magic
tech sky130A
magscale 1 2
timestamp 1733618896
<< viali >>
rect 1593 7497 1627 7531
rect 4169 7497 4203 7531
rect 5641 7497 5675 7531
rect 7757 7497 7791 7531
rect 9873 7497 9907 7531
rect 11989 7497 12023 7531
rect 14289 7497 14323 7531
rect 16221 7497 16255 7531
rect 18337 7497 18371 7531
rect 18705 7497 18739 7531
rect 20821 7497 20855 7531
rect 22569 7497 22603 7531
rect 23121 7497 23155 7531
rect 24869 7497 24903 7531
rect 27169 7497 27203 7531
rect 27537 7497 27571 7531
rect 29101 7497 29135 7531
rect 31033 7497 31067 7531
rect 33149 7497 33183 7531
rect 35265 7497 35299 7531
rect 37473 7497 37507 7531
rect 37841 7497 37875 7531
rect 40049 7497 40083 7531
rect 41613 7497 41647 7531
rect 43085 7497 43119 7531
rect 3893 7429 3927 7463
rect 18245 7429 18279 7463
rect 20361 7429 20395 7463
rect 27077 7429 27111 7463
rect 33057 7429 33091 7463
rect 1501 7361 1535 7395
rect 5549 7361 5583 7395
rect 7665 7361 7699 7395
rect 9781 7361 9815 7395
rect 11897 7361 11931 7395
rect 14197 7361 14231 7395
rect 16129 7361 16163 7395
rect 18889 7361 18923 7395
rect 20729 7361 20763 7395
rect 21005 7361 21039 7395
rect 22477 7361 22511 7395
rect 22937 7361 22971 7395
rect 24593 7361 24627 7395
rect 27721 7361 27755 7395
rect 28825 7361 28859 7395
rect 30941 7361 30975 7395
rect 35173 7361 35207 7395
rect 37381 7361 37415 7395
rect 38025 7361 38059 7395
rect 39957 7361 39991 7395
rect 41521 7361 41555 7395
rect 42809 7361 42843 7395
rect 22569 6885 22603 6919
rect 22753 6749 22787 6783
rect 24777 5865 24811 5899
rect 24961 5661 24995 5695
rect 16221 5321 16255 5355
rect 15945 5185 15979 5219
rect 16405 5185 16439 5219
rect 25421 3689 25455 3723
rect 27077 3689 27111 3723
rect 29009 3689 29043 3723
rect 33517 3689 33551 3723
rect 18153 3621 18187 3655
rect 18613 3621 18647 3655
rect 21465 3621 21499 3655
rect 25973 3621 26007 3655
rect 26525 3621 26559 3655
rect 27997 3621 28031 3655
rect 28273 3621 28307 3655
rect 18337 3485 18371 3519
rect 18429 3485 18463 3519
rect 18889 3485 18923 3519
rect 19441 3485 19475 3519
rect 19809 3485 19843 3519
rect 20085 3485 20119 3519
rect 20545 3485 20579 3519
rect 20821 3485 20855 3519
rect 21097 3485 21131 3519
rect 21373 3485 21407 3519
rect 21649 3485 21683 3519
rect 22477 3485 22511 3519
rect 22845 3485 22879 3519
rect 24225 3485 24259 3519
rect 24593 3485 24627 3519
rect 24869 3485 24903 3519
rect 25329 3485 25363 3519
rect 25605 3485 25639 3519
rect 25881 3485 25915 3519
rect 26157 3485 26191 3519
rect 26433 3485 26467 3519
rect 26709 3485 26743 3519
rect 26985 3485 27019 3519
rect 27261 3485 27295 3519
rect 27905 3485 27939 3519
rect 28181 3485 28215 3519
rect 28457 3485 28491 3519
rect 28733 3485 28767 3519
rect 29193 3485 29227 3519
rect 21833 3417 21867 3451
rect 32873 3417 32907 3451
rect 33425 3417 33459 3451
rect 18705 3349 18739 3383
rect 19257 3349 19291 3383
rect 19625 3349 19659 3383
rect 19901 3349 19935 3383
rect 20361 3349 20395 3383
rect 20637 3349 20671 3383
rect 20913 3349 20947 3383
rect 21189 3349 21223 3383
rect 21925 3349 21959 3383
rect 22293 3349 22327 3383
rect 22661 3349 22695 3383
rect 24041 3349 24075 3383
rect 24409 3349 24443 3383
rect 24685 3349 24719 3383
rect 25145 3349 25179 3383
rect 25697 3349 25731 3383
rect 26249 3349 26283 3383
rect 26801 3349 26835 3383
rect 27721 3349 27755 3383
rect 28549 3349 28583 3383
rect 32965 3349 32999 3383
rect 6745 3145 6779 3179
rect 14105 3145 14139 3179
rect 14657 3145 14691 3179
rect 15117 3145 15151 3179
rect 15393 3145 15427 3179
rect 15669 3145 15703 3179
rect 19165 3145 19199 3179
rect 19257 3145 19291 3179
rect 23397 3145 23431 3179
rect 29929 3145 29963 3179
rect 31585 3145 31619 3179
rect 32873 3145 32907 3179
rect 35633 3145 35667 3179
rect 38025 3145 38059 3179
rect 20177 3077 20211 3111
rect 20729 3077 20763 3111
rect 22385 3077 22419 3111
rect 22937 3077 22971 3111
rect 24041 3077 24075 3111
rect 25145 3077 25179 3111
rect 26249 3077 26283 3111
rect 27077 3077 27111 3111
rect 27629 3077 27663 3111
rect 28181 3077 28215 3111
rect 29837 3077 29871 3111
rect 31493 3077 31527 3111
rect 33885 3077 33919 3111
rect 34437 3077 34471 3111
rect 34989 3077 35023 3111
rect 35173 3077 35207 3111
rect 6561 3009 6595 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 14381 3009 14415 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 15209 3009 15243 3043
rect 15485 3009 15519 3043
rect 15945 3009 15979 3043
rect 16221 3009 16255 3043
rect 16497 3009 16531 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17509 3009 17543 3043
rect 17785 3009 17819 3043
rect 18061 3009 18095 3043
rect 18337 3009 18371 3043
rect 18613 3009 18647 3043
rect 18705 3009 18739 3043
rect 18981 3009 19015 3043
rect 19441 3009 19475 3043
rect 19625 3009 19659 3043
rect 21281 3009 21315 3043
rect 22201 3009 22235 3043
rect 23581 3009 23615 3043
rect 23857 3009 23891 3043
rect 24593 3009 24627 3043
rect 25697 3009 25731 3043
rect 28733 3009 28767 3043
rect 29285 3009 29319 3043
rect 30389 3009 30423 3043
rect 30941 3009 30975 3043
rect 32229 3009 32263 3043
rect 32781 3009 32815 3043
rect 33333 3009 33367 3043
rect 35357 3009 35391 3043
rect 35817 3009 35851 3043
rect 36093 3009 36127 3043
rect 36185 3009 36219 3043
rect 36461 3009 36495 3043
rect 37933 3009 37967 3043
rect 38209 3009 38243 3043
rect 39313 3009 39347 3043
rect 34161 2941 34195 2975
rect 13921 2873 13955 2907
rect 17049 2873 17083 2907
rect 18429 2873 18463 2907
rect 23673 2873 23707 2907
rect 36369 2873 36403 2907
rect 36645 2873 36679 2907
rect 37749 2873 37783 2907
rect 14565 2805 14599 2839
rect 15761 2805 15795 2839
rect 16037 2805 16071 2839
rect 16313 2805 16347 2839
rect 16773 2805 16807 2839
rect 17325 2805 17359 2839
rect 17601 2805 17635 2839
rect 17877 2805 17911 2839
rect 18153 2805 18187 2839
rect 18889 2805 18923 2839
rect 19717 2805 19751 2839
rect 20269 2805 20303 2839
rect 20821 2805 20855 2839
rect 21373 2805 21407 2839
rect 22017 2805 22051 2839
rect 22477 2805 22511 2839
rect 23029 2805 23063 2839
rect 24133 2805 24167 2839
rect 24685 2805 24719 2839
rect 25237 2805 25271 2839
rect 25789 2805 25823 2839
rect 26341 2805 26375 2839
rect 27169 2805 27203 2839
rect 27721 2805 27755 2839
rect 28273 2805 28307 2839
rect 29009 2805 29043 2839
rect 29377 2805 29411 2839
rect 30481 2805 30515 2839
rect 31033 2805 31067 2839
rect 32321 2805 32355 2839
rect 33425 2805 33459 2839
rect 34529 2805 34563 2839
rect 35449 2805 35483 2839
rect 35909 2805 35943 2839
rect 39129 2805 39163 2839
rect 5089 2601 5123 2635
rect 6193 2601 6227 2635
rect 8493 2601 8527 2635
rect 10793 2601 10827 2635
rect 11345 2601 11379 2635
rect 12817 2601 12851 2635
rect 14657 2601 14691 2635
rect 17509 2601 17543 2635
rect 18521 2601 18555 2635
rect 26249 2601 26283 2635
rect 26617 2601 26651 2635
rect 27721 2601 27755 2635
rect 29193 2601 29227 2635
rect 30849 2601 30883 2635
rect 31769 2601 31803 2635
rect 32321 2601 32355 2635
rect 34345 2601 34379 2635
rect 34897 2601 34931 2635
rect 35817 2601 35851 2635
rect 36185 2601 36219 2635
rect 37013 2601 37047 2635
rect 38025 2601 38059 2635
rect 38669 2601 38703 2635
rect 39865 2601 39899 2635
rect 40693 2601 40727 2635
rect 42441 2601 42475 2635
rect 5641 2533 5675 2567
rect 7665 2533 7699 2567
rect 9137 2533 9171 2567
rect 10241 2533 10275 2567
rect 10517 2533 10551 2567
rect 11069 2533 11103 2567
rect 11713 2533 11747 2567
rect 12265 2533 12299 2567
rect 14381 2533 14415 2567
rect 14933 2533 14967 2567
rect 16865 2533 16899 2567
rect 18061 2533 18095 2567
rect 23949 2533 23983 2567
rect 30389 2533 30423 2567
rect 36553 2533 36587 2567
rect 38945 2533 38979 2567
rect 39221 2533 39255 2567
rect 40141 2533 40175 2567
rect 40417 2533 40451 2567
rect 22661 2465 22695 2499
rect 25329 2465 25363 2499
rect 29009 2465 29043 2499
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 8033 2397 8067 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 8953 2397 8987 2431
rect 9229 2397 9263 2431
rect 9505 2397 9539 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 10885 2397 10919 2431
rect 11161 2397 11195 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13185 2397 13219 2431
rect 13461 2397 13495 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 14565 2397 14599 2431
rect 14841 2397 14875 2431
rect 15117 2397 15151 2431
rect 15209 2397 15243 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 16313 2397 16347 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 17233 2397 17267 2431
rect 17693 2397 17727 2431
rect 17785 2397 17819 2431
rect 18245 2397 18279 2431
rect 18337 2397 18371 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 20177 2397 20211 2431
rect 20729 2397 20763 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23489 2397 23523 2431
rect 24133 2397 24167 2431
rect 25053 2397 25087 2431
rect 26157 2397 26191 2431
rect 26801 2397 26835 2431
rect 29377 2397 29411 2431
rect 30205 2397 30239 2431
rect 30757 2397 30791 2431
rect 31953 2397 31987 2431
rect 33885 2397 33919 2431
rect 34529 2397 34563 2431
rect 35725 2397 35759 2431
rect 36001 2397 36035 2431
rect 36461 2397 36495 2431
rect 36737 2397 36771 2431
rect 36829 2397 36863 2431
rect 37289 2397 37323 2431
rect 37565 2397 37599 2431
rect 37841 2397 37875 2431
rect 38117 2397 38151 2431
rect 38577 2397 38611 2431
rect 38853 2397 38887 2431
rect 39129 2397 39163 2431
rect 39405 2397 39439 2431
rect 39681 2397 39715 2431
rect 40049 2397 40083 2431
rect 40325 2397 40359 2431
rect 40601 2397 40635 2431
rect 40877 2397 40911 2431
rect 42625 2397 42659 2431
rect 18705 2329 18739 2363
rect 19073 2329 19107 2363
rect 19993 2329 20027 2363
rect 20545 2329 20579 2363
rect 21097 2329 21131 2363
rect 21649 2329 21683 2363
rect 22385 2329 22419 2363
rect 24501 2329 24535 2363
rect 25605 2329 25639 2363
rect 27077 2329 27111 2363
rect 27629 2329 27663 2363
rect 28181 2329 28215 2363
rect 28733 2329 28767 2363
rect 29653 2329 29687 2363
rect 31309 2329 31343 2363
rect 32229 2329 32263 2363
rect 32781 2329 32815 2363
rect 33333 2329 33367 2363
rect 34805 2329 34839 2363
rect 35357 2329 35391 2363
rect 5365 2261 5399 2295
rect 5917 2261 5951 2295
rect 6561 2261 6595 2295
rect 6837 2261 6871 2295
rect 7113 2261 7147 2295
rect 7389 2261 7423 2295
rect 7941 2261 7975 2295
rect 8217 2261 8251 2295
rect 8769 2261 8803 2295
rect 9413 2261 9447 2295
rect 9689 2261 9723 2295
rect 9965 2261 9999 2295
rect 11989 2261 12023 2295
rect 12541 2261 12575 2295
rect 13093 2261 13127 2295
rect 13369 2261 13403 2295
rect 13645 2261 13679 2295
rect 13921 2261 13955 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 15669 2261 15703 2295
rect 15945 2261 15979 2295
rect 16221 2261 16255 2295
rect 16497 2261 16531 2295
rect 17141 2261 17175 2295
rect 17417 2261 17451 2295
rect 17969 2261 18003 2295
rect 19257 2261 19291 2295
rect 22017 2261 22051 2295
rect 23029 2261 23063 2295
rect 23581 2261 23615 2295
rect 24593 2261 24627 2295
rect 25697 2261 25731 2295
rect 27169 2261 27203 2295
rect 28273 2261 28307 2295
rect 29745 2261 29779 2295
rect 31401 2261 31435 2295
rect 32873 2261 32907 2295
rect 33425 2261 33459 2295
rect 33977 2261 34011 2295
rect 35449 2261 35483 2295
rect 36277 2261 36311 2295
rect 37473 2261 37507 2295
rect 37749 2261 37783 2295
rect 38301 2261 38335 2295
rect 38393 2261 38427 2295
rect 39497 2261 39531 2295
<< metal1 >>
rect 1104 7642 43675 7664
rect 1104 7590 11552 7642
rect 11604 7590 11616 7642
rect 11668 7590 11680 7642
rect 11732 7590 11744 7642
rect 11796 7590 11808 7642
rect 11860 7590 22155 7642
rect 22207 7590 22219 7642
rect 22271 7590 22283 7642
rect 22335 7590 22347 7642
rect 22399 7590 22411 7642
rect 22463 7590 32758 7642
rect 32810 7590 32822 7642
rect 32874 7590 32886 7642
rect 32938 7590 32950 7642
rect 33002 7590 33014 7642
rect 33066 7590 43361 7642
rect 43413 7590 43425 7642
rect 43477 7590 43489 7642
rect 43541 7590 43553 7642
rect 43605 7590 43617 7642
rect 43669 7590 43675 7642
rect 1104 7568 43675 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1581 7531 1639 7537
rect 1581 7528 1593 7531
rect 1176 7500 1593 7528
rect 1176 7488 1182 7500
rect 1581 7497 1593 7500
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 3476 7500 4169 7528
rect 3476 7488 3482 7500
rect 4157 7497 4169 7500
rect 4203 7497 4215 7531
rect 4157 7491 4215 7497
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 5408 7500 5641 7528
rect 5408 7488 5414 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7524 7500 7757 7528
rect 7524 7488 7530 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9732 7500 9873 7528
rect 9732 7488 9738 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 9861 7491 9919 7497
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 13872 7500 14289 7528
rect 13872 7488 13878 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15988 7500 16221 7528
rect 15988 7488 15994 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18104 7500 18337 7528
rect 18104 7488 18110 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7497 18751 7531
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 18693 7491 18751 7497
rect 20364 7500 20821 7528
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 18233 7463 18291 7469
rect 3927 7432 16574 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 6822 7392 6828 7404
rect 5583 7364 6828 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 9784 7256 9812 7355
rect 11900 7324 11928 7355
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16546 7392 16574 7432
rect 18233 7429 18245 7463
rect 18279 7460 18291 7463
rect 18708 7460 18736 7491
rect 20364 7469 20392 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 23109 7531 23167 7537
rect 23109 7497 23121 7531
rect 23155 7497 23167 7531
rect 23109 7491 23167 7497
rect 20349 7463 20407 7469
rect 18279 7432 18736 7460
rect 18800 7432 19840 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 18800 7392 18828 7432
rect 16546 7364 18828 7392
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 19812 7392 19840 7432
rect 20349 7429 20361 7463
rect 20395 7429 20407 7463
rect 23124 7460 23152 7491
rect 24854 7488 24860 7540
rect 24912 7488 24918 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 26568 7500 27169 7528
rect 26568 7488 26574 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 27157 7491 27215 7497
rect 27525 7531 27583 7537
rect 27525 7497 27537 7531
rect 27571 7497 27583 7531
rect 27525 7491 27583 7497
rect 20349 7423 20407 7429
rect 20456 7432 23152 7460
rect 27065 7463 27123 7469
rect 20456 7392 20484 7432
rect 27065 7429 27077 7463
rect 27111 7460 27123 7463
rect 27540 7460 27568 7491
rect 28810 7488 28816 7540
rect 28868 7528 28874 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 28868 7500 29101 7528
rect 28868 7488 28874 7500
rect 29089 7497 29101 7500
rect 29135 7497 29147 7531
rect 29089 7491 29147 7497
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 31021 7531 31079 7537
rect 31021 7528 31033 7531
rect 30800 7500 31033 7528
rect 30800 7488 30806 7500
rect 31021 7497 31033 7500
rect 31067 7497 31079 7531
rect 31021 7491 31079 7497
rect 33134 7488 33140 7540
rect 33192 7488 33198 7540
rect 34974 7488 34980 7540
rect 35032 7528 35038 7540
rect 35253 7531 35311 7537
rect 35253 7528 35265 7531
rect 35032 7500 35265 7528
rect 35032 7488 35038 7500
rect 35253 7497 35265 7500
rect 35299 7497 35311 7531
rect 35253 7491 35311 7497
rect 37182 7488 37188 7540
rect 37240 7528 37246 7540
rect 37461 7531 37519 7537
rect 37461 7528 37473 7531
rect 37240 7500 37473 7528
rect 37240 7488 37246 7500
rect 37461 7497 37473 7500
rect 37507 7497 37519 7531
rect 37461 7491 37519 7497
rect 37829 7531 37887 7537
rect 37829 7497 37841 7531
rect 37875 7497 37887 7531
rect 37829 7491 37887 7497
rect 27111 7432 27568 7460
rect 33045 7463 33103 7469
rect 27111 7429 27123 7432
rect 27065 7423 27123 7429
rect 33045 7429 33057 7463
rect 33091 7460 33103 7463
rect 37844 7460 37872 7491
rect 39298 7488 39304 7540
rect 39356 7528 39362 7540
rect 40037 7531 40095 7537
rect 40037 7528 40049 7531
rect 39356 7500 40049 7528
rect 39356 7488 39362 7500
rect 40037 7497 40049 7500
rect 40083 7497 40095 7531
rect 40037 7491 40095 7497
rect 41414 7488 41420 7540
rect 41472 7528 41478 7540
rect 41601 7531 41659 7537
rect 41601 7528 41613 7531
rect 41472 7500 41613 7528
rect 41472 7488 41478 7500
rect 41601 7497 41613 7500
rect 41647 7497 41659 7531
rect 41601 7491 41659 7497
rect 43073 7531 43131 7537
rect 43073 7497 43085 7531
rect 43119 7528 43131 7531
rect 43254 7528 43260 7540
rect 43119 7500 43260 7528
rect 43119 7497 43131 7500
rect 43073 7491 43131 7497
rect 43254 7488 43260 7500
rect 43312 7488 43318 7540
rect 33091 7432 37872 7460
rect 33091 7429 33103 7432
rect 33045 7423 33103 7429
rect 19812 7364 20484 7392
rect 20530 7352 20536 7404
rect 20588 7392 20594 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20588 7364 20729 7392
rect 20588 7352 20594 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20990 7352 20996 7404
rect 21048 7352 21054 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 22922 7352 22928 7404
rect 22980 7352 22986 7404
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7392 28871 7395
rect 29178 7392 29184 7404
rect 28859 7364 29184 7392
rect 28859 7361 28871 7364
rect 28813 7355 28871 7361
rect 20438 7324 20444 7336
rect 11900 7296 20444 7324
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 27724 7324 27752 7355
rect 29178 7352 29184 7364
rect 29236 7352 29242 7404
rect 30929 7395 30987 7401
rect 30929 7361 30941 7395
rect 30975 7392 30987 7395
rect 31754 7392 31760 7404
rect 30975 7364 31760 7392
rect 30975 7361 30987 7364
rect 30929 7355 30987 7361
rect 31754 7352 31760 7364
rect 31812 7352 31818 7404
rect 35161 7395 35219 7401
rect 35161 7361 35173 7395
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 33870 7324 33876 7336
rect 20640 7296 26234 7324
rect 27724 7296 33876 7324
rect 20640 7256 20668 7296
rect 9784 7228 20668 7256
rect 26206 7256 26234 7296
rect 33870 7284 33876 7296
rect 33928 7284 33934 7336
rect 35176 7324 35204 7355
rect 37366 7352 37372 7404
rect 37424 7352 37430 7404
rect 38013 7395 38071 7401
rect 38013 7361 38025 7395
rect 38059 7392 38071 7395
rect 38378 7392 38384 7404
rect 38059 7364 38384 7392
rect 38059 7361 38071 7364
rect 38013 7355 38071 7361
rect 38378 7352 38384 7364
rect 38436 7352 38442 7404
rect 39942 7352 39948 7404
rect 40000 7352 40006 7404
rect 41506 7352 41512 7404
rect 41564 7352 41570 7404
rect 42426 7352 42432 7404
rect 42484 7392 42490 7404
rect 42797 7395 42855 7401
rect 42797 7392 42809 7395
rect 42484 7364 42809 7392
rect 42484 7352 42490 7364
rect 42797 7361 42809 7364
rect 42843 7361 42855 7395
rect 42797 7355 42855 7361
rect 38654 7324 38660 7336
rect 35176 7296 38660 7324
rect 38654 7284 38660 7296
rect 38712 7284 38718 7336
rect 35710 7256 35716 7268
rect 26206 7228 35716 7256
rect 35710 7216 35716 7228
rect 35768 7216 35774 7268
rect 20530 7148 20536 7200
rect 20588 7188 20594 7200
rect 34790 7188 34796 7200
rect 20588 7160 34796 7188
rect 20588 7148 20594 7160
rect 34790 7148 34796 7160
rect 34848 7148 34854 7200
rect 1104 7098 43516 7120
rect 1104 7046 6251 7098
rect 6303 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 16854 7098
rect 16906 7046 16918 7098
rect 16970 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 27457 7098
rect 27509 7046 27521 7098
rect 27573 7046 27585 7098
rect 27637 7046 27649 7098
rect 27701 7046 27713 7098
rect 27765 7046 38060 7098
rect 38112 7046 38124 7098
rect 38176 7046 38188 7098
rect 38240 7046 38252 7098
rect 38304 7046 38316 7098
rect 38368 7046 43516 7098
rect 1104 7024 43516 7046
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 34422 6984 34428 6996
rect 7708 6956 34428 6984
rect 7708 6944 7714 6956
rect 34422 6944 34428 6956
rect 34480 6944 34486 6996
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 22557 6919 22615 6925
rect 22557 6916 22569 6919
rect 22520 6888 22569 6916
rect 22520 6876 22526 6888
rect 22557 6885 22569 6888
rect 22603 6885 22615 6919
rect 22557 6879 22615 6885
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6780 22799 6783
rect 23382 6780 23388 6792
rect 22787 6752 23388 6780
rect 22787 6749 22799 6752
rect 22741 6743 22799 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 1104 6554 43675 6576
rect 1104 6502 11552 6554
rect 11604 6502 11616 6554
rect 11668 6502 11680 6554
rect 11732 6502 11744 6554
rect 11796 6502 11808 6554
rect 11860 6502 22155 6554
rect 22207 6502 22219 6554
rect 22271 6502 22283 6554
rect 22335 6502 22347 6554
rect 22399 6502 22411 6554
rect 22463 6502 32758 6554
rect 32810 6502 32822 6554
rect 32874 6502 32886 6554
rect 32938 6502 32950 6554
rect 33002 6502 33014 6554
rect 33066 6502 43361 6554
rect 43413 6502 43425 6554
rect 43477 6502 43489 6554
rect 43541 6502 43553 6554
rect 43605 6502 43617 6554
rect 43669 6502 43675 6554
rect 1104 6480 43675 6502
rect 22922 6264 22928 6316
rect 22980 6304 22986 6316
rect 35986 6304 35992 6316
rect 22980 6276 35992 6304
rect 22980 6264 22986 6276
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 36630 6236 36636 6248
rect 18932 6208 36636 6236
rect 18932 6196 18938 6208
rect 36630 6196 36636 6208
rect 36688 6196 36694 6248
rect 1486 6128 1492 6180
rect 1544 6168 1550 6180
rect 33502 6168 33508 6180
rect 1544 6140 33508 6168
rect 1544 6128 1550 6140
rect 33502 6128 33508 6140
rect 33560 6128 33566 6180
rect 1104 6010 43516 6032
rect 1104 5958 6251 6010
rect 6303 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 16854 6010
rect 16906 5958 16918 6010
rect 16970 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 27457 6010
rect 27509 5958 27521 6010
rect 27573 5958 27585 6010
rect 27637 5958 27649 6010
rect 27701 5958 27713 6010
rect 27765 5958 38060 6010
rect 38112 5958 38124 6010
rect 38176 5958 38188 6010
rect 38240 5958 38252 6010
rect 38304 5958 38316 6010
rect 38368 5958 43516 6010
rect 1104 5936 43516 5958
rect 24578 5856 24584 5908
rect 24636 5896 24642 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 24636 5868 24777 5896
rect 24636 5856 24642 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5692 25007 5695
rect 37826 5692 37832 5704
rect 24995 5664 37832 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 1104 5466 43675 5488
rect 1104 5414 11552 5466
rect 11604 5414 11616 5466
rect 11668 5414 11680 5466
rect 11732 5414 11744 5466
rect 11796 5414 11808 5466
rect 11860 5414 22155 5466
rect 22207 5414 22219 5466
rect 22271 5414 22283 5466
rect 22335 5414 22347 5466
rect 22399 5414 22411 5466
rect 22463 5414 32758 5466
rect 32810 5414 32822 5466
rect 32874 5414 32886 5466
rect 32938 5414 32950 5466
rect 33002 5414 33014 5466
rect 33066 5414 43361 5466
rect 43413 5414 43425 5466
rect 43477 5414 43489 5466
rect 43541 5414 43553 5466
rect 43605 5414 43617 5466
rect 43669 5414 43675 5466
rect 1104 5392 43675 5414
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 16172 5324 16221 5352
rect 16172 5312 16178 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 16209 5315 16267 5321
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16393 5219 16451 5225
rect 16393 5216 16405 5219
rect 15979 5188 16405 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16393 5185 16405 5188
rect 16439 5216 16451 5219
rect 16439 5188 16528 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 16500 5160 16528 5188
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 1104 4922 43516 4944
rect 1104 4870 6251 4922
rect 6303 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 16854 4922
rect 16906 4870 16918 4922
rect 16970 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 27457 4922
rect 27509 4870 27521 4922
rect 27573 4870 27585 4922
rect 27637 4870 27649 4922
rect 27701 4870 27713 4922
rect 27765 4870 38060 4922
rect 38112 4870 38124 4922
rect 38176 4870 38188 4922
rect 38240 4870 38252 4922
rect 38304 4870 38316 4922
rect 38368 4870 43516 4922
rect 1104 4848 43516 4870
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 19426 4808 19432 4820
rect 10744 4780 19432 4808
rect 10744 4768 10750 4780
rect 19426 4768 19432 4780
rect 19484 4768 19490 4820
rect 8938 4700 8944 4752
rect 8996 4740 9002 4752
rect 24210 4740 24216 4752
rect 8996 4712 24216 4740
rect 8996 4700 9002 4712
rect 24210 4700 24216 4712
rect 24268 4700 24274 4752
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 23842 4672 23848 4684
rect 6788 4644 23848 4672
rect 6788 4632 6794 4644
rect 23842 4632 23848 4644
rect 23900 4632 23906 4684
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 22738 4604 22744 4616
rect 8812 4576 22744 4604
rect 8812 4564 8818 4576
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 15654 4496 15660 4548
rect 15712 4536 15718 4548
rect 33134 4536 33140 4548
rect 15712 4508 33140 4536
rect 15712 4496 15718 4508
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 28718 4468 28724 4480
rect 11020 4440 28724 4468
rect 11020 4428 11026 4440
rect 28718 4428 28724 4440
rect 28776 4428 28782 4480
rect 1104 4378 43675 4400
rect 1104 4326 11552 4378
rect 11604 4326 11616 4378
rect 11668 4326 11680 4378
rect 11732 4326 11744 4378
rect 11796 4326 11808 4378
rect 11860 4326 22155 4378
rect 22207 4326 22219 4378
rect 22271 4326 22283 4378
rect 22335 4326 22347 4378
rect 22399 4326 22411 4378
rect 22463 4326 32758 4378
rect 32810 4326 32822 4378
rect 32874 4326 32886 4378
rect 32938 4326 32950 4378
rect 33002 4326 33014 4378
rect 33066 4326 43361 4378
rect 43413 4326 43425 4378
rect 43477 4326 43489 4378
rect 43541 4326 43553 4378
rect 43605 4326 43617 4378
rect 43669 4326 43675 4378
rect 1104 4304 43675 4326
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 33962 4264 33968 4276
rect 15160 4236 33968 4264
rect 15160 4224 15166 4236
rect 33962 4224 33968 4236
rect 34020 4224 34026 4276
rect 14274 4156 14280 4208
rect 14332 4196 14338 4208
rect 36354 4196 36360 4208
rect 14332 4168 36360 4196
rect 14332 4156 14338 4168
rect 36354 4156 36360 4168
rect 36412 4156 36418 4208
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 24176 4032 28994 4060
rect 24176 4020 24182 4032
rect 17678 3952 17684 4004
rect 17736 3992 17742 4004
rect 25590 3992 25596 4004
rect 17736 3964 25596 3992
rect 17736 3952 17742 3964
rect 25590 3952 25596 3964
rect 25648 3952 25654 4004
rect 28966 3992 28994 4032
rect 30006 3992 30012 4004
rect 28966 3964 30012 3992
rect 30006 3952 30012 3964
rect 30064 3952 30070 4004
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 20070 3924 20076 3936
rect 11296 3896 20076 3924
rect 11296 3884 11302 3896
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 26418 3924 26424 3936
rect 22152 3896 26424 3924
rect 22152 3884 22158 3896
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 1104 3834 43516 3856
rect 1104 3782 6251 3834
rect 6303 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 16854 3834
rect 16906 3782 16918 3834
rect 16970 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 27457 3834
rect 27509 3782 27521 3834
rect 27573 3782 27585 3834
rect 27637 3782 27649 3834
rect 27701 3782 27713 3834
rect 27765 3782 38060 3834
rect 38112 3782 38124 3834
rect 38176 3782 38188 3834
rect 38240 3782 38252 3834
rect 38304 3782 38316 3834
rect 38368 3782 43516 3834
rect 1104 3760 43516 3782
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 20530 3720 20536 3732
rect 17460 3692 20536 3720
rect 17460 3680 17466 3692
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 21266 3680 21272 3732
rect 21324 3720 21330 3732
rect 25409 3723 25467 3729
rect 21324 3692 24900 3720
rect 21324 3680 21330 3692
rect 18141 3655 18199 3661
rect 18141 3621 18153 3655
rect 18187 3621 18199 3655
rect 18141 3615 18199 3621
rect 18601 3655 18659 3661
rect 18601 3621 18613 3655
rect 18647 3621 18659 3655
rect 18601 3615 18659 3621
rect 18156 3584 18184 3615
rect 18616 3584 18644 3615
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 20714 3652 20720 3664
rect 18840 3624 20720 3652
rect 18840 3612 18846 3624
rect 20714 3612 20720 3624
rect 20772 3612 20778 3664
rect 21453 3655 21511 3661
rect 21453 3621 21465 3655
rect 21499 3652 21511 3655
rect 22646 3652 22652 3664
rect 21499 3624 22652 3652
rect 21499 3621 21511 3624
rect 21453 3615 21511 3621
rect 22646 3612 22652 3624
rect 22704 3612 22710 3664
rect 24118 3584 24124 3596
rect 18156 3556 18460 3584
rect 18616 3556 24124 3584
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 18432 3525 18460 3556
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18104 3488 18337 3516
rect 18104 3476 18110 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 18656 3488 18889 3516
rect 18656 3476 18662 3488
rect 18877 3485 18889 3488
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 19794 3476 19800 3528
rect 19852 3476 19858 3528
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 20530 3476 20536 3528
rect 20588 3476 20594 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20680 3488 20821 3516
rect 20680 3476 20686 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 21085 3519 21143 3525
rect 21085 3516 21097 3519
rect 20956 3488 21097 3516
rect 20956 3476 20962 3488
rect 21085 3485 21097 3488
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 21361 3519 21419 3525
rect 21361 3485 21373 3519
rect 21407 3485 21419 3519
rect 21361 3479 21419 3485
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 21376 3448 21404 3479
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 21637 3519 21695 3525
rect 21637 3516 21649 3519
rect 21508 3488 21649 3516
rect 21508 3476 21514 3488
rect 21637 3485 21649 3488
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 22465 3519 22523 3525
rect 22465 3485 22477 3519
rect 22511 3485 22523 3519
rect 22465 3479 22523 3485
rect 17920 3420 21404 3448
rect 17920 3408 17926 3420
rect 21818 3408 21824 3460
rect 21876 3408 21882 3460
rect 22480 3448 22508 3479
rect 22830 3476 22836 3528
rect 22888 3476 22894 3528
rect 24210 3476 24216 3528
rect 24268 3476 24274 3528
rect 24872 3525 24900 3692
rect 25409 3689 25421 3723
rect 25455 3720 25467 3723
rect 26234 3720 26240 3732
rect 25455 3692 26240 3720
rect 25455 3689 25467 3692
rect 25409 3683 25467 3689
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 27065 3723 27123 3729
rect 27065 3689 27077 3723
rect 27111 3720 27123 3723
rect 28350 3720 28356 3732
rect 27111 3692 28356 3720
rect 27111 3689 27123 3692
rect 27065 3683 27123 3689
rect 28350 3680 28356 3692
rect 28408 3680 28414 3732
rect 28997 3723 29055 3729
rect 28997 3689 29009 3723
rect 29043 3720 29055 3723
rect 29178 3720 29184 3732
rect 29043 3692 29184 3720
rect 29043 3689 29055 3692
rect 28997 3683 29055 3689
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 33502 3680 33508 3732
rect 33560 3680 33566 3732
rect 25961 3655 26019 3661
rect 25961 3621 25973 3655
rect 26007 3652 26019 3655
rect 26513 3655 26571 3661
rect 26007 3624 26464 3652
rect 26007 3621 26019 3624
rect 25961 3615 26019 3621
rect 26436 3584 26464 3624
rect 26513 3621 26525 3655
rect 26559 3652 26571 3655
rect 27798 3652 27804 3664
rect 26559 3624 27804 3652
rect 26559 3621 26571 3624
rect 26513 3615 26571 3621
rect 27798 3612 27804 3624
rect 27856 3612 27862 3664
rect 27985 3655 28043 3661
rect 27985 3621 27997 3655
rect 28031 3621 28043 3655
rect 27985 3615 28043 3621
rect 28261 3655 28319 3661
rect 28261 3621 28273 3655
rect 28307 3652 28319 3655
rect 29730 3652 29736 3664
rect 28307 3624 29736 3652
rect 28307 3621 28319 3624
rect 28261 3615 28319 3621
rect 27614 3584 27620 3596
rect 26436 3556 27620 3584
rect 27614 3544 27620 3556
rect 27672 3544 27678 3596
rect 28000 3584 28028 3615
rect 29730 3612 29736 3624
rect 29788 3612 29794 3664
rect 29270 3584 29276 3596
rect 28000 3556 29276 3584
rect 29270 3544 29276 3556
rect 29328 3544 29334 3596
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 22922 3448 22928 3460
rect 22480 3420 22928 3448
rect 22922 3408 22928 3420
rect 22980 3408 22986 3460
rect 23106 3408 23112 3460
rect 23164 3448 23170 3460
rect 24596 3448 24624 3479
rect 25314 3476 25320 3528
rect 25372 3476 25378 3528
rect 25590 3476 25596 3528
rect 25648 3476 25654 3528
rect 25682 3476 25688 3528
rect 25740 3516 25746 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25740 3488 25881 3516
rect 25740 3476 25746 3488
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 25869 3479 25927 3485
rect 26142 3476 26148 3528
rect 26200 3476 26206 3528
rect 26418 3476 26424 3528
rect 26476 3476 26482 3528
rect 26694 3476 26700 3528
rect 26752 3476 26758 3528
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 27246 3476 27252 3528
rect 27304 3476 27310 3528
rect 27890 3476 27896 3528
rect 27948 3476 27954 3528
rect 28166 3476 28172 3528
rect 28224 3476 28230 3528
rect 28442 3476 28448 3528
rect 28500 3476 28506 3528
rect 28718 3476 28724 3528
rect 28776 3476 28782 3528
rect 29181 3519 29239 3525
rect 29181 3485 29193 3519
rect 29227 3516 29239 3519
rect 36262 3516 36268 3528
rect 29227 3488 36268 3516
rect 29227 3485 29239 3488
rect 29181 3479 29239 3485
rect 36262 3476 36268 3488
rect 36320 3476 36326 3528
rect 26326 3448 26332 3460
rect 23164 3420 24624 3448
rect 25700 3420 26332 3448
rect 23164 3408 23170 3420
rect 18690 3340 18696 3392
rect 18748 3340 18754 3392
rect 19245 3383 19303 3389
rect 19245 3349 19257 3383
rect 19291 3380 19303 3383
rect 19518 3380 19524 3392
rect 19291 3352 19524 3380
rect 19291 3349 19303 3352
rect 19245 3343 19303 3349
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 19610 3340 19616 3392
rect 19668 3340 19674 3392
rect 19886 3340 19892 3392
rect 19944 3340 19950 3392
rect 20346 3340 20352 3392
rect 20404 3340 20410 3392
rect 20622 3340 20628 3392
rect 20680 3340 20686 3392
rect 20898 3340 20904 3392
rect 20956 3340 20962 3392
rect 21174 3340 21180 3392
rect 21232 3340 21238 3392
rect 21634 3340 21640 3392
rect 21692 3380 21698 3392
rect 21913 3383 21971 3389
rect 21913 3380 21925 3383
rect 21692 3352 21925 3380
rect 21692 3340 21698 3352
rect 21913 3349 21925 3352
rect 21959 3349 21971 3383
rect 21913 3343 21971 3349
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 22554 3380 22560 3392
rect 22327 3352 22560 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 22649 3383 22707 3389
rect 22649 3349 22661 3383
rect 22695 3380 22707 3383
rect 23474 3380 23480 3392
rect 22695 3352 23480 3380
rect 22695 3349 22707 3352
rect 22649 3343 22707 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 24029 3383 24087 3389
rect 24029 3349 24041 3383
rect 24075 3380 24087 3383
rect 24302 3380 24308 3392
rect 24075 3352 24308 3380
rect 24075 3349 24087 3352
rect 24029 3343 24087 3349
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 24394 3340 24400 3392
rect 24452 3340 24458 3392
rect 24673 3383 24731 3389
rect 24673 3349 24685 3383
rect 24719 3380 24731 3383
rect 25038 3380 25044 3392
rect 24719 3352 25044 3380
rect 24719 3349 24731 3352
rect 24673 3343 24731 3349
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 25133 3383 25191 3389
rect 25133 3349 25145 3383
rect 25179 3380 25191 3383
rect 25314 3380 25320 3392
rect 25179 3352 25320 3380
rect 25179 3349 25191 3352
rect 25133 3343 25191 3349
rect 25314 3340 25320 3352
rect 25372 3340 25378 3392
rect 25700 3389 25728 3420
rect 26326 3408 26332 3420
rect 26384 3408 26390 3460
rect 28074 3448 28080 3460
rect 26804 3420 28080 3448
rect 25685 3383 25743 3389
rect 25685 3349 25697 3383
rect 25731 3349 25743 3383
rect 25685 3343 25743 3349
rect 26237 3383 26295 3389
rect 26237 3349 26249 3383
rect 26283 3380 26295 3383
rect 26418 3380 26424 3392
rect 26283 3352 26424 3380
rect 26283 3349 26295 3352
rect 26237 3343 26295 3349
rect 26418 3340 26424 3352
rect 26476 3340 26482 3392
rect 26804 3389 26832 3420
rect 28074 3408 28080 3420
rect 28132 3408 28138 3460
rect 28994 3448 29000 3460
rect 28460 3420 29000 3448
rect 26789 3383 26847 3389
rect 26789 3349 26801 3383
rect 26835 3349 26847 3383
rect 26789 3343 26847 3349
rect 27709 3383 27767 3389
rect 27709 3349 27721 3383
rect 27755 3380 27767 3383
rect 28460 3380 28488 3420
rect 28994 3408 29000 3420
rect 29052 3408 29058 3460
rect 32030 3408 32036 3460
rect 32088 3448 32094 3460
rect 32861 3451 32919 3457
rect 32861 3448 32873 3451
rect 32088 3420 32873 3448
rect 32088 3408 32094 3420
rect 32861 3417 32873 3420
rect 32907 3417 32919 3451
rect 32861 3411 32919 3417
rect 33410 3408 33416 3460
rect 33468 3408 33474 3460
rect 27755 3352 28488 3380
rect 27755 3349 27767 3352
rect 27709 3343 27767 3349
rect 28534 3340 28540 3392
rect 28592 3340 28598 3392
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 32953 3383 33011 3389
rect 32953 3380 32965 3383
rect 32732 3352 32965 3380
rect 32732 3340 32738 3352
rect 32953 3349 32965 3352
rect 32999 3349 33011 3383
rect 32953 3343 33011 3349
rect 34698 3340 34704 3392
rect 34756 3380 34762 3392
rect 35802 3380 35808 3392
rect 34756 3352 35808 3380
rect 34756 3340 34762 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 1104 3290 43675 3312
rect 1104 3238 11552 3290
rect 11604 3238 11616 3290
rect 11668 3238 11680 3290
rect 11732 3238 11744 3290
rect 11796 3238 11808 3290
rect 11860 3238 22155 3290
rect 22207 3238 22219 3290
rect 22271 3238 22283 3290
rect 22335 3238 22347 3290
rect 22399 3238 22411 3290
rect 22463 3238 32758 3290
rect 32810 3238 32822 3290
rect 32874 3238 32886 3290
rect 32938 3238 32950 3290
rect 33002 3238 33014 3290
rect 33066 3238 43361 3290
rect 43413 3238 43425 3290
rect 43477 3238 43489 3290
rect 43541 3238 43553 3290
rect 43605 3238 43617 3290
rect 43669 3238 43675 3290
rect 1104 3216 43675 3238
rect 6730 3136 6736 3188
rect 6788 3136 6794 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14182 3176 14188 3188
rect 14139 3148 14188 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14645 3179 14703 3185
rect 14645 3145 14657 3179
rect 14691 3145 14703 3179
rect 14645 3139 14703 3145
rect 14660 3108 14688 3139
rect 15102 3136 15108 3188
rect 15160 3136 15166 3188
rect 15378 3136 15384 3188
rect 15436 3136 15442 3188
rect 15654 3136 15660 3188
rect 15712 3136 15718 3188
rect 18690 3136 18696 3188
rect 18748 3136 18754 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 19076 3148 19165 3176
rect 14660 3080 14964 3108
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 14936 3049 14964 3080
rect 15010 3068 15016 3120
rect 15068 3108 15074 3120
rect 15068 3080 18644 3108
rect 15068 3068 15074 3080
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15194 3000 15200 3052
rect 15252 3000 15258 3052
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 15488 2972 15516 3003
rect 15930 3000 15936 3052
rect 15988 3000 15994 3052
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3040 16543 3043
rect 16574 3040 16580 3052
rect 16531 3012 16580 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 17218 3000 17224 3052
rect 17276 3000 17282 3052
rect 17494 3000 17500 3052
rect 17552 3000 17558 3052
rect 17678 3000 17684 3052
rect 17736 3000 17742 3052
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 18616 3049 18644 3080
rect 18708 3049 18736 3136
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 17696 2972 17724 3000
rect 14700 2944 15516 2972
rect 16546 2944 17724 2972
rect 18340 2972 18368 3003
rect 18966 3000 18972 3052
rect 19024 3000 19030 3052
rect 19076 3040 19104 3148
rect 19153 3145 19165 3148
rect 19199 3145 19211 3179
rect 19153 3139 19211 3145
rect 19242 3136 19248 3188
rect 19300 3136 19306 3188
rect 19518 3136 19524 3188
rect 19576 3136 19582 3188
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 19944 3148 20760 3176
rect 19944 3136 19950 3148
rect 19536 3108 19564 3136
rect 20165 3111 20223 3117
rect 20165 3108 20177 3111
rect 19536 3080 20177 3108
rect 20165 3077 20177 3080
rect 20211 3077 20223 3111
rect 20165 3071 20223 3077
rect 20346 3068 20352 3120
rect 20404 3068 20410 3120
rect 20732 3117 20760 3148
rect 21174 3136 21180 3188
rect 21232 3176 21238 3188
rect 21232 3148 22416 3176
rect 21232 3136 21238 3148
rect 22388 3117 22416 3148
rect 22554 3136 22560 3188
rect 22612 3136 22618 3188
rect 23385 3179 23443 3185
rect 23385 3145 23397 3179
rect 23431 3176 23443 3179
rect 23431 3148 24072 3176
rect 23431 3145 23443 3148
rect 23385 3139 23443 3145
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3077 20775 3111
rect 20717 3071 20775 3077
rect 22373 3111 22431 3117
rect 22373 3077 22385 3111
rect 22419 3077 22431 3111
rect 22572 3108 22600 3136
rect 24044 3117 24072 3148
rect 24394 3136 24400 3188
rect 24452 3176 24458 3188
rect 24452 3148 25176 3176
rect 24452 3136 24458 3148
rect 25148 3117 25176 3148
rect 25314 3136 25320 3188
rect 25372 3136 25378 3188
rect 26326 3136 26332 3188
rect 26384 3136 26390 3188
rect 26418 3136 26424 3188
rect 26476 3176 26482 3188
rect 26476 3148 27660 3176
rect 26476 3136 26482 3148
rect 22925 3111 22983 3117
rect 22925 3108 22937 3111
rect 22572 3080 22937 3108
rect 22373 3071 22431 3077
rect 22925 3077 22937 3080
rect 22971 3077 22983 3111
rect 22925 3071 22983 3077
rect 24029 3111 24087 3117
rect 24029 3077 24041 3111
rect 24075 3077 24087 3111
rect 24029 3071 24087 3077
rect 25133 3111 25191 3117
rect 25133 3077 25145 3111
rect 25179 3077 25191 3111
rect 25332 3108 25360 3136
rect 26237 3111 26295 3117
rect 26237 3108 26249 3111
rect 25332 3080 26249 3108
rect 25133 3071 25191 3077
rect 26237 3077 26249 3080
rect 26283 3077 26295 3111
rect 26344 3108 26372 3136
rect 27632 3117 27660 3148
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 28132 3148 28212 3176
rect 28132 3136 28138 3148
rect 28184 3117 28212 3148
rect 28534 3136 28540 3188
rect 28592 3136 28598 3188
rect 29086 3136 29092 3188
rect 29144 3176 29150 3188
rect 29917 3179 29975 3185
rect 29917 3176 29929 3179
rect 29144 3148 29929 3176
rect 29144 3136 29150 3148
rect 29917 3145 29929 3148
rect 29963 3145 29975 3179
rect 29917 3139 29975 3145
rect 30006 3136 30012 3188
rect 30064 3136 30070 3188
rect 30650 3136 30656 3188
rect 30708 3176 30714 3188
rect 31573 3179 31631 3185
rect 31573 3176 31585 3179
rect 30708 3148 31585 3176
rect 30708 3136 30714 3148
rect 31573 3145 31585 3148
rect 31619 3145 31631 3179
rect 31573 3139 31631 3145
rect 31846 3136 31852 3188
rect 31904 3176 31910 3188
rect 32861 3179 32919 3185
rect 32861 3176 32873 3179
rect 31904 3148 32873 3176
rect 31904 3136 31910 3148
rect 32861 3145 32873 3148
rect 32907 3145 32919 3179
rect 35621 3179 35679 3185
rect 35621 3176 35633 3179
rect 32861 3139 32919 3145
rect 34992 3148 35633 3176
rect 27065 3111 27123 3117
rect 27065 3108 27077 3111
rect 26344 3080 27077 3108
rect 26237 3071 26295 3077
rect 27065 3077 27077 3080
rect 27111 3077 27123 3111
rect 27065 3071 27123 3077
rect 27617 3111 27675 3117
rect 27617 3077 27629 3111
rect 27663 3077 27675 3111
rect 27617 3071 27675 3077
rect 28169 3111 28227 3117
rect 28169 3077 28181 3111
rect 28215 3077 28227 3111
rect 28552 3108 28580 3136
rect 29825 3111 29883 3117
rect 29825 3108 29837 3111
rect 28552 3080 29837 3108
rect 28169 3071 28227 3077
rect 29825 3077 29837 3080
rect 29871 3077 29883 3111
rect 30024 3108 30052 3136
rect 31481 3111 31539 3117
rect 31481 3108 31493 3111
rect 30024 3080 31493 3108
rect 29825 3071 29883 3077
rect 31481 3077 31493 3080
rect 31527 3077 31539 3111
rect 31481 3071 31539 3077
rect 33134 3068 33140 3120
rect 33192 3108 33198 3120
rect 33873 3111 33931 3117
rect 33873 3108 33885 3111
rect 33192 3080 33885 3108
rect 33192 3068 33198 3080
rect 33873 3077 33885 3080
rect 33919 3077 33931 3111
rect 33873 3071 33931 3077
rect 33962 3068 33968 3120
rect 34020 3108 34026 3120
rect 34992 3117 35020 3148
rect 35621 3145 35633 3148
rect 35667 3145 35679 3179
rect 35621 3139 35679 3145
rect 35802 3136 35808 3188
rect 35860 3176 35866 3188
rect 38013 3179 38071 3185
rect 38013 3176 38025 3179
rect 35860 3148 38025 3176
rect 35860 3136 35866 3148
rect 38013 3145 38025 3148
rect 38059 3145 38071 3179
rect 38013 3139 38071 3145
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 34020 3080 34437 3108
rect 34020 3068 34026 3080
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 34977 3111 35035 3117
rect 34977 3077 34989 3111
rect 35023 3077 35035 3111
rect 34977 3071 35035 3077
rect 35161 3111 35219 3117
rect 35161 3077 35173 3111
rect 35207 3077 35219 3111
rect 35161 3071 35219 3077
rect 19334 3040 19340 3052
rect 19076 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3009 19487 3043
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19429 3003 19487 3009
rect 19536 3012 19625 3040
rect 18874 2972 18880 2984
rect 18340 2944 18880 2972
rect 14700 2932 14706 2944
rect 13909 2907 13967 2913
rect 13909 2873 13921 2907
rect 13955 2904 13967 2907
rect 16546 2904 16574 2944
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19444 2972 19472 3003
rect 19116 2944 19472 2972
rect 19116 2932 19122 2944
rect 13955 2876 16574 2904
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 16666 2864 16672 2916
rect 16724 2904 16730 2916
rect 17037 2907 17095 2913
rect 17037 2904 17049 2907
rect 16724 2876 17049 2904
rect 16724 2864 16730 2876
rect 17037 2873 17049 2876
rect 17083 2873 17095 2907
rect 17037 2867 17095 2873
rect 18417 2907 18475 2913
rect 18417 2873 18429 2907
rect 18463 2904 18475 2907
rect 19536 2904 19564 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 20364 3040 20392 3068
rect 21269 3043 21327 3049
rect 21269 3040 21281 3043
rect 20364 3012 21281 3040
rect 19613 3003 19671 3009
rect 21269 3009 21281 3012
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22738 3040 22744 3052
rect 22235 3012 22744 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 23842 3000 23848 3052
rect 23900 3000 23906 3052
rect 24581 3043 24639 3049
rect 24581 3009 24593 3043
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 25685 3043 25743 3049
rect 25685 3009 25697 3043
rect 25731 3009 25743 3043
rect 25685 3003 25743 3009
rect 24596 2972 24624 3003
rect 22112 2944 23612 2972
rect 22112 2904 22140 2944
rect 18463 2876 19564 2904
rect 19628 2876 22140 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 14553 2839 14611 2845
rect 14553 2805 14565 2839
rect 14599 2836 14611 2839
rect 15010 2836 15016 2848
rect 14599 2808 15016 2836
rect 14599 2805 14611 2808
rect 14553 2799 14611 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15746 2796 15752 2848
rect 15804 2796 15810 2848
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 15896 2808 16037 2836
rect 15896 2796 15902 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16301 2839 16359 2845
rect 16301 2836 16313 2839
rect 16172 2808 16313 2836
rect 16172 2796 16178 2808
rect 16301 2805 16313 2808
rect 16347 2805 16359 2839
rect 16301 2799 16359 2805
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 16448 2808 16773 2836
rect 16448 2796 16454 2808
rect 16761 2805 16773 2808
rect 16807 2805 16819 2839
rect 16761 2799 16819 2805
rect 17310 2796 17316 2848
rect 17368 2796 17374 2848
rect 17586 2796 17592 2848
rect 17644 2796 17650 2848
rect 17862 2796 17868 2848
rect 17920 2796 17926 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 18322 2836 18328 2848
rect 18187 2808 18328 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 18877 2839 18935 2845
rect 18877 2805 18889 2839
rect 18923 2836 18935 2839
rect 19628 2836 19656 2876
rect 22186 2864 22192 2916
rect 22244 2904 22250 2916
rect 22244 2876 22508 2904
rect 22244 2864 22250 2876
rect 18923 2808 19656 2836
rect 18923 2805 18935 2808
rect 18877 2799 18935 2805
rect 19702 2796 19708 2848
rect 19760 2796 19766 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 20036 2808 20269 2836
rect 20036 2796 20042 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20257 2799 20315 2805
rect 20530 2796 20536 2848
rect 20588 2836 20594 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20588 2808 20821 2836
rect 20588 2796 20594 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 21140 2808 21373 2836
rect 21140 2796 21146 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21361 2799 21419 2805
rect 22005 2839 22063 2845
rect 22005 2805 22017 2839
rect 22051 2836 22063 2839
rect 22278 2836 22284 2848
rect 22051 2808 22284 2836
rect 22051 2805 22063 2808
rect 22005 2799 22063 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 22480 2845 22508 2876
rect 22465 2839 22523 2845
rect 22465 2805 22477 2839
rect 22511 2805 22523 2839
rect 22465 2799 22523 2805
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 23017 2839 23075 2845
rect 23017 2836 23029 2839
rect 22796 2808 23029 2836
rect 22796 2796 22802 2808
rect 23017 2805 23029 2808
rect 23063 2805 23075 2839
rect 23584 2836 23612 2944
rect 23676 2944 24624 2972
rect 25700 2972 25728 3003
rect 28718 3000 28724 3052
rect 28776 3000 28782 3052
rect 29270 3000 29276 3052
rect 29328 3000 29334 3052
rect 29362 3000 29368 3052
rect 29420 3040 29426 3052
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 29420 3012 30389 3040
rect 29420 3000 29426 3012
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30524 3012 30941 3040
rect 30524 3000 30530 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 31938 3000 31944 3052
rect 31996 3040 32002 3052
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 31996 3012 32229 3040
rect 31996 3000 32002 3012
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 32217 3003 32275 3009
rect 32766 3000 32772 3052
rect 32824 3000 32830 3052
rect 33321 3043 33379 3049
rect 33321 3009 33333 3043
rect 33367 3040 33379 3043
rect 33686 3040 33692 3052
rect 33367 3012 33692 3040
rect 33367 3009 33379 3012
rect 33321 3003 33379 3009
rect 33686 3000 33692 3012
rect 33744 3000 33750 3052
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 35176 3040 35204 3071
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 35492 3080 36124 3108
rect 35492 3068 35498 3080
rect 34572 3012 35204 3040
rect 35345 3043 35403 3049
rect 34572 3000 34578 3012
rect 35345 3009 35357 3043
rect 35391 3040 35403 3043
rect 35526 3040 35532 3052
rect 35391 3012 35532 3040
rect 35391 3009 35403 3012
rect 35345 3003 35403 3009
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 36096 3049 36124 3080
rect 36262 3068 36268 3120
rect 36320 3068 36326 3120
rect 35805 3043 35863 3049
rect 35805 3040 35817 3043
rect 35636 3012 35817 3040
rect 26602 2972 26608 2984
rect 25700 2944 26608 2972
rect 23676 2913 23704 2944
rect 26602 2932 26608 2944
rect 26660 2932 26666 2984
rect 27614 2932 27620 2984
rect 27672 2972 27678 2984
rect 27672 2944 27936 2972
rect 27672 2932 27678 2944
rect 23661 2907 23719 2913
rect 23661 2873 23673 2907
rect 23707 2873 23719 2907
rect 24854 2904 24860 2916
rect 23661 2867 23719 2873
rect 23768 2876 24860 2904
rect 23768 2836 23796 2876
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 25406 2864 25412 2916
rect 25464 2904 25470 2916
rect 26142 2904 26148 2916
rect 25464 2876 26148 2904
rect 25464 2864 25470 2876
rect 26142 2864 26148 2876
rect 26200 2864 26206 2916
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 27908 2904 27936 2944
rect 33042 2932 33048 2984
rect 33100 2972 33106 2984
rect 34149 2975 34207 2981
rect 34149 2972 34161 2975
rect 33100 2944 34161 2972
rect 33100 2932 33106 2944
rect 34149 2941 34161 2944
rect 34195 2941 34207 2975
rect 34149 2935 34207 2941
rect 34882 2932 34888 2984
rect 34940 2972 34946 2984
rect 35636 2972 35664 3012
rect 35805 3009 35817 3012
rect 35851 3009 35863 3043
rect 35805 3003 35863 3009
rect 36081 3043 36139 3049
rect 36081 3009 36093 3043
rect 36127 3009 36139 3043
rect 36081 3003 36139 3009
rect 36173 3043 36231 3049
rect 36173 3009 36185 3043
rect 36219 3009 36231 3043
rect 36173 3003 36231 3009
rect 34940 2944 35664 2972
rect 34940 2932 34946 2944
rect 35710 2932 35716 2984
rect 35768 2972 35774 2984
rect 36188 2972 36216 3003
rect 35768 2944 36216 2972
rect 36280 2972 36308 3068
rect 36446 3000 36452 3052
rect 36504 3000 36510 3052
rect 37642 3000 37648 3052
rect 37700 3040 37706 3052
rect 37921 3043 37979 3049
rect 37921 3040 37933 3043
rect 37700 3012 37933 3040
rect 37700 3000 37706 3012
rect 37921 3009 37933 3012
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38010 3000 38016 3052
rect 38068 3040 38074 3052
rect 38197 3043 38255 3049
rect 38197 3040 38209 3043
rect 38068 3012 38209 3040
rect 38068 3000 38074 3012
rect 38197 3009 38209 3012
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 39022 3000 39028 3052
rect 39080 3040 39086 3052
rect 39301 3043 39359 3049
rect 39301 3040 39313 3043
rect 39080 3012 39313 3040
rect 39080 3000 39086 3012
rect 39301 3009 39313 3012
rect 39347 3009 39359 3043
rect 39301 3003 39359 3009
rect 36280 2944 37780 2972
rect 35768 2932 35774 2944
rect 27982 2904 27988 2916
rect 26936 2876 27752 2904
rect 27908 2876 27988 2904
rect 26936 2864 26942 2876
rect 23584 2808 23796 2836
rect 23017 2799 23075 2805
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23900 2808 24133 2836
rect 23900 2796 23906 2808
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24121 2799 24179 2805
rect 24394 2796 24400 2848
rect 24452 2836 24458 2848
rect 24673 2839 24731 2845
rect 24673 2836 24685 2839
rect 24452 2808 24685 2836
rect 24452 2796 24458 2808
rect 24673 2805 24685 2808
rect 24719 2805 24731 2839
rect 24673 2799 24731 2805
rect 24946 2796 24952 2848
rect 25004 2836 25010 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 25004 2808 25237 2836
rect 25004 2796 25010 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 25498 2796 25504 2848
rect 25556 2836 25562 2848
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25556 2808 25789 2836
rect 25556 2796 25562 2808
rect 25777 2805 25789 2808
rect 25823 2805 25835 2839
rect 25777 2799 25835 2805
rect 25958 2796 25964 2848
rect 26016 2836 26022 2848
rect 26329 2839 26387 2845
rect 26329 2836 26341 2839
rect 26016 2808 26341 2836
rect 26016 2796 26022 2808
rect 26329 2805 26341 2808
rect 26375 2805 26387 2839
rect 26329 2799 26387 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 27724 2845 27752 2876
rect 27982 2864 27988 2876
rect 28040 2864 28046 2916
rect 28534 2864 28540 2916
rect 28592 2904 28598 2916
rect 28592 2876 29408 2904
rect 28592 2864 28598 2876
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 26568 2808 27169 2836
rect 26568 2796 26574 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 27157 2799 27215 2805
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 27798 2796 27804 2848
rect 27856 2836 27862 2848
rect 28261 2839 28319 2845
rect 28261 2836 28273 2839
rect 27856 2808 28273 2836
rect 27856 2796 27862 2808
rect 28261 2805 28273 2808
rect 28307 2805 28319 2839
rect 28261 2799 28319 2805
rect 28810 2796 28816 2848
rect 28868 2836 28874 2848
rect 29380 2845 29408 2876
rect 30190 2864 30196 2916
rect 30248 2904 30254 2916
rect 30248 2876 31064 2904
rect 30248 2864 30254 2876
rect 28997 2839 29055 2845
rect 28997 2836 29009 2839
rect 28868 2808 29009 2836
rect 28868 2796 28874 2808
rect 28997 2805 29009 2808
rect 29043 2805 29055 2839
rect 28997 2799 29055 2805
rect 29365 2839 29423 2845
rect 29365 2805 29377 2839
rect 29411 2805 29423 2839
rect 29365 2799 29423 2805
rect 29822 2796 29828 2848
rect 29880 2836 29886 2848
rect 31036 2845 31064 2876
rect 31294 2864 31300 2916
rect 31352 2904 31358 2916
rect 31352 2876 31754 2904
rect 31352 2864 31358 2876
rect 30469 2839 30527 2845
rect 30469 2836 30481 2839
rect 29880 2808 30481 2836
rect 29880 2796 29886 2808
rect 30469 2805 30481 2808
rect 30515 2805 30527 2839
rect 30469 2799 30527 2805
rect 31021 2839 31079 2845
rect 31021 2805 31033 2839
rect 31067 2805 31079 2839
rect 31726 2836 31754 2876
rect 32398 2864 32404 2916
rect 32456 2904 32462 2916
rect 32456 2876 33456 2904
rect 32456 2864 32462 2876
rect 33428 2845 33456 2876
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 33560 2876 34560 2904
rect 33560 2864 33566 2876
rect 34532 2845 34560 2876
rect 34606 2864 34612 2916
rect 34664 2904 34670 2916
rect 36170 2904 36176 2916
rect 34664 2876 36176 2904
rect 34664 2864 34670 2876
rect 36170 2864 36176 2876
rect 36228 2864 36234 2916
rect 36354 2864 36360 2916
rect 36412 2864 36418 2916
rect 36630 2864 36636 2916
rect 36688 2864 36694 2916
rect 37752 2913 37780 2944
rect 37737 2907 37795 2913
rect 37737 2873 37749 2907
rect 37783 2873 37795 2907
rect 37737 2867 37795 2873
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 31726 2808 32321 2836
rect 31021 2799 31079 2805
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 33413 2839 33471 2845
rect 33413 2805 33425 2839
rect 33459 2805 33471 2839
rect 33413 2799 33471 2805
rect 34517 2839 34575 2845
rect 34517 2805 34529 2839
rect 34563 2805 34575 2839
rect 34517 2799 34575 2805
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 35437 2839 35495 2845
rect 35437 2836 35449 2839
rect 34848 2808 35449 2836
rect 34848 2796 34854 2808
rect 35437 2805 35449 2808
rect 35483 2805 35495 2839
rect 35437 2799 35495 2805
rect 35894 2796 35900 2848
rect 35952 2796 35958 2848
rect 39117 2839 39175 2845
rect 39117 2805 39129 2839
rect 39163 2836 39175 2839
rect 40034 2836 40040 2848
rect 39163 2808 40040 2836
rect 39163 2805 39175 2808
rect 39117 2799 39175 2805
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 1104 2746 43516 2768
rect 1104 2694 6251 2746
rect 6303 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 16854 2746
rect 16906 2694 16918 2746
rect 16970 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 27457 2746
rect 27509 2694 27521 2746
rect 27573 2694 27585 2746
rect 27637 2694 27649 2746
rect 27701 2694 27713 2746
rect 27765 2694 38060 2746
rect 38112 2694 38124 2746
rect 38176 2694 38188 2746
rect 38240 2694 38252 2746
rect 38304 2694 38316 2746
rect 38368 2694 43516 2746
rect 1104 2672 43516 2694
rect 5074 2592 5080 2644
rect 5132 2592 5138 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 8481 2635 8539 2641
rect 6227 2604 8432 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 7466 2564 7472 2576
rect 5675 2536 7472 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7653 2567 7711 2573
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 8202 2564 8208 2576
rect 7699 2536 8208 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 8404 2564 8432 2604
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9306 2632 9312 2644
rect 8527 2604 9312 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 10778 2592 10784 2644
rect 10836 2592 10842 2644
rect 10962 2592 10968 2644
rect 11020 2592 11026 2644
rect 11330 2592 11336 2644
rect 11388 2592 11394 2644
rect 12710 2632 12716 2644
rect 11716 2604 12716 2632
rect 8938 2564 8944 2576
rect 8404 2536 8944 2564
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 9125 2567 9183 2573
rect 9125 2533 9137 2567
rect 9171 2533 9183 2567
rect 9125 2527 9183 2533
rect 10229 2567 10287 2573
rect 10229 2533 10241 2567
rect 10275 2564 10287 2567
rect 10410 2564 10416 2576
rect 10275 2536 10416 2564
rect 10275 2533 10287 2536
rect 10229 2527 10287 2533
rect 8110 2496 8116 2508
rect 7760 2468 8116 2496
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 5166 2388 5172 2440
rect 5224 2388 5230 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5626 2428 5632 2440
rect 5491 2400 5632 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5994 2388 6000 2440
rect 6052 2388 6058 2440
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 6917 2431 6975 2437
rect 6687 2400 6868 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 6380 2360 6408 2391
rect 6730 2360 6736 2372
rect 6380 2332 6736 2360
rect 6730 2320 6736 2332
rect 6788 2320 6794 2372
rect 6840 2360 6868 2400
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7098 2428 7104 2440
rect 6963 2400 7104 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7650 2428 7656 2440
rect 7515 2400 7656 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7006 2360 7012 2372
rect 6840 2332 7012 2360
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 7208 2360 7236 2391
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7760 2437 7788 2468
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 9140 2496 9168 2527
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 10980 2564 11008 2592
rect 10551 2536 11008 2564
rect 11057 2567 11115 2573
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 11422 2564 11428 2576
rect 11103 2536 11428 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 11716 2573 11744 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 12802 2592 12808 2644
rect 12860 2592 12866 2644
rect 13372 2604 13676 2632
rect 11701 2567 11759 2573
rect 11701 2533 11713 2567
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 12250 2524 12256 2576
rect 12308 2524 12314 2576
rect 13372 2564 13400 2604
rect 13648 2576 13676 2604
rect 14642 2592 14648 2644
rect 14700 2592 14706 2644
rect 15194 2632 15200 2644
rect 14752 2604 15200 2632
rect 12360 2536 13400 2564
rect 12158 2496 12164 2508
rect 9140 2468 12164 2496
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 12360 2496 12388 2536
rect 13446 2524 13452 2576
rect 13504 2524 13510 2576
rect 13630 2524 13636 2576
rect 13688 2524 13694 2576
rect 14369 2567 14427 2573
rect 14369 2533 14381 2567
rect 14415 2564 14427 2567
rect 14752 2564 14780 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17497 2635 17555 2641
rect 17497 2601 17509 2635
rect 17543 2632 17555 2635
rect 17543 2604 18000 2632
rect 17543 2601 17555 2604
rect 17497 2595 17555 2601
rect 14415 2536 14780 2564
rect 14921 2567 14979 2573
rect 14415 2533 14427 2536
rect 14369 2527 14427 2533
rect 14921 2533 14933 2567
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 13464 2496 13492 2524
rect 14458 2496 14464 2508
rect 12268 2468 12388 2496
rect 13004 2468 13492 2496
rect 13740 2468 14464 2496
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8478 2428 8484 2440
rect 8343 2400 8484 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 7558 2360 7564 2372
rect 7208 2332 7564 2360
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 8036 2360 8064 2391
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 8846 2428 8852 2440
rect 8619 2400 8852 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9398 2428 9404 2440
rect 9263 2400 9404 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9582 2428 9588 2440
rect 9539 2400 9588 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 9950 2428 9956 2440
rect 9815 2400 9956 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10226 2428 10232 2440
rect 10091 2400 10232 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10502 2428 10508 2440
rect 10367 2400 10508 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10778 2428 10784 2440
rect 10643 2400 10784 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11054 2428 11060 2440
rect 10919 2400 11060 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 11422 2428 11428 2440
rect 11195 2400 11428 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 11974 2428 11980 2440
rect 11839 2400 11980 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 8386 2360 8392 2372
rect 8036 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 8680 2332 9628 2360
rect 5350 2252 5356 2304
rect 5408 2252 5414 2304
rect 5902 2252 5908 2304
rect 5960 2252 5966 2304
rect 6546 2252 6552 2304
rect 6604 2252 6610 2304
rect 6825 2295 6883 2301
rect 6825 2261 6837 2295
rect 6871 2292 6883 2295
rect 6914 2292 6920 2304
rect 6871 2264 6920 2292
rect 6871 2261 6883 2264
rect 6825 2255 6883 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 7282 2292 7288 2304
rect 7147 2264 7288 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 7374 2252 7380 2304
rect 7432 2252 7438 2304
rect 7926 2252 7932 2304
rect 7984 2252 7990 2304
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8680 2292 8708 2332
rect 9600 2304 9628 2332
rect 9692 2332 10364 2360
rect 8251 2264 8708 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8754 2252 8760 2304
rect 8812 2252 8818 2304
rect 9398 2252 9404 2304
rect 9456 2252 9462 2304
rect 9582 2252 9588 2304
rect 9640 2252 9646 2304
rect 9692 2301 9720 2332
rect 9677 2295 9735 2301
rect 9677 2261 9689 2295
rect 9723 2261 9735 2295
rect 9677 2255 9735 2261
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10336 2292 10364 2332
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 11238 2360 11244 2372
rect 10468 2332 11244 2360
rect 10468 2320 10474 2332
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 12268 2360 12296 2468
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 13004 2360 13032 2468
rect 13170 2388 13176 2440
rect 13228 2388 13234 2440
rect 13740 2437 13768 2468
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 14936 2496 14964 2527
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 16114 2564 16120 2576
rect 15068 2536 16120 2564
rect 15068 2524 15074 2536
rect 16114 2524 16120 2536
rect 16172 2524 16178 2576
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 17678 2564 17684 2576
rect 16899 2536 17684 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 17678 2524 17684 2536
rect 17736 2524 17742 2576
rect 17310 2496 17316 2508
rect 14936 2468 15240 2496
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 11808 2332 12296 2360
rect 12406 2332 13032 2360
rect 13464 2360 13492 2391
rect 13814 2360 13820 2372
rect 13464 2332 13820 2360
rect 11808 2292 11836 2332
rect 10336 2264 11836 2292
rect 11977 2295 12035 2301
rect 11977 2261 11989 2295
rect 12023 2292 12035 2295
rect 12406 2292 12434 2332
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 14108 2360 14136 2391
rect 14550 2388 14556 2440
rect 14608 2388 14614 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 14734 2360 14740 2372
rect 14108 2332 14740 2360
rect 14734 2320 14740 2332
rect 14792 2320 14798 2372
rect 14844 2360 14872 2391
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15212 2437 15240 2468
rect 16960 2468 17316 2496
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 15746 2388 15752 2440
rect 15804 2388 15810 2440
rect 16022 2388 16028 2440
rect 16080 2388 16086 2440
rect 16298 2388 16304 2440
rect 16356 2388 16362 2440
rect 16666 2388 16672 2440
rect 16724 2388 16730 2440
rect 16960 2437 16988 2468
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17586 2428 17592 2440
rect 17267 2400 17592 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 17862 2428 17868 2440
rect 17819 2400 17868 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 15562 2360 15568 2372
rect 14844 2332 15568 2360
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 17310 2360 17316 2372
rect 15948 2332 17316 2360
rect 12023 2264 12434 2292
rect 12023 2261 12035 2264
rect 11977 2255 12035 2261
rect 12526 2252 12532 2304
rect 12584 2252 12590 2304
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 13354 2252 13360 2304
rect 13412 2252 13418 2304
rect 13630 2252 13636 2304
rect 13688 2252 13694 2304
rect 13906 2252 13912 2304
rect 13964 2252 13970 2304
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 15378 2252 15384 2304
rect 15436 2252 15442 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15838 2292 15844 2304
rect 15703 2264 15844 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 15948 2301 15976 2332
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 15933 2295 15991 2301
rect 15933 2261 15945 2295
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16390 2292 16396 2304
rect 16255 2264 16396 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16482 2252 16488 2304
rect 16540 2252 16546 2304
rect 17126 2252 17132 2304
rect 17184 2252 17190 2304
rect 17402 2252 17408 2304
rect 17460 2252 17466 2304
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 17696 2292 17724 2391
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 17972 2360 18000 2604
rect 18506 2592 18512 2644
rect 18564 2592 18570 2644
rect 18966 2592 18972 2644
rect 19024 2592 19030 2644
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 19392 2604 25452 2632
rect 19392 2592 19398 2604
rect 18049 2567 18107 2573
rect 18049 2533 18061 2567
rect 18095 2564 18107 2567
rect 18984 2564 19012 2592
rect 18095 2536 19012 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 21818 2564 21824 2576
rect 19300 2536 20208 2564
rect 19300 2524 19306 2536
rect 19150 2496 19156 2508
rect 18248 2468 19156 2496
rect 18248 2437 18276 2468
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 18322 2388 18328 2440
rect 18380 2388 18386 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 20180 2437 20208 2536
rect 20272 2536 21824 2564
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 18693 2363 18751 2369
rect 18693 2360 18705 2363
rect 17972 2332 18705 2360
rect 18693 2329 18705 2332
rect 18739 2329 18751 2363
rect 18693 2323 18751 2329
rect 19061 2363 19119 2369
rect 19061 2329 19073 2363
rect 19107 2360 19119 2363
rect 19334 2360 19340 2372
rect 19107 2332 19340 2360
rect 19107 2329 19119 2332
rect 19061 2323 19119 2329
rect 19334 2320 19340 2332
rect 19392 2320 19398 2372
rect 19981 2363 20039 2369
rect 19981 2329 19993 2363
rect 20027 2360 20039 2363
rect 20070 2360 20076 2372
rect 20027 2332 20076 2360
rect 20027 2329 20039 2332
rect 19981 2323 20039 2329
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 17644 2264 17724 2292
rect 17957 2295 18015 2301
rect 17644 2252 17650 2264
rect 17957 2261 17969 2295
rect 18003 2292 18015 2295
rect 18966 2292 18972 2304
rect 18003 2264 18972 2292
rect 18003 2261 18015 2264
rect 17957 2255 18015 2261
rect 18966 2252 18972 2264
rect 19024 2252 19030 2304
rect 19245 2295 19303 2301
rect 19245 2261 19257 2295
rect 19291 2292 19303 2295
rect 20272 2292 20300 2536
rect 21818 2524 21824 2536
rect 21876 2524 21882 2576
rect 23937 2567 23995 2573
rect 22066 2536 23888 2564
rect 22066 2496 22094 2536
rect 20824 2468 22094 2496
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20680 2400 20729 2428
rect 20680 2388 20686 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 20533 2363 20591 2369
rect 20533 2329 20545 2363
rect 20579 2329 20591 2363
rect 20533 2323 20591 2329
rect 19291 2264 20300 2292
rect 20548 2292 20576 2323
rect 20824 2304 20852 2468
rect 22554 2456 22560 2508
rect 22612 2496 22618 2508
rect 22649 2499 22707 2505
rect 22649 2496 22661 2499
rect 22612 2468 22661 2496
rect 22612 2456 22618 2468
rect 22649 2465 22661 2468
rect 22695 2465 22707 2499
rect 22649 2459 22707 2465
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 20956 2400 21281 2428
rect 20956 2388 20962 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21876 2400 22201 2428
rect 21876 2388 21882 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22336 2400 22937 2428
rect 22336 2388 22342 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23474 2388 23480 2440
rect 23532 2388 23538 2440
rect 23860 2428 23888 2536
rect 23937 2533 23949 2567
rect 23983 2533 23995 2567
rect 23937 2527 23995 2533
rect 23952 2496 23980 2527
rect 23952 2468 25084 2496
rect 23934 2428 23940 2440
rect 23860 2400 23940 2428
rect 23934 2388 23940 2400
rect 23992 2388 23998 2440
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24121 2431 24179 2437
rect 24121 2428 24133 2431
rect 24084 2400 24133 2428
rect 24084 2388 24090 2400
rect 24121 2397 24133 2400
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 25056 2437 25084 2468
rect 25314 2456 25320 2508
rect 25372 2456 25378 2508
rect 25424 2496 25452 2604
rect 26142 2592 26148 2644
rect 26200 2632 26206 2644
rect 26237 2635 26295 2641
rect 26237 2632 26249 2635
rect 26200 2604 26249 2632
rect 26200 2592 26206 2604
rect 26237 2601 26249 2604
rect 26283 2601 26295 2635
rect 26237 2595 26295 2601
rect 26602 2592 26608 2644
rect 26660 2592 26666 2644
rect 26786 2592 26792 2644
rect 26844 2632 26850 2644
rect 27709 2635 27767 2641
rect 27709 2632 27721 2635
rect 26844 2604 27721 2632
rect 26844 2592 26850 2604
rect 27709 2601 27721 2604
rect 27755 2601 27767 2635
rect 27709 2595 27767 2601
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 29181 2635 29239 2641
rect 29181 2632 29193 2635
rect 28776 2604 29193 2632
rect 28776 2592 28782 2604
rect 29181 2601 29193 2604
rect 29227 2601 29239 2635
rect 29181 2595 29239 2601
rect 29638 2592 29644 2644
rect 29696 2632 29702 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 29696 2604 30849 2632
rect 29696 2592 29702 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 31754 2592 31760 2644
rect 31812 2592 31818 2644
rect 32309 2635 32367 2641
rect 32309 2601 32321 2635
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 30377 2567 30435 2573
rect 30377 2564 30389 2567
rect 28960 2536 30389 2564
rect 28960 2524 28966 2536
rect 30377 2533 30389 2536
rect 30423 2533 30435 2567
rect 30377 2527 30435 2533
rect 31018 2524 31024 2576
rect 31076 2564 31082 2576
rect 32324 2564 32352 2595
rect 33410 2592 33416 2644
rect 33468 2632 33474 2644
rect 34333 2635 34391 2641
rect 34333 2632 34345 2635
rect 33468 2604 34345 2632
rect 33468 2592 33474 2604
rect 34333 2601 34345 2604
rect 34379 2601 34391 2635
rect 34333 2595 34391 2601
rect 34885 2635 34943 2641
rect 34885 2601 34897 2635
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 31076 2536 32352 2564
rect 31076 2524 31082 2536
rect 33318 2524 33324 2576
rect 33376 2564 33382 2576
rect 34900 2564 34928 2595
rect 35526 2592 35532 2644
rect 35584 2592 35590 2644
rect 35802 2592 35808 2644
rect 35860 2592 35866 2644
rect 35986 2592 35992 2644
rect 36044 2632 36050 2644
rect 36173 2635 36231 2641
rect 36173 2632 36185 2635
rect 36044 2604 36185 2632
rect 36044 2592 36050 2604
rect 36173 2601 36185 2604
rect 36219 2601 36231 2635
rect 36173 2595 36231 2601
rect 36998 2592 37004 2644
rect 37056 2592 37062 2644
rect 37826 2592 37832 2644
rect 37884 2632 37890 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 37884 2604 38025 2632
rect 37884 2592 37890 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 38378 2592 38384 2644
rect 38436 2592 38442 2644
rect 38654 2592 38660 2644
rect 38712 2592 38718 2644
rect 39853 2635 39911 2641
rect 39853 2601 39865 2635
rect 39899 2632 39911 2635
rect 39942 2632 39948 2644
rect 39899 2604 39948 2632
rect 39899 2601 39911 2604
rect 39853 2595 39911 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 40681 2635 40739 2641
rect 40681 2601 40693 2635
rect 40727 2632 40739 2635
rect 41506 2632 41512 2644
rect 40727 2604 41512 2632
rect 40727 2601 40739 2604
rect 40681 2595 40739 2601
rect 41506 2592 41512 2604
rect 41564 2592 41570 2644
rect 42426 2592 42432 2644
rect 42484 2592 42490 2644
rect 33376 2536 34928 2564
rect 35544 2564 35572 2592
rect 36541 2567 36599 2573
rect 36541 2564 36553 2567
rect 35544 2536 36553 2564
rect 33376 2524 33382 2536
rect 36541 2533 36553 2536
rect 36587 2533 36599 2567
rect 36541 2527 36599 2533
rect 37366 2524 37372 2576
rect 37424 2564 37430 2576
rect 38396 2564 38424 2592
rect 38933 2567 38991 2573
rect 38933 2564 38945 2567
rect 37424 2536 38148 2564
rect 38396 2536 38945 2564
rect 37424 2524 37430 2536
rect 25424 2468 27660 2496
rect 25041 2431 25099 2437
rect 24360 2400 24900 2428
rect 24360 2388 24366 2400
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21358 2360 21364 2372
rect 21131 2332 21364 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 21637 2363 21695 2369
rect 21637 2329 21649 2363
rect 21683 2360 21695 2363
rect 21910 2360 21916 2372
rect 21683 2332 21916 2360
rect 21683 2329 21695 2332
rect 21637 2323 21695 2329
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 22373 2363 22431 2369
rect 22373 2329 22385 2363
rect 22419 2360 22431 2363
rect 22646 2360 22652 2372
rect 22419 2332 22652 2360
rect 22419 2329 22431 2332
rect 22373 2323 22431 2329
rect 22646 2320 22652 2332
rect 22704 2320 22710 2372
rect 24489 2363 24547 2369
rect 24489 2360 24501 2363
rect 22940 2332 24501 2360
rect 20622 2292 20628 2304
rect 20548 2264 20628 2292
rect 19291 2261 19303 2264
rect 19245 2255 19303 2261
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 20806 2252 20812 2304
rect 20864 2252 20870 2304
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2292 22063 2295
rect 22940 2292 22968 2332
rect 24489 2329 24501 2332
rect 24535 2329 24547 2363
rect 24872 2360 24900 2400
rect 25041 2397 25053 2431
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 26145 2431 26203 2437
rect 26145 2428 26157 2431
rect 25188 2400 26157 2428
rect 25188 2388 25194 2400
rect 26145 2397 26157 2400
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26234 2388 26240 2440
rect 26292 2388 26298 2440
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26789 2431 26847 2437
rect 26789 2428 26801 2431
rect 26476 2400 26801 2428
rect 26476 2388 26482 2400
rect 26789 2397 26801 2400
rect 26835 2397 26847 2431
rect 27632 2428 27660 2468
rect 27706 2456 27712 2508
rect 27764 2496 27770 2508
rect 28997 2499 29055 2505
rect 28997 2496 29009 2499
rect 27764 2468 29009 2496
rect 27764 2456 27770 2468
rect 28997 2465 29009 2468
rect 29043 2465 29055 2499
rect 28997 2459 29055 2465
rect 29288 2468 30788 2496
rect 29288 2428 29316 2468
rect 27632 2400 29316 2428
rect 29365 2431 29423 2437
rect 26789 2391 26847 2397
rect 29365 2397 29377 2431
rect 29411 2428 29423 2431
rect 29454 2428 29460 2440
rect 29411 2400 29460 2428
rect 29411 2397 29423 2400
rect 29365 2391 29423 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 29730 2388 29736 2440
rect 29788 2428 29794 2440
rect 30760 2437 30788 2468
rect 31956 2468 33088 2496
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 29788 2400 30205 2428
rect 29788 2388 29794 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2397 30803 2431
rect 30745 2391 30803 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31956 2437 31984 2468
rect 31941 2431 31999 2437
rect 30892 2400 31432 2428
rect 30892 2388 30898 2400
rect 25593 2363 25651 2369
rect 25593 2360 25605 2363
rect 24872 2332 25605 2360
rect 24489 2323 24547 2329
rect 25593 2329 25605 2332
rect 25639 2329 25651 2363
rect 26252 2360 26280 2388
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 26252 2332 27077 2360
rect 25593 2323 25651 2329
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 27617 2363 27675 2369
rect 27617 2329 27629 2363
rect 27663 2360 27675 2363
rect 27798 2360 27804 2372
rect 27663 2332 27804 2360
rect 27663 2329 27675 2332
rect 27617 2323 27675 2329
rect 27798 2320 27804 2332
rect 27856 2320 27862 2372
rect 27890 2320 27896 2372
rect 27948 2360 27954 2372
rect 28169 2363 28227 2369
rect 28169 2360 28181 2363
rect 27948 2332 28181 2360
rect 27948 2320 27954 2332
rect 28169 2329 28181 2332
rect 28215 2329 28227 2363
rect 28169 2323 28227 2329
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28721 2363 28779 2369
rect 28721 2360 28733 2363
rect 28408 2332 28733 2360
rect 28408 2320 28414 2332
rect 28721 2329 28733 2332
rect 28767 2329 28779 2363
rect 28721 2323 28779 2329
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29641 2363 29699 2369
rect 29641 2360 29653 2363
rect 29052 2332 29653 2360
rect 29052 2320 29058 2332
rect 29641 2329 29653 2332
rect 29687 2329 29699 2363
rect 29641 2323 29699 2329
rect 29914 2320 29920 2372
rect 29972 2360 29978 2372
rect 31297 2363 31355 2369
rect 31297 2360 31309 2363
rect 29972 2332 31309 2360
rect 29972 2320 29978 2332
rect 31297 2329 31309 2332
rect 31343 2329 31355 2363
rect 31404 2360 31432 2400
rect 31941 2397 31953 2431
rect 31987 2397 31999 2431
rect 33060 2428 33088 2468
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 33192 2468 33916 2496
rect 33192 2456 33198 2468
rect 33888 2437 33916 2468
rect 34422 2456 34428 2508
rect 34480 2496 34486 2508
rect 34480 2468 36032 2496
rect 34480 2456 34486 2468
rect 33873 2431 33931 2437
rect 31941 2391 31999 2397
rect 32140 2400 32812 2428
rect 33060 2400 33824 2428
rect 32140 2360 32168 2400
rect 31404 2332 32168 2360
rect 31297 2323 31355 2329
rect 32214 2320 32220 2372
rect 32272 2320 32278 2372
rect 32784 2369 32812 2400
rect 32769 2363 32827 2369
rect 32769 2329 32781 2363
rect 32815 2329 32827 2363
rect 32769 2323 32827 2329
rect 33226 2320 33232 2372
rect 33284 2360 33290 2372
rect 33321 2363 33379 2369
rect 33321 2360 33333 2363
rect 33284 2332 33333 2360
rect 33284 2320 33290 2332
rect 33321 2329 33333 2332
rect 33367 2329 33379 2363
rect 33796 2360 33824 2400
rect 33873 2397 33885 2431
rect 33919 2397 33931 2431
rect 33873 2391 33931 2397
rect 34054 2388 34060 2440
rect 34112 2428 34118 2440
rect 34517 2431 34575 2437
rect 34517 2428 34529 2431
rect 34112 2400 34529 2428
rect 34112 2388 34118 2400
rect 34517 2397 34529 2400
rect 34563 2397 34575 2431
rect 34517 2391 34575 2397
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2428 35771 2431
rect 35894 2428 35900 2440
rect 35759 2400 35900 2428
rect 35759 2397 35771 2400
rect 35713 2391 35771 2397
rect 35894 2388 35900 2400
rect 35952 2388 35958 2440
rect 36004 2437 36032 2468
rect 36078 2456 36084 2508
rect 36136 2496 36142 2508
rect 36136 2468 36860 2496
rect 36136 2456 36142 2468
rect 35989 2431 36047 2437
rect 35989 2397 36001 2431
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36170 2388 36176 2440
rect 36228 2428 36234 2440
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 36228 2400 36461 2428
rect 36228 2388 36234 2400
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 36722 2388 36728 2440
rect 36780 2388 36786 2440
rect 36832 2437 36860 2468
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 36964 2468 37596 2496
rect 36964 2456 36970 2468
rect 37568 2437 37596 2468
rect 38120 2437 38148 2536
rect 38933 2533 38945 2536
rect 38979 2533 38991 2567
rect 38933 2527 38991 2533
rect 39209 2567 39267 2573
rect 39209 2533 39221 2567
rect 39255 2533 39267 2567
rect 39209 2527 39267 2533
rect 40129 2567 40187 2573
rect 40129 2533 40141 2567
rect 40175 2533 40187 2567
rect 40129 2527 40187 2533
rect 40405 2567 40463 2573
rect 40405 2533 40417 2567
rect 40451 2564 40463 2567
rect 40451 2536 42656 2564
rect 40451 2533 40463 2536
rect 40405 2527 40463 2533
rect 39224 2496 39252 2527
rect 38856 2468 39252 2496
rect 40144 2496 40172 2527
rect 40144 2468 40908 2496
rect 38856 2437 38884 2468
rect 36817 2431 36875 2437
rect 36817 2397 36829 2431
rect 36863 2397 36875 2431
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36817 2391 36875 2397
rect 37108 2400 37289 2428
rect 34698 2360 34704 2372
rect 33796 2332 34704 2360
rect 33321 2323 33379 2329
rect 34698 2320 34704 2332
rect 34756 2320 34762 2372
rect 34790 2320 34796 2372
rect 34848 2320 34854 2372
rect 35345 2363 35403 2369
rect 35345 2329 35357 2363
rect 35391 2360 35403 2363
rect 35391 2332 36308 2360
rect 35391 2329 35403 2332
rect 35345 2323 35403 2329
rect 22051 2264 22968 2292
rect 22051 2261 22063 2264
rect 22005 2255 22063 2261
rect 23014 2252 23020 2304
rect 23072 2252 23078 2304
rect 23290 2252 23296 2304
rect 23348 2292 23354 2304
rect 23569 2295 23627 2301
rect 23569 2292 23581 2295
rect 23348 2264 23581 2292
rect 23348 2252 23354 2264
rect 23569 2261 23581 2264
rect 23615 2261 23627 2295
rect 23569 2255 23627 2261
rect 23750 2252 23756 2304
rect 23808 2292 23814 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23808 2264 24593 2292
rect 23808 2252 23814 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 25685 2295 25743 2301
rect 25685 2292 25697 2295
rect 24728 2264 25697 2292
rect 24728 2252 24734 2264
rect 25685 2261 25697 2264
rect 25731 2261 25743 2295
rect 25685 2255 25743 2261
rect 26326 2252 26332 2304
rect 26384 2292 26390 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26384 2264 27169 2292
rect 26384 2252 26390 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27522 2252 27528 2304
rect 27580 2292 27586 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 27580 2264 28273 2292
rect 27580 2252 27586 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 28442 2252 28448 2304
rect 28500 2292 28506 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 28500 2264 29745 2292
rect 28500 2252 28506 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30098 2252 30104 2304
rect 30156 2292 30162 2304
rect 31389 2295 31447 2301
rect 31389 2292 31401 2295
rect 30156 2264 31401 2292
rect 30156 2252 30162 2264
rect 31389 2261 31401 2264
rect 31435 2261 31447 2295
rect 31389 2255 31447 2261
rect 32306 2252 32312 2304
rect 32364 2292 32370 2304
rect 32861 2295 32919 2301
rect 32861 2292 32873 2295
rect 32364 2264 32873 2292
rect 32364 2252 32370 2264
rect 32861 2261 32873 2264
rect 32907 2261 32919 2295
rect 32861 2255 32919 2261
rect 33410 2252 33416 2304
rect 33468 2252 33474 2304
rect 33962 2252 33968 2304
rect 34020 2252 34026 2304
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36280 2301 36308 2332
rect 36630 2320 36636 2372
rect 36688 2360 36694 2372
rect 37108 2360 37136 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 38841 2431 38899 2437
rect 38841 2397 38853 2431
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 36688 2332 37136 2360
rect 36688 2320 36694 2332
rect 37182 2320 37188 2372
rect 37240 2360 37246 2372
rect 37844 2360 37872 2391
rect 37240 2332 37872 2360
rect 38580 2360 38608 2391
rect 38930 2388 38936 2440
rect 38988 2428 38994 2440
rect 39117 2431 39175 2437
rect 39117 2428 39129 2431
rect 38988 2400 39129 2428
rect 38988 2388 38994 2400
rect 39117 2397 39129 2400
rect 39163 2397 39175 2431
rect 39117 2391 39175 2397
rect 39390 2388 39396 2440
rect 39448 2388 39454 2440
rect 39666 2388 39672 2440
rect 39724 2388 39730 2440
rect 40034 2388 40040 2440
rect 40092 2388 40098 2440
rect 40310 2388 40316 2440
rect 40368 2388 40374 2440
rect 40880 2437 40908 2468
rect 42628 2437 42656 2536
rect 40589 2431 40647 2437
rect 40589 2397 40601 2431
rect 40635 2397 40647 2431
rect 40589 2391 40647 2397
rect 40865 2431 40923 2437
rect 40865 2397 40877 2431
rect 40911 2397 40923 2431
rect 40865 2391 40923 2397
rect 42613 2431 42671 2437
rect 42613 2397 42625 2431
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 38580 2332 39528 2360
rect 37240 2320 37246 2332
rect 36265 2295 36323 2301
rect 36265 2261 36277 2295
rect 36311 2261 36323 2295
rect 36265 2255 36323 2261
rect 36354 2252 36360 2304
rect 36412 2292 36418 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 36412 2264 37473 2292
rect 36412 2252 36418 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37461 2255 37519 2261
rect 37734 2252 37740 2304
rect 37792 2252 37798 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38378 2252 38384 2304
rect 38436 2252 38442 2304
rect 39500 2301 39528 2332
rect 39942 2320 39948 2372
rect 40000 2360 40006 2372
rect 40604 2360 40632 2391
rect 40000 2332 40632 2360
rect 40000 2320 40006 2332
rect 39485 2295 39543 2301
rect 39485 2261 39497 2295
rect 39531 2261 39543 2295
rect 39485 2255 39543 2261
rect 1104 2202 43675 2224
rect 1104 2150 11552 2202
rect 11604 2150 11616 2202
rect 11668 2150 11680 2202
rect 11732 2150 11744 2202
rect 11796 2150 11808 2202
rect 11860 2150 22155 2202
rect 22207 2150 22219 2202
rect 22271 2150 22283 2202
rect 22335 2150 22347 2202
rect 22399 2150 22411 2202
rect 22463 2150 32758 2202
rect 32810 2150 32822 2202
rect 32874 2150 32886 2202
rect 32938 2150 32950 2202
rect 33002 2150 33014 2202
rect 33066 2150 43361 2202
rect 43413 2150 43425 2202
rect 43477 2150 43489 2202
rect 43541 2150 43553 2202
rect 43605 2150 43617 2202
rect 43669 2150 43675 2202
rect 1104 2128 43675 2150
rect 5902 2048 5908 2100
rect 5960 2048 5966 2100
rect 7926 2048 7932 2100
rect 7984 2088 7990 2100
rect 7984 2060 9904 2088
rect 7984 2048 7990 2060
rect 5920 1884 5948 2048
rect 6822 1980 6828 2032
rect 6880 2020 6886 2032
rect 9876 2020 9904 2060
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 13262 2088 13268 2100
rect 10008 2060 13268 2088
rect 10008 2048 10014 2060
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 13354 2048 13360 2100
rect 13412 2088 13418 2100
rect 15010 2088 15016 2100
rect 13412 2060 15016 2088
rect 13412 2048 13418 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 17402 2048 17408 2100
rect 17460 2088 17466 2100
rect 20806 2088 20812 2100
rect 17460 2060 20812 2088
rect 17460 2048 17466 2060
rect 20806 2048 20812 2060
rect 20864 2048 20870 2100
rect 22922 2088 22928 2100
rect 22066 2060 22928 2088
rect 22066 2020 22094 2060
rect 22922 2048 22928 2060
rect 22980 2048 22986 2100
rect 24854 2048 24860 2100
rect 24912 2088 24918 2100
rect 29914 2088 29920 2100
rect 24912 2060 29920 2088
rect 24912 2048 24918 2060
rect 29914 2048 29920 2060
rect 29972 2048 29978 2100
rect 31570 2048 31576 2100
rect 31628 2088 31634 2100
rect 33410 2088 33416 2100
rect 31628 2060 33416 2088
rect 31628 2048 31634 2060
rect 33410 2048 33416 2060
rect 33468 2048 33474 2100
rect 37458 2048 37464 2100
rect 37516 2088 37522 2100
rect 38378 2088 38384 2100
rect 37516 2060 38384 2088
rect 37516 2048 37522 2060
rect 38378 2048 38384 2060
rect 38436 2048 38442 2100
rect 6880 1992 9628 2020
rect 9876 1992 22094 2020
rect 6880 1980 6886 1992
rect 9600 1884 9628 1992
rect 23382 1980 23388 2032
rect 23440 2020 23446 2032
rect 37734 2020 37740 2032
rect 23440 1992 37740 2020
rect 23440 1980 23446 1992
rect 37734 1980 37740 1992
rect 37792 1980 37798 2032
rect 14274 1912 14280 1964
rect 14332 1952 14338 1964
rect 23106 1952 23112 1964
rect 14332 1924 23112 1952
rect 14332 1912 14338 1924
rect 23106 1912 23112 1924
rect 23164 1912 23170 1964
rect 24118 1912 24124 1964
rect 24176 1952 24182 1964
rect 25314 1952 25320 1964
rect 24176 1924 25320 1952
rect 24176 1912 24182 1924
rect 25314 1912 25320 1924
rect 25372 1912 25378 1964
rect 35434 1952 35440 1964
rect 26206 1924 35440 1952
rect 26206 1884 26234 1924
rect 35434 1912 35440 1924
rect 35492 1912 35498 1964
rect 36354 1912 36360 1964
rect 36412 1912 36418 1964
rect 36372 1884 36400 1912
rect 5920 1856 9352 1884
rect 9600 1856 26234 1884
rect 26344 1856 36400 1884
rect 7282 1776 7288 1828
rect 7340 1776 7346 1828
rect 9324 1816 9352 1856
rect 17586 1816 17592 1828
rect 9324 1788 17592 1816
rect 17586 1776 17592 1788
rect 17644 1776 17650 1828
rect 18046 1776 18052 1828
rect 18104 1776 18110 1828
rect 20990 1776 20996 1828
rect 21048 1816 21054 1828
rect 26344 1816 26372 1856
rect 21048 1788 26372 1816
rect 21048 1776 21054 1788
rect 33870 1776 33876 1828
rect 33928 1816 33934 1828
rect 38286 1816 38292 1828
rect 33928 1788 38292 1816
rect 33928 1776 33934 1788
rect 38286 1776 38292 1788
rect 38344 1776 38350 1828
rect 7300 1748 7328 1776
rect 7300 1720 9352 1748
rect 7374 1640 7380 1692
rect 7432 1640 7438 1692
rect 7466 1640 7472 1692
rect 7524 1640 7530 1692
rect 9324 1680 9352 1720
rect 9398 1708 9404 1760
rect 9456 1748 9462 1760
rect 12986 1748 12992 1760
rect 9456 1720 12992 1748
rect 9456 1708 9462 1720
rect 12986 1708 12992 1720
rect 13044 1708 13050 1760
rect 13906 1708 13912 1760
rect 13964 1748 13970 1760
rect 18064 1748 18092 1776
rect 29454 1748 29460 1760
rect 13964 1720 18092 1748
rect 26206 1720 29460 1748
rect 13964 1708 13970 1720
rect 9858 1680 9864 1692
rect 9324 1652 9864 1680
rect 9858 1640 9864 1652
rect 9916 1640 9922 1692
rect 12710 1640 12716 1692
rect 12768 1680 12774 1692
rect 26206 1680 26234 1720
rect 29454 1708 29460 1720
rect 29512 1708 29518 1760
rect 12768 1652 26234 1680
rect 12768 1640 12774 1652
rect 26418 1640 26424 1692
rect 26476 1640 26482 1692
rect 7392 1544 7420 1640
rect 7484 1612 7512 1640
rect 14918 1612 14924 1624
rect 7484 1584 14924 1612
rect 14918 1572 14924 1584
rect 14976 1572 14982 1624
rect 15102 1572 15108 1624
rect 15160 1612 15166 1624
rect 15654 1612 15660 1624
rect 15160 1584 15660 1612
rect 15160 1572 15166 1584
rect 15654 1572 15660 1584
rect 15712 1572 15718 1624
rect 16114 1572 16120 1624
rect 16172 1612 16178 1624
rect 26436 1612 26464 1640
rect 16172 1584 26464 1612
rect 16172 1572 16178 1584
rect 22830 1544 22836 1556
rect 7392 1516 22836 1544
rect 22830 1504 22836 1516
rect 22888 1504 22894 1556
rect 38746 1504 38752 1556
rect 38804 1544 38810 1556
rect 39666 1544 39672 1556
rect 38804 1516 39672 1544
rect 38804 1504 38810 1516
rect 39666 1504 39672 1516
rect 39724 1504 39730 1556
rect 5350 1436 5356 1488
rect 5408 1476 5414 1488
rect 10686 1476 10692 1488
rect 5408 1448 10692 1476
rect 5408 1436 5414 1448
rect 10686 1436 10692 1448
rect 10744 1436 10750 1488
rect 12526 1436 12532 1488
rect 12584 1476 12590 1488
rect 26694 1476 26700 1488
rect 12584 1448 26700 1476
rect 12584 1436 12590 1448
rect 26694 1436 26700 1448
rect 26752 1436 26758 1488
rect 32214 1436 32220 1488
rect 32272 1476 32278 1488
rect 33962 1476 33968 1488
rect 32272 1448 33968 1476
rect 32272 1436 32278 1448
rect 33962 1436 33968 1448
rect 34020 1436 34026 1488
rect 39390 1476 39396 1488
rect 38672 1448 39396 1476
rect 13262 1368 13268 1420
rect 13320 1408 13326 1420
rect 13320 1380 14504 1408
rect 13320 1368 13326 1380
rect 14476 1340 14504 1380
rect 14550 1368 14556 1420
rect 14608 1408 14614 1420
rect 15102 1408 15108 1420
rect 14608 1380 15108 1408
rect 14608 1368 14614 1380
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 19058 1408 19064 1420
rect 15212 1380 19064 1408
rect 15212 1340 15240 1380
rect 19058 1368 19064 1380
rect 19116 1368 19122 1420
rect 31202 1368 31208 1420
rect 31260 1408 31266 1420
rect 32306 1408 32312 1420
rect 31260 1380 32312 1408
rect 31260 1368 31266 1380
rect 32306 1368 32312 1380
rect 32364 1368 32370 1420
rect 35618 1368 35624 1420
rect 35676 1408 35682 1420
rect 36722 1408 36728 1420
rect 35676 1380 36728 1408
rect 35676 1368 35682 1380
rect 36722 1368 36728 1380
rect 36780 1368 36786 1420
rect 14476 1312 15240 1340
rect 18046 1300 18052 1352
rect 18104 1340 18110 1352
rect 21266 1340 21272 1352
rect 18104 1312 21272 1340
rect 18104 1300 18110 1312
rect 21266 1300 21272 1312
rect 21324 1300 21330 1352
rect 38562 1300 38568 1352
rect 38620 1340 38626 1352
rect 38672 1340 38700 1448
rect 39390 1436 39396 1448
rect 39448 1436 39454 1488
rect 39298 1368 39304 1420
rect 39356 1408 39362 1420
rect 40310 1408 40316 1420
rect 39356 1380 40316 1408
rect 39356 1368 39362 1380
rect 40310 1368 40316 1380
rect 40368 1368 40374 1420
rect 38620 1312 38700 1340
rect 38620 1300 38626 1312
rect 6546 1232 6552 1284
rect 6604 1272 6610 1284
rect 24026 1272 24032 1284
rect 6604 1244 24032 1272
rect 6604 1232 6610 1244
rect 24026 1232 24032 1244
rect 24084 1232 24090 1284
rect 16482 1164 16488 1216
rect 16540 1204 16546 1216
rect 33226 1204 33232 1216
rect 16540 1176 33232 1204
rect 16540 1164 16546 1176
rect 33226 1164 33232 1176
rect 33284 1164 33290 1216
rect 15010 1096 15016 1148
rect 15068 1136 15074 1148
rect 25682 1136 25688 1148
rect 15068 1108 25688 1136
rect 15068 1096 15074 1108
rect 25682 1096 25688 1108
rect 25740 1096 25746 1148
rect 9674 1028 9680 1080
rect 9732 1068 9738 1080
rect 21450 1068 21456 1080
rect 9732 1040 21456 1068
rect 9732 1028 9738 1040
rect 21450 1028 21456 1040
rect 21508 1028 21514 1080
rect 21818 1028 21824 1080
rect 21876 1028 21882 1080
rect 9858 960 9864 1012
rect 9916 1000 9922 1012
rect 21836 1000 21864 1028
rect 9916 972 21864 1000
rect 9916 960 9922 972
rect 15838 892 15844 944
rect 15896 932 15902 944
rect 33686 932 33692 944
rect 15896 904 33692 932
rect 15896 892 15902 904
rect 33686 892 33692 904
rect 33744 892 33750 944
<< via1 >>
rect 11552 7590 11604 7642
rect 11616 7590 11668 7642
rect 11680 7590 11732 7642
rect 11744 7590 11796 7642
rect 11808 7590 11860 7642
rect 22155 7590 22207 7642
rect 22219 7590 22271 7642
rect 22283 7590 22335 7642
rect 22347 7590 22399 7642
rect 22411 7590 22463 7642
rect 32758 7590 32810 7642
rect 32822 7590 32874 7642
rect 32886 7590 32938 7642
rect 32950 7590 33002 7642
rect 33014 7590 33066 7642
rect 43361 7590 43413 7642
rect 43425 7590 43477 7642
rect 43489 7590 43541 7642
rect 43553 7590 43605 7642
rect 43617 7590 43669 7642
rect 1124 7488 1176 7540
rect 3424 7488 3476 7540
rect 5356 7488 5408 7540
rect 7472 7488 7524 7540
rect 9680 7488 9732 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 13820 7488 13872 7540
rect 15936 7488 15988 7540
rect 18052 7488 18104 7540
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 6828 7352 6880 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 22560 7531 22612 7540
rect 22560 7497 22569 7531
rect 22569 7497 22603 7531
rect 22603 7497 22612 7531
rect 22560 7488 22612 7497
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 24860 7531 24912 7540
rect 24860 7497 24869 7531
rect 24869 7497 24903 7531
rect 24903 7497 24912 7531
rect 24860 7488 24912 7497
rect 26516 7488 26568 7540
rect 28816 7488 28868 7540
rect 30748 7488 30800 7540
rect 33140 7531 33192 7540
rect 33140 7497 33149 7531
rect 33149 7497 33183 7531
rect 33183 7497 33192 7531
rect 33140 7488 33192 7497
rect 34980 7488 35032 7540
rect 37188 7488 37240 7540
rect 39304 7488 39356 7540
rect 41420 7488 41472 7540
rect 43260 7488 43312 7540
rect 20536 7352 20588 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 20444 7284 20496 7336
rect 29184 7352 29236 7404
rect 31760 7352 31812 7404
rect 33876 7284 33928 7336
rect 37372 7395 37424 7404
rect 37372 7361 37381 7395
rect 37381 7361 37415 7395
rect 37415 7361 37424 7395
rect 37372 7352 37424 7361
rect 38384 7352 38436 7404
rect 39948 7395 40000 7404
rect 39948 7361 39957 7395
rect 39957 7361 39991 7395
rect 39991 7361 40000 7395
rect 39948 7352 40000 7361
rect 41512 7395 41564 7404
rect 41512 7361 41521 7395
rect 41521 7361 41555 7395
rect 41555 7361 41564 7395
rect 41512 7352 41564 7361
rect 42432 7352 42484 7404
rect 38660 7284 38712 7336
rect 35716 7216 35768 7268
rect 20536 7148 20588 7200
rect 34796 7148 34848 7200
rect 6251 7046 6303 7098
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 16854 7046 16906 7098
rect 16918 7046 16970 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 27457 7046 27509 7098
rect 27521 7046 27573 7098
rect 27585 7046 27637 7098
rect 27649 7046 27701 7098
rect 27713 7046 27765 7098
rect 38060 7046 38112 7098
rect 38124 7046 38176 7098
rect 38188 7046 38240 7098
rect 38252 7046 38304 7098
rect 38316 7046 38368 7098
rect 7656 6944 7708 6996
rect 34428 6944 34480 6996
rect 22468 6876 22520 6928
rect 23388 6740 23440 6792
rect 11552 6502 11604 6554
rect 11616 6502 11668 6554
rect 11680 6502 11732 6554
rect 11744 6502 11796 6554
rect 11808 6502 11860 6554
rect 22155 6502 22207 6554
rect 22219 6502 22271 6554
rect 22283 6502 22335 6554
rect 22347 6502 22399 6554
rect 22411 6502 22463 6554
rect 32758 6502 32810 6554
rect 32822 6502 32874 6554
rect 32886 6502 32938 6554
rect 32950 6502 33002 6554
rect 33014 6502 33066 6554
rect 43361 6502 43413 6554
rect 43425 6502 43477 6554
rect 43489 6502 43541 6554
rect 43553 6502 43605 6554
rect 43617 6502 43669 6554
rect 22928 6264 22980 6316
rect 35992 6264 36044 6316
rect 18880 6196 18932 6248
rect 36636 6196 36688 6248
rect 1492 6128 1544 6180
rect 33508 6128 33560 6180
rect 6251 5958 6303 6010
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 16854 5958 16906 6010
rect 16918 5958 16970 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 27457 5958 27509 6010
rect 27521 5958 27573 6010
rect 27585 5958 27637 6010
rect 27649 5958 27701 6010
rect 27713 5958 27765 6010
rect 38060 5958 38112 6010
rect 38124 5958 38176 6010
rect 38188 5958 38240 6010
rect 38252 5958 38304 6010
rect 38316 5958 38368 6010
rect 24584 5856 24636 5908
rect 37832 5652 37884 5704
rect 11552 5414 11604 5466
rect 11616 5414 11668 5466
rect 11680 5414 11732 5466
rect 11744 5414 11796 5466
rect 11808 5414 11860 5466
rect 22155 5414 22207 5466
rect 22219 5414 22271 5466
rect 22283 5414 22335 5466
rect 22347 5414 22399 5466
rect 22411 5414 22463 5466
rect 32758 5414 32810 5466
rect 32822 5414 32874 5466
rect 32886 5414 32938 5466
rect 32950 5414 33002 5466
rect 33014 5414 33066 5466
rect 43361 5414 43413 5466
rect 43425 5414 43477 5466
rect 43489 5414 43541 5466
rect 43553 5414 43605 5466
rect 43617 5414 43669 5466
rect 16120 5312 16172 5364
rect 16488 5108 16540 5160
rect 6251 4870 6303 4922
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 16854 4870 16906 4922
rect 16918 4870 16970 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 27457 4870 27509 4922
rect 27521 4870 27573 4922
rect 27585 4870 27637 4922
rect 27649 4870 27701 4922
rect 27713 4870 27765 4922
rect 38060 4870 38112 4922
rect 38124 4870 38176 4922
rect 38188 4870 38240 4922
rect 38252 4870 38304 4922
rect 38316 4870 38368 4922
rect 10692 4768 10744 4820
rect 19432 4768 19484 4820
rect 8944 4700 8996 4752
rect 24216 4700 24268 4752
rect 6736 4632 6788 4684
rect 23848 4632 23900 4684
rect 8760 4564 8812 4616
rect 22744 4564 22796 4616
rect 15660 4496 15712 4548
rect 33140 4496 33192 4548
rect 10968 4428 11020 4480
rect 28724 4428 28776 4480
rect 11552 4326 11604 4378
rect 11616 4326 11668 4378
rect 11680 4326 11732 4378
rect 11744 4326 11796 4378
rect 11808 4326 11860 4378
rect 22155 4326 22207 4378
rect 22219 4326 22271 4378
rect 22283 4326 22335 4378
rect 22347 4326 22399 4378
rect 22411 4326 22463 4378
rect 32758 4326 32810 4378
rect 32822 4326 32874 4378
rect 32886 4326 32938 4378
rect 32950 4326 33002 4378
rect 33014 4326 33066 4378
rect 43361 4326 43413 4378
rect 43425 4326 43477 4378
rect 43489 4326 43541 4378
rect 43553 4326 43605 4378
rect 43617 4326 43669 4378
rect 15108 4224 15160 4276
rect 33968 4224 34020 4276
rect 14280 4156 14332 4208
rect 36360 4156 36412 4208
rect 24124 4020 24176 4072
rect 17684 3952 17736 4004
rect 25596 3952 25648 4004
rect 30012 3952 30064 4004
rect 11244 3884 11296 3936
rect 20076 3884 20128 3936
rect 22100 3884 22152 3936
rect 26424 3884 26476 3936
rect 6251 3782 6303 3834
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 16854 3782 16906 3834
rect 16918 3782 16970 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 27457 3782 27509 3834
rect 27521 3782 27573 3834
rect 27585 3782 27637 3834
rect 27649 3782 27701 3834
rect 27713 3782 27765 3834
rect 38060 3782 38112 3834
rect 38124 3782 38176 3834
rect 38188 3782 38240 3834
rect 38252 3782 38304 3834
rect 38316 3782 38368 3834
rect 17408 3680 17460 3732
rect 20536 3680 20588 3732
rect 21272 3680 21324 3732
rect 18788 3612 18840 3664
rect 20720 3612 20772 3664
rect 22652 3612 22704 3664
rect 18052 3476 18104 3528
rect 24124 3544 24176 3596
rect 18604 3476 18656 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19800 3519 19852 3528
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 20628 3476 20680 3528
rect 20904 3476 20956 3528
rect 17868 3408 17920 3460
rect 21456 3476 21508 3528
rect 21824 3451 21876 3460
rect 21824 3417 21833 3451
rect 21833 3417 21867 3451
rect 21867 3417 21876 3451
rect 21824 3408 21876 3417
rect 22836 3519 22888 3528
rect 22836 3485 22845 3519
rect 22845 3485 22879 3519
rect 22879 3485 22888 3519
rect 22836 3476 22888 3485
rect 24216 3519 24268 3528
rect 24216 3485 24225 3519
rect 24225 3485 24259 3519
rect 24259 3485 24268 3519
rect 24216 3476 24268 3485
rect 26240 3680 26292 3732
rect 28356 3680 28408 3732
rect 29184 3680 29236 3732
rect 33508 3723 33560 3732
rect 33508 3689 33517 3723
rect 33517 3689 33551 3723
rect 33551 3689 33560 3723
rect 33508 3680 33560 3689
rect 27804 3612 27856 3664
rect 27620 3544 27672 3596
rect 29736 3612 29788 3664
rect 29276 3544 29328 3596
rect 22928 3408 22980 3460
rect 23112 3408 23164 3460
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 25596 3519 25648 3528
rect 25596 3485 25605 3519
rect 25605 3485 25639 3519
rect 25639 3485 25648 3519
rect 25596 3476 25648 3485
rect 25688 3476 25740 3528
rect 26148 3519 26200 3528
rect 26148 3485 26157 3519
rect 26157 3485 26191 3519
rect 26191 3485 26200 3519
rect 26148 3476 26200 3485
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 26700 3519 26752 3528
rect 26700 3485 26709 3519
rect 26709 3485 26743 3519
rect 26743 3485 26752 3519
rect 26700 3476 26752 3485
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 27252 3519 27304 3528
rect 27252 3485 27261 3519
rect 27261 3485 27295 3519
rect 27295 3485 27304 3519
rect 27252 3476 27304 3485
rect 27896 3519 27948 3528
rect 27896 3485 27905 3519
rect 27905 3485 27939 3519
rect 27939 3485 27948 3519
rect 27896 3476 27948 3485
rect 28172 3519 28224 3528
rect 28172 3485 28181 3519
rect 28181 3485 28215 3519
rect 28215 3485 28224 3519
rect 28172 3476 28224 3485
rect 28448 3519 28500 3528
rect 28448 3485 28457 3519
rect 28457 3485 28491 3519
rect 28491 3485 28500 3519
rect 28448 3476 28500 3485
rect 28724 3519 28776 3528
rect 28724 3485 28733 3519
rect 28733 3485 28767 3519
rect 28767 3485 28776 3519
rect 28724 3476 28776 3485
rect 36268 3476 36320 3528
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 19524 3340 19576 3392
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 19892 3383 19944 3392
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 20352 3383 20404 3392
rect 20352 3349 20361 3383
rect 20361 3349 20395 3383
rect 20395 3349 20404 3383
rect 20352 3340 20404 3349
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 20904 3340 20956 3349
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 21640 3340 21692 3392
rect 22560 3340 22612 3392
rect 23480 3340 23532 3392
rect 24308 3340 24360 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 25044 3340 25096 3392
rect 25320 3340 25372 3392
rect 26332 3408 26384 3460
rect 26424 3340 26476 3392
rect 28080 3408 28132 3460
rect 29000 3408 29052 3460
rect 32036 3408 32088 3460
rect 33416 3451 33468 3460
rect 33416 3417 33425 3451
rect 33425 3417 33459 3451
rect 33459 3417 33468 3451
rect 33416 3408 33468 3417
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 32680 3340 32732 3392
rect 34704 3340 34756 3392
rect 35808 3340 35860 3392
rect 11552 3238 11604 3290
rect 11616 3238 11668 3290
rect 11680 3238 11732 3290
rect 11744 3238 11796 3290
rect 11808 3238 11860 3290
rect 22155 3238 22207 3290
rect 22219 3238 22271 3290
rect 22283 3238 22335 3290
rect 22347 3238 22399 3290
rect 22411 3238 22463 3290
rect 32758 3238 32810 3290
rect 32822 3238 32874 3290
rect 32886 3238 32938 3290
rect 32950 3238 33002 3290
rect 33014 3238 33066 3290
rect 43361 3238 43413 3290
rect 43425 3238 43477 3290
rect 43489 3238 43541 3290
rect 43553 3238 43605 3290
rect 43617 3238 43669 3290
rect 6736 3179 6788 3188
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 14188 3136 14240 3188
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 18696 3136 18748 3188
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15016 3068 15068 3120
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 14648 2932 14700 2984
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16580 3000 16632 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17684 3000 17736 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 19248 3179 19300 3188
rect 19248 3145 19257 3179
rect 19257 3145 19291 3179
rect 19291 3145 19300 3179
rect 19248 3136 19300 3145
rect 19524 3136 19576 3188
rect 19892 3136 19944 3188
rect 20352 3068 20404 3120
rect 21180 3136 21232 3188
rect 22560 3136 22612 3188
rect 24400 3136 24452 3188
rect 25320 3136 25372 3188
rect 26332 3136 26384 3188
rect 26424 3136 26476 3188
rect 28080 3136 28132 3188
rect 28540 3136 28592 3188
rect 29092 3136 29144 3188
rect 30012 3136 30064 3188
rect 30656 3136 30708 3188
rect 31852 3136 31904 3188
rect 33140 3068 33192 3120
rect 33968 3068 34020 3120
rect 35808 3136 35860 3188
rect 19340 3000 19392 3052
rect 18880 2932 18932 2984
rect 19064 2932 19116 2984
rect 16672 2864 16724 2916
rect 22744 3000 22796 3052
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 23848 3043 23900 3052
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 15016 2796 15068 2848
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 15844 2796 15896 2848
rect 16120 2796 16172 2848
rect 16396 2796 16448 2848
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17592 2839 17644 2848
rect 17592 2805 17601 2839
rect 17601 2805 17635 2839
rect 17635 2805 17644 2839
rect 17592 2796 17644 2805
rect 17868 2839 17920 2848
rect 17868 2805 17877 2839
rect 17877 2805 17911 2839
rect 17911 2805 17920 2839
rect 17868 2796 17920 2805
rect 18328 2796 18380 2848
rect 22192 2864 22244 2916
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 19984 2796 20036 2848
rect 20536 2796 20588 2848
rect 21088 2796 21140 2848
rect 22284 2796 22336 2848
rect 22744 2796 22796 2848
rect 28724 3043 28776 3052
rect 28724 3009 28733 3043
rect 28733 3009 28767 3043
rect 28767 3009 28776 3043
rect 28724 3000 28776 3009
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 29368 3000 29420 3052
rect 30472 3000 30524 3052
rect 31944 3000 31996 3052
rect 32772 3043 32824 3052
rect 32772 3009 32781 3043
rect 32781 3009 32815 3043
rect 32815 3009 32824 3043
rect 32772 3000 32824 3009
rect 33692 3000 33744 3052
rect 34520 3000 34572 3052
rect 35440 3068 35492 3120
rect 35532 3000 35584 3052
rect 36268 3068 36320 3120
rect 26608 2932 26660 2984
rect 27620 2932 27672 2984
rect 24860 2864 24912 2916
rect 25412 2864 25464 2916
rect 26148 2864 26200 2916
rect 26884 2864 26936 2916
rect 33048 2932 33100 2984
rect 34888 2932 34940 2984
rect 35716 2932 35768 2984
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 37648 3000 37700 3052
rect 38016 3000 38068 3052
rect 39028 3000 39080 3052
rect 23848 2796 23900 2848
rect 24400 2796 24452 2848
rect 24952 2796 25004 2848
rect 25504 2796 25556 2848
rect 25964 2796 26016 2848
rect 26516 2796 26568 2848
rect 27988 2864 28040 2916
rect 28540 2864 28592 2916
rect 27804 2796 27856 2848
rect 28816 2796 28868 2848
rect 30196 2864 30248 2916
rect 29828 2796 29880 2848
rect 31300 2864 31352 2916
rect 32404 2864 32456 2916
rect 33508 2864 33560 2916
rect 34612 2864 34664 2916
rect 36176 2864 36228 2916
rect 36360 2907 36412 2916
rect 36360 2873 36369 2907
rect 36369 2873 36403 2907
rect 36403 2873 36412 2907
rect 36360 2864 36412 2873
rect 36636 2907 36688 2916
rect 36636 2873 36645 2907
rect 36645 2873 36679 2907
rect 36679 2873 36688 2907
rect 36636 2864 36688 2873
rect 34796 2796 34848 2848
rect 35900 2839 35952 2848
rect 35900 2805 35909 2839
rect 35909 2805 35943 2839
rect 35943 2805 35952 2839
rect 35900 2796 35952 2805
rect 40040 2796 40092 2848
rect 6251 2694 6303 2746
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 16854 2694 16906 2746
rect 16918 2694 16970 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 27457 2694 27509 2746
rect 27521 2694 27573 2746
rect 27585 2694 27637 2746
rect 27649 2694 27701 2746
rect 27713 2694 27765 2746
rect 38060 2694 38112 2746
rect 38124 2694 38176 2746
rect 38188 2694 38240 2746
rect 38252 2694 38304 2746
rect 38316 2694 38368 2746
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 7472 2524 7524 2576
rect 8208 2524 8260 2576
rect 9312 2592 9364 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 10968 2592 11020 2644
rect 11336 2635 11388 2644
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 8944 2524 8996 2576
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5632 2388 5684 2440
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6736 2320 6788 2372
rect 7104 2388 7156 2440
rect 7012 2320 7064 2372
rect 7656 2388 7708 2440
rect 8116 2456 8168 2508
rect 10416 2524 10468 2576
rect 11428 2524 11480 2576
rect 12716 2592 12768 2644
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 12256 2567 12308 2576
rect 12256 2533 12265 2567
rect 12265 2533 12299 2567
rect 12299 2533 12308 2567
rect 12256 2524 12308 2533
rect 14648 2635 14700 2644
rect 14648 2601 14657 2635
rect 14657 2601 14691 2635
rect 14691 2601 14700 2635
rect 14648 2592 14700 2601
rect 12164 2456 12216 2508
rect 13452 2524 13504 2576
rect 13636 2524 13688 2576
rect 15200 2592 15252 2644
rect 7564 2320 7616 2372
rect 8484 2388 8536 2440
rect 8852 2388 8904 2440
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 9404 2388 9456 2440
rect 9588 2388 9640 2440
rect 9956 2388 10008 2440
rect 10232 2388 10284 2440
rect 10508 2388 10560 2440
rect 10784 2388 10836 2440
rect 11060 2388 11112 2440
rect 11428 2388 11480 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11980 2388 12032 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 8392 2320 8444 2372
rect 5356 2295 5408 2304
rect 5356 2261 5365 2295
rect 5365 2261 5399 2295
rect 5399 2261 5408 2295
rect 5356 2252 5408 2261
rect 5908 2295 5960 2304
rect 5908 2261 5917 2295
rect 5917 2261 5951 2295
rect 5951 2261 5960 2295
rect 5908 2252 5960 2261
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 6920 2252 6972 2304
rect 7288 2252 7340 2304
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 9588 2252 9640 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10416 2320 10468 2372
rect 11244 2320 11296 2372
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 14464 2456 14516 2508
rect 15016 2524 15068 2576
rect 16120 2524 16172 2576
rect 17684 2524 17736 2576
rect 13820 2320 13872 2372
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 14740 2320 14792 2372
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17316 2456 17368 2508
rect 17592 2388 17644 2440
rect 15568 2320 15620 2372
rect 12532 2295 12584 2304
rect 12532 2261 12541 2295
rect 12541 2261 12575 2295
rect 12575 2261 12584 2295
rect 12532 2252 12584 2261
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 13912 2295 13964 2304
rect 13912 2261 13921 2295
rect 13921 2261 13955 2295
rect 13955 2261 13964 2295
rect 13912 2252 13964 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 15384 2295 15436 2304
rect 15384 2261 15393 2295
rect 15393 2261 15427 2295
rect 15427 2261 15436 2295
rect 15384 2252 15436 2261
rect 15844 2252 15896 2304
rect 17316 2320 17368 2372
rect 16396 2252 16448 2304
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 17132 2295 17184 2304
rect 17132 2261 17141 2295
rect 17141 2261 17175 2295
rect 17175 2261 17184 2295
rect 17132 2252 17184 2261
rect 17408 2295 17460 2304
rect 17408 2261 17417 2295
rect 17417 2261 17451 2295
rect 17451 2261 17460 2295
rect 17408 2252 17460 2261
rect 17592 2252 17644 2304
rect 17868 2388 17920 2440
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 18972 2592 19024 2644
rect 19340 2592 19392 2644
rect 19248 2524 19300 2576
rect 19156 2456 19208 2508
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19340 2320 19392 2372
rect 20076 2320 20128 2372
rect 18972 2252 19024 2304
rect 21824 2524 21876 2576
rect 20628 2388 20680 2440
rect 22560 2456 22612 2508
rect 20904 2388 20956 2440
rect 21824 2388 21876 2440
rect 22284 2388 22336 2440
rect 23480 2431 23532 2440
rect 23480 2397 23489 2431
rect 23489 2397 23523 2431
rect 23523 2397 23532 2431
rect 23480 2388 23532 2397
rect 23940 2388 23992 2440
rect 24032 2388 24084 2440
rect 24308 2388 24360 2440
rect 25320 2499 25372 2508
rect 25320 2465 25329 2499
rect 25329 2465 25363 2499
rect 25363 2465 25372 2499
rect 25320 2456 25372 2465
rect 26148 2592 26200 2644
rect 26608 2635 26660 2644
rect 26608 2601 26617 2635
rect 26617 2601 26651 2635
rect 26651 2601 26660 2635
rect 26608 2592 26660 2601
rect 26792 2592 26844 2644
rect 28724 2592 28776 2644
rect 29644 2592 29696 2644
rect 31760 2635 31812 2644
rect 31760 2601 31769 2635
rect 31769 2601 31803 2635
rect 31803 2601 31812 2635
rect 31760 2592 31812 2601
rect 28908 2524 28960 2576
rect 31024 2524 31076 2576
rect 33416 2592 33468 2644
rect 33324 2524 33376 2576
rect 35532 2592 35584 2644
rect 35808 2635 35860 2644
rect 35808 2601 35817 2635
rect 35817 2601 35851 2635
rect 35851 2601 35860 2635
rect 35808 2592 35860 2601
rect 35992 2592 36044 2644
rect 37004 2635 37056 2644
rect 37004 2601 37013 2635
rect 37013 2601 37047 2635
rect 37047 2601 37056 2635
rect 37004 2592 37056 2601
rect 37832 2592 37884 2644
rect 38384 2592 38436 2644
rect 38660 2635 38712 2644
rect 38660 2601 38669 2635
rect 38669 2601 38703 2635
rect 38703 2601 38712 2635
rect 38660 2592 38712 2601
rect 39948 2592 40000 2644
rect 41512 2592 41564 2644
rect 42432 2635 42484 2644
rect 42432 2601 42441 2635
rect 42441 2601 42475 2635
rect 42475 2601 42484 2635
rect 42432 2592 42484 2601
rect 37372 2524 37424 2576
rect 21364 2320 21416 2372
rect 21916 2320 21968 2372
rect 22652 2320 22704 2372
rect 20628 2252 20680 2304
rect 20812 2252 20864 2304
rect 25136 2388 25188 2440
rect 26240 2388 26292 2440
rect 26424 2388 26476 2440
rect 27712 2456 27764 2508
rect 29460 2388 29512 2440
rect 29736 2388 29788 2440
rect 30840 2388 30892 2440
rect 27804 2320 27856 2372
rect 27896 2320 27948 2372
rect 28356 2320 28408 2372
rect 29000 2320 29052 2372
rect 29920 2320 29972 2372
rect 33140 2456 33192 2508
rect 34428 2456 34480 2508
rect 32220 2363 32272 2372
rect 32220 2329 32229 2363
rect 32229 2329 32263 2363
rect 32263 2329 32272 2363
rect 32220 2320 32272 2329
rect 33232 2320 33284 2372
rect 34060 2388 34112 2440
rect 35900 2388 35952 2440
rect 36084 2456 36136 2508
rect 36176 2388 36228 2440
rect 36728 2431 36780 2440
rect 36728 2397 36737 2431
rect 36737 2397 36771 2431
rect 36771 2397 36780 2431
rect 36728 2388 36780 2397
rect 36912 2456 36964 2508
rect 34704 2320 34756 2372
rect 34796 2363 34848 2372
rect 34796 2329 34805 2363
rect 34805 2329 34839 2363
rect 34839 2329 34848 2363
rect 34796 2320 34848 2329
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 23296 2252 23348 2304
rect 23756 2252 23808 2304
rect 24676 2252 24728 2304
rect 26332 2252 26384 2304
rect 27528 2252 27580 2304
rect 28448 2252 28500 2304
rect 30104 2252 30156 2304
rect 32312 2252 32364 2304
rect 33416 2295 33468 2304
rect 33416 2261 33425 2295
rect 33425 2261 33459 2295
rect 33459 2261 33468 2295
rect 33416 2252 33468 2261
rect 33968 2295 34020 2304
rect 33968 2261 33977 2295
rect 33977 2261 34011 2295
rect 34011 2261 34020 2295
rect 33968 2252 34020 2261
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36636 2320 36688 2372
rect 37188 2320 37240 2372
rect 38936 2388 38988 2440
rect 39396 2431 39448 2440
rect 39396 2397 39405 2431
rect 39405 2397 39439 2431
rect 39439 2397 39448 2431
rect 39396 2388 39448 2397
rect 39672 2431 39724 2440
rect 39672 2397 39681 2431
rect 39681 2397 39715 2431
rect 39715 2397 39724 2431
rect 39672 2388 39724 2397
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 40316 2431 40368 2440
rect 40316 2397 40325 2431
rect 40325 2397 40359 2431
rect 40359 2397 40368 2431
rect 40316 2388 40368 2397
rect 36360 2252 36412 2304
rect 37740 2295 37792 2304
rect 37740 2261 37749 2295
rect 37749 2261 37783 2295
rect 37783 2261 37792 2295
rect 37740 2252 37792 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38384 2295 38436 2304
rect 38384 2261 38393 2295
rect 38393 2261 38427 2295
rect 38427 2261 38436 2295
rect 38384 2252 38436 2261
rect 39948 2320 40000 2372
rect 11552 2150 11604 2202
rect 11616 2150 11668 2202
rect 11680 2150 11732 2202
rect 11744 2150 11796 2202
rect 11808 2150 11860 2202
rect 22155 2150 22207 2202
rect 22219 2150 22271 2202
rect 22283 2150 22335 2202
rect 22347 2150 22399 2202
rect 22411 2150 22463 2202
rect 32758 2150 32810 2202
rect 32822 2150 32874 2202
rect 32886 2150 32938 2202
rect 32950 2150 33002 2202
rect 33014 2150 33066 2202
rect 43361 2150 43413 2202
rect 43425 2150 43477 2202
rect 43489 2150 43541 2202
rect 43553 2150 43605 2202
rect 43617 2150 43669 2202
rect 5908 2048 5960 2100
rect 7932 2048 7984 2100
rect 6828 1980 6880 2032
rect 9956 2048 10008 2100
rect 13268 2048 13320 2100
rect 13360 2048 13412 2100
rect 15016 2048 15068 2100
rect 17408 2048 17460 2100
rect 20812 2048 20864 2100
rect 22928 2048 22980 2100
rect 24860 2048 24912 2100
rect 29920 2048 29972 2100
rect 31576 2048 31628 2100
rect 33416 2048 33468 2100
rect 37464 2048 37516 2100
rect 38384 2048 38436 2100
rect 23388 1980 23440 2032
rect 37740 1980 37792 2032
rect 14280 1912 14332 1964
rect 23112 1912 23164 1964
rect 24124 1912 24176 1964
rect 25320 1912 25372 1964
rect 35440 1912 35492 1964
rect 36360 1912 36412 1964
rect 7288 1776 7340 1828
rect 17592 1776 17644 1828
rect 18052 1776 18104 1828
rect 20996 1776 21048 1828
rect 33876 1776 33928 1828
rect 38292 1776 38344 1828
rect 7380 1640 7432 1692
rect 7472 1640 7524 1692
rect 9404 1708 9456 1760
rect 12992 1708 13044 1760
rect 13912 1708 13964 1760
rect 9864 1640 9916 1692
rect 12716 1640 12768 1692
rect 29460 1708 29512 1760
rect 26424 1640 26476 1692
rect 14924 1572 14976 1624
rect 15108 1572 15160 1624
rect 15660 1572 15712 1624
rect 16120 1572 16172 1624
rect 22836 1504 22888 1556
rect 38752 1504 38804 1556
rect 39672 1504 39724 1556
rect 5356 1436 5408 1488
rect 10692 1436 10744 1488
rect 12532 1436 12584 1488
rect 26700 1436 26752 1488
rect 32220 1436 32272 1488
rect 33968 1436 34020 1488
rect 13268 1368 13320 1420
rect 14556 1368 14608 1420
rect 15108 1368 15160 1420
rect 19064 1368 19116 1420
rect 31208 1368 31260 1420
rect 32312 1368 32364 1420
rect 35624 1368 35676 1420
rect 36728 1368 36780 1420
rect 18052 1300 18104 1352
rect 21272 1300 21324 1352
rect 38568 1300 38620 1352
rect 39396 1436 39448 1488
rect 39304 1368 39356 1420
rect 40316 1368 40368 1420
rect 6552 1232 6604 1284
rect 24032 1232 24084 1284
rect 16488 1164 16540 1216
rect 33232 1164 33284 1216
rect 15016 1096 15068 1148
rect 25688 1096 25740 1148
rect 9680 1028 9732 1080
rect 21456 1028 21508 1080
rect 21824 1028 21876 1080
rect 9864 960 9916 1012
rect 15844 892 15896 944
rect 33692 892 33744 944
<< metal2 >>
rect 1122 9840 1178 10300
rect 3238 9840 3294 10300
rect 5354 9840 5410 10300
rect 7470 9840 7526 10300
rect 9586 9840 9642 10300
rect 11702 9840 11758 10300
rect 11808 9846 12020 9874
rect 1136 7546 1164 9840
rect 3252 9602 3280 9840
rect 3252 9574 3464 9602
rect 3436 7546 3464 9574
rect 5368 7546 5396 9840
rect 7484 7546 7512 9840
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 9600 7426 9628 9840
rect 11716 9738 11744 9840
rect 11808 9738 11836 9846
rect 11716 9710 11836 9738
rect 11552 7644 11860 7653
rect 11552 7642 11558 7644
rect 11614 7642 11638 7644
rect 11694 7642 11718 7644
rect 11774 7642 11798 7644
rect 11854 7642 11860 7644
rect 11614 7590 11616 7642
rect 11796 7590 11798 7642
rect 11552 7588 11558 7590
rect 11614 7588 11638 7590
rect 11694 7588 11718 7590
rect 11774 7588 11798 7590
rect 11854 7588 11860 7590
rect 11552 7579 11860 7588
rect 11992 7546 12020 9846
rect 13818 9840 13874 10300
rect 15934 9840 15990 10300
rect 18050 9840 18106 10300
rect 20166 9840 20222 10300
rect 20272 9846 20576 9874
rect 13832 7546 13860 9840
rect 15948 7546 15976 9840
rect 18064 7546 18092 9840
rect 20180 9738 20208 9840
rect 20272 9738 20300 9846
rect 20180 9710 20300 9738
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 9692 7426 9720 7482
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7656 7404 7708 7410
rect 9600 7398 9720 7426
rect 20548 7410 20576 9846
rect 22282 9840 22338 10300
rect 22388 9846 22600 9874
rect 22296 9738 22324 9840
rect 22388 9738 22416 9846
rect 22296 9710 22416 9738
rect 22155 7644 22463 7653
rect 22155 7642 22161 7644
rect 22217 7642 22241 7644
rect 22297 7642 22321 7644
rect 22377 7642 22401 7644
rect 22457 7642 22463 7644
rect 22217 7590 22219 7642
rect 22399 7590 22401 7642
rect 22155 7588 22161 7590
rect 22217 7588 22241 7590
rect 22297 7588 22321 7590
rect 22377 7588 22401 7590
rect 22457 7588 22463 7590
rect 22155 7579 22463 7588
rect 22572 7546 22600 9846
rect 24398 9840 24454 10300
rect 24504 9846 24808 9874
rect 24412 9738 24440 9840
rect 24504 9738 24532 9846
rect 24412 9710 24532 9738
rect 24780 8242 24808 9846
rect 26514 9840 26570 10300
rect 28630 9840 28686 10300
rect 30746 9840 30802 10300
rect 32862 9840 32918 10300
rect 34978 9840 35034 10300
rect 37094 9840 37150 10300
rect 39210 9840 39266 10300
rect 41326 9840 41382 10300
rect 43442 9840 43498 10300
rect 24780 8214 24900 8242
rect 24872 7546 24900 8214
rect 26528 7546 26556 9840
rect 28644 8514 28672 9840
rect 28644 8486 28856 8514
rect 28828 7546 28856 8486
rect 30760 7546 30788 9840
rect 32876 8242 32904 9840
rect 32876 8214 33180 8242
rect 32758 7644 33066 7653
rect 32758 7642 32764 7644
rect 32820 7642 32844 7644
rect 32900 7642 32924 7644
rect 32980 7642 33004 7644
rect 33060 7642 33066 7644
rect 32820 7590 32822 7642
rect 33002 7590 33004 7642
rect 32758 7588 32764 7590
rect 32820 7588 32844 7590
rect 32900 7588 32924 7590
rect 32980 7588 33004 7590
rect 33060 7588 33066 7590
rect 32758 7579 33066 7588
rect 33152 7546 33180 8214
rect 34992 7546 35020 9840
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 34980 7540 35032 7546
rect 37108 7528 37136 9840
rect 37188 7540 37240 7546
rect 37108 7500 37188 7528
rect 34980 7482 35032 7488
rect 39224 7528 39252 9840
rect 39304 7540 39356 7546
rect 39224 7500 39304 7528
rect 37188 7482 37240 7488
rect 39304 7482 39356 7488
rect 41340 7426 41368 9840
rect 43456 8242 43484 9840
rect 43272 8214 43484 8242
rect 43272 7546 43300 8214
rect 43361 7644 43669 7653
rect 43361 7642 43367 7644
rect 43423 7642 43447 7644
rect 43503 7642 43527 7644
rect 43583 7642 43607 7644
rect 43663 7642 43669 7644
rect 43423 7590 43425 7642
rect 43605 7590 43607 7642
rect 43361 7588 43367 7590
rect 43423 7588 43447 7590
rect 43503 7588 43527 7590
rect 43583 7588 43607 7590
rect 43663 7588 43669 7590
rect 43361 7579 43669 7588
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 43260 7540 43312 7546
rect 43260 7482 43312 7488
rect 41432 7426 41460 7482
rect 14188 7404 14240 7410
rect 7656 7346 7708 7352
rect 14188 7346 14240 7352
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 39948 7404 40000 7410
rect 41340 7398 41460 7426
rect 41512 7404 41564 7410
rect 39948 7346 40000 7352
rect 41512 7346 41564 7352
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 1504 6186 1532 7346
rect 6251 7100 6559 7109
rect 6251 7098 6257 7100
rect 6313 7098 6337 7100
rect 6393 7098 6417 7100
rect 6473 7098 6497 7100
rect 6553 7098 6559 7100
rect 6313 7046 6315 7098
rect 6495 7046 6497 7098
rect 6251 7044 6257 7046
rect 6313 7044 6337 7046
rect 6393 7044 6417 7046
rect 6473 7044 6497 7046
rect 6553 7044 6559 7046
rect 6251 7035 6559 7044
rect 1492 6180 1544 6186
rect 1492 6122 1544 6128
rect 6251 6012 6559 6021
rect 6251 6010 6257 6012
rect 6313 6010 6337 6012
rect 6393 6010 6417 6012
rect 6473 6010 6497 6012
rect 6553 6010 6559 6012
rect 6313 5958 6315 6010
rect 6495 5958 6497 6010
rect 6251 5956 6257 5958
rect 6313 5956 6337 5958
rect 6393 5956 6417 5958
rect 6473 5956 6497 5958
rect 6553 5956 6559 5958
rect 6251 5947 6559 5956
rect 6251 4924 6559 4933
rect 6251 4922 6257 4924
rect 6313 4922 6337 4924
rect 6393 4922 6417 4924
rect 6473 4922 6497 4924
rect 6553 4922 6559 4924
rect 6313 4870 6315 4922
rect 6495 4870 6497 4922
rect 6251 4868 6257 4870
rect 6313 4868 6337 4870
rect 6393 4868 6417 4870
rect 6473 4868 6497 4870
rect 6553 4868 6559 4870
rect 6251 4859 6559 4868
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6251 3836 6559 3845
rect 6251 3834 6257 3836
rect 6313 3834 6337 3836
rect 6393 3834 6417 3836
rect 6473 3834 6497 3836
rect 6553 3834 6559 3836
rect 6313 3782 6315 3834
rect 6495 3782 6497 3834
rect 6251 3780 6257 3782
rect 6313 3780 6337 3782
rect 6393 3780 6417 3782
rect 6473 3780 6497 3782
rect 6553 3780 6559 3782
rect 6251 3771 6559 3780
rect 6748 3194 6776 4626
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 5078 2952 5134 2961
rect 6564 2938 6592 2994
rect 6564 2910 6684 2938
rect 5078 2887 5134 2896
rect 5092 2650 5120 2887
rect 6251 2748 6559 2757
rect 6251 2746 6257 2748
rect 6313 2746 6337 2748
rect 6393 2746 6417 2748
rect 6473 2746 6497 2748
rect 6553 2746 6559 2748
rect 6313 2694 6315 2746
rect 6495 2694 6497 2746
rect 6251 2692 6257 2694
rect 6313 2692 6337 2694
rect 6393 2692 6417 2694
rect 6473 2692 6497 2694
rect 6553 2692 6559 2694
rect 6251 2683 6559 2692
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 4908 82 4936 2382
rect 5078 82 5134 160
rect 4908 54 5134 82
rect 5184 82 5212 2382
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5368 1494 5396 2246
rect 5356 1488 5408 1494
rect 5356 1430 5408 1436
rect 5644 160 5672 2382
rect 5354 82 5410 160
rect 5184 54 5410 82
rect 5078 -300 5134 54
rect 5354 -300 5410 54
rect 5630 -300 5686 160
rect 5736 82 5764 2382
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 2106 5948 2246
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 5906 82 5962 160
rect 5736 54 5962 82
rect 6012 82 6040 2382
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 1290 6592 2246
rect 6552 1284 6604 1290
rect 6552 1226 6604 1232
rect 6182 82 6238 160
rect 6012 54 6238 82
rect 5906 -300 5962 54
rect 6182 -300 6238 54
rect 6458 82 6514 160
rect 6656 82 6684 2910
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 160 6776 2314
rect 6840 2038 6868 7346
rect 7668 7002 7696 7346
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 11552 6556 11860 6565
rect 11552 6554 11558 6556
rect 11614 6554 11638 6556
rect 11694 6554 11718 6556
rect 11774 6554 11798 6556
rect 11854 6554 11860 6556
rect 11614 6502 11616 6554
rect 11796 6502 11798 6554
rect 11552 6500 11558 6502
rect 11614 6500 11638 6502
rect 11694 6500 11718 6502
rect 11774 6500 11798 6502
rect 11854 6500 11860 6502
rect 11552 6491 11860 6500
rect 11552 5468 11860 5477
rect 11552 5466 11558 5468
rect 11614 5466 11638 5468
rect 11694 5466 11718 5468
rect 11774 5466 11798 5468
rect 11854 5466 11860 5468
rect 11614 5414 11616 5466
rect 11796 5414 11798 5466
rect 11552 5412 11558 5414
rect 11614 5412 11638 5414
rect 11694 5412 11718 5414
rect 11774 5412 11798 5414
rect 11854 5412 11860 5414
rect 11552 5403 11860 5412
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8772 2774 8800 4558
rect 8404 2746 8800 2774
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 8208 2576 8260 2582
rect 8404 2530 8432 2746
rect 8956 2582 8984 4694
rect 9310 3496 9366 3505
rect 9310 3431 9366 3440
rect 9324 2650 9352 3431
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 8260 2524 8432 2530
rect 8208 2518 8432 2524
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 6932 921 6960 2246
rect 6918 912 6974 921
rect 6918 847 6974 856
rect 7024 160 7052 2314
rect 6458 54 6684 82
rect 6458 -300 6514 54
rect 6734 -300 6790 160
rect 7010 -300 7066 160
rect 7116 82 7144 2382
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7300 1834 7328 2246
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 7392 1698 7420 2246
rect 7484 1698 7512 2518
rect 8116 2508 8168 2514
rect 8220 2502 8432 2518
rect 8116 2450 8168 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7380 1692 7432 1698
rect 7380 1634 7432 1640
rect 7472 1692 7524 1698
rect 7472 1634 7524 1640
rect 7576 160 7604 2314
rect 7286 82 7342 160
rect 7116 54 7342 82
rect 7286 -300 7342 54
rect 7562 -300 7618 160
rect 7668 82 7696 2382
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 2106 7972 2246
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8128 160 8156 2450
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8944 2440 8996 2446
rect 9404 2440 9456 2446
rect 8996 2400 9260 2428
rect 8944 2382 8996 2388
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 160 8432 2314
rect 7838 82 7894 160
rect 7668 54 7894 82
rect 7838 -300 7894 54
rect 8114 -300 8170 160
rect 8390 -300 8446 160
rect 8496 82 8524 2382
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 1737 8800 2246
rect 8758 1728 8814 1737
rect 8758 1663 8814 1672
rect 8864 1306 8892 2382
rect 8864 1278 8984 1306
rect 8956 160 8984 1278
rect 9232 160 9260 2400
rect 9588 2440 9640 2446
rect 9456 2400 9536 2428
rect 9404 2382 9456 2388
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 1766 9444 2246
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 9508 160 9536 2400
rect 9956 2440 10008 2446
rect 9640 2400 9812 2428
rect 9588 2382 9640 2388
rect 9588 2304 9640 2310
rect 9640 2264 9720 2292
rect 9588 2246 9640 2252
rect 9692 1086 9720 2264
rect 9680 1080 9732 1086
rect 9680 1022 9732 1028
rect 9784 160 9812 2400
rect 10232 2440 10284 2446
rect 10008 2400 10088 2428
rect 9956 2382 10008 2388
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 2106 9996 2246
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 9864 1692 9916 1698
rect 9864 1634 9916 1640
rect 9876 1018 9904 1634
rect 9864 1012 9916 1018
rect 9864 954 9916 960
rect 10060 160 10088 2400
rect 10284 2400 10364 2428
rect 10232 2382 10284 2388
rect 10336 160 10364 2400
rect 10428 2378 10456 2518
rect 10508 2440 10560 2446
rect 10560 2400 10640 2428
rect 10508 2382 10560 2388
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10612 160 10640 2400
rect 10704 1494 10732 4762
rect 13450 4584 13506 4593
rect 13450 4519 13506 4528
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10782 3088 10838 3097
rect 10782 3023 10838 3032
rect 10796 2650 10824 3023
rect 10980 2650 11008 4422
rect 11552 4380 11860 4389
rect 11552 4378 11558 4380
rect 11614 4378 11638 4380
rect 11694 4378 11718 4380
rect 11774 4378 11798 4380
rect 11854 4378 11860 4380
rect 11614 4326 11616 4378
rect 11796 4326 11798 4378
rect 11552 4324 11558 4326
rect 11614 4324 11638 4326
rect 11694 4324 11718 4326
rect 11774 4324 11798 4326
rect 11854 4324 11860 4326
rect 11552 4315 11860 4324
rect 12990 4312 13046 4321
rect 12990 4247 13046 4256
rect 12806 4040 12862 4049
rect 12806 3975 12862 3984
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10784 2440 10836 2446
rect 11060 2440 11112 2446
rect 10836 2400 10916 2428
rect 10784 2382 10836 2388
rect 10692 1488 10744 1494
rect 10692 1430 10744 1436
rect 10888 160 10916 2400
rect 11112 2400 11192 2428
rect 11060 2382 11112 2388
rect 11164 160 11192 2400
rect 11256 2378 11284 3878
rect 11334 3632 11390 3641
rect 11334 3567 11390 3576
rect 11348 2650 11376 3567
rect 11552 3292 11860 3301
rect 11552 3290 11558 3292
rect 11614 3290 11638 3292
rect 11694 3290 11718 3292
rect 11774 3290 11798 3292
rect 11854 3290 11860 3292
rect 11614 3238 11616 3290
rect 11796 3238 11798 3290
rect 11552 3236 11558 3238
rect 11614 3236 11638 3238
rect 11694 3236 11718 3238
rect 11774 3236 11798 3238
rect 11854 3236 11860 3238
rect 11552 3227 11860 3236
rect 12254 3224 12310 3233
rect 12176 3182 12254 3210
rect 12176 2774 12204 3182
rect 12254 3159 12310 3168
rect 12176 2746 12296 2774
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 12268 2582 12296 2746
rect 12820 2650 12848 3975
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 11428 2576 11480 2582
rect 11348 2524 11428 2530
rect 11348 2518 11480 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 11348 2502 11468 2518
rect 12164 2508 12216 2514
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11348 2009 11376 2502
rect 12164 2450 12216 2456
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11520 2440 11572 2446
rect 11980 2440 12032 2446
rect 11572 2400 11928 2428
rect 11520 2382 11572 2388
rect 11334 2000 11390 2009
rect 11334 1935 11390 1944
rect 11440 160 11468 2382
rect 11552 2204 11860 2213
rect 11552 2202 11558 2204
rect 11614 2202 11638 2204
rect 11694 2202 11718 2204
rect 11774 2202 11798 2204
rect 11854 2202 11860 2204
rect 11614 2150 11616 2202
rect 11796 2150 11798 2202
rect 11552 2148 11558 2150
rect 11614 2148 11638 2150
rect 11694 2148 11718 2150
rect 11774 2148 11798 2150
rect 11854 2148 11860 2150
rect 11552 2139 11860 2148
rect 8666 82 8722 160
rect 8496 54 8722 82
rect 8666 -300 8722 54
rect 8942 -300 8998 160
rect 9218 -300 9274 160
rect 9494 -300 9550 160
rect 9770 -300 9826 160
rect 10046 -300 10102 160
rect 10322 -300 10378 160
rect 10598 -300 10654 160
rect 10874 -300 10930 160
rect 11150 -300 11206 160
rect 11426 -300 11482 160
rect 11702 82 11758 160
rect 11900 82 11928 2400
rect 11980 2382 12032 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11992 160 12020 2382
rect 11702 54 11928 82
rect 11702 -300 11758 54
rect 11978 -300 12034 160
rect 12084 82 12112 2382
rect 12176 2145 12204 2450
rect 12348 2440 12400 2446
rect 12624 2440 12676 2446
rect 12400 2400 12480 2428
rect 12348 2382 12400 2388
rect 12162 2136 12218 2145
rect 12162 2071 12218 2080
rect 12254 82 12310 160
rect 12084 54 12310 82
rect 12452 82 12480 2400
rect 12624 2382 12676 2388
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12544 1494 12572 2246
rect 12532 1488 12584 1494
rect 12532 1430 12584 1436
rect 12530 82 12586 160
rect 12452 54 12586 82
rect 12636 82 12664 2382
rect 12728 1698 12756 2586
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12716 1692 12768 1698
rect 12716 1634 12768 1640
rect 12806 82 12862 160
rect 12636 54 12862 82
rect 12912 82 12940 2382
rect 13004 1766 13032 4247
rect 13464 2582 13492 4519
rect 14200 3194 14228 7346
rect 16132 5370 16160 7346
rect 16854 7100 17162 7109
rect 16854 7098 16860 7100
rect 16916 7098 16940 7100
rect 16996 7098 17020 7100
rect 17076 7098 17100 7100
rect 17156 7098 17162 7100
rect 16916 7046 16918 7098
rect 17098 7046 17100 7098
rect 16854 7044 16860 7046
rect 16916 7044 16940 7046
rect 16996 7044 17020 7046
rect 17076 7044 17100 7046
rect 17156 7044 17162 7046
rect 16854 7035 17162 7044
rect 18892 6254 18920 7346
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20456 7188 20484 7278
rect 20536 7200 20588 7206
rect 20456 7160 20536 7188
rect 20536 7142 20588 7148
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 16854 6012 17162 6021
rect 16854 6010 16860 6012
rect 16916 6010 16940 6012
rect 16996 6010 17020 6012
rect 17076 6010 17100 6012
rect 17156 6010 17162 6012
rect 16916 5958 16918 6010
rect 17098 5958 17100 6010
rect 16854 5956 16860 5958
rect 16916 5956 16940 5958
rect 16996 5956 17020 5958
rect 17076 5956 17100 5958
rect 17156 5956 17162 5958
rect 16854 5947 17162 5956
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16488 5160 16540 5166
rect 16486 5128 16488 5137
rect 16540 5128 16542 5137
rect 16486 5063 16542 5072
rect 16854 4924 17162 4933
rect 16854 4922 16860 4924
rect 16916 4922 16940 4924
rect 16996 4922 17020 4924
rect 17076 4922 17100 4924
rect 17156 4922 17162 4924
rect 16916 4870 16918 4922
rect 17098 4870 17100 4922
rect 16854 4868 16860 4870
rect 16916 4868 16940 4870
rect 16996 4868 17020 4870
rect 17076 4868 17100 4870
rect 17156 4868 17162 4870
rect 16854 4859 17162 4868
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14292 3058 14320 4150
rect 15120 3194 15148 4218
rect 15672 3194 15700 4490
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 16854 3836 17162 3845
rect 16854 3834 16860 3836
rect 16916 3834 16940 3836
rect 16996 3834 17020 3836
rect 17076 3834 17100 3836
rect 17156 3834 17162 3836
rect 16916 3782 16918 3834
rect 17098 3782 17100 3834
rect 16854 3780 16860 3782
rect 16916 3780 16940 3782
rect 16996 3780 17020 3782
rect 17076 3780 17100 3782
rect 17156 3780 17162 3782
rect 16854 3771 17162 3780
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15016 3120 15068 3126
rect 15396 3097 15424 3130
rect 15016 3062 15068 3068
rect 15382 3088 15438 3097
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 13452 2576 13504 2582
rect 13636 2576 13688 2582
rect 13452 2518 13504 2524
rect 13634 2544 13636 2553
rect 13688 2544 13690 2553
rect 13634 2479 13690 2488
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 13096 1601 13124 2246
rect 13082 1592 13138 1601
rect 13082 1527 13138 1536
rect 13082 82 13138 160
rect 12912 54 13138 82
rect 13188 82 13216 2382
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13372 2106 13400 2246
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13280 1426 13308 2042
rect 13648 1873 13676 2246
rect 13634 1864 13690 1873
rect 13634 1799 13690 1808
rect 13268 1420 13320 1426
rect 13268 1362 13320 1368
rect 13358 82 13414 160
rect 13188 54 13414 82
rect 12254 -300 12310 54
rect 12530 -300 12586 54
rect 12806 -300 12862 54
rect 13082 -300 13138 54
rect 13358 -300 13414 54
rect 13634 82 13690 160
rect 13740 82 13768 2994
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13634 54 13768 82
rect 13832 82 13860 2314
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 13924 1766 13952 2246
rect 14292 1970 14320 2246
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 13912 1760 13964 1766
rect 13912 1702 13964 1708
rect 13910 82 13966 160
rect 13832 54 13966 82
rect 13634 -300 13690 54
rect 13910 -300 13966 54
rect 14186 82 14242 160
rect 14384 82 14412 2994
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14660 2650 14688 2926
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14476 160 14504 2450
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14568 1426 14596 2382
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14752 160 14780 2314
rect 14186 54 14412 82
rect 14186 -300 14242 54
rect 14462 -300 14518 160
rect 14738 -300 14794 160
rect 14844 82 14872 2994
rect 15028 2938 15056 3062
rect 15200 3052 15252 3058
rect 15382 3023 15438 3032
rect 15936 3052 15988 3058
rect 15200 2994 15252 3000
rect 15936 2994 15988 3000
rect 16212 3052 16264 3058
rect 16580 3052 16632 3058
rect 16264 3012 16344 3040
rect 16212 2994 16264 3000
rect 14936 2910 15056 2938
rect 14936 1630 14964 2910
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 2582 15056 2790
rect 15212 2650 15240 2994
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15764 2666 15792 2790
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15488 2638 15792 2666
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15488 2446 15516 2638
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15752 2440 15804 2446
rect 15856 2428 15884 2790
rect 15804 2400 15884 2428
rect 15752 2382 15804 2388
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 14924 1624 14976 1630
rect 14924 1566 14976 1572
rect 15028 1154 15056 2042
rect 15120 1630 15148 2382
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15108 1624 15160 1630
rect 15108 1566 15160 1572
rect 15120 1426 15240 1442
rect 15108 1420 15240 1426
rect 15160 1414 15240 1420
rect 15108 1362 15160 1368
rect 15016 1148 15068 1154
rect 15016 1090 15068 1096
rect 15014 82 15070 160
rect 14844 54 15070 82
rect 15212 82 15240 1414
rect 15396 1329 15424 2246
rect 15382 1320 15438 1329
rect 15382 1255 15438 1264
rect 15580 160 15608 2314
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15660 1624 15712 1630
rect 15660 1566 15712 1572
rect 15290 82 15346 160
rect 15212 54 15346 82
rect 15014 -300 15070 54
rect 15290 -300 15346 54
rect 15566 -300 15622 160
rect 15672 82 15700 1566
rect 15856 950 15884 2246
rect 15844 944 15896 950
rect 15844 886 15896 892
rect 15842 82 15898 160
rect 15672 54 15898 82
rect 15948 82 15976 2994
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 16132 2666 16160 2790
rect 16316 2774 16344 3012
rect 16948 3052 17000 3058
rect 16580 2994 16632 3000
rect 16776 3012 16948 3040
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16040 2638 16160 2666
rect 16224 2746 16344 2774
rect 16040 2446 16068 2638
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16132 1630 16160 2518
rect 16120 1624 16172 1630
rect 16120 1566 16172 1572
rect 16118 82 16174 160
rect 15948 54 16174 82
rect 16224 82 16252 2746
rect 16304 2440 16356 2446
rect 16408 2428 16436 2790
rect 16356 2400 16436 2428
rect 16304 2382 16356 2388
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16408 1193 16436 2246
rect 16500 1222 16528 2246
rect 16592 1442 16620 2994
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16684 2446 16712 2858
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16776 1442 16804 3012
rect 16948 2994 17000 3000
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 16854 2748 17162 2757
rect 16854 2746 16860 2748
rect 16916 2746 16940 2748
rect 16996 2746 17020 2748
rect 17076 2746 17100 2748
rect 17156 2746 17162 2748
rect 16916 2694 16918 2746
rect 17098 2694 17100 2746
rect 16854 2692 16860 2694
rect 16916 2692 16940 2694
rect 16996 2692 17020 2694
rect 17076 2692 17100 2694
rect 17156 2692 17162 2694
rect 16854 2683 17162 2692
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17144 1465 17172 2246
rect 17130 1456 17186 1465
rect 16592 1414 16712 1442
rect 16776 1414 16988 1442
rect 16488 1216 16540 1222
rect 16394 1184 16450 1193
rect 16488 1158 16540 1164
rect 16394 1119 16450 1128
rect 16684 160 16712 1414
rect 16960 160 16988 1414
rect 17130 1391 17186 1400
rect 17236 160 17264 2994
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17328 2514 17356 2790
rect 17420 2553 17448 3674
rect 17696 3058 17724 3946
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18052 3528 18104 3534
rect 17866 3496 17922 3505
rect 17866 3431 17868 3440
rect 17920 3431 17922 3440
rect 17972 3488 18052 3516
rect 17868 3402 17920 3408
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17406 2544 17462 2553
rect 17316 2508 17368 2514
rect 17406 2479 17462 2488
rect 17316 2450 17368 2456
rect 17314 2408 17370 2417
rect 17314 2343 17316 2352
rect 17368 2343 17370 2352
rect 17316 2314 17368 2320
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17420 2106 17448 2246
rect 17408 2100 17460 2106
rect 17408 2042 17460 2048
rect 17512 160 17540 2994
rect 17592 2848 17644 2854
rect 17592 2790 17644 2796
rect 17604 2446 17632 2790
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 1834 17632 2246
rect 17592 1828 17644 1834
rect 17592 1770 17644 1776
rect 17696 1057 17724 2518
rect 17682 1048 17738 1057
rect 17682 983 17738 992
rect 17788 160 17816 2994
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17880 2446 17908 2790
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 16394 82 16450 160
rect 16224 54 16450 82
rect 15842 -300 15898 54
rect 16118 -300 16174 54
rect 16394 -300 16450 54
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 -300 17278 160
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 17972 82 18000 3488
rect 18052 3470 18104 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18052 3052 18104 3058
rect 18104 3012 18276 3040
rect 18052 2994 18104 3000
rect 18052 1828 18104 1834
rect 18052 1770 18104 1776
rect 18064 1358 18092 1770
rect 18248 1442 18276 3012
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18510 2816 18566 2825
rect 18340 2446 18368 2790
rect 18510 2751 18566 2760
rect 18524 2650 18552 2751
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18248 1414 18368 1442
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 18340 160 18368 1414
rect 18616 160 18644 3470
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18708 3194 18736 3334
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18800 1737 18828 3606
rect 19444 3534 19472 4762
rect 20626 4312 20682 4321
rect 20626 4247 20682 4256
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 3534 20116 3878
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20548 3534 20576 3674
rect 20640 3534 20668 4247
rect 20720 3664 20772 3670
rect 20772 3624 20944 3652
rect 20720 3606 20772 3612
rect 20916 3534 20944 3624
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19536 3194 19564 3334
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 18786 1728 18842 1737
rect 18786 1663 18842 1672
rect 18892 160 18920 2926
rect 18984 2650 19012 2994
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18970 2408 19026 2417
rect 18970 2343 19026 2352
rect 18984 2310 19012 2343
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 19076 1426 19104 2926
rect 19260 2582 19288 3130
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2650 19380 2994
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 19168 160 19196 2450
rect 19628 2446 19656 3334
rect 19812 2961 19840 3470
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 19904 3194 19932 3334
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 20364 3126 20392 3334
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 19798 2952 19854 2961
rect 19798 2887 19854 2896
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19352 1170 19380 2314
rect 19444 2145 19472 2382
rect 19430 2136 19486 2145
rect 19430 2071 19486 2080
rect 19352 1142 19472 1170
rect 19444 160 19472 1142
rect 19720 160 19748 2790
rect 19996 160 20024 2790
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 18050 82 18106 160
rect 17972 54 18106 82
rect 18050 -300 18106 54
rect 18326 -300 18382 160
rect 18602 -300 18658 160
rect 18878 -300 18934 160
rect 19154 -300 19210 160
rect 19430 -300 19486 160
rect 19706 -300 19762 160
rect 19982 -300 20038 160
rect 20088 82 20116 2314
rect 20548 160 20576 2790
rect 20640 2446 20668 3334
rect 20916 2446 20944 3334
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20628 2304 20680 2310
rect 20812 2304 20864 2310
rect 20680 2264 20760 2292
rect 20628 2246 20680 2252
rect 20258 82 20314 160
rect 20088 54 20314 82
rect 20258 -300 20314 54
rect 20534 -300 20590 160
rect 20732 82 20760 2264
rect 20812 2246 20864 2252
rect 20824 2106 20852 2246
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 21008 1834 21036 7346
rect 22480 6934 22508 7346
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22155 6556 22463 6565
rect 22155 6554 22161 6556
rect 22217 6554 22241 6556
rect 22297 6554 22321 6556
rect 22377 6554 22401 6556
rect 22457 6554 22463 6556
rect 22217 6502 22219 6554
rect 22399 6502 22401 6554
rect 22155 6500 22161 6502
rect 22217 6500 22241 6502
rect 22297 6500 22321 6502
rect 22377 6500 22401 6502
rect 22457 6500 22463 6502
rect 22155 6491 22463 6500
rect 22940 6322 22968 7346
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 22155 5468 22463 5477
rect 22155 5466 22161 5468
rect 22217 5466 22241 5468
rect 22297 5466 22321 5468
rect 22377 5466 22401 5468
rect 22457 5466 22463 5468
rect 22217 5414 22219 5466
rect 22399 5414 22401 5466
rect 22155 5412 22161 5414
rect 22217 5412 22241 5414
rect 22297 5412 22321 5414
rect 22377 5412 22401 5414
rect 22457 5412 22463 5414
rect 22155 5403 22463 5412
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22155 4380 22463 4389
rect 22155 4378 22161 4380
rect 22217 4378 22241 4380
rect 22297 4378 22321 4380
rect 22377 4378 22401 4380
rect 22457 4378 22463 4380
rect 22217 4326 22219 4378
rect 22399 4326 22401 4378
rect 22155 4324 22161 4326
rect 22217 4324 22241 4326
rect 22297 4324 22321 4326
rect 22377 4324 22401 4326
rect 22457 4324 22463 4326
rect 22155 4315 22463 4324
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22112 3942 22140 3975
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21192 3194 21220 3334
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 20996 1828 21048 1834
rect 20996 1770 21048 1776
rect 21100 160 21128 2790
rect 21284 1358 21312 3674
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21272 1352 21324 1358
rect 21272 1294 21324 1300
rect 21376 160 21404 2314
rect 21468 1086 21496 3470
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21456 1080 21508 1086
rect 21456 1022 21508 1028
rect 21652 160 21680 3334
rect 21836 2582 21864 3402
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22155 3292 22463 3301
rect 22155 3290 22161 3292
rect 22217 3290 22241 3292
rect 22297 3290 22321 3292
rect 22377 3290 22401 3292
rect 22457 3290 22463 3292
rect 22217 3238 22219 3290
rect 22399 3238 22401 3290
rect 22155 3236 22161 3238
rect 22217 3236 22241 3238
rect 22297 3236 22321 3238
rect 22377 3236 22401 3238
rect 22457 3236 22463 3238
rect 22155 3227 22463 3236
rect 22572 3194 22600 3334
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 21824 2576 21876 2582
rect 21824 2518 21876 2524
rect 21824 2440 21876 2446
rect 22204 2394 22232 2858
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22296 2446 22324 2790
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 21824 2382 21876 2388
rect 21836 1086 21864 2382
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 22112 2366 22232 2394
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21824 1080 21876 1086
rect 21824 1022 21876 1028
rect 21928 160 21956 2314
rect 22112 2292 22140 2366
rect 22066 2264 22140 2292
rect 22066 2020 22094 2264
rect 22155 2204 22463 2213
rect 22155 2202 22161 2204
rect 22217 2202 22241 2204
rect 22297 2202 22321 2204
rect 22377 2202 22401 2204
rect 22457 2202 22463 2204
rect 22217 2150 22219 2202
rect 22399 2150 22401 2202
rect 22155 2148 22161 2150
rect 22217 2148 22241 2150
rect 22297 2148 22321 2150
rect 22377 2148 22401 2150
rect 22457 2148 22463 2150
rect 22155 2139 22463 2148
rect 22066 1992 22232 2020
rect 22204 160 22232 1992
rect 22572 1170 22600 2450
rect 22664 2378 22692 3606
rect 22756 3058 22784 4558
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 22480 1142 22600 1170
rect 22480 160 22508 1142
rect 22756 160 22784 2790
rect 22848 1562 22876 3470
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 22940 2106 22968 3402
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22928 2100 22980 2106
rect 22928 2042 22980 2048
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 23032 160 23060 2246
rect 23124 1970 23152 3402
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23112 1964 23164 1970
rect 23112 1906 23164 1912
rect 23308 160 23336 2246
rect 23400 2038 23428 6734
rect 24596 5914 24624 7346
rect 27457 7100 27765 7109
rect 27457 7098 27463 7100
rect 27519 7098 27543 7100
rect 27599 7098 27623 7100
rect 27679 7098 27703 7100
rect 27759 7098 27765 7100
rect 27519 7046 27521 7098
rect 27701 7046 27703 7098
rect 27457 7044 27463 7046
rect 27519 7044 27543 7046
rect 27599 7044 27623 7046
rect 27679 7044 27703 7046
rect 27759 7044 27765 7046
rect 27457 7035 27765 7044
rect 27457 6012 27765 6021
rect 27457 6010 27463 6012
rect 27519 6010 27543 6012
rect 27599 6010 27623 6012
rect 27679 6010 27703 6012
rect 27759 6010 27765 6012
rect 27519 5958 27521 6010
rect 27701 5958 27703 6010
rect 27457 5956 27463 5958
rect 27519 5956 27543 5958
rect 27599 5956 27623 5958
rect 27679 5956 27703 5958
rect 27759 5956 27765 5958
rect 27457 5947 27765 5956
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 27457 4924 27765 4933
rect 27457 4922 27463 4924
rect 27519 4922 27543 4924
rect 27599 4922 27623 4924
rect 27679 4922 27703 4924
rect 27759 4922 27765 4924
rect 27519 4870 27521 4922
rect 27701 4870 27703 4922
rect 27457 4868 27463 4870
rect 27519 4868 27543 4870
rect 27599 4868 27623 4870
rect 27679 4868 27703 4870
rect 27759 4868 27765 4870
rect 27457 4859 27765 4868
rect 24216 4752 24268 4758
rect 24216 4694 24268 4700
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2446 23520 3334
rect 23860 3058 23888 4626
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24136 3602 24164 4014
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24228 3534 24256 4694
rect 27250 4584 27306 4593
rect 27250 4519 27306 4528
rect 25596 4004 25648 4010
rect 25596 3946 25648 3952
rect 25608 3534 25636 3946
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 24216 3528 24268 3534
rect 25320 3528 25372 3534
rect 24216 3470 24268 3476
rect 25240 3488 25320 3516
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 25044 3392 25096 3398
rect 25096 3352 25176 3380
rect 25044 3334 25096 3340
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23584 2292 23612 2994
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23756 2304 23808 2310
rect 23492 2264 23612 2292
rect 23676 2264 23756 2292
rect 23388 2032 23440 2038
rect 23388 1974 23440 1980
rect 23492 921 23520 2264
rect 23676 1170 23704 2264
rect 23756 2246 23808 2252
rect 23584 1142 23704 1170
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 23584 160 23612 1142
rect 23860 160 23888 2790
rect 24320 2446 24348 3334
rect 24412 3194 24440 3334
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 23952 2145 23980 2382
rect 23938 2136 23994 2145
rect 23938 2071 23994 2080
rect 24044 1290 24072 2382
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24032 1284 24084 1290
rect 24032 1226 24084 1232
rect 24136 160 24164 1906
rect 24412 160 24440 2790
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 24688 160 24716 2246
rect 24872 2106 24900 2858
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 24860 2100 24912 2106
rect 24860 2042 24912 2048
rect 24964 160 24992 2790
rect 25148 2446 25176 3352
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25240 1873 25268 3488
rect 25320 3470 25372 3476
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25688 3528 25740 3534
rect 26148 3528 26200 3534
rect 25688 3470 25740 3476
rect 25884 3488 26148 3516
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25332 3194 25360 3334
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25412 2916 25464 2922
rect 25412 2858 25464 2864
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25332 1970 25360 2450
rect 25320 1964 25372 1970
rect 25320 1906 25372 1912
rect 25226 1864 25282 1873
rect 25226 1799 25282 1808
rect 20810 82 20866 160
rect 20732 54 20866 82
rect 20810 -300 20866 54
rect 21086 -300 21142 160
rect 21362 -300 21418 160
rect 21638 -300 21694 160
rect 21914 -300 21970 160
rect 22190 -300 22246 160
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 23018 -300 23074 160
rect 23294 -300 23350 160
rect 23570 -300 23626 160
rect 23846 -300 23902 160
rect 24122 -300 24178 160
rect 24398 -300 24454 160
rect 24674 -300 24730 160
rect 24950 -300 25006 160
rect 25226 82 25282 160
rect 25424 82 25452 2858
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25516 160 25544 2790
rect 25700 1154 25728 3470
rect 25884 1601 25912 3488
rect 26148 3470 26200 3476
rect 26054 2952 26110 2961
rect 26054 2887 26110 2896
rect 26148 2916 26200 2922
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 25870 1592 25926 1601
rect 25870 1527 25926 1536
rect 25688 1148 25740 1154
rect 25688 1090 25740 1096
rect 25226 54 25452 82
rect 25226 -300 25282 54
rect 25502 -300 25558 160
rect 25778 82 25834 160
rect 25976 82 26004 2790
rect 26068 1873 26096 2887
rect 26148 2858 26200 2864
rect 26160 2650 26188 2858
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 26252 2446 26280 3674
rect 26436 3534 26464 3878
rect 27264 3534 27292 4519
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 27894 4040 27950 4049
rect 27894 3975 27950 3984
rect 27457 3836 27765 3845
rect 27457 3834 27463 3836
rect 27519 3834 27543 3836
rect 27599 3834 27623 3836
rect 27679 3834 27703 3836
rect 27759 3834 27765 3836
rect 27519 3782 27521 3834
rect 27701 3782 27703 3834
rect 27457 3780 27463 3782
rect 27519 3780 27543 3782
rect 27599 3780 27623 3782
rect 27679 3780 27703 3782
rect 27759 3780 27765 3782
rect 27457 3771 27765 3780
rect 27804 3664 27856 3670
rect 27804 3606 27856 3612
rect 27620 3596 27672 3602
rect 27620 3538 27672 3544
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 26344 3194 26372 3402
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26436 3194 26464 3334
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26332 2304 26384 2310
rect 26332 2246 26384 2252
rect 26054 1864 26110 1873
rect 26054 1799 26110 1808
rect 26344 1442 26372 2246
rect 26436 1698 26464 2382
rect 26424 1692 26476 1698
rect 26424 1634 26476 1640
rect 26160 1414 26372 1442
rect 25778 54 26004 82
rect 26054 82 26110 160
rect 26160 82 26188 1414
rect 26054 54 26188 82
rect 26330 82 26386 160
rect 26528 82 26556 2790
rect 26620 2650 26648 2926
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26712 1494 26740 3470
rect 26988 3097 27016 3470
rect 26974 3088 27030 3097
rect 26974 3023 27030 3032
rect 27632 2990 27660 3538
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27816 2938 27844 3606
rect 27908 3534 27936 3975
rect 28356 3732 28408 3738
rect 28356 3674 28408 3680
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 28080 3460 28132 3466
rect 28080 3402 28132 3408
rect 28092 3194 28120 3402
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 26884 2916 26936 2922
rect 27816 2910 27936 2938
rect 26884 2858 26936 2864
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 26700 1488 26752 1494
rect 26700 1430 26752 1436
rect 26330 54 26556 82
rect 26606 82 26662 160
rect 26804 82 26832 2586
rect 26896 160 26924 2858
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27457 2748 27765 2757
rect 27457 2746 27463 2748
rect 27519 2746 27543 2748
rect 27599 2746 27623 2748
rect 27679 2746 27703 2748
rect 27759 2746 27765 2748
rect 27519 2694 27521 2746
rect 27701 2694 27703 2746
rect 27457 2692 27463 2694
rect 27519 2692 27543 2694
rect 27599 2692 27623 2694
rect 27679 2692 27703 2694
rect 27759 2692 27765 2694
rect 27457 2683 27765 2692
rect 27816 2632 27844 2790
rect 27632 2604 27844 2632
rect 27528 2304 27580 2310
rect 27356 2264 27528 2292
rect 26606 54 26832 82
rect 25778 -300 25834 54
rect 26054 -300 26110 54
rect 26330 -300 26386 54
rect 26606 -300 26662 54
rect 26882 -300 26938 160
rect 27158 82 27214 160
rect 27356 82 27384 2264
rect 27528 2246 27580 2252
rect 27632 2122 27660 2604
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 27540 2094 27660 2122
rect 27158 54 27384 82
rect 27434 82 27490 160
rect 27540 82 27568 2094
rect 27724 160 27752 2450
rect 27908 2378 27936 2910
rect 27988 2916 28040 2922
rect 28184 2904 28212 3470
rect 27988 2858 28040 2864
rect 28092 2876 28212 2904
rect 27804 2372 27856 2378
rect 27804 2314 27856 2320
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 27816 2258 27844 2314
rect 28000 2258 28028 2858
rect 28092 2281 28120 2876
rect 28170 2816 28226 2825
rect 28170 2751 28226 2760
rect 27816 2230 28028 2258
rect 28078 2272 28134 2281
rect 28078 2207 28134 2216
rect 27434 54 27568 82
rect 27158 -300 27214 54
rect 27434 -300 27490 54
rect 27710 -300 27766 160
rect 27986 82 28042 160
rect 28184 82 28212 2751
rect 28368 2378 28396 3674
rect 28446 3632 28502 3641
rect 28446 3567 28502 3576
rect 28460 3534 28488 3567
rect 28736 3534 28764 4422
rect 29196 3738 29224 7346
rect 30012 4004 30064 4010
rect 30012 3946 30064 3952
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29276 3596 29328 3602
rect 29276 3538 29328 3544
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 29000 3460 29052 3466
rect 29000 3402 29052 3408
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28552 3194 28580 3334
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28540 2916 28592 2922
rect 28540 2858 28592 2864
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28448 2304 28500 2310
rect 28448 2246 28500 2252
rect 27986 54 28212 82
rect 28262 82 28318 160
rect 28460 82 28488 2246
rect 28552 160 28580 2858
rect 28736 2650 28764 2994
rect 28816 2848 28868 2854
rect 28814 2816 28816 2825
rect 28868 2816 28870 2825
rect 28814 2751 28870 2760
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28920 1170 28948 2518
rect 29012 2378 29040 3402
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 28828 1142 28948 1170
rect 28828 160 28856 1142
rect 29104 160 29132 3130
rect 29288 3058 29316 3538
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 29380 2961 29408 2994
rect 29366 2952 29422 2961
rect 29366 2887 29422 2896
rect 29644 2644 29696 2650
rect 29380 2604 29644 2632
rect 29380 160 29408 2604
rect 29644 2586 29696 2592
rect 29748 2446 29776 3606
rect 30024 3194 30052 3946
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30196 2916 30248 2922
rect 30196 2858 30248 2864
rect 29828 2848 29880 2854
rect 29828 2790 29880 2796
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 29472 1766 29500 2382
rect 29460 1760 29512 1766
rect 29460 1702 29512 1708
rect 28262 54 28488 82
rect 27986 -300 28042 54
rect 28262 -300 28318 54
rect 28538 -300 28594 160
rect 28814 -300 28870 160
rect 29090 -300 29146 160
rect 29366 -300 29422 160
rect 29642 82 29698 160
rect 29840 82 29868 2790
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 2106 29960 2314
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 29920 2100 29972 2106
rect 29920 2042 29972 2048
rect 29642 54 29868 82
rect 29918 82 29974 160
rect 30116 82 30144 2246
rect 30208 160 30236 2858
rect 30484 2417 30512 2994
rect 30470 2408 30526 2417
rect 30470 2343 30526 2352
rect 29918 54 30144 82
rect 29642 -300 29698 54
rect 29918 -300 29974 54
rect 30194 -300 30250 160
rect 30470 82 30526 160
rect 30668 82 30696 3130
rect 31300 2916 31352 2922
rect 31300 2858 31352 2864
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 30840 2440 30892 2446
rect 31036 2394 31064 2518
rect 30840 2382 30892 2388
rect 30852 1465 30880 2382
rect 30944 2366 31064 2394
rect 30838 1456 30894 1465
rect 30838 1391 30894 1400
rect 30470 54 30696 82
rect 30746 82 30802 160
rect 30944 82 30972 2366
rect 31208 1420 31260 1426
rect 31208 1362 31260 1368
rect 30746 54 30972 82
rect 31022 82 31078 160
rect 31220 82 31248 1362
rect 31312 160 31340 2858
rect 31772 2650 31800 7346
rect 33876 7336 33928 7342
rect 33876 7278 33928 7284
rect 32758 6556 33066 6565
rect 32758 6554 32764 6556
rect 32820 6554 32844 6556
rect 32900 6554 32924 6556
rect 32980 6554 33004 6556
rect 33060 6554 33066 6556
rect 32820 6502 32822 6554
rect 33002 6502 33004 6554
rect 32758 6500 32764 6502
rect 32820 6500 32844 6502
rect 32900 6500 32924 6502
rect 32980 6500 33004 6502
rect 33060 6500 33066 6502
rect 32758 6491 33066 6500
rect 33508 6180 33560 6186
rect 33508 6122 33560 6128
rect 32758 5468 33066 5477
rect 32758 5466 32764 5468
rect 32820 5466 32844 5468
rect 32900 5466 32924 5468
rect 32980 5466 33004 5468
rect 33060 5466 33066 5468
rect 32820 5414 32822 5466
rect 33002 5414 33004 5466
rect 32758 5412 32764 5414
rect 32820 5412 32844 5414
rect 32900 5412 32924 5414
rect 32980 5412 33004 5414
rect 33060 5412 33066 5414
rect 32758 5403 33066 5412
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 32758 4380 33066 4389
rect 32758 4378 32764 4380
rect 32820 4378 32844 4380
rect 32900 4378 32924 4380
rect 32980 4378 33004 4380
rect 33060 4378 33066 4380
rect 32820 4326 32822 4378
rect 33002 4326 33004 4378
rect 32758 4324 32764 4326
rect 32820 4324 32844 4326
rect 32900 4324 32924 4326
rect 32980 4324 33004 4326
rect 33060 4324 33066 4326
rect 32758 4315 33066 4324
rect 32036 3460 32088 3466
rect 32036 3402 32088 3408
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31576 2100 31628 2106
rect 31576 2042 31628 2048
rect 31588 160 31616 2042
rect 31864 160 31892 3130
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 31956 1057 31984 2994
rect 32048 1329 32076 3402
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32232 2145 32260 2314
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 32218 2136 32274 2145
rect 32218 2071 32274 2080
rect 32220 1488 32272 1494
rect 32220 1430 32272 1436
rect 32034 1320 32090 1329
rect 32034 1255 32090 1264
rect 31942 1048 31998 1057
rect 31942 983 31998 992
rect 31022 54 31248 82
rect 30470 -300 30526 54
rect 30746 -300 30802 54
rect 31022 -300 31078 54
rect 31298 -300 31354 160
rect 31574 -300 31630 160
rect 31850 -300 31906 160
rect 32126 82 32182 160
rect 32232 82 32260 1430
rect 32324 1426 32352 2246
rect 32312 1420 32364 1426
rect 32312 1362 32364 1368
rect 32416 160 32444 2858
rect 32692 160 32720 3334
rect 32758 3292 33066 3301
rect 32758 3290 32764 3292
rect 32820 3290 32844 3292
rect 32900 3290 32924 3292
rect 32980 3290 33004 3292
rect 33060 3290 33066 3292
rect 32820 3238 32822 3290
rect 33002 3238 33004 3290
rect 32758 3236 32764 3238
rect 32820 3236 32844 3238
rect 32900 3236 32924 3238
rect 32980 3236 33004 3238
rect 33060 3236 33066 3238
rect 32758 3227 33066 3236
rect 33152 3126 33180 4490
rect 33520 3738 33548 6122
rect 33508 3732 33560 3738
rect 33508 3674 33560 3680
rect 33416 3460 33468 3466
rect 33416 3402 33468 3408
rect 33140 3120 33192 3126
rect 33140 3062 33192 3068
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32784 2825 32812 2994
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 32770 2816 32826 2825
rect 32770 2751 32826 2760
rect 33060 2394 33088 2926
rect 33428 2650 33456 3402
rect 33692 3052 33744 3058
rect 33692 2994 33744 3000
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33324 2576 33376 2582
rect 33138 2544 33194 2553
rect 33324 2518 33376 2524
rect 33138 2479 33140 2488
rect 33192 2479 33194 2488
rect 33140 2450 33192 2456
rect 33060 2366 33180 2394
rect 32758 2204 33066 2213
rect 32758 2202 32764 2204
rect 32820 2202 32844 2204
rect 32900 2202 32924 2204
rect 32980 2202 33004 2204
rect 33060 2202 33066 2204
rect 32820 2150 32822 2202
rect 33002 2150 33004 2202
rect 32758 2148 32764 2150
rect 32820 2148 32844 2150
rect 32900 2148 32924 2150
rect 32980 2148 33004 2150
rect 33060 2148 33066 2150
rect 32758 2139 33066 2148
rect 33152 2088 33180 2366
rect 33232 2372 33284 2378
rect 33232 2314 33284 2320
rect 33060 2060 33180 2088
rect 32126 54 32260 82
rect 32126 -300 32182 54
rect 32402 -300 32458 160
rect 32678 -300 32734 160
rect 32954 82 33010 160
rect 33060 82 33088 2060
rect 33244 1222 33272 2314
rect 33232 1216 33284 1222
rect 33232 1158 33284 1164
rect 32954 54 33088 82
rect 33230 82 33286 160
rect 33336 82 33364 2518
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 33428 2106 33456 2246
rect 33416 2100 33468 2106
rect 33416 2042 33468 2048
rect 33520 160 33548 2858
rect 33704 950 33732 2994
rect 33888 1834 33916 7278
rect 35716 7268 35768 7274
rect 35716 7210 35768 7216
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34440 5522 34468 6938
rect 34440 5494 34560 5522
rect 33968 4276 34020 4282
rect 33968 4218 34020 4224
rect 33980 3126 34008 4218
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 34532 3058 34560 5494
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 34612 2916 34664 2922
rect 34612 2858 34664 2864
rect 34428 2508 34480 2514
rect 34428 2450 34480 2456
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 33968 2304 34020 2310
rect 33968 2246 34020 2252
rect 33876 1828 33928 1834
rect 33876 1770 33928 1776
rect 33980 1494 34008 2246
rect 33968 1488 34020 1494
rect 33968 1430 34020 1436
rect 33692 944 33744 950
rect 33692 886 33744 892
rect 34072 218 34100 2382
rect 33980 190 34100 218
rect 33230 54 33364 82
rect 32954 -300 33010 54
rect 33230 -300 33286 54
rect 33506 -300 33562 160
rect 33782 82 33838 160
rect 33980 82 34008 190
rect 33782 54 34008 82
rect 33782 -300 33838 54
rect 34058 -300 34114 160
rect 34334 82 34390 160
rect 34440 82 34468 2450
rect 34624 160 34652 2858
rect 34716 2378 34744 3334
rect 34808 2854 34836 7142
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35728 3074 35756 7210
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35820 3194 35848 3334
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 34888 2984 34940 2990
rect 34888 2926 34940 2932
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 34808 1873 34836 2314
rect 34794 1864 34850 1873
rect 34794 1799 34850 1808
rect 34900 160 34928 2926
rect 35452 2774 35480 3062
rect 35532 3052 35584 3058
rect 35728 3046 35848 3074
rect 35532 2994 35584 3000
rect 35360 2746 35480 2774
rect 34334 54 34468 82
rect 34334 -300 34390 54
rect 34610 -300 34666 160
rect 34886 -300 34942 160
rect 35162 82 35218 160
rect 35360 82 35388 2746
rect 35544 2650 35572 2994
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35452 1970 35480 2246
rect 35440 1964 35492 1970
rect 35440 1906 35492 1912
rect 35624 1420 35676 1426
rect 35624 1362 35676 1368
rect 35162 54 35388 82
rect 35438 82 35494 160
rect 35636 82 35664 1362
rect 35728 160 35756 2926
rect 35820 2650 35848 3046
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 35912 2446 35940 2790
rect 36004 2650 36032 6258
rect 36636 6248 36688 6254
rect 36636 6190 36688 6196
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 36280 3126 36308 3470
rect 36268 3120 36320 3126
rect 36268 3062 36320 3068
rect 36372 2922 36400 4150
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36360 2916 36412 2922
rect 36360 2858 36412 2864
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 36084 2508 36136 2514
rect 36084 2450 36136 2456
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 36096 1306 36124 2450
rect 36188 2446 36216 2858
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 36372 1970 36400 2246
rect 36360 1964 36412 1970
rect 36360 1906 36412 1912
rect 36004 1278 36124 1306
rect 36004 160 36032 1278
rect 35438 54 35664 82
rect 35162 -300 35218 54
rect 35438 -300 35494 54
rect 35714 -300 35770 160
rect 35990 -300 36046 160
rect 36266 82 36322 160
rect 36464 82 36492 2994
rect 36648 2922 36676 6190
rect 36636 2916 36688 2922
rect 36636 2858 36688 2864
rect 37384 2774 37412 7346
rect 38060 7100 38368 7109
rect 38060 7098 38066 7100
rect 38122 7098 38146 7100
rect 38202 7098 38226 7100
rect 38282 7098 38306 7100
rect 38362 7098 38368 7100
rect 38122 7046 38124 7098
rect 38304 7046 38306 7098
rect 38060 7044 38066 7046
rect 38122 7044 38146 7046
rect 38202 7044 38226 7046
rect 38282 7044 38306 7046
rect 38362 7044 38368 7046
rect 38060 7035 38368 7044
rect 38060 6012 38368 6021
rect 38060 6010 38066 6012
rect 38122 6010 38146 6012
rect 38202 6010 38226 6012
rect 38282 6010 38306 6012
rect 38362 6010 38368 6012
rect 38122 5958 38124 6010
rect 38304 5958 38306 6010
rect 38060 5956 38066 5958
rect 38122 5956 38146 5958
rect 38202 5956 38226 5958
rect 38282 5956 38306 5958
rect 38362 5956 38368 5958
rect 38060 5947 38368 5956
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 37384 2746 37504 2774
rect 37002 2680 37058 2689
rect 37002 2615 37004 2624
rect 37056 2615 37058 2624
rect 37004 2586 37056 2592
rect 37372 2576 37424 2582
rect 37372 2518 37424 2524
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 36636 2372 36688 2378
rect 36636 2314 36688 2320
rect 36266 54 36492 82
rect 36542 82 36598 160
rect 36648 82 36676 2314
rect 36740 1426 36768 2382
rect 36728 1420 36780 1426
rect 36728 1362 36780 1368
rect 36924 1306 36952 2450
rect 36832 1278 36952 1306
rect 37108 2378 37228 2394
rect 37108 2372 37240 2378
rect 37108 2366 37188 2372
rect 36832 160 36860 1278
rect 37108 160 37136 2366
rect 37188 2314 37240 2320
rect 37384 160 37412 2518
rect 37476 2106 37504 2746
rect 37464 2100 37516 2106
rect 37464 2042 37516 2048
rect 37660 160 37688 2994
rect 37844 2650 37872 5646
rect 38060 4924 38368 4933
rect 38060 4922 38066 4924
rect 38122 4922 38146 4924
rect 38202 4922 38226 4924
rect 38282 4922 38306 4924
rect 38362 4922 38368 4924
rect 38122 4870 38124 4922
rect 38304 4870 38306 4922
rect 38060 4868 38066 4870
rect 38122 4868 38146 4870
rect 38202 4868 38226 4870
rect 38282 4868 38306 4870
rect 38362 4868 38368 4870
rect 38060 4859 38368 4868
rect 38060 3836 38368 3845
rect 38060 3834 38066 3836
rect 38122 3834 38146 3836
rect 38202 3834 38226 3836
rect 38282 3834 38306 3836
rect 38362 3834 38368 3836
rect 38122 3782 38124 3834
rect 38304 3782 38306 3834
rect 38060 3780 38066 3782
rect 38122 3780 38146 3782
rect 38202 3780 38226 3782
rect 38282 3780 38306 3782
rect 38362 3780 38368 3782
rect 38060 3771 38368 3780
rect 37936 3058 38056 3074
rect 37936 3052 38068 3058
rect 37936 3046 38016 3052
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 37740 2304 37792 2310
rect 37740 2246 37792 2252
rect 37752 2038 37780 2246
rect 37740 2032 37792 2038
rect 37740 1974 37792 1980
rect 37936 160 37964 3046
rect 38016 2994 38068 3000
rect 38060 2748 38368 2757
rect 38060 2746 38066 2748
rect 38122 2746 38146 2748
rect 38202 2746 38226 2748
rect 38282 2746 38306 2748
rect 38362 2746 38368 2748
rect 38122 2694 38124 2746
rect 38304 2694 38306 2746
rect 38060 2692 38066 2694
rect 38122 2692 38146 2694
rect 38202 2692 38226 2694
rect 38282 2692 38306 2694
rect 38362 2692 38368 2694
rect 38060 2683 38368 2692
rect 38396 2650 38424 7346
rect 38660 7336 38712 7342
rect 38660 7278 38712 7284
rect 38672 2650 38700 7278
rect 39028 3052 39080 3058
rect 39028 2994 39080 3000
rect 38384 2644 38436 2650
rect 38384 2586 38436 2592
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 38936 2440 38988 2446
rect 38936 2382 38988 2388
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38384 2304 38436 2310
rect 38384 2246 38436 2252
rect 38304 1834 38332 2246
rect 38396 2106 38424 2246
rect 38384 2100 38436 2106
rect 38384 2042 38436 2048
rect 38292 1828 38344 1834
rect 38292 1770 38344 1776
rect 38948 1714 38976 2382
rect 38396 1686 38976 1714
rect 36542 54 36676 82
rect 36266 -300 36322 54
rect 36542 -300 36598 54
rect 36818 -300 36874 160
rect 37094 -300 37150 160
rect 37370 -300 37426 160
rect 37646 -300 37702 160
rect 37922 -300 37978 160
rect 38198 82 38254 160
rect 38396 82 38424 1686
rect 38752 1556 38804 1562
rect 38752 1498 38804 1504
rect 38568 1352 38620 1358
rect 38568 1294 38620 1300
rect 38198 54 38424 82
rect 38474 82 38530 160
rect 38580 82 38608 1294
rect 38764 160 38792 1498
rect 39040 160 39068 2994
rect 39960 2650 39988 7346
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 40052 2446 40080 2790
rect 41524 2650 41552 7346
rect 42444 2650 42472 7346
rect 43361 6556 43669 6565
rect 43361 6554 43367 6556
rect 43423 6554 43447 6556
rect 43503 6554 43527 6556
rect 43583 6554 43607 6556
rect 43663 6554 43669 6556
rect 43423 6502 43425 6554
rect 43605 6502 43607 6554
rect 43361 6500 43367 6502
rect 43423 6500 43447 6502
rect 43503 6500 43527 6502
rect 43583 6500 43607 6502
rect 43663 6500 43669 6502
rect 43361 6491 43669 6500
rect 43361 5468 43669 5477
rect 43361 5466 43367 5468
rect 43423 5466 43447 5468
rect 43503 5466 43527 5468
rect 43583 5466 43607 5468
rect 43663 5466 43669 5468
rect 43423 5414 43425 5466
rect 43605 5414 43607 5466
rect 43361 5412 43367 5414
rect 43423 5412 43447 5414
rect 43503 5412 43527 5414
rect 43583 5412 43607 5414
rect 43663 5412 43669 5414
rect 43361 5403 43669 5412
rect 43361 4380 43669 4389
rect 43361 4378 43367 4380
rect 43423 4378 43447 4380
rect 43503 4378 43527 4380
rect 43583 4378 43607 4380
rect 43663 4378 43669 4380
rect 43423 4326 43425 4378
rect 43605 4326 43607 4378
rect 43361 4324 43367 4326
rect 43423 4324 43447 4326
rect 43503 4324 43527 4326
rect 43583 4324 43607 4326
rect 43663 4324 43669 4326
rect 43361 4315 43669 4324
rect 43361 3292 43669 3301
rect 43361 3290 43367 3292
rect 43423 3290 43447 3292
rect 43503 3290 43527 3292
rect 43583 3290 43607 3292
rect 43663 3290 43669 3292
rect 43423 3238 43425 3290
rect 43605 3238 43607 3290
rect 43361 3236 43367 3238
rect 43423 3236 43447 3238
rect 43503 3236 43527 3238
rect 43583 3236 43607 3238
rect 43663 3236 43669 3238
rect 43361 3227 43669 3236
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 42432 2644 42484 2650
rect 42432 2586 42484 2592
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39672 2440 39724 2446
rect 40040 2440 40092 2446
rect 39672 2382 39724 2388
rect 39408 1494 39436 2382
rect 39684 1562 39712 2382
rect 39868 2378 39988 2394
rect 40040 2382 40092 2388
rect 40316 2440 40368 2446
rect 40316 2382 40368 2388
rect 39868 2372 40000 2378
rect 39868 2366 39948 2372
rect 39672 1556 39724 1562
rect 39672 1498 39724 1504
rect 39396 1488 39448 1494
rect 39396 1430 39448 1436
rect 39304 1420 39356 1426
rect 39304 1362 39356 1368
rect 39316 160 39344 1362
rect 38474 54 38608 82
rect 38198 -300 38254 54
rect 38474 -300 38530 54
rect 38750 -300 38806 160
rect 39026 -300 39082 160
rect 39302 -300 39358 160
rect 39578 82 39634 160
rect 39868 82 39896 2366
rect 39948 2314 40000 2320
rect 40328 1426 40356 2382
rect 43361 2204 43669 2213
rect 43361 2202 43367 2204
rect 43423 2202 43447 2204
rect 43503 2202 43527 2204
rect 43583 2202 43607 2204
rect 43663 2202 43669 2204
rect 43423 2150 43425 2202
rect 43605 2150 43607 2202
rect 43361 2148 43367 2150
rect 43423 2148 43447 2150
rect 43503 2148 43527 2150
rect 43583 2148 43607 2150
rect 43663 2148 43669 2150
rect 43361 2139 43669 2148
rect 40316 1420 40368 1426
rect 40316 1362 40368 1368
rect 39578 54 39896 82
rect 39578 -300 39634 54
<< via2 >>
rect 11558 7642 11614 7644
rect 11638 7642 11694 7644
rect 11718 7642 11774 7644
rect 11798 7642 11854 7644
rect 11558 7590 11604 7642
rect 11604 7590 11614 7642
rect 11638 7590 11668 7642
rect 11668 7590 11680 7642
rect 11680 7590 11694 7642
rect 11718 7590 11732 7642
rect 11732 7590 11744 7642
rect 11744 7590 11774 7642
rect 11798 7590 11808 7642
rect 11808 7590 11854 7642
rect 11558 7588 11614 7590
rect 11638 7588 11694 7590
rect 11718 7588 11774 7590
rect 11798 7588 11854 7590
rect 22161 7642 22217 7644
rect 22241 7642 22297 7644
rect 22321 7642 22377 7644
rect 22401 7642 22457 7644
rect 22161 7590 22207 7642
rect 22207 7590 22217 7642
rect 22241 7590 22271 7642
rect 22271 7590 22283 7642
rect 22283 7590 22297 7642
rect 22321 7590 22335 7642
rect 22335 7590 22347 7642
rect 22347 7590 22377 7642
rect 22401 7590 22411 7642
rect 22411 7590 22457 7642
rect 22161 7588 22217 7590
rect 22241 7588 22297 7590
rect 22321 7588 22377 7590
rect 22401 7588 22457 7590
rect 32764 7642 32820 7644
rect 32844 7642 32900 7644
rect 32924 7642 32980 7644
rect 33004 7642 33060 7644
rect 32764 7590 32810 7642
rect 32810 7590 32820 7642
rect 32844 7590 32874 7642
rect 32874 7590 32886 7642
rect 32886 7590 32900 7642
rect 32924 7590 32938 7642
rect 32938 7590 32950 7642
rect 32950 7590 32980 7642
rect 33004 7590 33014 7642
rect 33014 7590 33060 7642
rect 32764 7588 32820 7590
rect 32844 7588 32900 7590
rect 32924 7588 32980 7590
rect 33004 7588 33060 7590
rect 43367 7642 43423 7644
rect 43447 7642 43503 7644
rect 43527 7642 43583 7644
rect 43607 7642 43663 7644
rect 43367 7590 43413 7642
rect 43413 7590 43423 7642
rect 43447 7590 43477 7642
rect 43477 7590 43489 7642
rect 43489 7590 43503 7642
rect 43527 7590 43541 7642
rect 43541 7590 43553 7642
rect 43553 7590 43583 7642
rect 43607 7590 43617 7642
rect 43617 7590 43663 7642
rect 43367 7588 43423 7590
rect 43447 7588 43503 7590
rect 43527 7588 43583 7590
rect 43607 7588 43663 7590
rect 6257 7098 6313 7100
rect 6337 7098 6393 7100
rect 6417 7098 6473 7100
rect 6497 7098 6553 7100
rect 6257 7046 6303 7098
rect 6303 7046 6313 7098
rect 6337 7046 6367 7098
rect 6367 7046 6379 7098
rect 6379 7046 6393 7098
rect 6417 7046 6431 7098
rect 6431 7046 6443 7098
rect 6443 7046 6473 7098
rect 6497 7046 6507 7098
rect 6507 7046 6553 7098
rect 6257 7044 6313 7046
rect 6337 7044 6393 7046
rect 6417 7044 6473 7046
rect 6497 7044 6553 7046
rect 6257 6010 6313 6012
rect 6337 6010 6393 6012
rect 6417 6010 6473 6012
rect 6497 6010 6553 6012
rect 6257 5958 6303 6010
rect 6303 5958 6313 6010
rect 6337 5958 6367 6010
rect 6367 5958 6379 6010
rect 6379 5958 6393 6010
rect 6417 5958 6431 6010
rect 6431 5958 6443 6010
rect 6443 5958 6473 6010
rect 6497 5958 6507 6010
rect 6507 5958 6553 6010
rect 6257 5956 6313 5958
rect 6337 5956 6393 5958
rect 6417 5956 6473 5958
rect 6497 5956 6553 5958
rect 6257 4922 6313 4924
rect 6337 4922 6393 4924
rect 6417 4922 6473 4924
rect 6497 4922 6553 4924
rect 6257 4870 6303 4922
rect 6303 4870 6313 4922
rect 6337 4870 6367 4922
rect 6367 4870 6379 4922
rect 6379 4870 6393 4922
rect 6417 4870 6431 4922
rect 6431 4870 6443 4922
rect 6443 4870 6473 4922
rect 6497 4870 6507 4922
rect 6507 4870 6553 4922
rect 6257 4868 6313 4870
rect 6337 4868 6393 4870
rect 6417 4868 6473 4870
rect 6497 4868 6553 4870
rect 6257 3834 6313 3836
rect 6337 3834 6393 3836
rect 6417 3834 6473 3836
rect 6497 3834 6553 3836
rect 6257 3782 6303 3834
rect 6303 3782 6313 3834
rect 6337 3782 6367 3834
rect 6367 3782 6379 3834
rect 6379 3782 6393 3834
rect 6417 3782 6431 3834
rect 6431 3782 6443 3834
rect 6443 3782 6473 3834
rect 6497 3782 6507 3834
rect 6507 3782 6553 3834
rect 6257 3780 6313 3782
rect 6337 3780 6393 3782
rect 6417 3780 6473 3782
rect 6497 3780 6553 3782
rect 5078 2896 5134 2952
rect 6257 2746 6313 2748
rect 6337 2746 6393 2748
rect 6417 2746 6473 2748
rect 6497 2746 6553 2748
rect 6257 2694 6303 2746
rect 6303 2694 6313 2746
rect 6337 2694 6367 2746
rect 6367 2694 6379 2746
rect 6379 2694 6393 2746
rect 6417 2694 6431 2746
rect 6431 2694 6443 2746
rect 6443 2694 6473 2746
rect 6497 2694 6507 2746
rect 6507 2694 6553 2746
rect 6257 2692 6313 2694
rect 6337 2692 6393 2694
rect 6417 2692 6473 2694
rect 6497 2692 6553 2694
rect 11558 6554 11614 6556
rect 11638 6554 11694 6556
rect 11718 6554 11774 6556
rect 11798 6554 11854 6556
rect 11558 6502 11604 6554
rect 11604 6502 11614 6554
rect 11638 6502 11668 6554
rect 11668 6502 11680 6554
rect 11680 6502 11694 6554
rect 11718 6502 11732 6554
rect 11732 6502 11744 6554
rect 11744 6502 11774 6554
rect 11798 6502 11808 6554
rect 11808 6502 11854 6554
rect 11558 6500 11614 6502
rect 11638 6500 11694 6502
rect 11718 6500 11774 6502
rect 11798 6500 11854 6502
rect 11558 5466 11614 5468
rect 11638 5466 11694 5468
rect 11718 5466 11774 5468
rect 11798 5466 11854 5468
rect 11558 5414 11604 5466
rect 11604 5414 11614 5466
rect 11638 5414 11668 5466
rect 11668 5414 11680 5466
rect 11680 5414 11694 5466
rect 11718 5414 11732 5466
rect 11732 5414 11744 5466
rect 11744 5414 11774 5466
rect 11798 5414 11808 5466
rect 11808 5414 11854 5466
rect 11558 5412 11614 5414
rect 11638 5412 11694 5414
rect 11718 5412 11774 5414
rect 11798 5412 11854 5414
rect 9310 3440 9366 3496
rect 6918 856 6974 912
rect 8758 1672 8814 1728
rect 13450 4528 13506 4584
rect 10782 3032 10838 3088
rect 11558 4378 11614 4380
rect 11638 4378 11694 4380
rect 11718 4378 11774 4380
rect 11798 4378 11854 4380
rect 11558 4326 11604 4378
rect 11604 4326 11614 4378
rect 11638 4326 11668 4378
rect 11668 4326 11680 4378
rect 11680 4326 11694 4378
rect 11718 4326 11732 4378
rect 11732 4326 11744 4378
rect 11744 4326 11774 4378
rect 11798 4326 11808 4378
rect 11808 4326 11854 4378
rect 11558 4324 11614 4326
rect 11638 4324 11694 4326
rect 11718 4324 11774 4326
rect 11798 4324 11854 4326
rect 12990 4256 13046 4312
rect 12806 3984 12862 4040
rect 11334 3576 11390 3632
rect 11558 3290 11614 3292
rect 11638 3290 11694 3292
rect 11718 3290 11774 3292
rect 11798 3290 11854 3292
rect 11558 3238 11604 3290
rect 11604 3238 11614 3290
rect 11638 3238 11668 3290
rect 11668 3238 11680 3290
rect 11680 3238 11694 3290
rect 11718 3238 11732 3290
rect 11732 3238 11744 3290
rect 11744 3238 11774 3290
rect 11798 3238 11808 3290
rect 11808 3238 11854 3290
rect 11558 3236 11614 3238
rect 11638 3236 11694 3238
rect 11718 3236 11774 3238
rect 11798 3236 11854 3238
rect 12254 3168 12310 3224
rect 11334 1944 11390 2000
rect 11558 2202 11614 2204
rect 11638 2202 11694 2204
rect 11718 2202 11774 2204
rect 11798 2202 11854 2204
rect 11558 2150 11604 2202
rect 11604 2150 11614 2202
rect 11638 2150 11668 2202
rect 11668 2150 11680 2202
rect 11680 2150 11694 2202
rect 11718 2150 11732 2202
rect 11732 2150 11744 2202
rect 11744 2150 11774 2202
rect 11798 2150 11808 2202
rect 11808 2150 11854 2202
rect 11558 2148 11614 2150
rect 11638 2148 11694 2150
rect 11718 2148 11774 2150
rect 11798 2148 11854 2150
rect 12162 2080 12218 2136
rect 16860 7098 16916 7100
rect 16940 7098 16996 7100
rect 17020 7098 17076 7100
rect 17100 7098 17156 7100
rect 16860 7046 16906 7098
rect 16906 7046 16916 7098
rect 16940 7046 16970 7098
rect 16970 7046 16982 7098
rect 16982 7046 16996 7098
rect 17020 7046 17034 7098
rect 17034 7046 17046 7098
rect 17046 7046 17076 7098
rect 17100 7046 17110 7098
rect 17110 7046 17156 7098
rect 16860 7044 16916 7046
rect 16940 7044 16996 7046
rect 17020 7044 17076 7046
rect 17100 7044 17156 7046
rect 16860 6010 16916 6012
rect 16940 6010 16996 6012
rect 17020 6010 17076 6012
rect 17100 6010 17156 6012
rect 16860 5958 16906 6010
rect 16906 5958 16916 6010
rect 16940 5958 16970 6010
rect 16970 5958 16982 6010
rect 16982 5958 16996 6010
rect 17020 5958 17034 6010
rect 17034 5958 17046 6010
rect 17046 5958 17076 6010
rect 17100 5958 17110 6010
rect 17110 5958 17156 6010
rect 16860 5956 16916 5958
rect 16940 5956 16996 5958
rect 17020 5956 17076 5958
rect 17100 5956 17156 5958
rect 16486 5108 16488 5128
rect 16488 5108 16540 5128
rect 16540 5108 16542 5128
rect 16486 5072 16542 5108
rect 16860 4922 16916 4924
rect 16940 4922 16996 4924
rect 17020 4922 17076 4924
rect 17100 4922 17156 4924
rect 16860 4870 16906 4922
rect 16906 4870 16916 4922
rect 16940 4870 16970 4922
rect 16970 4870 16982 4922
rect 16982 4870 16996 4922
rect 17020 4870 17034 4922
rect 17034 4870 17046 4922
rect 17046 4870 17076 4922
rect 17100 4870 17110 4922
rect 17110 4870 17156 4922
rect 16860 4868 16916 4870
rect 16940 4868 16996 4870
rect 17020 4868 17076 4870
rect 17100 4868 17156 4870
rect 16860 3834 16916 3836
rect 16940 3834 16996 3836
rect 17020 3834 17076 3836
rect 17100 3834 17156 3836
rect 16860 3782 16906 3834
rect 16906 3782 16916 3834
rect 16940 3782 16970 3834
rect 16970 3782 16982 3834
rect 16982 3782 16996 3834
rect 17020 3782 17034 3834
rect 17034 3782 17046 3834
rect 17046 3782 17076 3834
rect 17100 3782 17110 3834
rect 17110 3782 17156 3834
rect 16860 3780 16916 3782
rect 16940 3780 16996 3782
rect 17020 3780 17076 3782
rect 17100 3780 17156 3782
rect 13634 2524 13636 2544
rect 13636 2524 13688 2544
rect 13688 2524 13690 2544
rect 13634 2488 13690 2524
rect 13082 1536 13138 1592
rect 13634 1808 13690 1864
rect 15382 3032 15438 3088
rect 15382 1264 15438 1320
rect 16860 2746 16916 2748
rect 16940 2746 16996 2748
rect 17020 2746 17076 2748
rect 17100 2746 17156 2748
rect 16860 2694 16906 2746
rect 16906 2694 16916 2746
rect 16940 2694 16970 2746
rect 16970 2694 16982 2746
rect 16982 2694 16996 2746
rect 17020 2694 17034 2746
rect 17034 2694 17046 2746
rect 17046 2694 17076 2746
rect 17100 2694 17110 2746
rect 17110 2694 17156 2746
rect 16860 2692 16916 2694
rect 16940 2692 16996 2694
rect 17020 2692 17076 2694
rect 17100 2692 17156 2694
rect 16394 1128 16450 1184
rect 17130 1400 17186 1456
rect 17866 3460 17922 3496
rect 17866 3440 17868 3460
rect 17868 3440 17920 3460
rect 17920 3440 17922 3460
rect 17406 2488 17462 2544
rect 17314 2372 17370 2408
rect 17314 2352 17316 2372
rect 17316 2352 17368 2372
rect 17368 2352 17370 2372
rect 17682 992 17738 1048
rect 18510 2760 18566 2816
rect 20626 4256 20682 4312
rect 18786 1672 18842 1728
rect 18970 2352 19026 2408
rect 19798 2896 19854 2952
rect 19430 2080 19486 2136
rect 22161 6554 22217 6556
rect 22241 6554 22297 6556
rect 22321 6554 22377 6556
rect 22401 6554 22457 6556
rect 22161 6502 22207 6554
rect 22207 6502 22217 6554
rect 22241 6502 22271 6554
rect 22271 6502 22283 6554
rect 22283 6502 22297 6554
rect 22321 6502 22335 6554
rect 22335 6502 22347 6554
rect 22347 6502 22377 6554
rect 22401 6502 22411 6554
rect 22411 6502 22457 6554
rect 22161 6500 22217 6502
rect 22241 6500 22297 6502
rect 22321 6500 22377 6502
rect 22401 6500 22457 6502
rect 22161 5466 22217 5468
rect 22241 5466 22297 5468
rect 22321 5466 22377 5468
rect 22401 5466 22457 5468
rect 22161 5414 22207 5466
rect 22207 5414 22217 5466
rect 22241 5414 22271 5466
rect 22271 5414 22283 5466
rect 22283 5414 22297 5466
rect 22321 5414 22335 5466
rect 22335 5414 22347 5466
rect 22347 5414 22377 5466
rect 22401 5414 22411 5466
rect 22411 5414 22457 5466
rect 22161 5412 22217 5414
rect 22241 5412 22297 5414
rect 22321 5412 22377 5414
rect 22401 5412 22457 5414
rect 22161 4378 22217 4380
rect 22241 4378 22297 4380
rect 22321 4378 22377 4380
rect 22401 4378 22457 4380
rect 22161 4326 22207 4378
rect 22207 4326 22217 4378
rect 22241 4326 22271 4378
rect 22271 4326 22283 4378
rect 22283 4326 22297 4378
rect 22321 4326 22335 4378
rect 22335 4326 22347 4378
rect 22347 4326 22377 4378
rect 22401 4326 22411 4378
rect 22411 4326 22457 4378
rect 22161 4324 22217 4326
rect 22241 4324 22297 4326
rect 22321 4324 22377 4326
rect 22401 4324 22457 4326
rect 22098 3984 22154 4040
rect 22161 3290 22217 3292
rect 22241 3290 22297 3292
rect 22321 3290 22377 3292
rect 22401 3290 22457 3292
rect 22161 3238 22207 3290
rect 22207 3238 22217 3290
rect 22241 3238 22271 3290
rect 22271 3238 22283 3290
rect 22283 3238 22297 3290
rect 22321 3238 22335 3290
rect 22335 3238 22347 3290
rect 22347 3238 22377 3290
rect 22401 3238 22411 3290
rect 22411 3238 22457 3290
rect 22161 3236 22217 3238
rect 22241 3236 22297 3238
rect 22321 3236 22377 3238
rect 22401 3236 22457 3238
rect 22161 2202 22217 2204
rect 22241 2202 22297 2204
rect 22321 2202 22377 2204
rect 22401 2202 22457 2204
rect 22161 2150 22207 2202
rect 22207 2150 22217 2202
rect 22241 2150 22271 2202
rect 22271 2150 22283 2202
rect 22283 2150 22297 2202
rect 22321 2150 22335 2202
rect 22335 2150 22347 2202
rect 22347 2150 22377 2202
rect 22401 2150 22411 2202
rect 22411 2150 22457 2202
rect 22161 2148 22217 2150
rect 22241 2148 22297 2150
rect 22321 2148 22377 2150
rect 22401 2148 22457 2150
rect 27463 7098 27519 7100
rect 27543 7098 27599 7100
rect 27623 7098 27679 7100
rect 27703 7098 27759 7100
rect 27463 7046 27509 7098
rect 27509 7046 27519 7098
rect 27543 7046 27573 7098
rect 27573 7046 27585 7098
rect 27585 7046 27599 7098
rect 27623 7046 27637 7098
rect 27637 7046 27649 7098
rect 27649 7046 27679 7098
rect 27703 7046 27713 7098
rect 27713 7046 27759 7098
rect 27463 7044 27519 7046
rect 27543 7044 27599 7046
rect 27623 7044 27679 7046
rect 27703 7044 27759 7046
rect 27463 6010 27519 6012
rect 27543 6010 27599 6012
rect 27623 6010 27679 6012
rect 27703 6010 27759 6012
rect 27463 5958 27509 6010
rect 27509 5958 27519 6010
rect 27543 5958 27573 6010
rect 27573 5958 27585 6010
rect 27585 5958 27599 6010
rect 27623 5958 27637 6010
rect 27637 5958 27649 6010
rect 27649 5958 27679 6010
rect 27703 5958 27713 6010
rect 27713 5958 27759 6010
rect 27463 5956 27519 5958
rect 27543 5956 27599 5958
rect 27623 5956 27679 5958
rect 27703 5956 27759 5958
rect 27463 4922 27519 4924
rect 27543 4922 27599 4924
rect 27623 4922 27679 4924
rect 27703 4922 27759 4924
rect 27463 4870 27509 4922
rect 27509 4870 27519 4922
rect 27543 4870 27573 4922
rect 27573 4870 27585 4922
rect 27585 4870 27599 4922
rect 27623 4870 27637 4922
rect 27637 4870 27649 4922
rect 27649 4870 27679 4922
rect 27703 4870 27713 4922
rect 27713 4870 27759 4922
rect 27463 4868 27519 4870
rect 27543 4868 27599 4870
rect 27623 4868 27679 4870
rect 27703 4868 27759 4870
rect 27250 4528 27306 4584
rect 23478 856 23534 912
rect 23938 2080 23994 2136
rect 25226 1808 25282 1864
rect 26054 2896 26110 2952
rect 25870 1536 25926 1592
rect 27894 3984 27950 4040
rect 27463 3834 27519 3836
rect 27543 3834 27599 3836
rect 27623 3834 27679 3836
rect 27703 3834 27759 3836
rect 27463 3782 27509 3834
rect 27509 3782 27519 3834
rect 27543 3782 27573 3834
rect 27573 3782 27585 3834
rect 27585 3782 27599 3834
rect 27623 3782 27637 3834
rect 27637 3782 27649 3834
rect 27649 3782 27679 3834
rect 27703 3782 27713 3834
rect 27713 3782 27759 3834
rect 27463 3780 27519 3782
rect 27543 3780 27599 3782
rect 27623 3780 27679 3782
rect 27703 3780 27759 3782
rect 26054 1808 26110 1864
rect 26974 3032 27030 3088
rect 27463 2746 27519 2748
rect 27543 2746 27599 2748
rect 27623 2746 27679 2748
rect 27703 2746 27759 2748
rect 27463 2694 27509 2746
rect 27509 2694 27519 2746
rect 27543 2694 27573 2746
rect 27573 2694 27585 2746
rect 27585 2694 27599 2746
rect 27623 2694 27637 2746
rect 27637 2694 27649 2746
rect 27649 2694 27679 2746
rect 27703 2694 27713 2746
rect 27713 2694 27759 2746
rect 27463 2692 27519 2694
rect 27543 2692 27599 2694
rect 27623 2692 27679 2694
rect 27703 2692 27759 2694
rect 28170 2760 28226 2816
rect 28078 2216 28134 2272
rect 28446 3576 28502 3632
rect 28814 2796 28816 2816
rect 28816 2796 28868 2816
rect 28868 2796 28870 2816
rect 28814 2760 28870 2796
rect 29366 2896 29422 2952
rect 30470 2352 30526 2408
rect 30838 1400 30894 1456
rect 32764 6554 32820 6556
rect 32844 6554 32900 6556
rect 32924 6554 32980 6556
rect 33004 6554 33060 6556
rect 32764 6502 32810 6554
rect 32810 6502 32820 6554
rect 32844 6502 32874 6554
rect 32874 6502 32886 6554
rect 32886 6502 32900 6554
rect 32924 6502 32938 6554
rect 32938 6502 32950 6554
rect 32950 6502 32980 6554
rect 33004 6502 33014 6554
rect 33014 6502 33060 6554
rect 32764 6500 32820 6502
rect 32844 6500 32900 6502
rect 32924 6500 32980 6502
rect 33004 6500 33060 6502
rect 32764 5466 32820 5468
rect 32844 5466 32900 5468
rect 32924 5466 32980 5468
rect 33004 5466 33060 5468
rect 32764 5414 32810 5466
rect 32810 5414 32820 5466
rect 32844 5414 32874 5466
rect 32874 5414 32886 5466
rect 32886 5414 32900 5466
rect 32924 5414 32938 5466
rect 32938 5414 32950 5466
rect 32950 5414 32980 5466
rect 33004 5414 33014 5466
rect 33014 5414 33060 5466
rect 32764 5412 32820 5414
rect 32844 5412 32900 5414
rect 32924 5412 32980 5414
rect 33004 5412 33060 5414
rect 32764 4378 32820 4380
rect 32844 4378 32900 4380
rect 32924 4378 32980 4380
rect 33004 4378 33060 4380
rect 32764 4326 32810 4378
rect 32810 4326 32820 4378
rect 32844 4326 32874 4378
rect 32874 4326 32886 4378
rect 32886 4326 32900 4378
rect 32924 4326 32938 4378
rect 32938 4326 32950 4378
rect 32950 4326 32980 4378
rect 33004 4326 33014 4378
rect 33014 4326 33060 4378
rect 32764 4324 32820 4326
rect 32844 4324 32900 4326
rect 32924 4324 32980 4326
rect 33004 4324 33060 4326
rect 32218 2080 32274 2136
rect 32034 1264 32090 1320
rect 31942 992 31998 1048
rect 32764 3290 32820 3292
rect 32844 3290 32900 3292
rect 32924 3290 32980 3292
rect 33004 3290 33060 3292
rect 32764 3238 32810 3290
rect 32810 3238 32820 3290
rect 32844 3238 32874 3290
rect 32874 3238 32886 3290
rect 32886 3238 32900 3290
rect 32924 3238 32938 3290
rect 32938 3238 32950 3290
rect 32950 3238 32980 3290
rect 33004 3238 33014 3290
rect 33014 3238 33060 3290
rect 32764 3236 32820 3238
rect 32844 3236 32900 3238
rect 32924 3236 32980 3238
rect 33004 3236 33060 3238
rect 32770 2760 32826 2816
rect 33138 2508 33194 2544
rect 33138 2488 33140 2508
rect 33140 2488 33192 2508
rect 33192 2488 33194 2508
rect 32764 2202 32820 2204
rect 32844 2202 32900 2204
rect 32924 2202 32980 2204
rect 33004 2202 33060 2204
rect 32764 2150 32810 2202
rect 32810 2150 32820 2202
rect 32844 2150 32874 2202
rect 32874 2150 32886 2202
rect 32886 2150 32900 2202
rect 32924 2150 32938 2202
rect 32938 2150 32950 2202
rect 32950 2150 32980 2202
rect 33004 2150 33014 2202
rect 33014 2150 33060 2202
rect 32764 2148 32820 2150
rect 32844 2148 32900 2150
rect 32924 2148 32980 2150
rect 33004 2148 33060 2150
rect 34794 1808 34850 1864
rect 38066 7098 38122 7100
rect 38146 7098 38202 7100
rect 38226 7098 38282 7100
rect 38306 7098 38362 7100
rect 38066 7046 38112 7098
rect 38112 7046 38122 7098
rect 38146 7046 38176 7098
rect 38176 7046 38188 7098
rect 38188 7046 38202 7098
rect 38226 7046 38240 7098
rect 38240 7046 38252 7098
rect 38252 7046 38282 7098
rect 38306 7046 38316 7098
rect 38316 7046 38362 7098
rect 38066 7044 38122 7046
rect 38146 7044 38202 7046
rect 38226 7044 38282 7046
rect 38306 7044 38362 7046
rect 38066 6010 38122 6012
rect 38146 6010 38202 6012
rect 38226 6010 38282 6012
rect 38306 6010 38362 6012
rect 38066 5958 38112 6010
rect 38112 5958 38122 6010
rect 38146 5958 38176 6010
rect 38176 5958 38188 6010
rect 38188 5958 38202 6010
rect 38226 5958 38240 6010
rect 38240 5958 38252 6010
rect 38252 5958 38282 6010
rect 38306 5958 38316 6010
rect 38316 5958 38362 6010
rect 38066 5956 38122 5958
rect 38146 5956 38202 5958
rect 38226 5956 38282 5958
rect 38306 5956 38362 5958
rect 37002 2644 37058 2680
rect 37002 2624 37004 2644
rect 37004 2624 37056 2644
rect 37056 2624 37058 2644
rect 38066 4922 38122 4924
rect 38146 4922 38202 4924
rect 38226 4922 38282 4924
rect 38306 4922 38362 4924
rect 38066 4870 38112 4922
rect 38112 4870 38122 4922
rect 38146 4870 38176 4922
rect 38176 4870 38188 4922
rect 38188 4870 38202 4922
rect 38226 4870 38240 4922
rect 38240 4870 38252 4922
rect 38252 4870 38282 4922
rect 38306 4870 38316 4922
rect 38316 4870 38362 4922
rect 38066 4868 38122 4870
rect 38146 4868 38202 4870
rect 38226 4868 38282 4870
rect 38306 4868 38362 4870
rect 38066 3834 38122 3836
rect 38146 3834 38202 3836
rect 38226 3834 38282 3836
rect 38306 3834 38362 3836
rect 38066 3782 38112 3834
rect 38112 3782 38122 3834
rect 38146 3782 38176 3834
rect 38176 3782 38188 3834
rect 38188 3782 38202 3834
rect 38226 3782 38240 3834
rect 38240 3782 38252 3834
rect 38252 3782 38282 3834
rect 38306 3782 38316 3834
rect 38316 3782 38362 3834
rect 38066 3780 38122 3782
rect 38146 3780 38202 3782
rect 38226 3780 38282 3782
rect 38306 3780 38362 3782
rect 38066 2746 38122 2748
rect 38146 2746 38202 2748
rect 38226 2746 38282 2748
rect 38306 2746 38362 2748
rect 38066 2694 38112 2746
rect 38112 2694 38122 2746
rect 38146 2694 38176 2746
rect 38176 2694 38188 2746
rect 38188 2694 38202 2746
rect 38226 2694 38240 2746
rect 38240 2694 38252 2746
rect 38252 2694 38282 2746
rect 38306 2694 38316 2746
rect 38316 2694 38362 2746
rect 38066 2692 38122 2694
rect 38146 2692 38202 2694
rect 38226 2692 38282 2694
rect 38306 2692 38362 2694
rect 43367 6554 43423 6556
rect 43447 6554 43503 6556
rect 43527 6554 43583 6556
rect 43607 6554 43663 6556
rect 43367 6502 43413 6554
rect 43413 6502 43423 6554
rect 43447 6502 43477 6554
rect 43477 6502 43489 6554
rect 43489 6502 43503 6554
rect 43527 6502 43541 6554
rect 43541 6502 43553 6554
rect 43553 6502 43583 6554
rect 43607 6502 43617 6554
rect 43617 6502 43663 6554
rect 43367 6500 43423 6502
rect 43447 6500 43503 6502
rect 43527 6500 43583 6502
rect 43607 6500 43663 6502
rect 43367 5466 43423 5468
rect 43447 5466 43503 5468
rect 43527 5466 43583 5468
rect 43607 5466 43663 5468
rect 43367 5414 43413 5466
rect 43413 5414 43423 5466
rect 43447 5414 43477 5466
rect 43477 5414 43489 5466
rect 43489 5414 43503 5466
rect 43527 5414 43541 5466
rect 43541 5414 43553 5466
rect 43553 5414 43583 5466
rect 43607 5414 43617 5466
rect 43617 5414 43663 5466
rect 43367 5412 43423 5414
rect 43447 5412 43503 5414
rect 43527 5412 43583 5414
rect 43607 5412 43663 5414
rect 43367 4378 43423 4380
rect 43447 4378 43503 4380
rect 43527 4378 43583 4380
rect 43607 4378 43663 4380
rect 43367 4326 43413 4378
rect 43413 4326 43423 4378
rect 43447 4326 43477 4378
rect 43477 4326 43489 4378
rect 43489 4326 43503 4378
rect 43527 4326 43541 4378
rect 43541 4326 43553 4378
rect 43553 4326 43583 4378
rect 43607 4326 43617 4378
rect 43617 4326 43663 4378
rect 43367 4324 43423 4326
rect 43447 4324 43503 4326
rect 43527 4324 43583 4326
rect 43607 4324 43663 4326
rect 43367 3290 43423 3292
rect 43447 3290 43503 3292
rect 43527 3290 43583 3292
rect 43607 3290 43663 3292
rect 43367 3238 43413 3290
rect 43413 3238 43423 3290
rect 43447 3238 43477 3290
rect 43477 3238 43489 3290
rect 43489 3238 43503 3290
rect 43527 3238 43541 3290
rect 43541 3238 43553 3290
rect 43553 3238 43583 3290
rect 43607 3238 43617 3290
rect 43617 3238 43663 3290
rect 43367 3236 43423 3238
rect 43447 3236 43503 3238
rect 43527 3236 43583 3238
rect 43607 3236 43663 3238
rect 43367 2202 43423 2204
rect 43447 2202 43503 2204
rect 43527 2202 43583 2204
rect 43607 2202 43663 2204
rect 43367 2150 43413 2202
rect 43413 2150 43423 2202
rect 43447 2150 43477 2202
rect 43477 2150 43489 2202
rect 43489 2150 43503 2202
rect 43527 2150 43541 2202
rect 43541 2150 43553 2202
rect 43553 2150 43583 2202
rect 43607 2150 43617 2202
rect 43617 2150 43663 2202
rect 43367 2148 43423 2150
rect 43447 2148 43503 2150
rect 43527 2148 43583 2150
rect 43607 2148 43663 2150
<< metal3 >>
rect 11548 7648 11864 7649
rect 11548 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11864 7648
rect 11548 7583 11864 7584
rect 22151 7648 22467 7649
rect 22151 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22467 7648
rect 22151 7583 22467 7584
rect 32754 7648 33070 7649
rect 32754 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33070 7648
rect 32754 7583 33070 7584
rect 43357 7648 43673 7649
rect 43357 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43673 7648
rect 43357 7583 43673 7584
rect 6247 7104 6563 7105
rect 6247 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6563 7104
rect 6247 7039 6563 7040
rect 16850 7104 17166 7105
rect 16850 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17166 7104
rect 16850 7039 17166 7040
rect 27453 7104 27769 7105
rect 27453 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27769 7104
rect 27453 7039 27769 7040
rect 38056 7104 38372 7105
rect 38056 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38372 7104
rect 38056 7039 38372 7040
rect 11548 6560 11864 6561
rect 11548 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11864 6560
rect 11548 6495 11864 6496
rect 22151 6560 22467 6561
rect 22151 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22467 6560
rect 22151 6495 22467 6496
rect 32754 6560 33070 6561
rect 32754 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33070 6560
rect 32754 6495 33070 6496
rect 43357 6560 43673 6561
rect 43357 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43673 6560
rect 43357 6495 43673 6496
rect 6247 6016 6563 6017
rect 6247 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6563 6016
rect 6247 5951 6563 5952
rect 16850 6016 17166 6017
rect 16850 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17166 6016
rect 16850 5951 17166 5952
rect 27453 6016 27769 6017
rect 27453 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27769 6016
rect 27453 5951 27769 5952
rect 38056 6016 38372 6017
rect 38056 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38372 6016
rect 38056 5951 38372 5952
rect 11548 5472 11864 5473
rect 11548 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11864 5472
rect 11548 5407 11864 5408
rect 22151 5472 22467 5473
rect 22151 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22467 5472
rect 22151 5407 22467 5408
rect 32754 5472 33070 5473
rect 32754 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33070 5472
rect 32754 5407 33070 5408
rect 43357 5472 43673 5473
rect 43357 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43673 5472
rect 43357 5407 43673 5408
rect 16481 5130 16547 5133
rect 36486 5130 36492 5132
rect 16481 5128 36492 5130
rect 16481 5072 16486 5128
rect 16542 5072 36492 5128
rect 16481 5070 36492 5072
rect 16481 5067 16547 5070
rect 36486 5068 36492 5070
rect 36556 5068 36562 5132
rect 6247 4928 6563 4929
rect 6247 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6563 4928
rect 6247 4863 6563 4864
rect 16850 4928 17166 4929
rect 16850 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17166 4928
rect 16850 4863 17166 4864
rect 27453 4928 27769 4929
rect 27453 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27769 4928
rect 27453 4863 27769 4864
rect 38056 4928 38372 4929
rect 38056 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38372 4928
rect 38056 4863 38372 4864
rect 13445 4586 13511 4589
rect 27245 4586 27311 4589
rect 13445 4584 27311 4586
rect 13445 4528 13450 4584
rect 13506 4528 27250 4584
rect 27306 4528 27311 4584
rect 13445 4526 27311 4528
rect 13445 4523 13511 4526
rect 27245 4523 27311 4526
rect 11548 4384 11864 4385
rect 11548 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11864 4384
rect 11548 4319 11864 4320
rect 22151 4384 22467 4385
rect 22151 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22467 4384
rect 22151 4319 22467 4320
rect 32754 4384 33070 4385
rect 32754 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33070 4384
rect 32754 4319 33070 4320
rect 43357 4384 43673 4385
rect 43357 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43673 4384
rect 43357 4319 43673 4320
rect 12985 4314 13051 4317
rect 20621 4314 20687 4317
rect 12985 4312 20687 4314
rect 12985 4256 12990 4312
rect 13046 4256 20626 4312
rect 20682 4256 20687 4312
rect 12985 4254 20687 4256
rect 12985 4251 13051 4254
rect 20621 4251 20687 4254
rect 12801 4042 12867 4045
rect 22093 4042 22159 4045
rect 27889 4042 27955 4045
rect 12801 4040 22159 4042
rect 12801 3984 12806 4040
rect 12862 3984 22098 4040
rect 22154 3984 22159 4040
rect 12801 3982 22159 3984
rect 12801 3979 12867 3982
rect 22093 3979 22159 3982
rect 26190 4040 27955 4042
rect 26190 3984 27894 4040
rect 27950 3984 27955 4040
rect 26190 3982 27955 3984
rect 6247 3840 6563 3841
rect 6247 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6563 3840
rect 6247 3775 6563 3776
rect 16850 3840 17166 3841
rect 16850 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17166 3840
rect 16850 3775 17166 3776
rect 26190 3770 26250 3982
rect 27889 3979 27955 3982
rect 27453 3840 27769 3841
rect 27453 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27769 3840
rect 27453 3775 27769 3776
rect 38056 3840 38372 3841
rect 38056 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38372 3840
rect 38056 3775 38372 3776
rect 21406 3710 26250 3770
rect 11329 3634 11395 3637
rect 21406 3634 21466 3710
rect 28441 3634 28507 3637
rect 11329 3632 21466 3634
rect 11329 3576 11334 3632
rect 11390 3576 21466 3632
rect 11329 3574 21466 3576
rect 21958 3632 28507 3634
rect 21958 3576 28446 3632
rect 28502 3576 28507 3632
rect 21958 3574 28507 3576
rect 11329 3571 11395 3574
rect 9305 3498 9371 3501
rect 17861 3498 17927 3501
rect 9305 3496 17927 3498
rect 9305 3440 9310 3496
rect 9366 3440 17866 3496
rect 17922 3440 17927 3496
rect 9305 3438 17927 3440
rect 9305 3435 9371 3438
rect 17861 3435 17927 3438
rect 21958 3362 22018 3574
rect 28441 3571 28507 3574
rect 12022 3302 22018 3362
rect 11548 3296 11864 3297
rect 11548 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11864 3296
rect 11548 3231 11864 3232
rect 10777 3090 10843 3093
rect 12022 3090 12082 3302
rect 22151 3296 22467 3297
rect 22151 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22467 3296
rect 22151 3231 22467 3232
rect 32754 3296 33070 3297
rect 32754 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33070 3296
rect 32754 3231 33070 3232
rect 43357 3296 43673 3297
rect 43357 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43673 3296
rect 43357 3231 43673 3232
rect 12249 3226 12315 3229
rect 12249 3224 21466 3226
rect 12249 3168 12254 3224
rect 12310 3168 21466 3224
rect 12249 3166 21466 3168
rect 12249 3163 12315 3166
rect 10777 3088 12082 3090
rect 10777 3032 10782 3088
rect 10838 3032 12082 3088
rect 10777 3030 12082 3032
rect 15377 3090 15443 3093
rect 21406 3090 21466 3166
rect 26969 3090 27035 3093
rect 15377 3088 21282 3090
rect 15377 3032 15382 3088
rect 15438 3032 21282 3088
rect 15377 3030 21282 3032
rect 21406 3088 27035 3090
rect 21406 3032 26974 3088
rect 27030 3032 27035 3088
rect 21406 3030 27035 3032
rect 10777 3027 10843 3030
rect 15377 3027 15443 3030
rect 5073 2954 5139 2957
rect 19793 2954 19859 2957
rect 5073 2952 19859 2954
rect 5073 2896 5078 2952
rect 5134 2896 19798 2952
rect 19854 2896 19859 2952
rect 5073 2894 19859 2896
rect 21222 2954 21282 3030
rect 26969 3027 27035 3030
rect 26049 2954 26115 2957
rect 29361 2954 29427 2957
rect 21222 2952 26115 2954
rect 21222 2896 26054 2952
rect 26110 2896 26115 2952
rect 21222 2894 26115 2896
rect 5073 2891 5139 2894
rect 19793 2891 19859 2894
rect 26049 2891 26115 2894
rect 26190 2952 29427 2954
rect 26190 2896 29366 2952
rect 29422 2896 29427 2952
rect 26190 2894 29427 2896
rect 18505 2818 18571 2821
rect 26190 2818 26250 2894
rect 29361 2891 29427 2894
rect 18505 2816 26250 2818
rect 18505 2760 18510 2816
rect 18566 2760 26250 2816
rect 18505 2758 26250 2760
rect 28165 2818 28231 2821
rect 28809 2818 28875 2821
rect 28165 2816 28875 2818
rect 28165 2760 28170 2816
rect 28226 2760 28814 2816
rect 28870 2760 28875 2816
rect 28165 2758 28875 2760
rect 18505 2755 18571 2758
rect 28165 2755 28231 2758
rect 28809 2755 28875 2758
rect 30414 2756 30420 2820
rect 30484 2818 30490 2820
rect 32765 2818 32831 2821
rect 30484 2816 32831 2818
rect 30484 2760 32770 2816
rect 32826 2760 32831 2816
rect 30484 2758 32831 2760
rect 30484 2756 30490 2758
rect 32765 2755 32831 2758
rect 6247 2752 6563 2753
rect 6247 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6563 2752
rect 6247 2687 6563 2688
rect 16850 2752 17166 2753
rect 16850 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17166 2752
rect 16850 2687 17166 2688
rect 27453 2752 27769 2753
rect 27453 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27769 2752
rect 27453 2687 27769 2688
rect 38056 2752 38372 2753
rect 38056 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38372 2752
rect 38056 2687 38372 2688
rect 36486 2620 36492 2684
rect 36556 2682 36562 2684
rect 36997 2682 37063 2685
rect 36556 2680 37063 2682
rect 36556 2624 37002 2680
rect 37058 2624 37063 2680
rect 36556 2622 37063 2624
rect 36556 2620 36562 2622
rect 36997 2619 37063 2622
rect 13629 2546 13695 2549
rect 17401 2546 17467 2549
rect 33133 2546 33199 2549
rect 13629 2544 17467 2546
rect 13629 2488 13634 2544
rect 13690 2488 17406 2544
rect 17462 2488 17467 2544
rect 13629 2486 17467 2488
rect 13629 2483 13695 2486
rect 17401 2483 17467 2486
rect 18830 2544 33199 2546
rect 18830 2488 33138 2544
rect 33194 2488 33199 2544
rect 18830 2486 33199 2488
rect 17309 2410 17375 2413
rect 18830 2410 18890 2486
rect 33133 2483 33199 2486
rect 17309 2408 18890 2410
rect 17309 2352 17314 2408
rect 17370 2352 18890 2408
rect 17309 2350 18890 2352
rect 18965 2410 19031 2413
rect 30465 2410 30531 2413
rect 18965 2408 30531 2410
rect 18965 2352 18970 2408
rect 19026 2352 30470 2408
rect 30526 2352 30531 2408
rect 18965 2350 30531 2352
rect 17309 2347 17375 2350
rect 18965 2347 19031 2350
rect 30465 2347 30531 2350
rect 28073 2274 28139 2277
rect 22694 2272 28139 2274
rect 22694 2216 28078 2272
rect 28134 2216 28139 2272
rect 22694 2214 28139 2216
rect 11548 2208 11864 2209
rect 11548 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11864 2208
rect 11548 2143 11864 2144
rect 22151 2208 22467 2209
rect 22151 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22467 2208
rect 22151 2143 22467 2144
rect 12157 2138 12223 2141
rect 19425 2138 19491 2141
rect 12157 2136 19491 2138
rect 12157 2080 12162 2136
rect 12218 2080 19430 2136
rect 19486 2080 19491 2136
rect 12157 2078 19491 2080
rect 12157 2075 12223 2078
rect 19425 2075 19491 2078
rect 11329 2002 11395 2005
rect 22694 2002 22754 2214
rect 28073 2211 28139 2214
rect 32754 2208 33070 2209
rect 32754 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33070 2208
rect 32754 2143 33070 2144
rect 43357 2208 43673 2209
rect 43357 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43673 2208
rect 43357 2143 43673 2144
rect 23933 2138 23999 2141
rect 32213 2138 32279 2141
rect 23933 2136 32279 2138
rect 23933 2080 23938 2136
rect 23994 2080 32218 2136
rect 32274 2080 32279 2136
rect 23933 2078 32279 2080
rect 23933 2075 23999 2078
rect 32213 2075 32279 2078
rect 11329 2000 22754 2002
rect 11329 1944 11334 2000
rect 11390 1944 22754 2000
rect 11329 1942 22754 1944
rect 11329 1939 11395 1942
rect 13629 1866 13695 1869
rect 25221 1866 25287 1869
rect 13629 1864 25287 1866
rect 13629 1808 13634 1864
rect 13690 1808 25226 1864
rect 25282 1808 25287 1864
rect 13629 1806 25287 1808
rect 13629 1803 13695 1806
rect 25221 1803 25287 1806
rect 26049 1866 26115 1869
rect 34789 1866 34855 1869
rect 26049 1864 34855 1866
rect 26049 1808 26054 1864
rect 26110 1808 34794 1864
rect 34850 1808 34855 1864
rect 26049 1806 34855 1808
rect 26049 1803 26115 1806
rect 34789 1803 34855 1806
rect 8753 1730 8819 1733
rect 18781 1730 18847 1733
rect 8753 1728 18847 1730
rect 8753 1672 8758 1728
rect 8814 1672 18786 1728
rect 18842 1672 18847 1728
rect 8753 1670 18847 1672
rect 8753 1667 8819 1670
rect 18781 1667 18847 1670
rect 13077 1594 13143 1597
rect 25865 1594 25931 1597
rect 13077 1592 25931 1594
rect 13077 1536 13082 1592
rect 13138 1536 25870 1592
rect 25926 1536 25931 1592
rect 13077 1534 25931 1536
rect 13077 1531 13143 1534
rect 25865 1531 25931 1534
rect 17125 1458 17191 1461
rect 30833 1458 30899 1461
rect 17125 1456 30899 1458
rect 17125 1400 17130 1456
rect 17186 1400 30838 1456
rect 30894 1400 30899 1456
rect 17125 1398 30899 1400
rect 17125 1395 17191 1398
rect 30833 1395 30899 1398
rect 15377 1322 15443 1325
rect 32029 1322 32095 1325
rect 15377 1320 32095 1322
rect 15377 1264 15382 1320
rect 15438 1264 32034 1320
rect 32090 1264 32095 1320
rect 15377 1262 32095 1264
rect 15377 1259 15443 1262
rect 32029 1259 32095 1262
rect 16389 1186 16455 1189
rect 30414 1186 30420 1188
rect 16389 1184 30420 1186
rect 16389 1128 16394 1184
rect 16450 1128 30420 1184
rect 16389 1126 30420 1128
rect 16389 1123 16455 1126
rect 30414 1124 30420 1126
rect 30484 1124 30490 1188
rect 17677 1050 17743 1053
rect 31937 1050 32003 1053
rect 17677 1048 32003 1050
rect 17677 992 17682 1048
rect 17738 992 31942 1048
rect 31998 992 32003 1048
rect 17677 990 32003 992
rect 17677 987 17743 990
rect 31937 987 32003 990
rect 6913 914 6979 917
rect 23473 914 23539 917
rect 6913 912 23539 914
rect 6913 856 6918 912
rect 6974 856 23478 912
rect 23534 856 23539 912
rect 6913 854 23539 856
rect 6913 851 6979 854
rect 23473 851 23539 854
<< via3 >>
rect 11554 7644 11618 7648
rect 11554 7588 11558 7644
rect 11558 7588 11614 7644
rect 11614 7588 11618 7644
rect 11554 7584 11618 7588
rect 11634 7644 11698 7648
rect 11634 7588 11638 7644
rect 11638 7588 11694 7644
rect 11694 7588 11698 7644
rect 11634 7584 11698 7588
rect 11714 7644 11778 7648
rect 11714 7588 11718 7644
rect 11718 7588 11774 7644
rect 11774 7588 11778 7644
rect 11714 7584 11778 7588
rect 11794 7644 11858 7648
rect 11794 7588 11798 7644
rect 11798 7588 11854 7644
rect 11854 7588 11858 7644
rect 11794 7584 11858 7588
rect 22157 7644 22221 7648
rect 22157 7588 22161 7644
rect 22161 7588 22217 7644
rect 22217 7588 22221 7644
rect 22157 7584 22221 7588
rect 22237 7644 22301 7648
rect 22237 7588 22241 7644
rect 22241 7588 22297 7644
rect 22297 7588 22301 7644
rect 22237 7584 22301 7588
rect 22317 7644 22381 7648
rect 22317 7588 22321 7644
rect 22321 7588 22377 7644
rect 22377 7588 22381 7644
rect 22317 7584 22381 7588
rect 22397 7644 22461 7648
rect 22397 7588 22401 7644
rect 22401 7588 22457 7644
rect 22457 7588 22461 7644
rect 22397 7584 22461 7588
rect 32760 7644 32824 7648
rect 32760 7588 32764 7644
rect 32764 7588 32820 7644
rect 32820 7588 32824 7644
rect 32760 7584 32824 7588
rect 32840 7644 32904 7648
rect 32840 7588 32844 7644
rect 32844 7588 32900 7644
rect 32900 7588 32904 7644
rect 32840 7584 32904 7588
rect 32920 7644 32984 7648
rect 32920 7588 32924 7644
rect 32924 7588 32980 7644
rect 32980 7588 32984 7644
rect 32920 7584 32984 7588
rect 33000 7644 33064 7648
rect 33000 7588 33004 7644
rect 33004 7588 33060 7644
rect 33060 7588 33064 7644
rect 33000 7584 33064 7588
rect 43363 7644 43427 7648
rect 43363 7588 43367 7644
rect 43367 7588 43423 7644
rect 43423 7588 43427 7644
rect 43363 7584 43427 7588
rect 43443 7644 43507 7648
rect 43443 7588 43447 7644
rect 43447 7588 43503 7644
rect 43503 7588 43507 7644
rect 43443 7584 43507 7588
rect 43523 7644 43587 7648
rect 43523 7588 43527 7644
rect 43527 7588 43583 7644
rect 43583 7588 43587 7644
rect 43523 7584 43587 7588
rect 43603 7644 43667 7648
rect 43603 7588 43607 7644
rect 43607 7588 43663 7644
rect 43663 7588 43667 7644
rect 43603 7584 43667 7588
rect 6253 7100 6317 7104
rect 6253 7044 6257 7100
rect 6257 7044 6313 7100
rect 6313 7044 6317 7100
rect 6253 7040 6317 7044
rect 6333 7100 6397 7104
rect 6333 7044 6337 7100
rect 6337 7044 6393 7100
rect 6393 7044 6397 7100
rect 6333 7040 6397 7044
rect 6413 7100 6477 7104
rect 6413 7044 6417 7100
rect 6417 7044 6473 7100
rect 6473 7044 6477 7100
rect 6413 7040 6477 7044
rect 6493 7100 6557 7104
rect 6493 7044 6497 7100
rect 6497 7044 6553 7100
rect 6553 7044 6557 7100
rect 6493 7040 6557 7044
rect 16856 7100 16920 7104
rect 16856 7044 16860 7100
rect 16860 7044 16916 7100
rect 16916 7044 16920 7100
rect 16856 7040 16920 7044
rect 16936 7100 17000 7104
rect 16936 7044 16940 7100
rect 16940 7044 16996 7100
rect 16996 7044 17000 7100
rect 16936 7040 17000 7044
rect 17016 7100 17080 7104
rect 17016 7044 17020 7100
rect 17020 7044 17076 7100
rect 17076 7044 17080 7100
rect 17016 7040 17080 7044
rect 17096 7100 17160 7104
rect 17096 7044 17100 7100
rect 17100 7044 17156 7100
rect 17156 7044 17160 7100
rect 17096 7040 17160 7044
rect 27459 7100 27523 7104
rect 27459 7044 27463 7100
rect 27463 7044 27519 7100
rect 27519 7044 27523 7100
rect 27459 7040 27523 7044
rect 27539 7100 27603 7104
rect 27539 7044 27543 7100
rect 27543 7044 27599 7100
rect 27599 7044 27603 7100
rect 27539 7040 27603 7044
rect 27619 7100 27683 7104
rect 27619 7044 27623 7100
rect 27623 7044 27679 7100
rect 27679 7044 27683 7100
rect 27619 7040 27683 7044
rect 27699 7100 27763 7104
rect 27699 7044 27703 7100
rect 27703 7044 27759 7100
rect 27759 7044 27763 7100
rect 27699 7040 27763 7044
rect 38062 7100 38126 7104
rect 38062 7044 38066 7100
rect 38066 7044 38122 7100
rect 38122 7044 38126 7100
rect 38062 7040 38126 7044
rect 38142 7100 38206 7104
rect 38142 7044 38146 7100
rect 38146 7044 38202 7100
rect 38202 7044 38206 7100
rect 38142 7040 38206 7044
rect 38222 7100 38286 7104
rect 38222 7044 38226 7100
rect 38226 7044 38282 7100
rect 38282 7044 38286 7100
rect 38222 7040 38286 7044
rect 38302 7100 38366 7104
rect 38302 7044 38306 7100
rect 38306 7044 38362 7100
rect 38362 7044 38366 7100
rect 38302 7040 38366 7044
rect 11554 6556 11618 6560
rect 11554 6500 11558 6556
rect 11558 6500 11614 6556
rect 11614 6500 11618 6556
rect 11554 6496 11618 6500
rect 11634 6556 11698 6560
rect 11634 6500 11638 6556
rect 11638 6500 11694 6556
rect 11694 6500 11698 6556
rect 11634 6496 11698 6500
rect 11714 6556 11778 6560
rect 11714 6500 11718 6556
rect 11718 6500 11774 6556
rect 11774 6500 11778 6556
rect 11714 6496 11778 6500
rect 11794 6556 11858 6560
rect 11794 6500 11798 6556
rect 11798 6500 11854 6556
rect 11854 6500 11858 6556
rect 11794 6496 11858 6500
rect 22157 6556 22221 6560
rect 22157 6500 22161 6556
rect 22161 6500 22217 6556
rect 22217 6500 22221 6556
rect 22157 6496 22221 6500
rect 22237 6556 22301 6560
rect 22237 6500 22241 6556
rect 22241 6500 22297 6556
rect 22297 6500 22301 6556
rect 22237 6496 22301 6500
rect 22317 6556 22381 6560
rect 22317 6500 22321 6556
rect 22321 6500 22377 6556
rect 22377 6500 22381 6556
rect 22317 6496 22381 6500
rect 22397 6556 22461 6560
rect 22397 6500 22401 6556
rect 22401 6500 22457 6556
rect 22457 6500 22461 6556
rect 22397 6496 22461 6500
rect 32760 6556 32824 6560
rect 32760 6500 32764 6556
rect 32764 6500 32820 6556
rect 32820 6500 32824 6556
rect 32760 6496 32824 6500
rect 32840 6556 32904 6560
rect 32840 6500 32844 6556
rect 32844 6500 32900 6556
rect 32900 6500 32904 6556
rect 32840 6496 32904 6500
rect 32920 6556 32984 6560
rect 32920 6500 32924 6556
rect 32924 6500 32980 6556
rect 32980 6500 32984 6556
rect 32920 6496 32984 6500
rect 33000 6556 33064 6560
rect 33000 6500 33004 6556
rect 33004 6500 33060 6556
rect 33060 6500 33064 6556
rect 33000 6496 33064 6500
rect 43363 6556 43427 6560
rect 43363 6500 43367 6556
rect 43367 6500 43423 6556
rect 43423 6500 43427 6556
rect 43363 6496 43427 6500
rect 43443 6556 43507 6560
rect 43443 6500 43447 6556
rect 43447 6500 43503 6556
rect 43503 6500 43507 6556
rect 43443 6496 43507 6500
rect 43523 6556 43587 6560
rect 43523 6500 43527 6556
rect 43527 6500 43583 6556
rect 43583 6500 43587 6556
rect 43523 6496 43587 6500
rect 43603 6556 43667 6560
rect 43603 6500 43607 6556
rect 43607 6500 43663 6556
rect 43663 6500 43667 6556
rect 43603 6496 43667 6500
rect 6253 6012 6317 6016
rect 6253 5956 6257 6012
rect 6257 5956 6313 6012
rect 6313 5956 6317 6012
rect 6253 5952 6317 5956
rect 6333 6012 6397 6016
rect 6333 5956 6337 6012
rect 6337 5956 6393 6012
rect 6393 5956 6397 6012
rect 6333 5952 6397 5956
rect 6413 6012 6477 6016
rect 6413 5956 6417 6012
rect 6417 5956 6473 6012
rect 6473 5956 6477 6012
rect 6413 5952 6477 5956
rect 6493 6012 6557 6016
rect 6493 5956 6497 6012
rect 6497 5956 6553 6012
rect 6553 5956 6557 6012
rect 6493 5952 6557 5956
rect 16856 6012 16920 6016
rect 16856 5956 16860 6012
rect 16860 5956 16916 6012
rect 16916 5956 16920 6012
rect 16856 5952 16920 5956
rect 16936 6012 17000 6016
rect 16936 5956 16940 6012
rect 16940 5956 16996 6012
rect 16996 5956 17000 6012
rect 16936 5952 17000 5956
rect 17016 6012 17080 6016
rect 17016 5956 17020 6012
rect 17020 5956 17076 6012
rect 17076 5956 17080 6012
rect 17016 5952 17080 5956
rect 17096 6012 17160 6016
rect 17096 5956 17100 6012
rect 17100 5956 17156 6012
rect 17156 5956 17160 6012
rect 17096 5952 17160 5956
rect 27459 6012 27523 6016
rect 27459 5956 27463 6012
rect 27463 5956 27519 6012
rect 27519 5956 27523 6012
rect 27459 5952 27523 5956
rect 27539 6012 27603 6016
rect 27539 5956 27543 6012
rect 27543 5956 27599 6012
rect 27599 5956 27603 6012
rect 27539 5952 27603 5956
rect 27619 6012 27683 6016
rect 27619 5956 27623 6012
rect 27623 5956 27679 6012
rect 27679 5956 27683 6012
rect 27619 5952 27683 5956
rect 27699 6012 27763 6016
rect 27699 5956 27703 6012
rect 27703 5956 27759 6012
rect 27759 5956 27763 6012
rect 27699 5952 27763 5956
rect 38062 6012 38126 6016
rect 38062 5956 38066 6012
rect 38066 5956 38122 6012
rect 38122 5956 38126 6012
rect 38062 5952 38126 5956
rect 38142 6012 38206 6016
rect 38142 5956 38146 6012
rect 38146 5956 38202 6012
rect 38202 5956 38206 6012
rect 38142 5952 38206 5956
rect 38222 6012 38286 6016
rect 38222 5956 38226 6012
rect 38226 5956 38282 6012
rect 38282 5956 38286 6012
rect 38222 5952 38286 5956
rect 38302 6012 38366 6016
rect 38302 5956 38306 6012
rect 38306 5956 38362 6012
rect 38362 5956 38366 6012
rect 38302 5952 38366 5956
rect 11554 5468 11618 5472
rect 11554 5412 11558 5468
rect 11558 5412 11614 5468
rect 11614 5412 11618 5468
rect 11554 5408 11618 5412
rect 11634 5468 11698 5472
rect 11634 5412 11638 5468
rect 11638 5412 11694 5468
rect 11694 5412 11698 5468
rect 11634 5408 11698 5412
rect 11714 5468 11778 5472
rect 11714 5412 11718 5468
rect 11718 5412 11774 5468
rect 11774 5412 11778 5468
rect 11714 5408 11778 5412
rect 11794 5468 11858 5472
rect 11794 5412 11798 5468
rect 11798 5412 11854 5468
rect 11854 5412 11858 5468
rect 11794 5408 11858 5412
rect 22157 5468 22221 5472
rect 22157 5412 22161 5468
rect 22161 5412 22217 5468
rect 22217 5412 22221 5468
rect 22157 5408 22221 5412
rect 22237 5468 22301 5472
rect 22237 5412 22241 5468
rect 22241 5412 22297 5468
rect 22297 5412 22301 5468
rect 22237 5408 22301 5412
rect 22317 5468 22381 5472
rect 22317 5412 22321 5468
rect 22321 5412 22377 5468
rect 22377 5412 22381 5468
rect 22317 5408 22381 5412
rect 22397 5468 22461 5472
rect 22397 5412 22401 5468
rect 22401 5412 22457 5468
rect 22457 5412 22461 5468
rect 22397 5408 22461 5412
rect 32760 5468 32824 5472
rect 32760 5412 32764 5468
rect 32764 5412 32820 5468
rect 32820 5412 32824 5468
rect 32760 5408 32824 5412
rect 32840 5468 32904 5472
rect 32840 5412 32844 5468
rect 32844 5412 32900 5468
rect 32900 5412 32904 5468
rect 32840 5408 32904 5412
rect 32920 5468 32984 5472
rect 32920 5412 32924 5468
rect 32924 5412 32980 5468
rect 32980 5412 32984 5468
rect 32920 5408 32984 5412
rect 33000 5468 33064 5472
rect 33000 5412 33004 5468
rect 33004 5412 33060 5468
rect 33060 5412 33064 5468
rect 33000 5408 33064 5412
rect 43363 5468 43427 5472
rect 43363 5412 43367 5468
rect 43367 5412 43423 5468
rect 43423 5412 43427 5468
rect 43363 5408 43427 5412
rect 43443 5468 43507 5472
rect 43443 5412 43447 5468
rect 43447 5412 43503 5468
rect 43503 5412 43507 5468
rect 43443 5408 43507 5412
rect 43523 5468 43587 5472
rect 43523 5412 43527 5468
rect 43527 5412 43583 5468
rect 43583 5412 43587 5468
rect 43523 5408 43587 5412
rect 43603 5468 43667 5472
rect 43603 5412 43607 5468
rect 43607 5412 43663 5468
rect 43663 5412 43667 5468
rect 43603 5408 43667 5412
rect 36492 5068 36556 5132
rect 6253 4924 6317 4928
rect 6253 4868 6257 4924
rect 6257 4868 6313 4924
rect 6313 4868 6317 4924
rect 6253 4864 6317 4868
rect 6333 4924 6397 4928
rect 6333 4868 6337 4924
rect 6337 4868 6393 4924
rect 6393 4868 6397 4924
rect 6333 4864 6397 4868
rect 6413 4924 6477 4928
rect 6413 4868 6417 4924
rect 6417 4868 6473 4924
rect 6473 4868 6477 4924
rect 6413 4864 6477 4868
rect 6493 4924 6557 4928
rect 6493 4868 6497 4924
rect 6497 4868 6553 4924
rect 6553 4868 6557 4924
rect 6493 4864 6557 4868
rect 16856 4924 16920 4928
rect 16856 4868 16860 4924
rect 16860 4868 16916 4924
rect 16916 4868 16920 4924
rect 16856 4864 16920 4868
rect 16936 4924 17000 4928
rect 16936 4868 16940 4924
rect 16940 4868 16996 4924
rect 16996 4868 17000 4924
rect 16936 4864 17000 4868
rect 17016 4924 17080 4928
rect 17016 4868 17020 4924
rect 17020 4868 17076 4924
rect 17076 4868 17080 4924
rect 17016 4864 17080 4868
rect 17096 4924 17160 4928
rect 17096 4868 17100 4924
rect 17100 4868 17156 4924
rect 17156 4868 17160 4924
rect 17096 4864 17160 4868
rect 27459 4924 27523 4928
rect 27459 4868 27463 4924
rect 27463 4868 27519 4924
rect 27519 4868 27523 4924
rect 27459 4864 27523 4868
rect 27539 4924 27603 4928
rect 27539 4868 27543 4924
rect 27543 4868 27599 4924
rect 27599 4868 27603 4924
rect 27539 4864 27603 4868
rect 27619 4924 27683 4928
rect 27619 4868 27623 4924
rect 27623 4868 27679 4924
rect 27679 4868 27683 4924
rect 27619 4864 27683 4868
rect 27699 4924 27763 4928
rect 27699 4868 27703 4924
rect 27703 4868 27759 4924
rect 27759 4868 27763 4924
rect 27699 4864 27763 4868
rect 38062 4924 38126 4928
rect 38062 4868 38066 4924
rect 38066 4868 38122 4924
rect 38122 4868 38126 4924
rect 38062 4864 38126 4868
rect 38142 4924 38206 4928
rect 38142 4868 38146 4924
rect 38146 4868 38202 4924
rect 38202 4868 38206 4924
rect 38142 4864 38206 4868
rect 38222 4924 38286 4928
rect 38222 4868 38226 4924
rect 38226 4868 38282 4924
rect 38282 4868 38286 4924
rect 38222 4864 38286 4868
rect 38302 4924 38366 4928
rect 38302 4868 38306 4924
rect 38306 4868 38362 4924
rect 38362 4868 38366 4924
rect 38302 4864 38366 4868
rect 11554 4380 11618 4384
rect 11554 4324 11558 4380
rect 11558 4324 11614 4380
rect 11614 4324 11618 4380
rect 11554 4320 11618 4324
rect 11634 4380 11698 4384
rect 11634 4324 11638 4380
rect 11638 4324 11694 4380
rect 11694 4324 11698 4380
rect 11634 4320 11698 4324
rect 11714 4380 11778 4384
rect 11714 4324 11718 4380
rect 11718 4324 11774 4380
rect 11774 4324 11778 4380
rect 11714 4320 11778 4324
rect 11794 4380 11858 4384
rect 11794 4324 11798 4380
rect 11798 4324 11854 4380
rect 11854 4324 11858 4380
rect 11794 4320 11858 4324
rect 22157 4380 22221 4384
rect 22157 4324 22161 4380
rect 22161 4324 22217 4380
rect 22217 4324 22221 4380
rect 22157 4320 22221 4324
rect 22237 4380 22301 4384
rect 22237 4324 22241 4380
rect 22241 4324 22297 4380
rect 22297 4324 22301 4380
rect 22237 4320 22301 4324
rect 22317 4380 22381 4384
rect 22317 4324 22321 4380
rect 22321 4324 22377 4380
rect 22377 4324 22381 4380
rect 22317 4320 22381 4324
rect 22397 4380 22461 4384
rect 22397 4324 22401 4380
rect 22401 4324 22457 4380
rect 22457 4324 22461 4380
rect 22397 4320 22461 4324
rect 32760 4380 32824 4384
rect 32760 4324 32764 4380
rect 32764 4324 32820 4380
rect 32820 4324 32824 4380
rect 32760 4320 32824 4324
rect 32840 4380 32904 4384
rect 32840 4324 32844 4380
rect 32844 4324 32900 4380
rect 32900 4324 32904 4380
rect 32840 4320 32904 4324
rect 32920 4380 32984 4384
rect 32920 4324 32924 4380
rect 32924 4324 32980 4380
rect 32980 4324 32984 4380
rect 32920 4320 32984 4324
rect 33000 4380 33064 4384
rect 33000 4324 33004 4380
rect 33004 4324 33060 4380
rect 33060 4324 33064 4380
rect 33000 4320 33064 4324
rect 43363 4380 43427 4384
rect 43363 4324 43367 4380
rect 43367 4324 43423 4380
rect 43423 4324 43427 4380
rect 43363 4320 43427 4324
rect 43443 4380 43507 4384
rect 43443 4324 43447 4380
rect 43447 4324 43503 4380
rect 43503 4324 43507 4380
rect 43443 4320 43507 4324
rect 43523 4380 43587 4384
rect 43523 4324 43527 4380
rect 43527 4324 43583 4380
rect 43583 4324 43587 4380
rect 43523 4320 43587 4324
rect 43603 4380 43667 4384
rect 43603 4324 43607 4380
rect 43607 4324 43663 4380
rect 43663 4324 43667 4380
rect 43603 4320 43667 4324
rect 6253 3836 6317 3840
rect 6253 3780 6257 3836
rect 6257 3780 6313 3836
rect 6313 3780 6317 3836
rect 6253 3776 6317 3780
rect 6333 3836 6397 3840
rect 6333 3780 6337 3836
rect 6337 3780 6393 3836
rect 6393 3780 6397 3836
rect 6333 3776 6397 3780
rect 6413 3836 6477 3840
rect 6413 3780 6417 3836
rect 6417 3780 6473 3836
rect 6473 3780 6477 3836
rect 6413 3776 6477 3780
rect 6493 3836 6557 3840
rect 6493 3780 6497 3836
rect 6497 3780 6553 3836
rect 6553 3780 6557 3836
rect 6493 3776 6557 3780
rect 16856 3836 16920 3840
rect 16856 3780 16860 3836
rect 16860 3780 16916 3836
rect 16916 3780 16920 3836
rect 16856 3776 16920 3780
rect 16936 3836 17000 3840
rect 16936 3780 16940 3836
rect 16940 3780 16996 3836
rect 16996 3780 17000 3836
rect 16936 3776 17000 3780
rect 17016 3836 17080 3840
rect 17016 3780 17020 3836
rect 17020 3780 17076 3836
rect 17076 3780 17080 3836
rect 17016 3776 17080 3780
rect 17096 3836 17160 3840
rect 17096 3780 17100 3836
rect 17100 3780 17156 3836
rect 17156 3780 17160 3836
rect 17096 3776 17160 3780
rect 27459 3836 27523 3840
rect 27459 3780 27463 3836
rect 27463 3780 27519 3836
rect 27519 3780 27523 3836
rect 27459 3776 27523 3780
rect 27539 3836 27603 3840
rect 27539 3780 27543 3836
rect 27543 3780 27599 3836
rect 27599 3780 27603 3836
rect 27539 3776 27603 3780
rect 27619 3836 27683 3840
rect 27619 3780 27623 3836
rect 27623 3780 27679 3836
rect 27679 3780 27683 3836
rect 27619 3776 27683 3780
rect 27699 3836 27763 3840
rect 27699 3780 27703 3836
rect 27703 3780 27759 3836
rect 27759 3780 27763 3836
rect 27699 3776 27763 3780
rect 38062 3836 38126 3840
rect 38062 3780 38066 3836
rect 38066 3780 38122 3836
rect 38122 3780 38126 3836
rect 38062 3776 38126 3780
rect 38142 3836 38206 3840
rect 38142 3780 38146 3836
rect 38146 3780 38202 3836
rect 38202 3780 38206 3836
rect 38142 3776 38206 3780
rect 38222 3836 38286 3840
rect 38222 3780 38226 3836
rect 38226 3780 38282 3836
rect 38282 3780 38286 3836
rect 38222 3776 38286 3780
rect 38302 3836 38366 3840
rect 38302 3780 38306 3836
rect 38306 3780 38362 3836
rect 38362 3780 38366 3836
rect 38302 3776 38366 3780
rect 11554 3292 11618 3296
rect 11554 3236 11558 3292
rect 11558 3236 11614 3292
rect 11614 3236 11618 3292
rect 11554 3232 11618 3236
rect 11634 3292 11698 3296
rect 11634 3236 11638 3292
rect 11638 3236 11694 3292
rect 11694 3236 11698 3292
rect 11634 3232 11698 3236
rect 11714 3292 11778 3296
rect 11714 3236 11718 3292
rect 11718 3236 11774 3292
rect 11774 3236 11778 3292
rect 11714 3232 11778 3236
rect 11794 3292 11858 3296
rect 11794 3236 11798 3292
rect 11798 3236 11854 3292
rect 11854 3236 11858 3292
rect 11794 3232 11858 3236
rect 22157 3292 22221 3296
rect 22157 3236 22161 3292
rect 22161 3236 22217 3292
rect 22217 3236 22221 3292
rect 22157 3232 22221 3236
rect 22237 3292 22301 3296
rect 22237 3236 22241 3292
rect 22241 3236 22297 3292
rect 22297 3236 22301 3292
rect 22237 3232 22301 3236
rect 22317 3292 22381 3296
rect 22317 3236 22321 3292
rect 22321 3236 22377 3292
rect 22377 3236 22381 3292
rect 22317 3232 22381 3236
rect 22397 3292 22461 3296
rect 22397 3236 22401 3292
rect 22401 3236 22457 3292
rect 22457 3236 22461 3292
rect 22397 3232 22461 3236
rect 32760 3292 32824 3296
rect 32760 3236 32764 3292
rect 32764 3236 32820 3292
rect 32820 3236 32824 3292
rect 32760 3232 32824 3236
rect 32840 3292 32904 3296
rect 32840 3236 32844 3292
rect 32844 3236 32900 3292
rect 32900 3236 32904 3292
rect 32840 3232 32904 3236
rect 32920 3292 32984 3296
rect 32920 3236 32924 3292
rect 32924 3236 32980 3292
rect 32980 3236 32984 3292
rect 32920 3232 32984 3236
rect 33000 3292 33064 3296
rect 33000 3236 33004 3292
rect 33004 3236 33060 3292
rect 33060 3236 33064 3292
rect 33000 3232 33064 3236
rect 43363 3292 43427 3296
rect 43363 3236 43367 3292
rect 43367 3236 43423 3292
rect 43423 3236 43427 3292
rect 43363 3232 43427 3236
rect 43443 3292 43507 3296
rect 43443 3236 43447 3292
rect 43447 3236 43503 3292
rect 43503 3236 43507 3292
rect 43443 3232 43507 3236
rect 43523 3292 43587 3296
rect 43523 3236 43527 3292
rect 43527 3236 43583 3292
rect 43583 3236 43587 3292
rect 43523 3232 43587 3236
rect 43603 3292 43667 3296
rect 43603 3236 43607 3292
rect 43607 3236 43663 3292
rect 43663 3236 43667 3292
rect 43603 3232 43667 3236
rect 30420 2756 30484 2820
rect 6253 2748 6317 2752
rect 6253 2692 6257 2748
rect 6257 2692 6313 2748
rect 6313 2692 6317 2748
rect 6253 2688 6317 2692
rect 6333 2748 6397 2752
rect 6333 2692 6337 2748
rect 6337 2692 6393 2748
rect 6393 2692 6397 2748
rect 6333 2688 6397 2692
rect 6413 2748 6477 2752
rect 6413 2692 6417 2748
rect 6417 2692 6473 2748
rect 6473 2692 6477 2748
rect 6413 2688 6477 2692
rect 6493 2748 6557 2752
rect 6493 2692 6497 2748
rect 6497 2692 6553 2748
rect 6553 2692 6557 2748
rect 6493 2688 6557 2692
rect 16856 2748 16920 2752
rect 16856 2692 16860 2748
rect 16860 2692 16916 2748
rect 16916 2692 16920 2748
rect 16856 2688 16920 2692
rect 16936 2748 17000 2752
rect 16936 2692 16940 2748
rect 16940 2692 16996 2748
rect 16996 2692 17000 2748
rect 16936 2688 17000 2692
rect 17016 2748 17080 2752
rect 17016 2692 17020 2748
rect 17020 2692 17076 2748
rect 17076 2692 17080 2748
rect 17016 2688 17080 2692
rect 17096 2748 17160 2752
rect 17096 2692 17100 2748
rect 17100 2692 17156 2748
rect 17156 2692 17160 2748
rect 17096 2688 17160 2692
rect 27459 2748 27523 2752
rect 27459 2692 27463 2748
rect 27463 2692 27519 2748
rect 27519 2692 27523 2748
rect 27459 2688 27523 2692
rect 27539 2748 27603 2752
rect 27539 2692 27543 2748
rect 27543 2692 27599 2748
rect 27599 2692 27603 2748
rect 27539 2688 27603 2692
rect 27619 2748 27683 2752
rect 27619 2692 27623 2748
rect 27623 2692 27679 2748
rect 27679 2692 27683 2748
rect 27619 2688 27683 2692
rect 27699 2748 27763 2752
rect 27699 2692 27703 2748
rect 27703 2692 27759 2748
rect 27759 2692 27763 2748
rect 27699 2688 27763 2692
rect 38062 2748 38126 2752
rect 38062 2692 38066 2748
rect 38066 2692 38122 2748
rect 38122 2692 38126 2748
rect 38062 2688 38126 2692
rect 38142 2748 38206 2752
rect 38142 2692 38146 2748
rect 38146 2692 38202 2748
rect 38202 2692 38206 2748
rect 38142 2688 38206 2692
rect 38222 2748 38286 2752
rect 38222 2692 38226 2748
rect 38226 2692 38282 2748
rect 38282 2692 38286 2748
rect 38222 2688 38286 2692
rect 38302 2748 38366 2752
rect 38302 2692 38306 2748
rect 38306 2692 38362 2748
rect 38362 2692 38366 2748
rect 38302 2688 38366 2692
rect 36492 2620 36556 2684
rect 11554 2204 11618 2208
rect 11554 2148 11558 2204
rect 11558 2148 11614 2204
rect 11614 2148 11618 2204
rect 11554 2144 11618 2148
rect 11634 2204 11698 2208
rect 11634 2148 11638 2204
rect 11638 2148 11694 2204
rect 11694 2148 11698 2204
rect 11634 2144 11698 2148
rect 11714 2204 11778 2208
rect 11714 2148 11718 2204
rect 11718 2148 11774 2204
rect 11774 2148 11778 2204
rect 11714 2144 11778 2148
rect 11794 2204 11858 2208
rect 11794 2148 11798 2204
rect 11798 2148 11854 2204
rect 11854 2148 11858 2204
rect 11794 2144 11858 2148
rect 22157 2204 22221 2208
rect 22157 2148 22161 2204
rect 22161 2148 22217 2204
rect 22217 2148 22221 2204
rect 22157 2144 22221 2148
rect 22237 2204 22301 2208
rect 22237 2148 22241 2204
rect 22241 2148 22297 2204
rect 22297 2148 22301 2204
rect 22237 2144 22301 2148
rect 22317 2204 22381 2208
rect 22317 2148 22321 2204
rect 22321 2148 22377 2204
rect 22377 2148 22381 2204
rect 22317 2144 22381 2148
rect 22397 2204 22461 2208
rect 22397 2148 22401 2204
rect 22401 2148 22457 2204
rect 22457 2148 22461 2204
rect 22397 2144 22461 2148
rect 32760 2204 32824 2208
rect 32760 2148 32764 2204
rect 32764 2148 32820 2204
rect 32820 2148 32824 2204
rect 32760 2144 32824 2148
rect 32840 2204 32904 2208
rect 32840 2148 32844 2204
rect 32844 2148 32900 2204
rect 32900 2148 32904 2204
rect 32840 2144 32904 2148
rect 32920 2204 32984 2208
rect 32920 2148 32924 2204
rect 32924 2148 32980 2204
rect 32980 2148 32984 2204
rect 32920 2144 32984 2148
rect 33000 2204 33064 2208
rect 33000 2148 33004 2204
rect 33004 2148 33060 2204
rect 33060 2148 33064 2204
rect 33000 2144 33064 2148
rect 43363 2204 43427 2208
rect 43363 2148 43367 2204
rect 43367 2148 43423 2204
rect 43423 2148 43427 2204
rect 43363 2144 43427 2148
rect 43443 2204 43507 2208
rect 43443 2148 43447 2204
rect 43447 2148 43503 2204
rect 43503 2148 43507 2204
rect 43443 2144 43507 2148
rect 43523 2204 43587 2208
rect 43523 2148 43527 2204
rect 43527 2148 43583 2204
rect 43583 2148 43587 2204
rect 43523 2144 43587 2148
rect 43603 2204 43667 2208
rect 43603 2148 43607 2204
rect 43607 2148 43663 2204
rect 43663 2148 43667 2204
rect 43603 2144 43667 2148
rect 30420 1124 30484 1188
<< metal4 >>
rect 6245 7104 6565 7664
rect 6245 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6565 7104
rect 6245 6016 6565 7040
rect 6245 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6565 6016
rect 6245 4928 6565 5952
rect 6245 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6565 4928
rect 6245 3840 6565 4864
rect 6245 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6565 3840
rect 6245 2752 6565 3776
rect 6245 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6565 2752
rect 6245 2128 6565 2688
rect 11546 7648 11866 7664
rect 11546 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11866 7648
rect 11546 6560 11866 7584
rect 11546 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11866 6560
rect 11546 5472 11866 6496
rect 11546 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11866 5472
rect 11546 4384 11866 5408
rect 11546 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11866 4384
rect 11546 3296 11866 4320
rect 11546 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11866 3296
rect 11546 2208 11866 3232
rect 11546 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11866 2208
rect 11546 2128 11866 2144
rect 16848 7104 17168 7664
rect 16848 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17168 7104
rect 16848 6016 17168 7040
rect 16848 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17168 6016
rect 16848 4928 17168 5952
rect 16848 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17168 4928
rect 16848 3840 17168 4864
rect 16848 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17168 3840
rect 16848 2752 17168 3776
rect 16848 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17168 2752
rect 16848 2128 17168 2688
rect 22149 7648 22469 7664
rect 22149 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22469 7648
rect 22149 6560 22469 7584
rect 22149 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22469 6560
rect 22149 5472 22469 6496
rect 22149 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22469 5472
rect 22149 4384 22469 5408
rect 22149 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22469 4384
rect 22149 3296 22469 4320
rect 22149 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22469 3296
rect 22149 2208 22469 3232
rect 22149 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22469 2208
rect 22149 2128 22469 2144
rect 27451 7104 27771 7664
rect 27451 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27771 7104
rect 27451 6016 27771 7040
rect 27451 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27771 6016
rect 27451 4928 27771 5952
rect 27451 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27771 4928
rect 27451 3840 27771 4864
rect 27451 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27771 3840
rect 27451 2752 27771 3776
rect 32752 7648 33072 7664
rect 32752 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33072 7648
rect 32752 6560 33072 7584
rect 32752 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33072 6560
rect 32752 5472 33072 6496
rect 32752 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33072 5472
rect 32752 4384 33072 5408
rect 38054 7104 38374 7664
rect 38054 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38374 7104
rect 38054 6016 38374 7040
rect 38054 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38374 6016
rect 36491 5132 36557 5133
rect 36491 5068 36492 5132
rect 36556 5068 36557 5132
rect 36491 5067 36557 5068
rect 32752 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33072 4384
rect 32752 3296 33072 4320
rect 32752 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33072 3296
rect 30419 2820 30485 2821
rect 30419 2756 30420 2820
rect 30484 2756 30485 2820
rect 30419 2755 30485 2756
rect 27451 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27771 2752
rect 27451 2128 27771 2688
rect 30422 1189 30482 2755
rect 32752 2208 33072 3232
rect 36494 2685 36554 5067
rect 38054 4928 38374 5952
rect 38054 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38374 4928
rect 38054 3840 38374 4864
rect 38054 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38374 3840
rect 38054 2752 38374 3776
rect 38054 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38374 2752
rect 36491 2684 36557 2685
rect 36491 2620 36492 2684
rect 36556 2620 36557 2684
rect 36491 2619 36557 2620
rect 32752 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33072 2208
rect 32752 2128 33072 2144
rect 38054 2128 38374 2688
rect 43355 7648 43675 7664
rect 43355 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43675 7648
rect 43355 6560 43675 7584
rect 43355 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43675 6560
rect 43355 5472 43675 6496
rect 43355 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43675 5472
rect 43355 4384 43675 5408
rect 43355 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43675 4384
rect 43355 3296 43675 4320
rect 43355 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43675 3296
rect 43355 2208 43675 3232
rect 43355 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43675 2208
rect 43355 2128 43675 2144
rect 30419 1188 30485 1189
rect 30419 1124 30420 1188
rect 30484 1124 30485 1188
rect 30419 1123 30485 1124
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 24748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 37812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 23368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform 1 0 25392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 25668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 25944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _49_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _50_
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _51_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _52_
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _53_
timestamp 1688980957
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _54_
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _55_
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _56_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _57_
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _58_
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _59_
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _60_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _61_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _62_
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _63_
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _64_
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _65_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _66_
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _67_
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _68_
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _69_
timestamp 1688980957
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _70_
timestamp 1688980957
transform 1 0 35236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_452 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42688 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_86
timestamp 1688980957
transform 1 0 9016 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_98
timestamp 1688980957
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_140
timestamp 1688980957
transform 1 0 13984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1688980957
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_387
timestamp 1688980957
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_397
timestamp 1688980957
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_404 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38272 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_412
timestamp 1688980957
transform 1 0 39008 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_416
timestamp 1688980957
transform 1 0 39376 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_428
timestamp 1688980957
transform 1 0 40480 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_440
timestamp 1688980957
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_200
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_207
timestamp 1688980957
transform 1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_237
timestamp 1688980957
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_259
timestamp 1688980957
transform 1 0 24932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_285
timestamp 1688980957
transform 1 0 27324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_341
timestamp 1688980957
transform 1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_354
timestamp 1688980957
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1688980957
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_457
timestamp 1688980957
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_157
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_162
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_457
timestamp 1688980957
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_260
timestamp 1688980957
transform 1 0 25024 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_272
timestamp 1688980957
transform 1 0 26128 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_284
timestamp 1688980957
transform 1 0 27232 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_296
timestamp 1688980957
transform 1 0 28336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_236
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_76
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_122
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_134
timestamp 1688980957
transform 1 0 13432 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_147
timestamp 1688980957
transform 1 0 14628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_194
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_197
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_240
timestamp 1688980957
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_260
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_272
timestamp 1688980957
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_298
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_306
timestamp 1688980957
transform 1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_309
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_321
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_345
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_352
timestamp 1688980957
transform 1 0 33488 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_365
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_375
timestamp 1688980957
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_387
timestamp 1688980957
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_402
timestamp 1688980957
transform 1 0 38088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_414
timestamp 1688980957
transform 1 0 39192 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_427
timestamp 1688980957
transform 1 0 40388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_435
timestamp 1688980957
transform 1 0 41124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_444
timestamp 1688980957
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 35972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 37996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 35880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 36800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 28704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 30820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 32936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 35052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 41400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 42688 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 11776 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 22356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 22816 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 23368 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 23920 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 24472 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 21712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 22264 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 22264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 25024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 28612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 25576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 26128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 32752 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 33764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 32660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 34058 -300 34114 160 0 FreeSans 224 90 0 0 Ci
port 0 nsew signal input
flabel metal2 s 34334 -300 34390 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 37094 -300 37150 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 37370 -300 37426 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 37646 -300 37702 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 37922 -300 37978 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 38198 -300 38254 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 38474 -300 38530 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 38750 -300 38806 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 39026 -300 39082 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 39302 -300 39358 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 39578 -300 39634 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 34610 -300 34666 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 34886 -300 34942 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 35162 -300 35218 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 35438 -300 35494 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 35714 -300 35770 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 35990 -300 36046 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 36266 -300 36322 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 36542 -300 36598 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 36818 -300 36874 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 3238 9840 3294 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 24398 9840 24454 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 26514 9840 26570 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 28630 9840 28686 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 30746 9840 30802 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 32862 9840 32918 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 34978 9840 35034 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 37094 9840 37150 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 39210 9840 39266 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 41326 9840 41382 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 43442 9840 43498 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 5354 9840 5410 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 7470 9840 7526 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 9586 9840 9642 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 11702 9840 11758 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 13818 9840 13874 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 15934 9840 15990 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 18050 9840 18106 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 20166 9840 20222 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 22282 9840 22338 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5078 -300 5134 160 0 FreeSans 224 90 0 0 N1END[0]
port 41 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 N1END[1]
port 42 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 N1END[2]
port 43 nsew signal input
flabel metal2 s 5906 -300 5962 160 0 FreeSans 224 90 0 0 N1END[3]
port 44 nsew signal input
flabel metal2 s 8390 -300 8446 160 0 FreeSans 224 90 0 0 N2END[0]
port 45 nsew signal input
flabel metal2 s 8666 -300 8722 160 0 FreeSans 224 90 0 0 N2END[1]
port 46 nsew signal input
flabel metal2 s 8942 -300 8998 160 0 FreeSans 224 90 0 0 N2END[2]
port 47 nsew signal input
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 N2END[3]
port 48 nsew signal input
flabel metal2 s 9494 -300 9550 160 0 FreeSans 224 90 0 0 N2END[4]
port 49 nsew signal input
flabel metal2 s 9770 -300 9826 160 0 FreeSans 224 90 0 0 N2END[5]
port 50 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 N2END[6]
port 51 nsew signal input
flabel metal2 s 10322 -300 10378 160 0 FreeSans 224 90 0 0 N2END[7]
port 52 nsew signal input
flabel metal2 s 6182 -300 6238 160 0 FreeSans 224 90 0 0 N2MID[0]
port 53 nsew signal input
flabel metal2 s 6458 -300 6514 160 0 FreeSans 224 90 0 0 N2MID[1]
port 54 nsew signal input
flabel metal2 s 6734 -300 6790 160 0 FreeSans 224 90 0 0 N2MID[2]
port 55 nsew signal input
flabel metal2 s 7010 -300 7066 160 0 FreeSans 224 90 0 0 N2MID[3]
port 56 nsew signal input
flabel metal2 s 7286 -300 7342 160 0 FreeSans 224 90 0 0 N2MID[4]
port 57 nsew signal input
flabel metal2 s 7562 -300 7618 160 0 FreeSans 224 90 0 0 N2MID[5]
port 58 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 N2MID[6]
port 59 nsew signal input
flabel metal2 s 8114 -300 8170 160 0 FreeSans 224 90 0 0 N2MID[7]
port 60 nsew signal input
flabel metal2 s 10598 -300 10654 160 0 FreeSans 224 90 0 0 N4END[0]
port 61 nsew signal input
flabel metal2 s 13358 -300 13414 160 0 FreeSans 224 90 0 0 N4END[10]
port 62 nsew signal input
flabel metal2 s 13634 -300 13690 160 0 FreeSans 224 90 0 0 N4END[11]
port 63 nsew signal input
flabel metal2 s 13910 -300 13966 160 0 FreeSans 224 90 0 0 N4END[12]
port 64 nsew signal input
flabel metal2 s 14186 -300 14242 160 0 FreeSans 224 90 0 0 N4END[13]
port 65 nsew signal input
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 N4END[14]
port 66 nsew signal input
flabel metal2 s 14738 -300 14794 160 0 FreeSans 224 90 0 0 N4END[15]
port 67 nsew signal input
flabel metal2 s 10874 -300 10930 160 0 FreeSans 224 90 0 0 N4END[1]
port 68 nsew signal input
flabel metal2 s 11150 -300 11206 160 0 FreeSans 224 90 0 0 N4END[2]
port 69 nsew signal input
flabel metal2 s 11426 -300 11482 160 0 FreeSans 224 90 0 0 N4END[3]
port 70 nsew signal input
flabel metal2 s 11702 -300 11758 160 0 FreeSans 224 90 0 0 N4END[4]
port 71 nsew signal input
flabel metal2 s 11978 -300 12034 160 0 FreeSans 224 90 0 0 N4END[5]
port 72 nsew signal input
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 N4END[6]
port 73 nsew signal input
flabel metal2 s 12530 -300 12586 160 0 FreeSans 224 90 0 0 N4END[7]
port 74 nsew signal input
flabel metal2 s 12806 -300 12862 160 0 FreeSans 224 90 0 0 N4END[8]
port 75 nsew signal input
flabel metal2 s 13082 -300 13138 160 0 FreeSans 224 90 0 0 N4END[9]
port 76 nsew signal input
flabel metal2 s 15014 -300 15070 160 0 FreeSans 224 90 0 0 NN4END[0]
port 77 nsew signal input
flabel metal2 s 17774 -300 17830 160 0 FreeSans 224 90 0 0 NN4END[10]
port 78 nsew signal input
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 NN4END[11]
port 79 nsew signal input
flabel metal2 s 18326 -300 18382 160 0 FreeSans 224 90 0 0 NN4END[12]
port 80 nsew signal input
flabel metal2 s 18602 -300 18658 160 0 FreeSans 224 90 0 0 NN4END[13]
port 81 nsew signal input
flabel metal2 s 18878 -300 18934 160 0 FreeSans 224 90 0 0 NN4END[14]
port 82 nsew signal input
flabel metal2 s 19154 -300 19210 160 0 FreeSans 224 90 0 0 NN4END[15]
port 83 nsew signal input
flabel metal2 s 15290 -300 15346 160 0 FreeSans 224 90 0 0 NN4END[1]
port 84 nsew signal input
flabel metal2 s 15566 -300 15622 160 0 FreeSans 224 90 0 0 NN4END[2]
port 85 nsew signal input
flabel metal2 s 15842 -300 15898 160 0 FreeSans 224 90 0 0 NN4END[3]
port 86 nsew signal input
flabel metal2 s 16118 -300 16174 160 0 FreeSans 224 90 0 0 NN4END[4]
port 87 nsew signal input
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 NN4END[5]
port 88 nsew signal input
flabel metal2 s 16670 -300 16726 160 0 FreeSans 224 90 0 0 NN4END[6]
port 89 nsew signal input
flabel metal2 s 16946 -300 17002 160 0 FreeSans 224 90 0 0 NN4END[7]
port 90 nsew signal input
flabel metal2 s 17222 -300 17278 160 0 FreeSans 224 90 0 0 NN4END[8]
port 91 nsew signal input
flabel metal2 s 17498 -300 17554 160 0 FreeSans 224 90 0 0 NN4END[9]
port 92 nsew signal input
flabel metal2 s 19430 -300 19486 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 93 nsew signal tristate
flabel metal2 s 19706 -300 19762 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 94 nsew signal tristate
flabel metal2 s 19982 -300 20038 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 95 nsew signal tristate
flabel metal2 s 20258 -300 20314 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 96 nsew signal tristate
flabel metal2 s 22742 -300 22798 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 97 nsew signal tristate
flabel metal2 s 23018 -300 23074 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 98 nsew signal tristate
flabel metal2 s 23294 -300 23350 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 99 nsew signal tristate
flabel metal2 s 23570 -300 23626 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 100 nsew signal tristate
flabel metal2 s 23846 -300 23902 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 101 nsew signal tristate
flabel metal2 s 24122 -300 24178 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 102 nsew signal tristate
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 103 nsew signal tristate
flabel metal2 s 24674 -300 24730 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 104 nsew signal tristate
flabel metal2 s 20534 -300 20590 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 105 nsew signal tristate
flabel metal2 s 20810 -300 20866 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 106 nsew signal tristate
flabel metal2 s 21086 -300 21142 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 107 nsew signal tristate
flabel metal2 s 21362 -300 21418 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 108 nsew signal tristate
flabel metal2 s 21638 -300 21694 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 109 nsew signal tristate
flabel metal2 s 21914 -300 21970 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 110 nsew signal tristate
flabel metal2 s 22190 -300 22246 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 111 nsew signal tristate
flabel metal2 s 22466 -300 22522 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 112 nsew signal tristate
flabel metal2 s 24950 -300 25006 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 113 nsew signal tristate
flabel metal2 s 27710 -300 27766 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 114 nsew signal tristate
flabel metal2 s 27986 -300 28042 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 115 nsew signal tristate
flabel metal2 s 28262 -300 28318 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 116 nsew signal tristate
flabel metal2 s 28538 -300 28594 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 117 nsew signal tristate
flabel metal2 s 28814 -300 28870 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 118 nsew signal tristate
flabel metal2 s 29090 -300 29146 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 119 nsew signal tristate
flabel metal2 s 25226 -300 25282 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 120 nsew signal tristate
flabel metal2 s 25502 -300 25558 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 121 nsew signal tristate
flabel metal2 s 25778 -300 25834 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 122 nsew signal tristate
flabel metal2 s 26054 -300 26110 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 123 nsew signal tristate
flabel metal2 s 26330 -300 26386 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 124 nsew signal tristate
flabel metal2 s 26606 -300 26662 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 125 nsew signal tristate
flabel metal2 s 26882 -300 26938 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 126 nsew signal tristate
flabel metal2 s 27158 -300 27214 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 127 nsew signal tristate
flabel metal2 s 27434 -300 27490 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 128 nsew signal tristate
flabel metal2 s 29366 -300 29422 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 129 nsew signal tristate
flabel metal2 s 32126 -300 32182 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 130 nsew signal tristate
flabel metal2 s 32402 -300 32458 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 131 nsew signal tristate
flabel metal2 s 32678 -300 32734 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 132 nsew signal tristate
flabel metal2 s 32954 -300 33010 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 133 nsew signal tristate
flabel metal2 s 33230 -300 33286 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 134 nsew signal tristate
flabel metal2 s 33506 -300 33562 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 135 nsew signal tristate
flabel metal2 s 29642 -300 29698 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 136 nsew signal tristate
flabel metal2 s 29918 -300 29974 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 137 nsew signal tristate
flabel metal2 s 30194 -300 30250 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 138 nsew signal tristate
flabel metal2 s 30470 -300 30526 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 139 nsew signal tristate
flabel metal2 s 30746 -300 30802 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 140 nsew signal tristate
flabel metal2 s 31022 -300 31078 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 141 nsew signal tristate
flabel metal2 s 31298 -300 31354 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 142 nsew signal tristate
flabel metal2 s 31574 -300 31630 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 143 nsew signal tristate
flabel metal2 s 31850 -300 31906 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 144 nsew signal tristate
flabel metal2 s 33782 -300 33838 160 0 FreeSans 224 90 0 0 UserCLK
port 145 nsew signal input
flabel metal2 s 1122 9840 1178 10300 0 FreeSans 224 90 0 0 UserCLKo
port 146 nsew signal tristate
flabel metal4 s 6245 2128 6565 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 16848 2128 17168 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 27451 2128 27771 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 38054 2128 38374 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 11546 2128 11866 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 22149 2128 22469 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 32752 2128 33072 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 43355 2128 43675 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
rlabel metal1 22310 7072 22310 7072 0 vccd1
rlabel via1 22389 7616 22389 7616 0 vssd1
rlabel metal2 34415 68 34415 68 0 FrameStrobe[0]
rlabel metal2 37122 1231 37122 1231 0 FrameStrobe[10]
rlabel metal2 37398 1316 37398 1316 0 FrameStrobe[11]
rlabel metal1 37812 3026 37812 3026 0 FrameStrobe[12]
rlabel metal2 37996 3060 37996 3060 0 FrameStrobe[13]
rlabel metal2 38325 68 38325 68 0 FrameStrobe[14]
rlabel metal2 38555 68 38555 68 0 FrameStrobe[15]
rlabel metal2 38778 806 38778 806 0 FrameStrobe[16]
rlabel metal1 39192 3026 39192 3026 0 FrameStrobe[17]
rlabel metal2 39330 738 39330 738 0 FrameStrobe[18]
rlabel metal2 39751 68 39751 68 0 FrameStrobe[19]
rlabel metal1 36340 2414 36340 2414 0 FrameStrobe[1]
rlabel metal1 35282 2958 35282 2958 0 FrameStrobe[2]
rlabel metal2 35289 68 35289 68 0 FrameStrobe[3]
rlabel metal2 35565 68 35565 68 0 FrameStrobe[4]
rlabel metal1 35972 2958 35972 2958 0 FrameStrobe[5]
rlabel metal2 36018 687 36018 687 0 FrameStrobe[6]
rlabel metal2 36393 68 36393 68 0 FrameStrobe[7]
rlabel metal2 36623 68 36623 68 0 FrameStrobe[8]
rlabel metal2 36846 687 36846 687 0 FrameStrobe[9]
rlabel metal2 3266 9717 3266 9717 0 FrameStrobe_O[0]
rlabel metal2 24426 9785 24426 9785 0 FrameStrobe_O[10]
rlabel metal2 26542 8680 26542 8680 0 FrameStrobe_O[11]
rlabel metal2 28658 9173 28658 9173 0 FrameStrobe_O[12]
rlabel metal2 30774 8680 30774 8680 0 FrameStrobe_O[13]
rlabel metal2 32890 9037 32890 9037 0 FrameStrobe_O[14]
rlabel metal2 35006 8680 35006 8680 0 FrameStrobe_O[15]
rlabel metal2 37122 8680 37122 8680 0 FrameStrobe_O[16]
rlabel metal2 39238 8680 39238 8680 0 FrameStrobe_O[17]
rlabel metal2 41446 7463 41446 7463 0 FrameStrobe_O[18]
rlabel metal1 43194 7514 43194 7514 0 FrameStrobe_O[19]
rlabel metal2 5382 8680 5382 8680 0 FrameStrobe_O[1]
rlabel metal2 7498 8680 7498 8680 0 FrameStrobe_O[2]
rlabel metal2 9614 8629 9614 8629 0 FrameStrobe_O[3]
rlabel metal2 11730 9785 11730 9785 0 FrameStrobe_O[4]
rlabel metal2 13846 8680 13846 8680 0 FrameStrobe_O[5]
rlabel metal2 15962 8680 15962 8680 0 FrameStrobe_O[6]
rlabel metal2 18078 8680 18078 8680 0 FrameStrobe_O[7]
rlabel metal2 20194 9785 20194 9785 0 FrameStrobe_O[8]
rlabel metal2 22310 9785 22310 9785 0 FrameStrobe_O[9]
rlabel metal2 5007 68 5007 68 0 N1END[0]
rlabel metal2 5283 68 5283 68 0 N1END[1]
rlabel metal2 5658 1248 5658 1248 0 N1END[2]
rlabel metal2 5835 68 5835 68 0 N1END[3]
rlabel metal2 8418 1214 8418 1214 0 N2END[0]
rlabel metal2 8595 68 8595 68 0 N2END[1]
rlabel metal2 8970 687 8970 687 0 N2END[2]
rlabel metal2 9246 1248 9246 1248 0 N2END[3]
rlabel metal2 9522 1248 9522 1248 0 N2END[4]
rlabel metal2 9798 1248 9798 1248 0 N2END[5]
rlabel metal2 10074 1248 10074 1248 0 N2END[6]
rlabel metal2 10350 1248 10350 1248 0 N2END[7]
rlabel metal2 6111 68 6111 68 0 N2MID[0]
rlabel metal2 6624 2924 6624 2924 0 N2MID[1]
rlabel metal2 6762 1214 6762 1214 0 N2MID[2]
rlabel metal2 7038 1214 7038 1214 0 N2MID[3]
rlabel metal2 7215 68 7215 68 0 N2MID[4]
rlabel metal2 7590 1214 7590 1214 0 N2MID[5]
rlabel metal2 7767 68 7767 68 0 N2MID[6]
rlabel metal2 8142 1282 8142 1282 0 N2MID[7]
rlabel metal2 10626 1248 10626 1248 0 N4END[0]
rlabel metal2 13287 68 13287 68 0 N4END[10]
rlabel metal2 13715 68 13715 68 0 N4END[11]
rlabel metal2 13885 68 13885 68 0 N4END[12]
rlabel metal2 14313 68 14313 68 0 N4END[13]
rlabel metal2 14490 1282 14490 1282 0 N4END[14]
rlabel metal2 14766 1214 14766 1214 0 N4END[15]
rlabel metal2 10902 1248 10902 1248 0 N4END[1]
rlabel metal2 11178 1248 11178 1248 0 N4END[2]
rlabel metal2 11454 1248 11454 1248 0 N4END[3]
rlabel metal2 11829 68 11829 68 0 N4END[4]
rlabel metal2 12006 1248 12006 1248 0 N4END[5]
rlabel metal2 12183 68 12183 68 0 N4END[6]
rlabel metal2 12505 68 12505 68 0 N4END[7]
rlabel metal2 12735 68 12735 68 0 N4END[8]
rlabel metal2 13011 68 13011 68 0 N4END[9]
rlabel metal2 14943 68 14943 68 0 NN4END[0]
rlabel metal2 17802 1554 17802 1554 0 NN4END[10]
rlabel metal2 18032 3502 18032 3502 0 NN4END[11]
rlabel metal2 18170 3026 18170 3026 0 NN4END[12]
rlabel metal1 18768 3502 18768 3502 0 NN4END[13]
rlabel metal1 18630 2958 18630 2958 0 NN4END[14]
rlabel metal2 19182 1282 19182 1282 0 NN4END[15]
rlabel metal2 15265 68 15265 68 0 NN4END[1]
rlabel metal2 15594 1214 15594 1214 0 NN4END[2]
rlabel metal2 15771 68 15771 68 0 NN4END[3]
rlabel metal2 16047 68 16047 68 0 NN4END[4]
rlabel metal2 16284 3026 16284 3026 0 NN4END[5]
rlabel metal1 16560 3026 16560 3026 0 NN4END[6]
rlabel metal2 16882 3026 16882 3026 0 NN4END[7]
rlabel metal2 17250 1554 17250 1554 0 NN4END[8]
rlabel metal2 17526 1554 17526 1554 0 NN4END[9]
rlabel metal2 19458 619 19458 619 0 S1BEG[0]
rlabel metal2 19734 1452 19734 1452 0 S1BEG[1]
rlabel metal1 20148 2822 20148 2822 0 S1BEG[2]
rlabel metal2 20187 68 20187 68 0 S1BEG[3]
rlabel metal2 22770 1452 22770 1452 0 S2BEG[0]
rlabel metal2 23046 1180 23046 1180 0 S2BEG[1]
rlabel metal2 23322 1180 23322 1180 0 S2BEG[2]
rlabel metal2 23598 619 23598 619 0 S2BEG[3]
rlabel metal2 23874 1452 23874 1452 0 S2BEG[4]
rlabel metal2 24150 1010 24150 1010 0 S2BEG[5]
rlabel metal2 24426 1452 24426 1452 0 S2BEG[6]
rlabel metal2 24702 1180 24702 1180 0 S2BEG[7]
rlabel metal1 20700 2822 20700 2822 0 S2BEGb[0]
rlabel metal2 20785 68 20785 68 0 S2BEGb[1]
rlabel metal1 21252 2822 21252 2822 0 S2BEGb[2]
rlabel metal2 21390 1214 21390 1214 0 S2BEGb[3]
rlabel metal1 21804 3366 21804 3366 0 S2BEGb[4]
rlabel metal2 21942 1214 21942 1214 0 S2BEGb[5]
rlabel metal2 22218 1044 22218 1044 0 S2BEGb[6]
rlabel metal2 22494 619 22494 619 0 S2BEGb[7]
rlabel metal2 24978 1452 24978 1452 0 S4BEG[0]
rlabel metal2 27738 1282 27738 1282 0 S4BEG[10]
rlabel metal2 28113 68 28113 68 0 S4BEG[11]
rlabel metal2 28389 68 28389 68 0 S4BEG[12]
rlabel metal2 28566 1486 28566 1486 0 S4BEG[13]
rlabel metal2 28842 619 28842 619 0 S4BEG[14]
rlabel metal2 29118 1622 29118 1622 0 S4BEG[15]
rlabel metal2 25353 68 25353 68 0 S4BEG[1]
rlabel metal2 25530 1452 25530 1452 0 S4BEG[2]
rlabel metal2 25905 68 25905 68 0 S4BEG[3]
rlabel metal2 26135 68 26135 68 0 S4BEG[4]
rlabel metal2 26457 68 26457 68 0 S4BEG[5]
rlabel metal2 26733 68 26733 68 0 S4BEG[6]
rlabel metal2 26910 1486 26910 1486 0 S4BEG[7]
rlabel metal2 27285 68 27285 68 0 S4BEG[8]
rlabel metal2 27515 68 27515 68 0 S4BEG[9]
rlabel metal2 29394 1350 29394 1350 0 SS4BEG[0]
rlabel metal2 32207 68 32207 68 0 SS4BEG[10]
rlabel metal1 32936 2890 32936 2890 0 SS4BEG[11]
rlabel metal1 32844 3366 32844 3366 0 SS4BEG[12]
rlabel metal2 33035 68 33035 68 0 SS4BEG[13]
rlabel metal2 33311 68 33311 68 0 SS4BEG[14]
rlabel metal1 34040 2890 34040 2890 0 SS4BEG[15]
rlabel metal2 29769 68 29769 68 0 SS4BEG[1]
rlabel metal2 30045 68 30045 68 0 SS4BEG[2]
rlabel metal2 30222 1486 30222 1486 0 SS4BEG[3]
rlabel metal2 30597 68 30597 68 0 SS4BEG[4]
rlabel metal2 30873 68 30873 68 0 SS4BEG[5]
rlabel metal2 31149 68 31149 68 0 SS4BEG[6]
rlabel metal2 31326 1486 31326 1486 0 SS4BEG[7]
rlabel metal2 31602 1078 31602 1078 0 SS4BEG[8]
rlabel metal1 32384 3162 32384 3162 0 SS4BEG[9]
rlabel metal2 33909 68 33909 68 0 UserCLK
rlabel metal2 1150 8680 1150 8680 0 UserCLKo
rlabel metal2 22954 6834 22954 6834 0 net1
rlabel metal1 40894 2448 40894 2448 0 net10
rlabel metal2 23506 2890 23506 2890 0 net100
rlabel metal1 23736 2346 23736 2346 0 net101
rlabel metal1 24058 3128 24058 3128 0 net102
rlabel metal1 25070 2448 25070 2448 0 net103
rlabel metal1 24610 2992 24610 2992 0 net104
rlabel metal1 25254 2346 25254 2346 0 net105
rlabel metal1 20746 3128 20746 3128 0 net106
rlabel metal1 20194 2482 20194 2482 0 net107
rlabel metal1 20838 3026 20838 3026 0 net108
rlabel metal1 20700 2414 20700 2414 0 net109
rlabel metal1 42642 2482 42642 2482 0 net11
rlabel metal1 19780 2278 19780 2278 0 net110
rlabel metal1 21114 2414 21114 2414 0 net111
rlabel metal1 22402 3128 22402 3128 0 net112
rlabel metal1 22540 2346 22540 2346 0 net113
rlabel metal1 25162 3128 25162 3128 0 net114
rlabel metal1 28566 2346 28566 2346 0 net115
rlabel metal1 28980 2618 28980 2618 0 net116
rlabel metal1 29348 2346 29348 2346 0 net117
rlabel metal2 29302 3298 29302 3298 0 net118
rlabel metal1 29992 2414 29992 2414 0 net119
rlabel metal1 35834 2346 35834 2346 0 net12
rlabel metal1 29210 3094 29210 3094 0 net120
rlabel metal1 25668 2414 25668 2414 0 net121
rlabel metal1 25714 2992 25714 2992 0 net122
rlabel metal1 25346 3128 25346 3128 0 net123
rlabel metal1 26680 2346 26680 2346 0 net124
rlabel metal1 25714 3400 25714 3400 0 net125
rlabel metal1 27738 2346 27738 2346 0 net126
rlabel metal1 27646 3128 27646 3128 0 net127
rlabel metal1 28060 2346 28060 2346 0 net128
rlabel metal1 28198 3128 28198 3128 0 net129
rlabel metal1 35006 3128 35006 3128 0 net13
rlabel metal1 25438 2550 25438 2550 0 net130
rlabel metal3 18860 2448 18860 2448 0 net131
rlabel metal2 15870 1598 15870 1598 0 net132
rlabel metal2 15410 1785 15410 1785 0 net133
rlabel metal2 15686 3842 15686 3842 0 net134
rlabel metal3 21252 2992 21252 2992 0 net135
rlabel metal2 15134 3706 15134 3706 0 net136
rlabel metal3 22379 2788 22379 2788 0 net137
rlabel metal2 24886 2482 24886 2482 0 net138
rlabel metal2 30498 2703 30498 2703 0 net139
rlabel metal1 35834 2414 35834 2414 0 net14
rlabel metal1 18630 3604 18630 3604 0 net140
rlabel metal2 23966 2261 23966 2261 0 net141
rlabel metal2 30866 1921 30866 1921 0 net142
rlabel metal2 17710 1785 17710 1785 0 net143
rlabel metal2 16514 1734 16514 1734 0 net144
rlabel metal4 30452 1972 30452 1972 0 net145
rlabel metal2 1518 6766 1518 6766 0 net146
rlabel metal1 36064 2550 36064 2550 0 net15
rlabel metal2 14306 3604 14306 3604 0 net16
rlabel metal1 16468 5202 16468 5202 0 net17
rlabel metal2 18906 6800 18906 6800 0 net18
rlabel metal1 26358 1836 26358 1836 0 net19
rlabel metal1 37950 2618 37950 2618 0 net2
rlabel metal2 23414 4386 23414 4386 0 net20
rlabel metal2 19826 3213 19826 3213 0 net21
rlabel metal2 19458 4148 19458 4148 0 net22
rlabel metal1 18630 3060 18630 3060 0 net23
rlabel metal2 17618 2040 17618 2040 0 net24
rlabel metal1 21574 3502 21574 3502 0 net25
rlabel via2 17894 3451 17894 3451 0 net26
rlabel metal2 18814 2669 18814 2669 0 net27
rlabel metal2 19458 2261 19458 2261 0 net28
rlabel metal2 20654 3893 20654 3893 0 net29
rlabel metal1 27738 7344 27738 7344 0 net3
rlabel metal1 18998 3706 18998 3706 0 net30
rlabel metal1 19274 2958 19274 2958 0 net31
rlabel metal2 20102 3706 20102 3706 0 net32
rlabel metal2 24242 4114 24242 4114 0 net33
rlabel metal2 6762 3910 6762 3910 0 net34
rlabel metal2 24058 1836 24058 1836 0 net35
rlabel metal2 23506 1581 23506 1581 0 net36
rlabel metal1 21850 1020 21850 1020 0 net37
rlabel metal2 22862 2516 22862 2516 0 net38
rlabel metal2 22770 3808 22770 3808 0 net39
rlabel metal1 37766 2924 37766 2924 0 net4
rlabel metal2 22954 2754 22954 2754 0 net40
rlabel metal2 28750 3978 28750 3978 0 net41
rlabel metal2 25714 2312 25714 2312 0 net42
rlabel metal1 17710 2992 17710 2992 0 net43
rlabel metal2 25254 2669 25254 2669 0 net44
rlabel metal1 14812 2822 14812 2822 0 net45
rlabel metal1 23092 3706 23092 3706 0 net46
rlabel metal2 23138 2686 23138 2686 0 net47
rlabel metal3 21988 3468 21988 3468 0 net48
rlabel metal3 22724 2108 22724 2108 0 net49
rlabel metal1 34270 2346 34270 2346 0 net5
rlabel metal3 21436 3672 21436 3672 0 net50
rlabel metal1 26220 1700 26220 1700 0 net51
rlabel metal2 27278 4029 27278 4029 0 net52
rlabel metal3 21436 3128 21436 3128 0 net53
rlabel metal2 26726 2482 26726 2482 0 net54
rlabel metal2 22126 3961 22126 3961 0 net55
rlabel metal2 25898 2533 25898 2533 0 net56
rlabel metal1 14950 3060 14950 3060 0 net57
rlabel metal1 17434 2414 17434 2414 0 net58
rlabel metal1 18446 3536 18446 3536 0 net59
rlabel metal1 38686 2550 38686 2550 0 net6
rlabel metal1 17848 2414 17848 2414 0 net60
rlabel metal1 18722 3094 18722 3094 0 net61
rlabel metal1 18262 2822 18262 2822 0 net62
rlabel metal1 18538 2550 18538 2550 0 net63
rlabel metal1 14582 2550 14582 2550 0 net64
rlabel metal1 15088 2958 15088 2958 0 net65
rlabel metal1 15226 2448 15226 2448 0 net66
rlabel metal2 15640 2652 15640 2652 0 net67
rlabel metal1 15962 2822 15962 2822 0 net68
rlabel metal1 16238 2822 16238 2822 0 net69
rlabel metal1 38870 2448 38870 2448 0 net7
rlabel metal1 16606 2822 16606 2822 0 net70
rlabel metal1 16882 2890 16882 2890 0 net71
rlabel metal1 17158 2482 17158 2482 0 net72
rlabel metal1 33902 2618 33902 2618 0 net73
rlabel metal1 18814 7412 18814 7412 0 net74
rlabel metal1 24702 5882 24702 5882 0 net75
rlabel metal1 27324 7446 27324 7446 0 net76
rlabel metal1 29118 3706 29118 3706 0 net77
rlabel metal1 31372 7378 31372 7378 0 net78
rlabel metal1 35466 7446 35466 7446 0 net79
rlabel metal1 38594 2380 38594 2380 0 net8
rlabel metal1 36938 7310 36938 7310 0 net80
rlabel metal2 38410 2176 38410 2176 0 net81
rlabel metal1 39928 2618 39928 2618 0 net82
rlabel metal2 41538 4998 41538 4998 0 net83
rlabel metal1 42642 7378 42642 7378 0 net84
rlabel metal1 6210 7378 6210 7378 0 net85
rlabel metal2 7682 7174 7682 7174 0 net86
rlabel metal1 20654 7276 20654 7276 0 net87
rlabel metal2 20470 7242 20470 7242 0 net88
rlabel metal1 14168 3162 14168 3162 0 net89
rlabel metal1 39606 2822 39606 2822 0 net9
rlabel metal1 16192 5338 16192 5338 0 net90
rlabel metal1 18492 7446 18492 7446 0 net91
rlabel metal1 20378 7480 20378 7480 0 net92
rlabel metal1 22540 6902 22540 6902 0 net93
rlabel metal1 18354 2346 18354 2346 0 net94
rlabel metal1 19596 3026 19596 3026 0 net95
rlabel metal1 19872 3094 19872 3094 0 net96
rlabel metal2 19642 2890 19642 2890 0 net97
rlabel metal1 22770 3094 22770 3094 0 net98
rlabel metal1 22632 2414 22632 2414 0 net99
<< properties >>
string FIXED_BBOX 0 0 44700 10000
<< end >>
