magic
tech sky130A
magscale 1 2
timestamp 1734825407
<< obsli1 >>
rect 1104 1071 108836 86513
<< obsm1 >>
rect 290 76 108864 87644
<< metal2 >>
rect 54956 0 54984 800
<< obsm2 >>
rect 296 856 108858 87650
rect 296 70 54900 856
rect 55040 70 108858 856
<< metal3 >>
rect 0 84358 800 84418
rect 0 83406 800 83466
rect 0 82454 800 82514
rect 0 81502 800 81562
rect 0 80550 800 80610
rect 0 79598 800 79658
rect 0 78646 800 78706
rect 0 77694 800 77754
rect 0 76742 800 76802
rect 0 75790 800 75850
rect 0 74838 800 74898
rect 0 73886 800 73946
rect 0 72934 800 72994
rect 0 71982 800 72042
rect 0 71030 800 71090
rect 0 70078 800 70138
rect 0 69126 800 69186
rect 0 68174 800 68234
rect 0 67222 800 67282
rect 0 66270 800 66330
rect 0 65318 800 65378
rect 0 64366 800 64426
rect 0 63414 800 63474
rect 0 62462 800 62522
rect 0 61510 800 61570
rect 0 60558 800 60618
rect 0 59606 800 59666
rect 0 58654 800 58714
rect 0 57702 800 57762
rect 0 56750 800 56810
rect 0 55798 800 55858
rect 0 54846 800 54906
rect 0 53894 800 53954
rect 0 52942 800 53002
rect 0 51990 800 52050
rect 0 51038 800 51098
rect 0 50086 800 50146
rect 0 49134 800 49194
rect 0 48182 800 48242
rect 0 47230 800 47290
rect 0 46278 800 46338
rect 0 45326 800 45386
rect 0 44374 800 44434
rect 0 43422 800 43482
rect 0 42470 800 42530
rect 0 41518 800 41578
rect 0 40566 800 40626
rect 0 39614 800 39674
rect 0 38662 800 38722
rect 0 37710 800 37770
rect 0 36758 800 36818
rect 0 35806 800 35866
rect 0 34854 800 34914
rect 0 33902 800 33962
rect 0 32950 800 33010
rect 0 31998 800 32058
rect 0 31046 800 31106
rect 0 30094 800 30154
rect 0 29142 800 29202
rect 0 28190 800 28250
rect 0 27238 800 27298
rect 0 26286 800 26346
rect 0 25334 800 25394
rect 0 24382 800 24442
rect 0 23430 800 23490
rect 0 22478 800 22538
rect 0 21526 800 21586
rect 0 20574 800 20634
rect 0 19622 800 19682
rect 0 18670 800 18730
rect 0 17718 800 17778
rect 0 16766 800 16826
rect 0 15814 800 15874
rect 0 14862 800 14922
rect 0 13910 800 13970
rect 0 12958 800 13018
rect 0 12006 800 12066
rect 0 11054 800 11114
rect 0 10102 800 10162
rect 0 9150 800 9210
rect 0 8198 800 8258
rect 0 7246 800 7306
rect 0 6294 800 6354
rect 0 5342 800 5402
rect 0 4390 800 4450
rect 0 3438 800 3498
<< obsm3 >>
rect 790 84498 108862 86529
rect 880 84278 108862 84498
rect 790 83546 108862 84278
rect 880 83326 108862 83546
rect 790 82594 108862 83326
rect 880 82374 108862 82594
rect 790 81642 108862 82374
rect 880 81422 108862 81642
rect 790 80690 108862 81422
rect 880 80470 108862 80690
rect 790 79738 108862 80470
rect 880 79518 108862 79738
rect 790 78786 108862 79518
rect 880 78566 108862 78786
rect 790 77834 108862 78566
rect 880 77614 108862 77834
rect 790 76882 108862 77614
rect 880 76662 108862 76882
rect 790 75930 108862 76662
rect 880 75710 108862 75930
rect 790 74978 108862 75710
rect 880 74758 108862 74978
rect 790 74026 108862 74758
rect 880 73806 108862 74026
rect 790 73074 108862 73806
rect 880 72854 108862 73074
rect 790 72122 108862 72854
rect 880 71902 108862 72122
rect 790 71170 108862 71902
rect 880 70950 108862 71170
rect 790 70218 108862 70950
rect 880 69998 108862 70218
rect 790 69266 108862 69998
rect 880 69046 108862 69266
rect 790 68314 108862 69046
rect 880 68094 108862 68314
rect 790 67362 108862 68094
rect 880 67142 108862 67362
rect 790 66410 108862 67142
rect 880 66190 108862 66410
rect 790 65458 108862 66190
rect 880 65238 108862 65458
rect 790 64506 108862 65238
rect 880 64286 108862 64506
rect 790 63554 108862 64286
rect 880 63334 108862 63554
rect 790 62602 108862 63334
rect 880 62382 108862 62602
rect 790 61650 108862 62382
rect 880 61430 108862 61650
rect 790 60698 108862 61430
rect 880 60478 108862 60698
rect 790 59746 108862 60478
rect 880 59526 108862 59746
rect 790 58794 108862 59526
rect 880 58574 108862 58794
rect 790 57842 108862 58574
rect 880 57622 108862 57842
rect 790 56890 108862 57622
rect 880 56670 108862 56890
rect 790 55938 108862 56670
rect 880 55718 108862 55938
rect 790 54986 108862 55718
rect 880 54766 108862 54986
rect 790 54034 108862 54766
rect 880 53814 108862 54034
rect 790 53082 108862 53814
rect 880 52862 108862 53082
rect 790 52130 108862 52862
rect 880 51910 108862 52130
rect 790 51178 108862 51910
rect 880 50958 108862 51178
rect 790 50226 108862 50958
rect 880 50006 108862 50226
rect 790 49274 108862 50006
rect 880 49054 108862 49274
rect 790 48322 108862 49054
rect 880 48102 108862 48322
rect 790 47370 108862 48102
rect 880 47150 108862 47370
rect 790 46418 108862 47150
rect 880 46198 108862 46418
rect 790 45466 108862 46198
rect 880 45246 108862 45466
rect 790 44514 108862 45246
rect 880 44294 108862 44514
rect 790 43562 108862 44294
rect 880 43342 108862 43562
rect 790 42610 108862 43342
rect 880 42390 108862 42610
rect 790 41658 108862 42390
rect 880 41438 108862 41658
rect 790 40706 108862 41438
rect 880 40486 108862 40706
rect 790 39754 108862 40486
rect 880 39534 108862 39754
rect 790 38802 108862 39534
rect 880 38582 108862 38802
rect 790 37850 108862 38582
rect 880 37630 108862 37850
rect 790 36898 108862 37630
rect 880 36678 108862 36898
rect 790 35946 108862 36678
rect 880 35726 108862 35946
rect 790 34994 108862 35726
rect 880 34774 108862 34994
rect 790 34042 108862 34774
rect 880 33822 108862 34042
rect 790 33090 108862 33822
rect 880 32870 108862 33090
rect 790 32138 108862 32870
rect 880 31918 108862 32138
rect 790 31186 108862 31918
rect 880 30966 108862 31186
rect 790 30234 108862 30966
rect 880 30014 108862 30234
rect 790 29282 108862 30014
rect 880 29062 108862 29282
rect 790 28330 108862 29062
rect 880 28110 108862 28330
rect 790 27378 108862 28110
rect 880 27158 108862 27378
rect 790 26426 108862 27158
rect 880 26206 108862 26426
rect 790 25474 108862 26206
rect 880 25254 108862 25474
rect 790 24522 108862 25254
rect 880 24302 108862 24522
rect 790 23570 108862 24302
rect 880 23350 108862 23570
rect 790 22618 108862 23350
rect 880 22398 108862 22618
rect 790 21666 108862 22398
rect 880 21446 108862 21666
rect 790 20714 108862 21446
rect 880 20494 108862 20714
rect 790 19762 108862 20494
rect 880 19542 108862 19762
rect 790 18810 108862 19542
rect 880 18590 108862 18810
rect 790 17858 108862 18590
rect 880 17638 108862 17858
rect 790 16906 108862 17638
rect 880 16686 108862 16906
rect 790 15954 108862 16686
rect 880 15734 108862 15954
rect 790 15002 108862 15734
rect 880 14782 108862 15002
rect 790 14050 108862 14782
rect 880 13830 108862 14050
rect 790 13098 108862 13830
rect 880 12878 108862 13098
rect 790 12146 108862 12878
rect 880 11926 108862 12146
rect 790 11194 108862 11926
rect 880 10974 108862 11194
rect 790 10242 108862 10974
rect 880 10022 108862 10242
rect 790 9290 108862 10022
rect 880 9070 108862 9290
rect 790 8338 108862 9070
rect 880 8118 108862 8338
rect 790 7386 108862 8118
rect 880 7166 108862 7386
rect 790 6434 108862 7166
rect 880 6214 108862 6434
rect 790 5482 108862 6214
rect 880 5262 108862 5482
rect 790 4530 108862 5262
rect 880 4310 108862 4530
rect 790 3578 108862 4310
rect 880 3358 108862 3578
rect 790 307 108862 3358
<< metal4 >>
rect -1076 -1092 -756 88676
rect -416 -432 -96 88016
rect 2944 -1092 3264 88676
rect 3604 -1092 3924 88676
rect 4544 -1092 4864 88676
rect 5204 -1092 5524 88676
rect 6144 -1092 6464 88676
rect 6804 -1092 7124 88676
rect 7744 -1092 8064 88676
rect 8404 -1092 8724 88676
rect 9344 -1092 9664 88676
rect 10004 85496 10324 88676
rect 10944 85496 11264 88676
rect 11604 85496 11924 88676
rect 12544 85496 12864 88676
rect 13204 85496 13524 88676
rect 14144 85496 14464 88676
rect 14804 85496 15124 88676
rect 15744 85496 16064 88676
rect 16404 85496 16724 88676
rect 17344 85496 17664 88676
rect 18004 85496 18324 88676
rect 18944 85496 19264 88676
rect 19604 85496 19924 88676
rect 20544 85496 20864 88676
rect 21204 85496 21524 88676
rect 22144 85496 22464 88676
rect 22804 85496 23124 88676
rect 23744 85496 24064 88676
rect 24404 85496 24724 88676
rect 25344 85496 25664 88676
rect 26004 85496 26324 88676
rect 26944 85496 27264 88676
rect 27604 85496 27924 88676
rect 28544 85496 28864 88676
rect 29204 85496 29524 88676
rect 30144 85496 30464 88676
rect 30804 85496 31124 88676
rect 31744 85496 32064 88676
rect 32404 85496 32724 88676
rect 33344 85496 33664 88676
rect 34004 85496 34324 88676
rect 34944 85496 35264 88676
rect 35604 85496 35924 88676
rect 36544 85496 36864 88676
rect 37204 85496 37524 88676
rect 38144 85496 38464 88676
rect 38804 85496 39124 88676
rect 39744 85620 40064 88676
rect 40404 85496 40724 88676
rect 41344 85620 41664 88676
rect 42004 85496 42324 88676
rect 42944 85496 43264 88676
rect 43604 85620 43924 88676
rect 44544 85496 44864 88676
rect 45204 85620 45524 88676
rect 46144 85620 46464 88676
rect 46804 85496 47124 88676
rect 47744 85620 48064 88676
rect 48404 85496 48724 88676
rect 49344 85496 49664 88676
rect 50004 85620 50324 88676
rect 50944 85620 51264 88676
rect 51604 85496 51924 88676
rect 52544 85620 52864 88676
rect 53204 85496 53524 88676
rect 54144 85496 54464 88676
rect 54804 85496 55124 88676
rect 55744 85496 56064 88676
rect 56404 85620 56724 88676
rect 57344 85620 57664 88676
rect 58004 85496 58324 88676
rect 58944 85620 59264 88676
rect 59604 85496 59924 88676
rect 60544 85496 60864 88676
rect 61204 85620 61524 88676
rect 62144 85496 62464 88676
rect 62804 85496 63124 88676
rect 63744 85620 64064 88676
rect 64404 85496 64724 88676
rect 65344 85496 65664 88676
rect 66004 85620 66324 88676
rect 66944 85496 67264 88676
rect 67604 85620 67924 88676
rect 68544 85620 68864 88676
rect 69204 85496 69524 88676
rect 70144 85620 70464 88676
rect 70804 85496 71124 88676
rect 71744 85496 72064 88676
rect 72404 85620 72724 88676
rect 73344 85496 73664 88676
rect 74004 85620 74324 88676
rect 74944 85620 75264 88676
rect 75604 85496 75924 88676
rect 76544 85496 76864 88676
rect 77204 85620 77524 88676
rect 78144 85496 78464 88676
rect 78804 85620 79124 88676
rect 79744 85496 80064 88676
rect 80404 85496 80724 88676
rect 81344 85496 81664 88676
rect 82004 85496 82324 88676
rect 82944 85496 83264 88676
rect 83604 85496 83924 88676
rect 84544 85496 84864 88676
rect 85204 85496 85524 88676
rect 86144 85496 86464 88676
rect 86804 85496 87124 88676
rect 87744 85496 88064 88676
rect 88404 85496 88724 88676
rect 89344 85496 89664 88676
rect 90004 85496 90324 88676
rect 90944 85496 91264 88676
rect 91604 85620 91924 88676
rect 92544 85496 92864 88676
rect 93204 85496 93524 88676
rect 94144 85496 94464 88676
rect 94804 85496 95124 88676
rect 95744 85496 96064 88676
rect 96404 85496 96724 88676
rect 97344 85496 97664 88676
rect 98004 85496 98324 88676
rect 98944 85496 99264 88676
rect 99604 85496 99924 88676
rect 100544 85496 100864 88676
rect 101204 85496 101524 88676
rect 102144 85620 102464 88676
rect 102804 85496 103124 88676
rect 103744 85496 104064 88676
rect 104404 85496 104724 88676
rect 105344 85496 105664 88676
rect 106004 85496 106324 88676
rect 106944 85496 107264 88676
rect 107604 85496 107924 88676
rect 108544 85496 108864 88676
rect 10004 -1092 10324 2004
rect 10944 -1092 11264 2004
rect 11604 -1092 11924 2004
rect 12544 -1092 12864 2004
rect 13204 -1092 13524 2004
rect 14144 -1092 14464 2004
rect 14804 -1092 15124 2004
rect 15744 -1092 16064 2004
rect 16404 -1092 16724 2004
rect 17344 -1092 17664 2004
rect 18004 -1092 18324 1880
rect 18944 -1092 19264 2004
rect 19604 -1092 19924 2004
rect 20544 -1092 20864 2004
rect 21204 -1092 21524 2004
rect 22144 -1092 22464 2004
rect 22804 -1092 23124 2004
rect 23744 -1092 24064 2004
rect 24404 -1092 24724 2004
rect 25344 -1092 25664 2004
rect 26004 -1092 26324 2004
rect 26944 -1092 27264 2004
rect 27604 -1092 27924 1880
rect 28544 -1092 28864 1880
rect 29204 -1092 29524 2004
rect 30144 -1092 30464 2004
rect 30804 -1092 31124 1880
rect 31744 -1092 32064 1880
rect 32404 -1092 32724 2004
rect 33344 -1092 33664 1880
rect 34004 -1092 34324 2004
rect 34944 -1092 35264 2004
rect 35604 -1092 35924 1880
rect 36544 -1092 36864 2004
rect 37204 -1092 37524 1880
rect 38144 -1092 38464 1880
rect 38804 -1092 39124 1880
rect 39744 -1092 40064 1880
rect 40404 -1092 40724 1880
rect 41344 -1092 41664 1880
rect 42004 -1092 42324 1880
rect 42944 -1092 43264 2004
rect 43604 -1092 43924 1880
rect 44544 -1092 44864 2004
rect 45204 -1092 45524 1880
rect 46144 -1092 46464 1880
rect 46804 -1092 47124 2004
rect 47744 -1092 48064 1880
rect 48404 -1092 48724 1880
rect 49344 -1092 49664 1880
rect 50004 -1092 50324 1880
rect 50944 -1092 51264 1880
rect 51604 -1092 51924 2004
rect 52544 -1092 52864 1880
rect 53204 -1092 53524 1880
rect 54144 -1092 54464 1880
rect 54804 -1092 55124 1880
rect 55744 -1092 56064 2004
rect 56404 -1092 56724 1880
rect 57344 -1092 57664 1880
rect 58004 -1092 58324 1880
rect 58944 -1092 59264 1880
rect 59604 -1092 59924 1880
rect 60544 -1092 60864 2004
rect 61204 -1092 61524 1880
rect 62144 -1092 62464 2004
rect 62804 -1092 63124 1880
rect 63744 -1092 64064 1880
rect 64404 -1092 64724 2004
rect 65344 -1092 65664 1880
rect 66004 -1092 66324 1880
rect 66944 -1092 67264 1880
rect 67604 -1092 67924 1880
rect 68544 -1092 68864 1880
rect 69204 -1092 69524 2004
rect 70144 -1092 70464 2004
rect 70804 -1092 71124 2004
rect 71744 -1092 72064 2004
rect 72404 -1092 72724 1880
rect 73344 -1092 73664 2004
rect 74004 -1092 74324 1880
rect 74944 -1092 75264 1880
rect 75604 -1092 75924 2004
rect 76544 -1092 76864 2004
rect 77204 -1092 77524 1880
rect 78144 -1092 78464 2004
rect 78804 -1092 79124 1880
rect 79744 -1092 80064 2004
rect 80404 -1092 80724 2004
rect 81344 -1092 81664 2004
rect 82004 -1092 82324 2004
rect 82944 -1092 83264 2004
rect 83604 -1092 83924 2004
rect 84544 -1092 84864 2004
rect 85204 -1092 85524 2004
rect 86144 -1092 86464 2004
rect 86804 -1092 87124 2004
rect 87744 -1092 88064 2004
rect 88404 -1092 88724 2004
rect 89344 -1092 89664 2004
rect 90004 -1092 90324 2004
rect 90944 -1092 91264 2004
rect 91604 -1092 91924 2004
rect 92544 -1092 92864 2004
rect 93204 -1092 93524 2004
rect 94144 -1092 94464 2004
rect 94804 -1092 95124 1880
rect 95744 -1092 96064 2004
rect 96404 -1092 96724 2004
rect 97344 -1092 97664 2004
rect 98004 -1092 98324 2004
rect 98944 -1092 99264 2004
rect 99604 -1092 99924 2004
rect 100544 -1092 100864 2004
rect 101204 -1092 101524 2004
rect 102144 -1092 102464 2004
rect 102804 -1092 103124 2004
rect 103744 -1092 104064 2004
rect 104404 -1092 104724 2004
rect 105344 -1092 105664 2004
rect 106004 -1092 106324 2004
rect 106944 -1092 107264 2004
rect 107604 -1092 107924 2004
rect 108544 -1092 108864 2004
rect 110036 -432 110356 88016
rect 110696 -1092 111016 88676
<< obsm4 >>
rect 795 443 2864 86189
rect 3344 443 3524 86189
rect 4004 443 4464 86189
rect 4944 443 5124 86189
rect 5604 443 6064 86189
rect 6544 443 6724 86189
rect 7204 443 7664 86189
rect 8144 443 8324 86189
rect 8804 443 9264 86189
rect 9744 85416 9924 86189
rect 10404 85416 10864 86189
rect 11344 85416 11524 86189
rect 12004 85416 12464 86189
rect 12944 85416 13124 86189
rect 13604 85416 14064 86189
rect 14544 85416 14724 86189
rect 15204 85416 15664 86189
rect 16144 85416 16324 86189
rect 16804 85416 17264 86189
rect 17744 85416 17924 86189
rect 18404 85416 18864 86189
rect 19344 85416 19524 86189
rect 20004 85416 20464 86189
rect 20944 85416 21124 86189
rect 21604 85416 22064 86189
rect 22544 85416 22724 86189
rect 23204 85416 23664 86189
rect 24144 85416 24324 86189
rect 24804 85416 25264 86189
rect 25744 85416 25924 86189
rect 26404 85416 26864 86189
rect 27344 85416 27524 86189
rect 28004 85416 28464 86189
rect 28944 85416 29124 86189
rect 29604 85416 30064 86189
rect 30544 85416 30724 86189
rect 31204 85416 31664 86189
rect 32144 85416 32324 86189
rect 32804 85416 33264 86189
rect 33744 85416 33924 86189
rect 34404 85416 34864 86189
rect 35344 85416 35524 86189
rect 36004 85416 36464 86189
rect 36944 85416 37124 86189
rect 37604 85416 38064 86189
rect 38544 85416 38724 86189
rect 39204 85540 39664 86189
rect 40144 85540 40324 86189
rect 39204 85416 40324 85540
rect 40804 85540 41264 86189
rect 41744 85540 41924 86189
rect 40804 85416 41924 85540
rect 42404 85416 42864 86189
rect 43344 85540 43524 86189
rect 44004 85540 44464 86189
rect 43344 85416 44464 85540
rect 44944 85540 45124 86189
rect 45604 85540 46064 86189
rect 46544 85540 46724 86189
rect 44944 85416 46724 85540
rect 47204 85540 47664 86189
rect 48144 85540 48324 86189
rect 47204 85416 48324 85540
rect 48804 85416 49264 86189
rect 49744 85540 49924 86189
rect 50404 85540 50864 86189
rect 51344 85540 51524 86189
rect 49744 85416 51524 85540
rect 52004 85540 52464 86189
rect 52944 85540 53124 86189
rect 52004 85416 53124 85540
rect 53604 85416 54064 86189
rect 54544 85416 54724 86189
rect 55204 85416 55664 86189
rect 56144 85540 56324 86189
rect 56804 85540 57264 86189
rect 57744 85540 57924 86189
rect 56144 85416 57924 85540
rect 58404 85540 58864 86189
rect 59344 85540 59524 86189
rect 58404 85416 59524 85540
rect 60004 85416 60464 86189
rect 60944 85540 61124 86189
rect 61604 85540 62064 86189
rect 60944 85416 62064 85540
rect 62544 85416 62724 86189
rect 63204 85540 63664 86189
rect 64144 85540 64324 86189
rect 63204 85416 64324 85540
rect 64804 85416 65264 86189
rect 65744 85540 65924 86189
rect 66404 85540 66864 86189
rect 65744 85416 66864 85540
rect 67344 85540 67524 86189
rect 68004 85540 68464 86189
rect 68944 85540 69124 86189
rect 67344 85416 69124 85540
rect 69604 85540 70064 86189
rect 70544 85540 70724 86189
rect 69604 85416 70724 85540
rect 71204 85416 71664 86189
rect 72144 85540 72324 86189
rect 72804 85540 73264 86189
rect 72144 85416 73264 85540
rect 73744 85540 73924 86189
rect 74404 85540 74864 86189
rect 75344 85540 75524 86189
rect 73744 85416 75524 85540
rect 76004 85416 76464 86189
rect 76944 85540 77124 86189
rect 77604 85540 78064 86189
rect 76944 85416 78064 85540
rect 78544 85540 78724 86189
rect 79204 85540 79664 86189
rect 78544 85416 79664 85540
rect 80144 85416 80324 86189
rect 80804 85416 81264 86189
rect 81744 85416 81924 86189
rect 82404 85416 82864 86189
rect 83344 85416 83524 86189
rect 84004 85416 84464 86189
rect 84944 85416 85124 86189
rect 85604 85416 86064 86189
rect 86544 85416 86724 86189
rect 87204 85416 87664 86189
rect 88144 85416 88324 86189
rect 88804 85416 89264 86189
rect 89744 85416 89924 86189
rect 90404 85416 90864 86189
rect 91344 85540 91524 86189
rect 92004 85540 92464 86189
rect 91344 85416 92464 85540
rect 92944 85416 93124 86189
rect 93604 85416 94064 86189
rect 94544 85416 94724 86189
rect 95204 85416 95664 86189
rect 96144 85416 96324 86189
rect 96804 85416 97264 86189
rect 97744 85416 97924 86189
rect 98404 85416 98864 86189
rect 99344 85416 99524 86189
rect 100004 85416 100464 86189
rect 100944 85416 101124 86189
rect 101604 85540 102064 86189
rect 102544 85540 102724 86189
rect 101604 85416 102724 85540
rect 103204 85416 103664 86189
rect 104144 85416 104324 86189
rect 104804 85416 105264 86189
rect 105744 85416 105924 86189
rect 106404 85416 106864 86189
rect 107344 85416 107524 86189
rect 9744 2084 107832 85416
rect 9744 443 9924 2084
rect 10404 443 10864 2084
rect 11344 443 11524 2084
rect 12004 443 12464 2084
rect 12944 443 13124 2084
rect 13604 443 14064 2084
rect 14544 443 14724 2084
rect 15204 443 15664 2084
rect 16144 443 16324 2084
rect 16804 443 17264 2084
rect 17744 1960 18864 2084
rect 17744 443 17924 1960
rect 18404 443 18864 1960
rect 19344 443 19524 2084
rect 20004 443 20464 2084
rect 20944 443 21124 2084
rect 21604 443 22064 2084
rect 22544 443 22724 2084
rect 23204 443 23664 2084
rect 24144 443 24324 2084
rect 24804 443 25264 2084
rect 25744 443 25924 2084
rect 26404 443 26864 2084
rect 27344 1960 29124 2084
rect 27344 443 27524 1960
rect 28004 443 28464 1960
rect 28944 443 29124 1960
rect 29604 443 30064 2084
rect 30544 1960 32324 2084
rect 30544 443 30724 1960
rect 31204 443 31664 1960
rect 32144 443 32324 1960
rect 32804 1960 33924 2084
rect 32804 443 33264 1960
rect 33744 443 33924 1960
rect 34404 443 34864 2084
rect 35344 1960 36464 2084
rect 35344 443 35524 1960
rect 36004 443 36464 1960
rect 36944 1960 42864 2084
rect 36944 443 37124 1960
rect 37604 443 38064 1960
rect 38544 443 38724 1960
rect 39204 443 39664 1960
rect 40144 443 40324 1960
rect 40804 443 41264 1960
rect 41744 443 41924 1960
rect 42404 443 42864 1960
rect 43344 1960 44464 2084
rect 43344 443 43524 1960
rect 44004 443 44464 1960
rect 44944 1960 46724 2084
rect 44944 443 45124 1960
rect 45604 443 46064 1960
rect 46544 443 46724 1960
rect 47204 1960 51524 2084
rect 47204 443 47664 1960
rect 48144 443 48324 1960
rect 48804 443 49264 1960
rect 49744 443 49924 1960
rect 50404 443 50864 1960
rect 51344 443 51524 1960
rect 52004 1960 55664 2084
rect 52004 443 52464 1960
rect 52944 443 53124 1960
rect 53604 443 54064 1960
rect 54544 443 54724 1960
rect 55204 443 55664 1960
rect 56144 1960 60464 2084
rect 56144 443 56324 1960
rect 56804 443 57264 1960
rect 57744 443 57924 1960
rect 58404 443 58864 1960
rect 59344 443 59524 1960
rect 60004 443 60464 1960
rect 60944 1960 62064 2084
rect 60944 443 61124 1960
rect 61604 443 62064 1960
rect 62544 1960 64324 2084
rect 62544 443 62724 1960
rect 63204 443 63664 1960
rect 64144 443 64324 1960
rect 64804 1960 69124 2084
rect 64804 443 65264 1960
rect 65744 443 65924 1960
rect 66404 443 66864 1960
rect 67344 443 67524 1960
rect 68004 443 68464 1960
rect 68944 443 69124 1960
rect 69604 443 70064 2084
rect 70544 443 70724 2084
rect 71204 443 71664 2084
rect 72144 1960 73264 2084
rect 72144 443 72324 1960
rect 72804 443 73264 1960
rect 73744 1960 75524 2084
rect 73744 443 73924 1960
rect 74404 443 74864 1960
rect 75344 443 75524 1960
rect 76004 443 76464 2084
rect 76944 1960 78064 2084
rect 76944 443 77124 1960
rect 77604 443 78064 1960
rect 78544 1960 79664 2084
rect 78544 443 78724 1960
rect 79204 443 79664 1960
rect 80144 443 80324 2084
rect 80804 443 81264 2084
rect 81744 443 81924 2084
rect 82404 443 82864 2084
rect 83344 443 83524 2084
rect 84004 443 84464 2084
rect 84944 443 85124 2084
rect 85604 443 86064 2084
rect 86544 443 86724 2084
rect 87204 443 87664 2084
rect 88144 443 88324 2084
rect 88804 443 89264 2084
rect 89744 443 89924 2084
rect 90404 443 90864 2084
rect 91344 443 91524 2084
rect 92004 443 92464 2084
rect 92944 443 93124 2084
rect 93604 443 94064 2084
rect 94544 1960 95664 2084
rect 94544 443 94724 1960
rect 95204 443 95664 1960
rect 96144 443 96324 2084
rect 96804 443 97264 2084
rect 97744 443 97924 2084
rect 98404 443 98864 2084
rect 99344 443 99524 2084
rect 100004 443 100464 2084
rect 100944 443 101124 2084
rect 101604 443 102064 2084
rect 102544 443 102724 2084
rect 103204 443 103664 2084
rect 104144 443 104324 2084
rect 104804 443 105264 2084
rect 105744 443 105924 2084
rect 106404 443 106864 2084
rect 107344 443 107524 2084
<< metal5 >>
rect -1076 88356 111016 88676
rect -416 87696 110356 88016
rect -1076 82588 111016 82908
rect -1076 81928 111016 82248
rect -1076 6588 111016 6908
rect -1076 5928 111016 6248
rect -416 -432 110356 -112
rect -1076 -1092 111016 -772
<< labels >>
rlabel metal3 s 0 22478 800 22538 6 C0
port 1 nsew signal input
rlabel metal3 s 0 23430 800 23490 6 C1
port 2 nsew signal input
rlabel metal3 s 0 24382 800 24442 6 C2
port 3 nsew signal input
rlabel metal3 s 0 25334 800 25394 6 C3
port 4 nsew signal input
rlabel metal3 s 0 60558 800 60618 6 C4
port 5 nsew signal input
rlabel metal3 s 0 61510 800 61570 6 C5
port 6 nsew signal input
rlabel metal2 s 54956 0 54984 800 6 clk
port 7 nsew signal input
rlabel metal3 s 0 18670 800 18730 6 rd_addr[0]
port 8 nsew signal input
rlabel metal3 s 0 19622 800 19682 6 rd_addr[1]
port 9 nsew signal input
rlabel metal3 s 0 20574 800 20634 6 rd_addr[2]
port 10 nsew signal input
rlabel metal3 s 0 21526 800 21586 6 rd_addr[3]
port 11 nsew signal input
rlabel metal3 s 0 26286 800 26346 6 rd_addr[4]
port 12 nsew signal input
rlabel metal3 s 0 27238 800 27298 6 rd_addr[5]
port 13 nsew signal input
rlabel metal3 s 0 35806 800 35866 6 rd_addr[6]
port 14 nsew signal input
rlabel metal3 s 0 36758 800 36818 6 rd_addr[7]
port 15 nsew signal input
rlabel metal3 s 0 17718 800 17778 6 rd_data[0]
port 16 nsew signal output
rlabel metal3 s 0 8198 800 8258 6 rd_data[10]
port 17 nsew signal output
rlabel metal3 s 0 7246 800 7306 6 rd_data[11]
port 18 nsew signal output
rlabel metal3 s 0 3438 800 3498 6 rd_data[12]
port 19 nsew signal output
rlabel metal3 s 0 4390 800 4450 6 rd_data[13]
port 20 nsew signal output
rlabel metal3 s 0 5342 800 5402 6 rd_data[14]
port 21 nsew signal output
rlabel metal3 s 0 6294 800 6354 6 rd_data[15]
port 22 nsew signal output
rlabel metal3 s 0 45326 800 45386 6 rd_data[16]
port 23 nsew signal output
rlabel metal3 s 0 46278 800 46338 6 rd_data[17]
port 24 nsew signal output
rlabel metal3 s 0 47230 800 47290 6 rd_data[18]
port 25 nsew signal output
rlabel metal3 s 0 48182 800 48242 6 rd_data[19]
port 26 nsew signal output
rlabel metal3 s 0 16766 800 16826 6 rd_data[1]
port 27 nsew signal output
rlabel metal3 s 0 49134 800 49194 6 rd_data[20]
port 28 nsew signal output
rlabel metal3 s 0 50086 800 50146 6 rd_data[21]
port 29 nsew signal output
rlabel metal3 s 0 51038 800 51098 6 rd_data[22]
port 30 nsew signal output
rlabel metal3 s 0 51990 800 52050 6 rd_data[23]
port 31 nsew signal output
rlabel metal3 s 0 52942 800 53002 6 rd_data[24]
port 32 nsew signal output
rlabel metal3 s 0 53894 800 53954 6 rd_data[25]
port 33 nsew signal output
rlabel metal3 s 0 54846 800 54906 6 rd_data[26]
port 34 nsew signal output
rlabel metal3 s 0 55798 800 55858 6 rd_data[27]
port 35 nsew signal output
rlabel metal3 s 0 56750 800 56810 6 rd_data[28]
port 36 nsew signal output
rlabel metal3 s 0 57702 800 57762 6 rd_data[29]
port 37 nsew signal output
rlabel metal3 s 0 15814 800 15874 6 rd_data[2]
port 38 nsew signal output
rlabel metal3 s 0 58654 800 58714 6 rd_data[30]
port 39 nsew signal output
rlabel metal3 s 0 59606 800 59666 6 rd_data[31]
port 40 nsew signal output
rlabel metal3 s 0 14862 800 14922 6 rd_data[3]
port 41 nsew signal output
rlabel metal3 s 0 13910 800 13970 6 rd_data[4]
port 42 nsew signal output
rlabel metal3 s 0 12958 800 13018 6 rd_data[5]
port 43 nsew signal output
rlabel metal3 s 0 12006 800 12066 6 rd_data[6]
port 44 nsew signal output
rlabel metal3 s 0 11054 800 11114 6 rd_data[7]
port 45 nsew signal output
rlabel metal3 s 0 10102 800 10162 6 rd_data[8]
port 46 nsew signal output
rlabel metal3 s 0 9150 800 9210 6 rd_data[9]
port 47 nsew signal output
rlabel metal4 s -416 -432 -96 88016 4 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -416 -432 110356 -112 8 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -416 87696 110356 88016 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 110036 -432 110356 88016 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 3604 -1092 3924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 5204 -1092 5524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 6804 -1092 7124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 8404 -1092 8724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 10004 -1092 10324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 10004 85496 10324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 11604 -1092 11924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 11604 85496 11924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 13204 -1092 13524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 13204 85496 13524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 14804 -1092 15124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 14804 85496 15124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 16404 -1092 16724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 16404 85496 16724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 18004 -1092 18324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 18004 85496 18324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 19604 -1092 19924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 19604 85496 19924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 21204 -1092 21524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 21204 85496 21524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 22804 -1092 23124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 22804 85496 23124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 24404 -1092 24724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 24404 85496 24724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 26004 -1092 26324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 26004 85496 26324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 27604 -1092 27924 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 27604 85496 27924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 29204 -1092 29524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 29204 85496 29524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 30804 -1092 31124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 30804 85496 31124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 32404 -1092 32724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 32404 85496 32724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 34004 -1092 34324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 34004 85496 34324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 35604 -1092 35924 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 35604 85496 35924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 37204 -1092 37524 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 37204 85496 37524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 38804 -1092 39124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 38804 85496 39124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 40404 -1092 40724 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 40404 85496 40724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 42004 -1092 42324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 42004 85496 42324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 43604 -1092 43924 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 43604 85620 43924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 45204 -1092 45524 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 45204 85620 45524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 46804 -1092 47124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 46804 85496 47124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 48404 -1092 48724 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 48404 85496 48724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 50004 -1092 50324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 50004 85620 50324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 51604 -1092 51924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 51604 85496 51924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 53204 -1092 53524 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 53204 85496 53524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 54804 -1092 55124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 54804 85496 55124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 56404 -1092 56724 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 56404 85620 56724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 58004 -1092 58324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 58004 85496 58324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 59604 -1092 59924 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 59604 85496 59924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 61204 -1092 61524 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 61204 85620 61524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 62804 -1092 63124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 62804 85496 63124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 64404 -1092 64724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 64404 85496 64724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 66004 -1092 66324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 66004 85620 66324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 67604 -1092 67924 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 67604 85620 67924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 69204 -1092 69524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 69204 85496 69524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 70804 -1092 71124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 70804 85496 71124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 72404 -1092 72724 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 72404 85620 72724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 74004 -1092 74324 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 74004 85620 74324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 75604 -1092 75924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 75604 85496 75924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 77204 -1092 77524 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 77204 85620 77524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 78804 -1092 79124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 78804 85620 79124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 80404 -1092 80724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 80404 85496 80724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 82004 -1092 82324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 82004 85496 82324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 83604 -1092 83924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 83604 85496 83924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 85204 -1092 85524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 85204 85496 85524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 86804 -1092 87124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 86804 85496 87124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 88404 -1092 88724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 88404 85496 88724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 90004 -1092 90324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 90004 85496 90324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 91604 -1092 91924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 91604 85620 91924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 93204 -1092 93524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 93204 85496 93524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 94804 -1092 95124 1880 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 94804 85496 95124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 96404 -1092 96724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 96404 85496 96724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 98004 -1092 98324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 98004 85496 98324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 99604 -1092 99924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 99604 85496 99924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 101204 -1092 101524 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 101204 85496 101524 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 102804 -1092 103124 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 102804 85496 103124 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 104404 -1092 104724 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 104404 85496 104724 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 106004 -1092 106324 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 106004 85496 106324 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 107604 -1092 107924 2004 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 107604 85496 107924 88676 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -1076 6588 111016 6908 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -1076 82588 111016 82908 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s -1076 -1092 -756 88676 4 vssd1
port 49 nsew ground bidirectional
rlabel metal5 s -1076 -1092 111016 -772 8 vssd1
port 49 nsew ground bidirectional
rlabel metal5 s -1076 88356 111016 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 110696 -1092 111016 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 2944 -1092 3264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 4544 -1092 4864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 6144 -1092 6464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 7744 -1092 8064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 9344 -1092 9664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 10944 -1092 11264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 10944 85496 11264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 12544 -1092 12864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 12544 85496 12864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 14144 -1092 14464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 14144 85496 14464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 15744 -1092 16064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 15744 85496 16064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 17344 -1092 17664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 17344 85496 17664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 18944 -1092 19264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 18944 85496 19264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 20544 -1092 20864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 20544 85496 20864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 22144 -1092 22464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 22144 85496 22464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 23744 -1092 24064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 23744 85496 24064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 25344 -1092 25664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 25344 85496 25664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 26944 -1092 27264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 26944 85496 27264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 28544 -1092 28864 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 28544 85496 28864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 30144 -1092 30464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 30144 85496 30464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 31744 -1092 32064 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 31744 85496 32064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 33344 -1092 33664 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 33344 85496 33664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 34944 -1092 35264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 34944 85496 35264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 36544 -1092 36864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 36544 85496 36864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 38144 -1092 38464 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 38144 85496 38464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 39744 -1092 40064 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 39744 85620 40064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 41344 -1092 41664 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 41344 85620 41664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 42944 -1092 43264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 42944 85496 43264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 44544 -1092 44864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 44544 85496 44864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 46144 -1092 46464 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 46144 85620 46464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 47744 -1092 48064 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 47744 85620 48064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 49344 -1092 49664 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 49344 85496 49664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 50944 -1092 51264 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 50944 85620 51264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 52544 -1092 52864 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 52544 85620 52864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 54144 -1092 54464 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 54144 85496 54464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 55744 -1092 56064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 55744 85496 56064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 57344 -1092 57664 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 57344 85620 57664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 58944 -1092 59264 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 58944 85620 59264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 60544 -1092 60864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 60544 85496 60864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 62144 -1092 62464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 62144 85496 62464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 63744 -1092 64064 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 63744 85620 64064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 65344 -1092 65664 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 65344 85496 65664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 66944 -1092 67264 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 66944 85496 67264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 68544 -1092 68864 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 68544 85620 68864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 70144 -1092 70464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 70144 85620 70464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 71744 -1092 72064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 71744 85496 72064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 73344 -1092 73664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 73344 85496 73664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 74944 -1092 75264 1880 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 74944 85620 75264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 76544 -1092 76864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 76544 85496 76864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 78144 -1092 78464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 78144 85496 78464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 79744 -1092 80064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 79744 85496 80064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 81344 -1092 81664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 81344 85496 81664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 82944 -1092 83264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 82944 85496 83264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 84544 -1092 84864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 84544 85496 84864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 86144 -1092 86464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 86144 85496 86464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 87744 -1092 88064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 87744 85496 88064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 89344 -1092 89664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 89344 85496 89664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 90944 -1092 91264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 90944 85496 91264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 92544 -1092 92864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 92544 85496 92864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 94144 -1092 94464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 94144 85496 94464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 95744 -1092 96064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 95744 85496 96064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 97344 -1092 97664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 97344 85496 97664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 98944 -1092 99264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 98944 85496 99264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 100544 -1092 100864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 100544 85496 100864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 102144 -1092 102464 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 102144 85620 102464 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 103744 -1092 104064 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 103744 85496 104064 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 105344 -1092 105664 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 105344 85496 105664 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 106944 -1092 107264 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 106944 85496 107264 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 108544 -1092 108864 2004 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 108544 85496 108864 88676 6 vssd1
port 49 nsew ground bidirectional
rlabel metal5 s -1076 5928 111016 6248 6 vssd1
port 49 nsew ground bidirectional
rlabel metal5 s -1076 81928 111016 82248 6 vssd1
port 49 nsew ground bidirectional
rlabel metal3 s 0 62462 800 62522 6 wr_addr[0]
port 50 nsew signal input
rlabel metal3 s 0 63414 800 63474 6 wr_addr[1]
port 51 nsew signal input
rlabel metal3 s 0 64366 800 64426 6 wr_addr[2]
port 52 nsew signal input
rlabel metal3 s 0 65318 800 65378 6 wr_addr[3]
port 53 nsew signal input
rlabel metal3 s 0 66270 800 66330 6 wr_addr[4]
port 54 nsew signal input
rlabel metal3 s 0 67222 800 67282 6 wr_addr[5]
port 55 nsew signal input
rlabel metal3 s 0 68174 800 68234 6 wr_addr[6]
port 56 nsew signal input
rlabel metal3 s 0 69126 800 69186 6 wr_addr[7]
port 57 nsew signal input
rlabel metal3 s 0 37710 800 37770 6 wr_data[0]
port 58 nsew signal input
rlabel metal3 s 0 28190 800 28250 6 wr_data[10]
port 59 nsew signal input
rlabel metal3 s 0 29142 800 29202 6 wr_data[11]
port 60 nsew signal input
rlabel metal3 s 0 30094 800 30154 6 wr_data[12]
port 61 nsew signal input
rlabel metal3 s 0 31046 800 31106 6 wr_data[13]
port 62 nsew signal input
rlabel metal3 s 0 43422 800 43482 6 wr_data[14]
port 63 nsew signal input
rlabel metal3 s 0 44374 800 44434 6 wr_data[15]
port 64 nsew signal input
rlabel metal3 s 0 70078 800 70138 6 wr_data[16]
port 65 nsew signal input
rlabel metal3 s 0 71030 800 71090 6 wr_data[17]
port 66 nsew signal input
rlabel metal3 s 0 71982 800 72042 6 wr_data[18]
port 67 nsew signal input
rlabel metal3 s 0 72934 800 72994 6 wr_data[19]
port 68 nsew signal input
rlabel metal3 s 0 38662 800 38722 6 wr_data[1]
port 69 nsew signal input
rlabel metal3 s 0 73886 800 73946 6 wr_data[20]
port 70 nsew signal input
rlabel metal3 s 0 74838 800 74898 6 wr_data[21]
port 71 nsew signal input
rlabel metal3 s 0 75790 800 75850 6 wr_data[22]
port 72 nsew signal input
rlabel metal3 s 0 76742 800 76802 6 wr_data[23]
port 73 nsew signal input
rlabel metal3 s 0 77694 800 77754 6 wr_data[24]
port 74 nsew signal input
rlabel metal3 s 0 78646 800 78706 6 wr_data[25]
port 75 nsew signal input
rlabel metal3 s 0 79598 800 79658 6 wr_data[26]
port 76 nsew signal input
rlabel metal3 s 0 80550 800 80610 6 wr_data[27]
port 77 nsew signal input
rlabel metal3 s 0 81502 800 81562 6 wr_data[28]
port 78 nsew signal input
rlabel metal3 s 0 82454 800 82514 6 wr_data[29]
port 79 nsew signal input
rlabel metal3 s 0 39614 800 39674 6 wr_data[2]
port 80 nsew signal input
rlabel metal3 s 0 83406 800 83466 6 wr_data[30]
port 81 nsew signal input
rlabel metal3 s 0 84358 800 84418 6 wr_data[31]
port 82 nsew signal input
rlabel metal3 s 0 40566 800 40626 6 wr_data[3]
port 83 nsew signal input
rlabel metal3 s 0 41518 800 41578 6 wr_data[4]
port 84 nsew signal input
rlabel metal3 s 0 42470 800 42530 6 wr_data[5]
port 85 nsew signal input
rlabel metal3 s 0 31998 800 32058 6 wr_data[6]
port 86 nsew signal input
rlabel metal3 s 0 32950 800 33010 6 wr_data[7]
port 87 nsew signal input
rlabel metal3 s 0 33902 800 33962 6 wr_data[8]
port 88 nsew signal input
rlabel metal3 s 0 34854 800 34914 6 wr_data[9]
port 89 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 88000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12083696
string GDS_FILE /home/asma/open_eFPGA_v2/openlane/BRAM/runs/24_12_21_23_54/results/signoff/BlockRAM_1KB.magic.gds
string GDS_START 9636152
<< end >>

