magic
tech sky130A
magscale 1 2
timestamp 1733616291
<< obsli1 >>
rect 1104 1071 24564 43537
<< obsm1 >>
rect 14 416 25654 44328
<< metal2 >>
rect 110 44540 166 45000
rect 386 44540 442 45000
rect 662 44540 718 45000
rect 938 44540 994 45000
rect 1214 44540 1270 45000
rect 1490 44540 1546 45000
rect 1766 44540 1822 45000
rect 2042 44540 2098 45000
rect 2318 44540 2374 45000
rect 2594 44540 2650 45000
rect 2870 44540 2926 45000
rect 3146 44540 3202 45000
rect 3422 44540 3478 45000
rect 3698 44540 3754 45000
rect 3974 44540 4030 45000
rect 4250 44540 4306 45000
rect 4526 44540 4582 45000
rect 4802 44540 4858 45000
rect 5078 44540 5134 45000
rect 5354 44540 5410 45000
rect 5630 44540 5686 45000
rect 5906 44540 5962 45000
rect 6182 44540 6238 45000
rect 6458 44540 6514 45000
rect 6734 44540 6790 45000
rect 7010 44540 7066 45000
rect 7286 44540 7342 45000
rect 7562 44540 7618 45000
rect 7838 44540 7894 45000
rect 8114 44540 8170 45000
rect 8390 44540 8446 45000
rect 8666 44540 8722 45000
rect 8942 44540 8998 45000
rect 9218 44540 9274 45000
rect 9494 44540 9550 45000
rect 9770 44540 9826 45000
rect 10046 44540 10102 45000
rect 10322 44540 10378 45000
rect 10598 44540 10654 45000
rect 10874 44540 10930 45000
rect 11150 44540 11206 45000
rect 11426 44540 11482 45000
rect 11702 44540 11758 45000
rect 11978 44540 12034 45000
rect 12254 44540 12310 45000
rect 12530 44540 12586 45000
rect 12806 44540 12862 45000
rect 13082 44540 13138 45000
rect 13358 44540 13414 45000
rect 13634 44540 13690 45000
rect 13910 44540 13966 45000
rect 14186 44540 14242 45000
rect 14462 44540 14518 45000
rect 14738 44540 14794 45000
rect 15014 44540 15070 45000
rect 15290 44540 15346 45000
rect 15566 44540 15622 45000
rect 15842 44540 15898 45000
rect 16118 44540 16174 45000
rect 16394 44540 16450 45000
rect 16670 44540 16726 45000
rect 16946 44540 17002 45000
rect 17222 44540 17278 45000
rect 17498 44540 17554 45000
rect 17774 44540 17830 45000
rect 18050 44540 18106 45000
rect 18326 44540 18382 45000
rect 18602 44540 18658 45000
rect 18878 44540 18934 45000
rect 19154 44540 19210 45000
rect 19430 44540 19486 45000
rect 19706 44540 19762 45000
rect 19982 44540 20038 45000
rect 20258 44540 20314 45000
rect 20534 44540 20590 45000
rect 20810 44540 20866 45000
rect 21086 44540 21142 45000
rect 21362 44540 21418 45000
rect 21638 44540 21694 45000
rect 21914 44540 21970 45000
rect 22190 44540 22246 45000
rect 22466 44540 22522 45000
rect 22742 44540 22798 45000
rect 23018 44540 23074 45000
rect 23294 44540 23350 45000
rect 23570 44540 23626 45000
rect 23846 44540 23902 45000
rect 24122 44540 24178 45000
rect 24398 44540 24454 45000
rect 24674 44540 24730 45000
rect 24950 44540 25006 45000
rect 25226 44540 25282 45000
rect 25502 44540 25558 45000
rect 110 -300 166 160
rect 386 -300 442 160
rect 662 -300 718 160
rect 938 -300 994 160
rect 1214 -300 1270 160
rect 1490 -300 1546 160
rect 1766 -300 1822 160
rect 2042 -300 2098 160
rect 2318 -300 2374 160
rect 2594 -300 2650 160
rect 2870 -300 2926 160
rect 3146 -300 3202 160
rect 3422 -300 3478 160
rect 3698 -300 3754 160
rect 3974 -300 4030 160
rect 4250 -300 4306 160
rect 4526 -300 4582 160
rect 4802 -300 4858 160
rect 5078 -300 5134 160
rect 5354 -300 5410 160
rect 5630 -300 5686 160
rect 5906 -300 5962 160
rect 6182 -300 6238 160
rect 6458 -300 6514 160
rect 6734 -300 6790 160
rect 7010 -300 7066 160
rect 7286 -300 7342 160
rect 7562 -300 7618 160
rect 7838 -300 7894 160
rect 8114 -300 8170 160
rect 8390 -300 8446 160
rect 8666 -300 8722 160
rect 8942 -300 8998 160
rect 9218 -300 9274 160
rect 9494 -300 9550 160
rect 9770 -300 9826 160
rect 10046 -300 10102 160
rect 10322 -300 10378 160
rect 10598 -300 10654 160
rect 10874 -300 10930 160
rect 11150 -300 11206 160
rect 11426 -300 11482 160
rect 11702 -300 11758 160
rect 11978 -300 12034 160
rect 12254 -300 12310 160
rect 12530 -300 12586 160
rect 12806 -300 12862 160
rect 13082 -300 13138 160
rect 13358 -300 13414 160
rect 13634 -300 13690 160
rect 13910 -300 13966 160
rect 14186 -300 14242 160
rect 14462 -300 14518 160
rect 14738 -300 14794 160
rect 15014 -300 15070 160
rect 15290 -300 15346 160
rect 15566 -300 15622 160
rect 15842 -300 15898 160
rect 16118 -300 16174 160
rect 16394 -300 16450 160
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 -300 17278 160
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 18050 -300 18106 160
rect 18326 -300 18382 160
rect 18602 -300 18658 160
rect 18878 -300 18934 160
rect 19154 -300 19210 160
rect 19430 -300 19486 160
rect 19706 -300 19762 160
rect 19982 -300 20038 160
rect 20258 -300 20314 160
rect 20534 -300 20590 160
rect 20810 -300 20866 160
rect 21086 -300 21142 160
rect 21362 -300 21418 160
rect 21638 -300 21694 160
rect 21914 -300 21970 160
rect 22190 -300 22246 160
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 23018 -300 23074 160
rect 23294 -300 23350 160
rect 23570 -300 23626 160
rect 23846 -300 23902 160
rect 24122 -300 24178 160
rect 24398 -300 24454 160
rect 24674 -300 24730 160
rect 24950 -300 25006 160
rect 25226 -300 25282 160
rect 25502 -300 25558 160
<< obsm2 >>
rect 20 44484 54 44540
rect 222 44484 330 44540
rect 498 44484 606 44540
rect 774 44484 882 44540
rect 1050 44484 1158 44540
rect 1326 44484 1434 44540
rect 1602 44484 1710 44540
rect 1878 44484 1986 44540
rect 2154 44484 2262 44540
rect 2430 44484 2538 44540
rect 2706 44484 2814 44540
rect 2982 44484 3090 44540
rect 3258 44484 3366 44540
rect 3534 44484 3642 44540
rect 3810 44484 3918 44540
rect 4086 44484 4194 44540
rect 4362 44484 4470 44540
rect 4638 44484 4746 44540
rect 4914 44484 5022 44540
rect 5190 44484 5298 44540
rect 5466 44484 5574 44540
rect 5742 44484 5850 44540
rect 6018 44484 6126 44540
rect 6294 44484 6402 44540
rect 6570 44484 6678 44540
rect 6846 44484 6954 44540
rect 7122 44484 7230 44540
rect 7398 44484 7506 44540
rect 7674 44484 7782 44540
rect 7950 44484 8058 44540
rect 8226 44484 8334 44540
rect 8502 44484 8610 44540
rect 8778 44484 8886 44540
rect 9054 44484 9162 44540
rect 9330 44484 9438 44540
rect 9606 44484 9714 44540
rect 9882 44484 9990 44540
rect 10158 44484 10266 44540
rect 10434 44484 10542 44540
rect 10710 44484 10818 44540
rect 10986 44484 11094 44540
rect 11262 44484 11370 44540
rect 11538 44484 11646 44540
rect 11814 44484 11922 44540
rect 12090 44484 12198 44540
rect 12366 44484 12474 44540
rect 12642 44484 12750 44540
rect 12918 44484 13026 44540
rect 13194 44484 13302 44540
rect 13470 44484 13578 44540
rect 13746 44484 13854 44540
rect 14022 44484 14130 44540
rect 14298 44484 14406 44540
rect 14574 44484 14682 44540
rect 14850 44484 14958 44540
rect 15126 44484 15234 44540
rect 15402 44484 15510 44540
rect 15678 44484 15786 44540
rect 15954 44484 16062 44540
rect 16230 44484 16338 44540
rect 16506 44484 16614 44540
rect 16782 44484 16890 44540
rect 17058 44484 17166 44540
rect 17334 44484 17442 44540
rect 17610 44484 17718 44540
rect 17886 44484 17994 44540
rect 18162 44484 18270 44540
rect 18438 44484 18546 44540
rect 18714 44484 18822 44540
rect 18990 44484 19098 44540
rect 19266 44484 19374 44540
rect 19542 44484 19650 44540
rect 19818 44484 19926 44540
rect 20094 44484 20202 44540
rect 20370 44484 20478 44540
rect 20646 44484 20754 44540
rect 20922 44484 21030 44540
rect 21198 44484 21306 44540
rect 21474 44484 21582 44540
rect 21750 44484 21858 44540
rect 22026 44484 22134 44540
rect 22302 44484 22410 44540
rect 22578 44484 22686 44540
rect 22854 44484 22962 44540
rect 23130 44484 23238 44540
rect 23406 44484 23514 44540
rect 23682 44484 23790 44540
rect 23958 44484 24066 44540
rect 24234 44484 24342 44540
rect 24510 44484 24618 44540
rect 24786 44484 24894 44540
rect 25062 44484 25170 44540
rect 25338 44484 25446 44540
rect 25614 44484 25648 44540
rect 20 216 25648 44484
rect 20 54 54 216
rect 222 54 330 216
rect 498 54 606 216
rect 774 54 882 216
rect 1050 54 1158 216
rect 1326 54 1434 216
rect 1602 54 1710 216
rect 1878 54 1986 216
rect 2154 54 2262 216
rect 2430 54 2538 216
rect 2706 54 2814 216
rect 2982 54 3090 216
rect 3258 54 3366 216
rect 3534 54 3642 216
rect 3810 54 3918 216
rect 4086 54 4194 216
rect 4362 54 4470 216
rect 4638 54 4746 216
rect 4914 54 5022 216
rect 5190 54 5298 216
rect 5466 54 5574 216
rect 5742 54 5850 216
rect 6018 54 6126 216
rect 6294 54 6402 216
rect 6570 54 6678 216
rect 6846 54 6954 216
rect 7122 54 7230 216
rect 7398 54 7506 216
rect 7674 54 7782 216
rect 7950 54 8058 216
rect 8226 54 8334 216
rect 8502 54 8610 216
rect 8778 54 8886 216
rect 9054 54 9162 216
rect 9330 54 9438 216
rect 9606 54 9714 216
rect 9882 54 9990 216
rect 10158 54 10266 216
rect 10434 54 10542 216
rect 10710 54 10818 216
rect 10986 54 11094 216
rect 11262 54 11370 216
rect 11538 54 11646 216
rect 11814 54 11922 216
rect 12090 54 12198 216
rect 12366 54 12474 216
rect 12642 54 12750 216
rect 12918 54 13026 216
rect 13194 54 13302 216
rect 13470 54 13578 216
rect 13746 54 13854 216
rect 14022 54 14130 216
rect 14298 54 14406 216
rect 14574 54 14682 216
rect 14850 54 14958 216
rect 15126 54 15234 216
rect 15402 54 15510 216
rect 15678 54 15786 216
rect 15954 54 16062 216
rect 16230 54 16338 216
rect 16506 54 16614 216
rect 16782 54 16890 216
rect 17058 54 17166 216
rect 17334 54 17442 216
rect 17610 54 17718 216
rect 17886 54 17994 216
rect 18162 54 18270 216
rect 18438 54 18546 216
rect 18714 54 18822 216
rect 18990 54 19098 216
rect 19266 54 19374 216
rect 19542 54 19650 216
rect 19818 54 19926 216
rect 20094 54 20202 216
rect 20370 54 20478 216
rect 20646 54 20754 216
rect 20922 54 21030 216
rect 21198 54 21306 216
rect 21474 54 21582 216
rect 21750 54 21858 216
rect 22026 54 22134 216
rect 22302 54 22410 216
rect 22578 54 22686 216
rect 22854 54 22962 216
rect 23130 54 23238 216
rect 23406 54 23514 216
rect 23682 54 23790 216
rect 23958 54 24066 216
rect 24234 54 24342 216
rect 24510 54 24618 216
rect 24786 54 24894 216
rect 25062 54 25170 216
rect 25338 54 25446 216
rect 25614 54 25648 216
<< metal3 >>
rect 25540 43528 26000 43648
rect 25540 42984 26000 43104
rect 25540 42440 26000 42560
rect 25540 41896 26000 42016
rect 25540 41352 26000 41472
rect 25540 40808 26000 40928
rect 25540 40264 26000 40384
rect 25540 39720 26000 39840
rect -300 39448 160 39568
rect -300 39176 160 39296
rect 25540 39176 26000 39296
rect -300 38904 160 39024
rect -300 38632 160 38752
rect 25540 38632 26000 38752
rect -300 38360 160 38480
rect -300 38088 160 38208
rect 25540 38088 26000 38208
rect -300 37816 160 37936
rect -300 37544 160 37664
rect 25540 37544 26000 37664
rect -300 37272 160 37392
rect -300 37000 160 37120
rect 25540 37000 26000 37120
rect -300 36728 160 36848
rect -300 36456 160 36576
rect 25540 36456 26000 36576
rect -300 36184 160 36304
rect -300 35912 160 36032
rect 25540 35912 26000 36032
rect -300 35640 160 35760
rect -300 35368 160 35488
rect 25540 35368 26000 35488
rect -300 35096 160 35216
rect -300 34824 160 34944
rect 25540 34824 26000 34944
rect -300 34552 160 34672
rect -300 34280 160 34400
rect 25540 34280 26000 34400
rect -300 34008 160 34128
rect -300 33736 160 33856
rect 25540 33736 26000 33856
rect -300 33464 160 33584
rect -300 33192 160 33312
rect 25540 33192 26000 33312
rect -300 32920 160 33040
rect -300 32648 160 32768
rect 25540 32648 26000 32768
rect -300 32376 160 32496
rect -300 32104 160 32224
rect 25540 32104 26000 32224
rect -300 31832 160 31952
rect -300 31560 160 31680
rect 25540 31560 26000 31680
rect -300 31288 160 31408
rect -300 31016 160 31136
rect 25540 31016 26000 31136
rect -300 30744 160 30864
rect -300 30472 160 30592
rect 25540 30472 26000 30592
rect -300 30200 160 30320
rect -300 29928 160 30048
rect 25540 29928 26000 30048
rect -300 29656 160 29776
rect -300 29384 160 29504
rect 25540 29384 26000 29504
rect -300 29112 160 29232
rect -300 28840 160 28960
rect 25540 28840 26000 28960
rect -300 28568 160 28688
rect -300 28296 160 28416
rect 25540 28296 26000 28416
rect -300 28024 160 28144
rect -300 27752 160 27872
rect 25540 27752 26000 27872
rect -300 27480 160 27600
rect -300 27208 160 27328
rect 25540 27208 26000 27328
rect -300 26936 160 27056
rect -300 26664 160 26784
rect 25540 26664 26000 26784
rect -300 26392 160 26512
rect -300 26120 160 26240
rect 25540 26120 26000 26240
rect -300 25848 160 25968
rect -300 25576 160 25696
rect 25540 25576 26000 25696
rect -300 25304 160 25424
rect -300 25032 160 25152
rect 25540 25032 26000 25152
rect -300 24760 160 24880
rect -300 24488 160 24608
rect 25540 24488 26000 24608
rect -300 24216 160 24336
rect -300 23944 160 24064
rect 25540 23944 26000 24064
rect -300 23672 160 23792
rect -300 23400 160 23520
rect 25540 23400 26000 23520
rect -300 23128 160 23248
rect -300 22856 160 22976
rect 25540 22856 26000 22976
rect -300 22584 160 22704
rect -300 22312 160 22432
rect 25540 22312 26000 22432
rect -300 22040 160 22160
rect -300 21768 160 21888
rect 25540 21768 26000 21888
rect -300 21496 160 21616
rect -300 21224 160 21344
rect 25540 21224 26000 21344
rect -300 20952 160 21072
rect -300 20680 160 20800
rect 25540 20680 26000 20800
rect -300 20408 160 20528
rect -300 20136 160 20256
rect 25540 20136 26000 20256
rect -300 19864 160 19984
rect -300 19592 160 19712
rect 25540 19592 26000 19712
rect -300 19320 160 19440
rect -300 19048 160 19168
rect 25540 19048 26000 19168
rect -300 18776 160 18896
rect -300 18504 160 18624
rect 25540 18504 26000 18624
rect -300 18232 160 18352
rect -300 17960 160 18080
rect 25540 17960 26000 18080
rect -300 17688 160 17808
rect -300 17416 160 17536
rect 25540 17416 26000 17536
rect -300 17144 160 17264
rect -300 16872 160 16992
rect 25540 16872 26000 16992
rect -300 16600 160 16720
rect -300 16328 160 16448
rect 25540 16328 26000 16448
rect -300 16056 160 16176
rect -300 15784 160 15904
rect 25540 15784 26000 15904
rect -300 15512 160 15632
rect -300 15240 160 15360
rect 25540 15240 26000 15360
rect -300 14968 160 15088
rect -300 14696 160 14816
rect 25540 14696 26000 14816
rect -300 14424 160 14544
rect -300 14152 160 14272
rect 25540 14152 26000 14272
rect -300 13880 160 14000
rect -300 13608 160 13728
rect 25540 13608 26000 13728
rect -300 13336 160 13456
rect -300 13064 160 13184
rect 25540 13064 26000 13184
rect -300 12792 160 12912
rect -300 12520 160 12640
rect 25540 12520 26000 12640
rect -300 12248 160 12368
rect -300 11976 160 12096
rect 25540 11976 26000 12096
rect -300 11704 160 11824
rect -300 11432 160 11552
rect 25540 11432 26000 11552
rect -300 11160 160 11280
rect -300 10888 160 11008
rect 25540 10888 26000 11008
rect -300 10616 160 10736
rect -300 10344 160 10464
rect 25540 10344 26000 10464
rect -300 10072 160 10192
rect -300 9800 160 9920
rect 25540 9800 26000 9920
rect -300 9528 160 9648
rect -300 9256 160 9376
rect 25540 9256 26000 9376
rect -300 8984 160 9104
rect -300 8712 160 8832
rect 25540 8712 26000 8832
rect -300 8440 160 8560
rect -300 8168 160 8288
rect 25540 8168 26000 8288
rect -300 7896 160 8016
rect -300 7624 160 7744
rect 25540 7624 26000 7744
rect -300 7352 160 7472
rect -300 7080 160 7200
rect 25540 7080 26000 7200
rect -300 6808 160 6928
rect -300 6536 160 6656
rect 25540 6536 26000 6656
rect -300 6264 160 6384
rect -300 5992 160 6112
rect 25540 5992 26000 6112
rect -300 5720 160 5840
rect -300 5448 160 5568
rect 25540 5448 26000 5568
rect -300 5176 160 5296
rect -300 4904 160 5024
rect 25540 4904 26000 5024
rect 25540 4360 26000 4480
rect 25540 3816 26000 3936
rect 25540 3272 26000 3392
rect 25540 2728 26000 2848
rect 25540 2184 26000 2304
rect 25540 1640 26000 1760
rect 25540 1096 26000 1216
rect 25540 552 26000 672
<< obsm3 >>
rect 160 43728 25540 43757
rect 160 43448 25460 43728
rect 160 43184 25540 43448
rect 160 42904 25460 43184
rect 160 42640 25540 42904
rect 160 42360 25460 42640
rect 160 42096 25540 42360
rect 160 41816 25460 42096
rect 160 41552 25540 41816
rect 160 41272 25460 41552
rect 160 41008 25540 41272
rect 160 40728 25460 41008
rect 160 40464 25540 40728
rect 160 40184 25460 40464
rect 160 39920 25540 40184
rect 160 39648 25460 39920
rect 240 39640 25460 39648
rect 240 39376 25540 39640
rect 240 39096 25460 39376
rect 240 38832 25540 39096
rect 240 38552 25460 38832
rect 240 38288 25540 38552
rect 240 38008 25460 38288
rect 240 37744 25540 38008
rect 240 37464 25460 37744
rect 240 37200 25540 37464
rect 240 36920 25460 37200
rect 240 36656 25540 36920
rect 240 36376 25460 36656
rect 240 36112 25540 36376
rect 240 35832 25460 36112
rect 240 35568 25540 35832
rect 240 35288 25460 35568
rect 240 35024 25540 35288
rect 240 34744 25460 35024
rect 240 34480 25540 34744
rect 240 34200 25460 34480
rect 240 33936 25540 34200
rect 240 33656 25460 33936
rect 240 33392 25540 33656
rect 240 33112 25460 33392
rect 240 32848 25540 33112
rect 240 32568 25460 32848
rect 240 32304 25540 32568
rect 240 32024 25460 32304
rect 240 31760 25540 32024
rect 240 31480 25460 31760
rect 240 31216 25540 31480
rect 240 30936 25460 31216
rect 240 30672 25540 30936
rect 240 30392 25460 30672
rect 240 30128 25540 30392
rect 240 29848 25460 30128
rect 240 29584 25540 29848
rect 240 29304 25460 29584
rect 240 29040 25540 29304
rect 240 28760 25460 29040
rect 240 28496 25540 28760
rect 240 28216 25460 28496
rect 240 27952 25540 28216
rect 240 27672 25460 27952
rect 240 27408 25540 27672
rect 240 27128 25460 27408
rect 240 26864 25540 27128
rect 240 26584 25460 26864
rect 240 26320 25540 26584
rect 240 26040 25460 26320
rect 240 25776 25540 26040
rect 240 25496 25460 25776
rect 240 25232 25540 25496
rect 240 24952 25460 25232
rect 240 24688 25540 24952
rect 240 24408 25460 24688
rect 240 24144 25540 24408
rect 240 23864 25460 24144
rect 240 23600 25540 23864
rect 240 23320 25460 23600
rect 240 23056 25540 23320
rect 240 22776 25460 23056
rect 240 22512 25540 22776
rect 240 22232 25460 22512
rect 240 21968 25540 22232
rect 240 21688 25460 21968
rect 240 21424 25540 21688
rect 240 21144 25460 21424
rect 240 20880 25540 21144
rect 240 20600 25460 20880
rect 240 20336 25540 20600
rect 240 20056 25460 20336
rect 240 19792 25540 20056
rect 240 19512 25460 19792
rect 240 19248 25540 19512
rect 240 18968 25460 19248
rect 240 18704 25540 18968
rect 240 18424 25460 18704
rect 240 18160 25540 18424
rect 240 17880 25460 18160
rect 240 17616 25540 17880
rect 240 17336 25460 17616
rect 240 17072 25540 17336
rect 240 16792 25460 17072
rect 240 16528 25540 16792
rect 240 16248 25460 16528
rect 240 15984 25540 16248
rect 240 15704 25460 15984
rect 240 15440 25540 15704
rect 240 15160 25460 15440
rect 240 14896 25540 15160
rect 240 14616 25460 14896
rect 240 14352 25540 14616
rect 240 14072 25460 14352
rect 240 13808 25540 14072
rect 240 13528 25460 13808
rect 240 13264 25540 13528
rect 240 12984 25460 13264
rect 240 12720 25540 12984
rect 240 12440 25460 12720
rect 240 12176 25540 12440
rect 240 11896 25460 12176
rect 240 11632 25540 11896
rect 240 11352 25460 11632
rect 240 11088 25540 11352
rect 240 10808 25460 11088
rect 240 10544 25540 10808
rect 240 10264 25460 10544
rect 240 10000 25540 10264
rect 240 9720 25460 10000
rect 240 9456 25540 9720
rect 240 9176 25460 9456
rect 240 8912 25540 9176
rect 240 8632 25460 8912
rect 240 8368 25540 8632
rect 240 8088 25460 8368
rect 240 7824 25540 8088
rect 240 7544 25460 7824
rect 240 7280 25540 7544
rect 240 7000 25460 7280
rect 240 6736 25540 7000
rect 240 6456 25460 6736
rect 240 6192 25540 6456
rect 240 5912 25460 6192
rect 240 5648 25540 5912
rect 240 5368 25460 5648
rect 240 5104 25540 5368
rect 240 4824 25460 5104
rect 160 4560 25540 4824
rect 160 4280 25460 4560
rect 160 4016 25540 4280
rect 160 3736 25460 4016
rect 160 3472 25540 3736
rect 160 3192 25460 3472
rect 160 2928 25540 3192
rect 160 2648 25460 2928
rect 160 2384 25540 2648
rect 160 2104 25460 2384
rect 160 1840 25540 2104
rect 160 1560 25460 1840
rect 160 1296 25540 1560
rect 160 1016 25460 1296
rect 160 752 25540 1016
rect 160 472 25460 752
rect 160 443 25540 472
<< metal4 >>
rect 3876 1040 4196 43568
rect 6808 1040 7128 43568
rect 9741 1040 10061 43568
rect 12673 1040 12993 43568
rect 15606 1040 15926 43568
rect 18538 1040 18858 43568
rect 21471 1040 21791 43568
rect 24403 1040 24723 43568
<< obsm4 >>
rect 611 960 3796 43213
rect 4276 960 6728 43213
rect 7208 960 9661 43213
rect 10141 960 12593 43213
rect 13073 960 15526 43213
rect 16006 960 18458 43213
rect 18938 960 21391 43213
rect 21871 960 22757 43213
rect 611 443 22757 960
<< labels >>
rlabel metal3 s 25540 9256 26000 9376 6 Config_accessC_bit0
port 1 nsew signal output
rlabel metal3 s 25540 9800 26000 9920 6 Config_accessC_bit1
port 2 nsew signal output
rlabel metal3 s 25540 10344 26000 10464 6 Config_accessC_bit2
port 3 nsew signal output
rlabel metal3 s 25540 10888 26000 11008 6 Config_accessC_bit3
port 4 nsew signal output
rlabel metal3 s -300 17960 160 18080 4 E1END[0]
port 5 nsew signal input
rlabel metal3 s -300 18232 160 18352 4 E1END[1]
port 6 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 E1END[2]
port 7 nsew signal input
rlabel metal3 s -300 18776 160 18896 4 E1END[3]
port 8 nsew signal input
rlabel metal3 s -300 21224 160 21344 4 E2END[0]
port 9 nsew signal input
rlabel metal3 s -300 21496 160 21616 4 E2END[1]
port 10 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 E2END[2]
port 11 nsew signal input
rlabel metal3 s -300 22040 160 22160 4 E2END[3]
port 12 nsew signal input
rlabel metal3 s -300 22312 160 22432 4 E2END[4]
port 13 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 E2END[5]
port 14 nsew signal input
rlabel metal3 s -300 22856 160 22976 4 E2END[6]
port 15 nsew signal input
rlabel metal3 s -300 23128 160 23248 4 E2END[7]
port 16 nsew signal input
rlabel metal3 s -300 19048 160 19168 4 E2MID[0]
port 17 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 E2MID[1]
port 18 nsew signal input
rlabel metal3 s -300 19592 160 19712 4 E2MID[2]
port 19 nsew signal input
rlabel metal3 s -300 19864 160 19984 4 E2MID[3]
port 20 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 E2MID[4]
port 21 nsew signal input
rlabel metal3 s -300 20408 160 20528 4 E2MID[5]
port 22 nsew signal input
rlabel metal3 s -300 20680 160 20800 4 E2MID[6]
port 23 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 E2MID[7]
port 24 nsew signal input
rlabel metal3 s -300 27752 160 27872 4 E6END[0]
port 25 nsew signal input
rlabel metal3 s -300 30472 160 30592 4 E6END[10]
port 26 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 E6END[11]
port 27 nsew signal input
rlabel metal3 s -300 28024 160 28144 4 E6END[1]
port 28 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 E6END[2]
port 29 nsew signal input
rlabel metal3 s -300 28568 160 28688 4 E6END[3]
port 30 nsew signal input
rlabel metal3 s -300 28840 160 28960 4 E6END[4]
port 31 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 E6END[5]
port 32 nsew signal input
rlabel metal3 s -300 29384 160 29504 4 E6END[6]
port 33 nsew signal input
rlabel metal3 s -300 29656 160 29776 4 E6END[7]
port 34 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 E6END[8]
port 35 nsew signal input
rlabel metal3 s -300 30200 160 30320 4 E6END[9]
port 36 nsew signal input
rlabel metal3 s -300 23400 160 23520 4 EE4END[0]
port 37 nsew signal input
rlabel metal3 s -300 26120 160 26240 4 EE4END[10]
port 38 nsew signal input
rlabel metal3 s -300 26392 160 26512 4 EE4END[11]
port 39 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 EE4END[12]
port 40 nsew signal input
rlabel metal3 s -300 26936 160 27056 4 EE4END[13]
port 41 nsew signal input
rlabel metal3 s -300 27208 160 27328 4 EE4END[14]
port 42 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 EE4END[15]
port 43 nsew signal input
rlabel metal3 s -300 23672 160 23792 4 EE4END[1]
port 44 nsew signal input
rlabel metal3 s -300 23944 160 24064 4 EE4END[2]
port 45 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 EE4END[3]
port 46 nsew signal input
rlabel metal3 s -300 24488 160 24608 4 EE4END[4]
port 47 nsew signal input
rlabel metal3 s -300 24760 160 24880 4 EE4END[5]
port 48 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 EE4END[6]
port 49 nsew signal input
rlabel metal3 s -300 25304 160 25424 4 EE4END[7]
port 50 nsew signal input
rlabel metal3 s -300 25576 160 25696 4 EE4END[8]
port 51 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 EE4END[9]
port 52 nsew signal input
rlabel metal3 s 25540 15784 26000 15904 6 FAB2RAM_A0_O0
port 53 nsew signal output
rlabel metal3 s 25540 16328 26000 16448 6 FAB2RAM_A0_O1
port 54 nsew signal output
rlabel metal3 s 25540 16872 26000 16992 6 FAB2RAM_A0_O2
port 55 nsew signal output
rlabel metal3 s 25540 17416 26000 17536 6 FAB2RAM_A0_O3
port 56 nsew signal output
rlabel metal3 s 25540 13608 26000 13728 6 FAB2RAM_A1_O0
port 57 nsew signal output
rlabel metal3 s 25540 14152 26000 14272 6 FAB2RAM_A1_O1
port 58 nsew signal output
rlabel metal3 s 25540 14696 26000 14816 6 FAB2RAM_A1_O2
port 59 nsew signal output
rlabel metal3 s 25540 15240 26000 15360 6 FAB2RAM_A1_O3
port 60 nsew signal output
rlabel metal3 s 25540 11432 26000 11552 6 FAB2RAM_C_O0
port 61 nsew signal output
rlabel metal3 s 25540 11976 26000 12096 6 FAB2RAM_C_O1
port 62 nsew signal output
rlabel metal3 s 25540 12520 26000 12640 6 FAB2RAM_C_O2
port 63 nsew signal output
rlabel metal3 s 25540 13064 26000 13184 6 FAB2RAM_C_O3
port 64 nsew signal output
rlabel metal3 s 25540 24488 26000 24608 6 FAB2RAM_D0_O0
port 65 nsew signal output
rlabel metal3 s 25540 25032 26000 25152 6 FAB2RAM_D0_O1
port 66 nsew signal output
rlabel metal3 s 25540 25576 26000 25696 6 FAB2RAM_D0_O2
port 67 nsew signal output
rlabel metal3 s 25540 26120 26000 26240 6 FAB2RAM_D0_O3
port 68 nsew signal output
rlabel metal3 s 25540 22312 26000 22432 6 FAB2RAM_D1_O0
port 69 nsew signal output
rlabel metal3 s 25540 22856 26000 22976 6 FAB2RAM_D1_O1
port 70 nsew signal output
rlabel metal3 s 25540 23400 26000 23520 6 FAB2RAM_D1_O2
port 71 nsew signal output
rlabel metal3 s 25540 23944 26000 24064 6 FAB2RAM_D1_O3
port 72 nsew signal output
rlabel metal3 s 25540 20136 26000 20256 6 FAB2RAM_D2_O0
port 73 nsew signal output
rlabel metal3 s 25540 20680 26000 20800 6 FAB2RAM_D2_O1
port 74 nsew signal output
rlabel metal3 s 25540 21224 26000 21344 6 FAB2RAM_D2_O2
port 75 nsew signal output
rlabel metal3 s 25540 21768 26000 21888 6 FAB2RAM_D2_O3
port 76 nsew signal output
rlabel metal3 s 25540 17960 26000 18080 6 FAB2RAM_D3_O0
port 77 nsew signal output
rlabel metal3 s 25540 18504 26000 18624 6 FAB2RAM_D3_O1
port 78 nsew signal output
rlabel metal3 s 25540 19048 26000 19168 6 FAB2RAM_D3_O2
port 79 nsew signal output
rlabel metal3 s 25540 19592 26000 19712 6 FAB2RAM_D3_O3
port 80 nsew signal output
rlabel metal3 s -300 31016 160 31136 4 FrameData[0]
port 81 nsew signal input
rlabel metal3 s -300 33736 160 33856 4 FrameData[10]
port 82 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 FrameData[11]
port 83 nsew signal input
rlabel metal3 s -300 34280 160 34400 4 FrameData[12]
port 84 nsew signal input
rlabel metal3 s -300 34552 160 34672 4 FrameData[13]
port 85 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 FrameData[14]
port 86 nsew signal input
rlabel metal3 s -300 35096 160 35216 4 FrameData[15]
port 87 nsew signal input
rlabel metal3 s -300 35368 160 35488 4 FrameData[16]
port 88 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 FrameData[17]
port 89 nsew signal input
rlabel metal3 s -300 35912 160 36032 4 FrameData[18]
port 90 nsew signal input
rlabel metal3 s -300 36184 160 36304 4 FrameData[19]
port 91 nsew signal input
rlabel metal3 s -300 31288 160 31408 4 FrameData[1]
port 92 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 FrameData[20]
port 93 nsew signal input
rlabel metal3 s -300 36728 160 36848 4 FrameData[21]
port 94 nsew signal input
rlabel metal3 s -300 37000 160 37120 4 FrameData[22]
port 95 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 FrameData[23]
port 96 nsew signal input
rlabel metal3 s -300 37544 160 37664 4 FrameData[24]
port 97 nsew signal input
rlabel metal3 s -300 37816 160 37936 4 FrameData[25]
port 98 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 FrameData[26]
port 99 nsew signal input
rlabel metal3 s -300 38360 160 38480 4 FrameData[27]
port 100 nsew signal input
rlabel metal3 s -300 38632 160 38752 4 FrameData[28]
port 101 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 FrameData[29]
port 102 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 FrameData[2]
port 103 nsew signal input
rlabel metal3 s -300 39176 160 39296 4 FrameData[30]
port 104 nsew signal input
rlabel metal3 s -300 39448 160 39568 4 FrameData[31]
port 105 nsew signal input
rlabel metal3 s -300 31832 160 31952 4 FrameData[3]
port 106 nsew signal input
rlabel metal3 s -300 32104 160 32224 4 FrameData[4]
port 107 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 FrameData[5]
port 108 nsew signal input
rlabel metal3 s -300 32648 160 32768 4 FrameData[6]
port 109 nsew signal input
rlabel metal3 s -300 32920 160 33040 4 FrameData[7]
port 110 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 FrameData[8]
port 111 nsew signal input
rlabel metal3 s -300 33464 160 33584 4 FrameData[9]
port 112 nsew signal input
rlabel metal3 s 25540 26664 26000 26784 6 FrameData_O[0]
port 113 nsew signal output
rlabel metal3 s 25540 32104 26000 32224 6 FrameData_O[10]
port 114 nsew signal output
rlabel metal3 s 25540 32648 26000 32768 6 FrameData_O[11]
port 115 nsew signal output
rlabel metal3 s 25540 33192 26000 33312 6 FrameData_O[12]
port 116 nsew signal output
rlabel metal3 s 25540 33736 26000 33856 6 FrameData_O[13]
port 117 nsew signal output
rlabel metal3 s 25540 34280 26000 34400 6 FrameData_O[14]
port 118 nsew signal output
rlabel metal3 s 25540 34824 26000 34944 6 FrameData_O[15]
port 119 nsew signal output
rlabel metal3 s 25540 35368 26000 35488 6 FrameData_O[16]
port 120 nsew signal output
rlabel metal3 s 25540 35912 26000 36032 6 FrameData_O[17]
port 121 nsew signal output
rlabel metal3 s 25540 36456 26000 36576 6 FrameData_O[18]
port 122 nsew signal output
rlabel metal3 s 25540 37000 26000 37120 6 FrameData_O[19]
port 123 nsew signal output
rlabel metal3 s 25540 27208 26000 27328 6 FrameData_O[1]
port 124 nsew signal output
rlabel metal3 s 25540 37544 26000 37664 6 FrameData_O[20]
port 125 nsew signal output
rlabel metal3 s 25540 38088 26000 38208 6 FrameData_O[21]
port 126 nsew signal output
rlabel metal3 s 25540 38632 26000 38752 6 FrameData_O[22]
port 127 nsew signal output
rlabel metal3 s 25540 39176 26000 39296 6 FrameData_O[23]
port 128 nsew signal output
rlabel metal3 s 25540 39720 26000 39840 6 FrameData_O[24]
port 129 nsew signal output
rlabel metal3 s 25540 40264 26000 40384 6 FrameData_O[25]
port 130 nsew signal output
rlabel metal3 s 25540 40808 26000 40928 6 FrameData_O[26]
port 131 nsew signal output
rlabel metal3 s 25540 41352 26000 41472 6 FrameData_O[27]
port 132 nsew signal output
rlabel metal3 s 25540 41896 26000 42016 6 FrameData_O[28]
port 133 nsew signal output
rlabel metal3 s 25540 42440 26000 42560 6 FrameData_O[29]
port 134 nsew signal output
rlabel metal3 s 25540 27752 26000 27872 6 FrameData_O[2]
port 135 nsew signal output
rlabel metal3 s 25540 42984 26000 43104 6 FrameData_O[30]
port 136 nsew signal output
rlabel metal3 s 25540 43528 26000 43648 6 FrameData_O[31]
port 137 nsew signal output
rlabel metal3 s 25540 28296 26000 28416 6 FrameData_O[3]
port 138 nsew signal output
rlabel metal3 s 25540 28840 26000 28960 6 FrameData_O[4]
port 139 nsew signal output
rlabel metal3 s 25540 29384 26000 29504 6 FrameData_O[5]
port 140 nsew signal output
rlabel metal3 s 25540 29928 26000 30048 6 FrameData_O[6]
port 141 nsew signal output
rlabel metal3 s 25540 30472 26000 30592 6 FrameData_O[7]
port 142 nsew signal output
rlabel metal3 s 25540 31016 26000 31136 6 FrameData_O[8]
port 143 nsew signal output
rlabel metal3 s 25540 31560 26000 31680 6 FrameData_O[9]
port 144 nsew signal output
rlabel metal2 s 20258 -300 20314 160 8 FrameStrobe[0]
port 145 nsew signal input
rlabel metal2 s 23018 -300 23074 160 8 FrameStrobe[10]
port 146 nsew signal input
rlabel metal2 s 23294 -300 23350 160 8 FrameStrobe[11]
port 147 nsew signal input
rlabel metal2 s 23570 -300 23626 160 8 FrameStrobe[12]
port 148 nsew signal input
rlabel metal2 s 23846 -300 23902 160 8 FrameStrobe[13]
port 149 nsew signal input
rlabel metal2 s 24122 -300 24178 160 8 FrameStrobe[14]
port 150 nsew signal input
rlabel metal2 s 24398 -300 24454 160 8 FrameStrobe[15]
port 151 nsew signal input
rlabel metal2 s 24674 -300 24730 160 8 FrameStrobe[16]
port 152 nsew signal input
rlabel metal2 s 24950 -300 25006 160 8 FrameStrobe[17]
port 153 nsew signal input
rlabel metal2 s 25226 -300 25282 160 8 FrameStrobe[18]
port 154 nsew signal input
rlabel metal2 s 25502 -300 25558 160 8 FrameStrobe[19]
port 155 nsew signal input
rlabel metal2 s 20534 -300 20590 160 8 FrameStrobe[1]
port 156 nsew signal input
rlabel metal2 s 20810 -300 20866 160 8 FrameStrobe[2]
port 157 nsew signal input
rlabel metal2 s 21086 -300 21142 160 8 FrameStrobe[3]
port 158 nsew signal input
rlabel metal2 s 21362 -300 21418 160 8 FrameStrobe[4]
port 159 nsew signal input
rlabel metal2 s 21638 -300 21694 160 8 FrameStrobe[5]
port 160 nsew signal input
rlabel metal2 s 21914 -300 21970 160 8 FrameStrobe[6]
port 161 nsew signal input
rlabel metal2 s 22190 -300 22246 160 8 FrameStrobe[7]
port 162 nsew signal input
rlabel metal2 s 22466 -300 22522 160 8 FrameStrobe[8]
port 163 nsew signal input
rlabel metal2 s 22742 -300 22798 160 8 FrameStrobe[9]
port 164 nsew signal input
rlabel metal2 s 20258 44540 20314 45000 6 FrameStrobe_O[0]
port 165 nsew signal output
rlabel metal2 s 23018 44540 23074 45000 6 FrameStrobe_O[10]
port 166 nsew signal output
rlabel metal2 s 23294 44540 23350 45000 6 FrameStrobe_O[11]
port 167 nsew signal output
rlabel metal2 s 23570 44540 23626 45000 6 FrameStrobe_O[12]
port 168 nsew signal output
rlabel metal2 s 23846 44540 23902 45000 6 FrameStrobe_O[13]
port 169 nsew signal output
rlabel metal2 s 24122 44540 24178 45000 6 FrameStrobe_O[14]
port 170 nsew signal output
rlabel metal2 s 24398 44540 24454 45000 6 FrameStrobe_O[15]
port 171 nsew signal output
rlabel metal2 s 24674 44540 24730 45000 6 FrameStrobe_O[16]
port 172 nsew signal output
rlabel metal2 s 24950 44540 25006 45000 6 FrameStrobe_O[17]
port 173 nsew signal output
rlabel metal2 s 25226 44540 25282 45000 6 FrameStrobe_O[18]
port 174 nsew signal output
rlabel metal2 s 25502 44540 25558 45000 6 FrameStrobe_O[19]
port 175 nsew signal output
rlabel metal2 s 20534 44540 20590 45000 6 FrameStrobe_O[1]
port 176 nsew signal output
rlabel metal2 s 20810 44540 20866 45000 6 FrameStrobe_O[2]
port 177 nsew signal output
rlabel metal2 s 21086 44540 21142 45000 6 FrameStrobe_O[3]
port 178 nsew signal output
rlabel metal2 s 21362 44540 21418 45000 6 FrameStrobe_O[4]
port 179 nsew signal output
rlabel metal2 s 21638 44540 21694 45000 6 FrameStrobe_O[5]
port 180 nsew signal output
rlabel metal2 s 21914 44540 21970 45000 6 FrameStrobe_O[6]
port 181 nsew signal output
rlabel metal2 s 22190 44540 22246 45000 6 FrameStrobe_O[7]
port 182 nsew signal output
rlabel metal2 s 22466 44540 22522 45000 6 FrameStrobe_O[8]
port 183 nsew signal output
rlabel metal2 s 22742 44540 22798 45000 6 FrameStrobe_O[9]
port 184 nsew signal output
rlabel metal2 s 110 44540 166 45000 6 N1BEG[0]
port 185 nsew signal output
rlabel metal2 s 386 44540 442 45000 6 N1BEG[1]
port 186 nsew signal output
rlabel metal2 s 662 44540 718 45000 6 N1BEG[2]
port 187 nsew signal output
rlabel metal2 s 938 44540 994 45000 6 N1BEG[3]
port 188 nsew signal output
rlabel metal2 s 110 -300 166 160 8 N1END[0]
port 189 nsew signal input
rlabel metal2 s 386 -300 442 160 8 N1END[1]
port 190 nsew signal input
rlabel metal2 s 662 -300 718 160 8 N1END[2]
port 191 nsew signal input
rlabel metal2 s 938 -300 994 160 8 N1END[3]
port 192 nsew signal input
rlabel metal2 s 1214 44540 1270 45000 6 N2BEG[0]
port 193 nsew signal output
rlabel metal2 s 1490 44540 1546 45000 6 N2BEG[1]
port 194 nsew signal output
rlabel metal2 s 1766 44540 1822 45000 6 N2BEG[2]
port 195 nsew signal output
rlabel metal2 s 2042 44540 2098 45000 6 N2BEG[3]
port 196 nsew signal output
rlabel metal2 s 2318 44540 2374 45000 6 N2BEG[4]
port 197 nsew signal output
rlabel metal2 s 2594 44540 2650 45000 6 N2BEG[5]
port 198 nsew signal output
rlabel metal2 s 2870 44540 2926 45000 6 N2BEG[6]
port 199 nsew signal output
rlabel metal2 s 3146 44540 3202 45000 6 N2BEG[7]
port 200 nsew signal output
rlabel metal2 s 3422 44540 3478 45000 6 N2BEGb[0]
port 201 nsew signal output
rlabel metal2 s 3698 44540 3754 45000 6 N2BEGb[1]
port 202 nsew signal output
rlabel metal2 s 3974 44540 4030 45000 6 N2BEGb[2]
port 203 nsew signal output
rlabel metal2 s 4250 44540 4306 45000 6 N2BEGb[3]
port 204 nsew signal output
rlabel metal2 s 4526 44540 4582 45000 6 N2BEGb[4]
port 205 nsew signal output
rlabel metal2 s 4802 44540 4858 45000 6 N2BEGb[5]
port 206 nsew signal output
rlabel metal2 s 5078 44540 5134 45000 6 N2BEGb[6]
port 207 nsew signal output
rlabel metal2 s 5354 44540 5410 45000 6 N2BEGb[7]
port 208 nsew signal output
rlabel metal2 s 3422 -300 3478 160 8 N2END[0]
port 209 nsew signal input
rlabel metal2 s 3698 -300 3754 160 8 N2END[1]
port 210 nsew signal input
rlabel metal2 s 3974 -300 4030 160 8 N2END[2]
port 211 nsew signal input
rlabel metal2 s 4250 -300 4306 160 8 N2END[3]
port 212 nsew signal input
rlabel metal2 s 4526 -300 4582 160 8 N2END[4]
port 213 nsew signal input
rlabel metal2 s 4802 -300 4858 160 8 N2END[5]
port 214 nsew signal input
rlabel metal2 s 5078 -300 5134 160 8 N2END[6]
port 215 nsew signal input
rlabel metal2 s 5354 -300 5410 160 8 N2END[7]
port 216 nsew signal input
rlabel metal2 s 1214 -300 1270 160 8 N2MID[0]
port 217 nsew signal input
rlabel metal2 s 1490 -300 1546 160 8 N2MID[1]
port 218 nsew signal input
rlabel metal2 s 1766 -300 1822 160 8 N2MID[2]
port 219 nsew signal input
rlabel metal2 s 2042 -300 2098 160 8 N2MID[3]
port 220 nsew signal input
rlabel metal2 s 2318 -300 2374 160 8 N2MID[4]
port 221 nsew signal input
rlabel metal2 s 2594 -300 2650 160 8 N2MID[5]
port 222 nsew signal input
rlabel metal2 s 2870 -300 2926 160 8 N2MID[6]
port 223 nsew signal input
rlabel metal2 s 3146 -300 3202 160 8 N2MID[7]
port 224 nsew signal input
rlabel metal2 s 5630 44540 5686 45000 6 N4BEG[0]
port 225 nsew signal output
rlabel metal2 s 8390 44540 8446 45000 6 N4BEG[10]
port 226 nsew signal output
rlabel metal2 s 8666 44540 8722 45000 6 N4BEG[11]
port 227 nsew signal output
rlabel metal2 s 8942 44540 8998 45000 6 N4BEG[12]
port 228 nsew signal output
rlabel metal2 s 9218 44540 9274 45000 6 N4BEG[13]
port 229 nsew signal output
rlabel metal2 s 9494 44540 9550 45000 6 N4BEG[14]
port 230 nsew signal output
rlabel metal2 s 9770 44540 9826 45000 6 N4BEG[15]
port 231 nsew signal output
rlabel metal2 s 5906 44540 5962 45000 6 N4BEG[1]
port 232 nsew signal output
rlabel metal2 s 6182 44540 6238 45000 6 N4BEG[2]
port 233 nsew signal output
rlabel metal2 s 6458 44540 6514 45000 6 N4BEG[3]
port 234 nsew signal output
rlabel metal2 s 6734 44540 6790 45000 6 N4BEG[4]
port 235 nsew signal output
rlabel metal2 s 7010 44540 7066 45000 6 N4BEG[5]
port 236 nsew signal output
rlabel metal2 s 7286 44540 7342 45000 6 N4BEG[6]
port 237 nsew signal output
rlabel metal2 s 7562 44540 7618 45000 6 N4BEG[7]
port 238 nsew signal output
rlabel metal2 s 7838 44540 7894 45000 6 N4BEG[8]
port 239 nsew signal output
rlabel metal2 s 8114 44540 8170 45000 6 N4BEG[9]
port 240 nsew signal output
rlabel metal2 s 5630 -300 5686 160 8 N4END[0]
port 241 nsew signal input
rlabel metal2 s 8390 -300 8446 160 8 N4END[10]
port 242 nsew signal input
rlabel metal2 s 8666 -300 8722 160 8 N4END[11]
port 243 nsew signal input
rlabel metal2 s 8942 -300 8998 160 8 N4END[12]
port 244 nsew signal input
rlabel metal2 s 9218 -300 9274 160 8 N4END[13]
port 245 nsew signal input
rlabel metal2 s 9494 -300 9550 160 8 N4END[14]
port 246 nsew signal input
rlabel metal2 s 9770 -300 9826 160 8 N4END[15]
port 247 nsew signal input
rlabel metal2 s 5906 -300 5962 160 8 N4END[1]
port 248 nsew signal input
rlabel metal2 s 6182 -300 6238 160 8 N4END[2]
port 249 nsew signal input
rlabel metal2 s 6458 -300 6514 160 8 N4END[3]
port 250 nsew signal input
rlabel metal2 s 6734 -300 6790 160 8 N4END[4]
port 251 nsew signal input
rlabel metal2 s 7010 -300 7066 160 8 N4END[5]
port 252 nsew signal input
rlabel metal2 s 7286 -300 7342 160 8 N4END[6]
port 253 nsew signal input
rlabel metal2 s 7562 -300 7618 160 8 N4END[7]
port 254 nsew signal input
rlabel metal2 s 7838 -300 7894 160 8 N4END[8]
port 255 nsew signal input
rlabel metal2 s 8114 -300 8170 160 8 N4END[9]
port 256 nsew signal input
rlabel metal3 s 25540 7080 26000 7200 6 RAM2FAB_D0_I0
port 257 nsew signal input
rlabel metal3 s 25540 7624 26000 7744 6 RAM2FAB_D0_I1
port 258 nsew signal input
rlabel metal3 s 25540 8168 26000 8288 6 RAM2FAB_D0_I2
port 259 nsew signal input
rlabel metal3 s 25540 8712 26000 8832 6 RAM2FAB_D0_I3
port 260 nsew signal input
rlabel metal3 s 25540 4904 26000 5024 6 RAM2FAB_D1_I0
port 261 nsew signal input
rlabel metal3 s 25540 5448 26000 5568 6 RAM2FAB_D1_I1
port 262 nsew signal input
rlabel metal3 s 25540 5992 26000 6112 6 RAM2FAB_D1_I2
port 263 nsew signal input
rlabel metal3 s 25540 6536 26000 6656 6 RAM2FAB_D1_I3
port 264 nsew signal input
rlabel metal3 s 25540 2728 26000 2848 6 RAM2FAB_D2_I0
port 265 nsew signal input
rlabel metal3 s 25540 3272 26000 3392 6 RAM2FAB_D2_I1
port 266 nsew signal input
rlabel metal3 s 25540 3816 26000 3936 6 RAM2FAB_D2_I2
port 267 nsew signal input
rlabel metal3 s 25540 4360 26000 4480 6 RAM2FAB_D2_I3
port 268 nsew signal input
rlabel metal3 s 25540 552 26000 672 6 RAM2FAB_D3_I0
port 269 nsew signal input
rlabel metal3 s 25540 1096 26000 1216 6 RAM2FAB_D3_I1
port 270 nsew signal input
rlabel metal3 s 25540 1640 26000 1760 6 RAM2FAB_D3_I2
port 271 nsew signal input
rlabel metal3 s 25540 2184 26000 2304 6 RAM2FAB_D3_I3
port 272 nsew signal input
rlabel metal2 s 10046 -300 10102 160 8 S1BEG[0]
port 273 nsew signal output
rlabel metal2 s 10322 -300 10378 160 8 S1BEG[1]
port 274 nsew signal output
rlabel metal2 s 10598 -300 10654 160 8 S1BEG[2]
port 275 nsew signal output
rlabel metal2 s 10874 -300 10930 160 8 S1BEG[3]
port 276 nsew signal output
rlabel metal2 s 10046 44540 10102 45000 6 S1END[0]
port 277 nsew signal input
rlabel metal2 s 10322 44540 10378 45000 6 S1END[1]
port 278 nsew signal input
rlabel metal2 s 10598 44540 10654 45000 6 S1END[2]
port 279 nsew signal input
rlabel metal2 s 10874 44540 10930 45000 6 S1END[3]
port 280 nsew signal input
rlabel metal2 s 13358 -300 13414 160 8 S2BEG[0]
port 281 nsew signal output
rlabel metal2 s 13634 -300 13690 160 8 S2BEG[1]
port 282 nsew signal output
rlabel metal2 s 13910 -300 13966 160 8 S2BEG[2]
port 283 nsew signal output
rlabel metal2 s 14186 -300 14242 160 8 S2BEG[3]
port 284 nsew signal output
rlabel metal2 s 14462 -300 14518 160 8 S2BEG[4]
port 285 nsew signal output
rlabel metal2 s 14738 -300 14794 160 8 S2BEG[5]
port 286 nsew signal output
rlabel metal2 s 15014 -300 15070 160 8 S2BEG[6]
port 287 nsew signal output
rlabel metal2 s 15290 -300 15346 160 8 S2BEG[7]
port 288 nsew signal output
rlabel metal2 s 11150 -300 11206 160 8 S2BEGb[0]
port 289 nsew signal output
rlabel metal2 s 11426 -300 11482 160 8 S2BEGb[1]
port 290 nsew signal output
rlabel metal2 s 11702 -300 11758 160 8 S2BEGb[2]
port 291 nsew signal output
rlabel metal2 s 11978 -300 12034 160 8 S2BEGb[3]
port 292 nsew signal output
rlabel metal2 s 12254 -300 12310 160 8 S2BEGb[4]
port 293 nsew signal output
rlabel metal2 s 12530 -300 12586 160 8 S2BEGb[5]
port 294 nsew signal output
rlabel metal2 s 12806 -300 12862 160 8 S2BEGb[6]
port 295 nsew signal output
rlabel metal2 s 13082 -300 13138 160 8 S2BEGb[7]
port 296 nsew signal output
rlabel metal2 s 11150 44540 11206 45000 6 S2END[0]
port 297 nsew signal input
rlabel metal2 s 11426 44540 11482 45000 6 S2END[1]
port 298 nsew signal input
rlabel metal2 s 11702 44540 11758 45000 6 S2END[2]
port 299 nsew signal input
rlabel metal2 s 11978 44540 12034 45000 6 S2END[3]
port 300 nsew signal input
rlabel metal2 s 12254 44540 12310 45000 6 S2END[4]
port 301 nsew signal input
rlabel metal2 s 12530 44540 12586 45000 6 S2END[5]
port 302 nsew signal input
rlabel metal2 s 12806 44540 12862 45000 6 S2END[6]
port 303 nsew signal input
rlabel metal2 s 13082 44540 13138 45000 6 S2END[7]
port 304 nsew signal input
rlabel metal2 s 13358 44540 13414 45000 6 S2MID[0]
port 305 nsew signal input
rlabel metal2 s 13634 44540 13690 45000 6 S2MID[1]
port 306 nsew signal input
rlabel metal2 s 13910 44540 13966 45000 6 S2MID[2]
port 307 nsew signal input
rlabel metal2 s 14186 44540 14242 45000 6 S2MID[3]
port 308 nsew signal input
rlabel metal2 s 14462 44540 14518 45000 6 S2MID[4]
port 309 nsew signal input
rlabel metal2 s 14738 44540 14794 45000 6 S2MID[5]
port 310 nsew signal input
rlabel metal2 s 15014 44540 15070 45000 6 S2MID[6]
port 311 nsew signal input
rlabel metal2 s 15290 44540 15346 45000 6 S2MID[7]
port 312 nsew signal input
rlabel metal2 s 15566 -300 15622 160 8 S4BEG[0]
port 313 nsew signal output
rlabel metal2 s 18326 -300 18382 160 8 S4BEG[10]
port 314 nsew signal output
rlabel metal2 s 18602 -300 18658 160 8 S4BEG[11]
port 315 nsew signal output
rlabel metal2 s 18878 -300 18934 160 8 S4BEG[12]
port 316 nsew signal output
rlabel metal2 s 19154 -300 19210 160 8 S4BEG[13]
port 317 nsew signal output
rlabel metal2 s 19430 -300 19486 160 8 S4BEG[14]
port 318 nsew signal output
rlabel metal2 s 19706 -300 19762 160 8 S4BEG[15]
port 319 nsew signal output
rlabel metal2 s 15842 -300 15898 160 8 S4BEG[1]
port 320 nsew signal output
rlabel metal2 s 16118 -300 16174 160 8 S4BEG[2]
port 321 nsew signal output
rlabel metal2 s 16394 -300 16450 160 8 S4BEG[3]
port 322 nsew signal output
rlabel metal2 s 16670 -300 16726 160 8 S4BEG[4]
port 323 nsew signal output
rlabel metal2 s 16946 -300 17002 160 8 S4BEG[5]
port 324 nsew signal output
rlabel metal2 s 17222 -300 17278 160 8 S4BEG[6]
port 325 nsew signal output
rlabel metal2 s 17498 -300 17554 160 8 S4BEG[7]
port 326 nsew signal output
rlabel metal2 s 17774 -300 17830 160 8 S4BEG[8]
port 327 nsew signal output
rlabel metal2 s 18050 -300 18106 160 8 S4BEG[9]
port 328 nsew signal output
rlabel metal2 s 15566 44540 15622 45000 6 S4END[0]
port 329 nsew signal input
rlabel metal2 s 18326 44540 18382 45000 6 S4END[10]
port 330 nsew signal input
rlabel metal2 s 18602 44540 18658 45000 6 S4END[11]
port 331 nsew signal input
rlabel metal2 s 18878 44540 18934 45000 6 S4END[12]
port 332 nsew signal input
rlabel metal2 s 19154 44540 19210 45000 6 S4END[13]
port 333 nsew signal input
rlabel metal2 s 19430 44540 19486 45000 6 S4END[14]
port 334 nsew signal input
rlabel metal2 s 19706 44540 19762 45000 6 S4END[15]
port 335 nsew signal input
rlabel metal2 s 15842 44540 15898 45000 6 S4END[1]
port 336 nsew signal input
rlabel metal2 s 16118 44540 16174 45000 6 S4END[2]
port 337 nsew signal input
rlabel metal2 s 16394 44540 16450 45000 6 S4END[3]
port 338 nsew signal input
rlabel metal2 s 16670 44540 16726 45000 6 S4END[4]
port 339 nsew signal input
rlabel metal2 s 16946 44540 17002 45000 6 S4END[5]
port 340 nsew signal input
rlabel metal2 s 17222 44540 17278 45000 6 S4END[6]
port 341 nsew signal input
rlabel metal2 s 17498 44540 17554 45000 6 S4END[7]
port 342 nsew signal input
rlabel metal2 s 17774 44540 17830 45000 6 S4END[8]
port 343 nsew signal input
rlabel metal2 s 18050 44540 18106 45000 6 S4END[9]
port 344 nsew signal input
rlabel metal2 s 19982 -300 20038 160 8 UserCLK
port 345 nsew signal input
rlabel metal2 s 19982 44540 20038 45000 6 UserCLKo
port 346 nsew signal output
rlabel metal4 s 6808 1040 7128 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 12673 1040 12993 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 18538 1040 18858 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 24403 1040 24723 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 3876 1040 4196 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 9741 1040 10061 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 15606 1040 15926 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 21471 1040 21791 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal3 s -300 4904 160 5024 4 W1BEG[0]
port 349 nsew signal output
rlabel metal3 s -300 5176 160 5296 4 W1BEG[1]
port 350 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 W1BEG[2]
port 351 nsew signal output
rlabel metal3 s -300 5720 160 5840 4 W1BEG[3]
port 352 nsew signal output
rlabel metal3 s -300 5992 160 6112 4 W2BEG[0]
port 353 nsew signal output
rlabel metal3 s -300 6264 160 6384 4 W2BEG[1]
port 354 nsew signal output
rlabel metal3 s -300 6536 160 6656 4 W2BEG[2]
port 355 nsew signal output
rlabel metal3 s -300 6808 160 6928 4 W2BEG[3]
port 356 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 W2BEG[4]
port 357 nsew signal output
rlabel metal3 s -300 7352 160 7472 4 W2BEG[5]
port 358 nsew signal output
rlabel metal3 s -300 7624 160 7744 4 W2BEG[6]
port 359 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 W2BEG[7]
port 360 nsew signal output
rlabel metal3 s -300 8168 160 8288 4 W2BEGb[0]
port 361 nsew signal output
rlabel metal3 s -300 8440 160 8560 4 W2BEGb[1]
port 362 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 W2BEGb[2]
port 363 nsew signal output
rlabel metal3 s -300 8984 160 9104 4 W2BEGb[3]
port 364 nsew signal output
rlabel metal3 s -300 9256 160 9376 4 W2BEGb[4]
port 365 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 W2BEGb[5]
port 366 nsew signal output
rlabel metal3 s -300 9800 160 9920 4 W2BEGb[6]
port 367 nsew signal output
rlabel metal3 s -300 10072 160 10192 4 W2BEGb[7]
port 368 nsew signal output
rlabel metal3 s -300 14696 160 14816 4 W6BEG[0]
port 369 nsew signal output
rlabel metal3 s -300 17416 160 17536 4 W6BEG[10]
port 370 nsew signal output
rlabel metal3 s -300 17688 160 17808 4 W6BEG[11]
port 371 nsew signal output
rlabel metal3 s -300 14968 160 15088 4 W6BEG[1]
port 372 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 W6BEG[2]
port 373 nsew signal output
rlabel metal3 s -300 15512 160 15632 4 W6BEG[3]
port 374 nsew signal output
rlabel metal3 s -300 15784 160 15904 4 W6BEG[4]
port 375 nsew signal output
rlabel metal3 s -300 16056 160 16176 4 W6BEG[5]
port 376 nsew signal output
rlabel metal3 s -300 16328 160 16448 4 W6BEG[6]
port 377 nsew signal output
rlabel metal3 s -300 16600 160 16720 4 W6BEG[7]
port 378 nsew signal output
rlabel metal3 s -300 16872 160 16992 4 W6BEG[8]
port 379 nsew signal output
rlabel metal3 s -300 17144 160 17264 4 W6BEG[9]
port 380 nsew signal output
rlabel metal3 s -300 10344 160 10464 4 WW4BEG[0]
port 381 nsew signal output
rlabel metal3 s -300 13064 160 13184 4 WW4BEG[10]
port 382 nsew signal output
rlabel metal3 s -300 13336 160 13456 4 WW4BEG[11]
port 383 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 WW4BEG[12]
port 384 nsew signal output
rlabel metal3 s -300 13880 160 14000 4 WW4BEG[13]
port 385 nsew signal output
rlabel metal3 s -300 14152 160 14272 4 WW4BEG[14]
port 386 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 WW4BEG[15]
port 387 nsew signal output
rlabel metal3 s -300 10616 160 10736 4 WW4BEG[1]
port 388 nsew signal output
rlabel metal3 s -300 10888 160 11008 4 WW4BEG[2]
port 389 nsew signal output
rlabel metal3 s -300 11160 160 11280 4 WW4BEG[3]
port 390 nsew signal output
rlabel metal3 s -300 11432 160 11552 4 WW4BEG[4]
port 391 nsew signal output
rlabel metal3 s -300 11704 160 11824 4 WW4BEG[5]
port 392 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 WW4BEG[6]
port 393 nsew signal output
rlabel metal3 s -300 12248 160 12368 4 WW4BEG[7]
port 394 nsew signal output
rlabel metal3 s -300 12520 160 12640 4 WW4BEG[8]
port 395 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 WW4BEG[9]
port 396 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 25700 44700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4100600
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/RAM_IO/runs/24_12_08_00_02/results/signoff/RAM_IO.magic.gds
string GDS_START 173598
<< end >>

