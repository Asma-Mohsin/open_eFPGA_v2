// This is the unpowered netlist.
module W_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire A_I;
 wire A_O;
 wire A_Q;
 wire A_T;
 wire B_I;
 wire B_O;
 wire B_Q;
 wire B_T;
 wire \ConfigBits[0] ;
 wire \ConfigBits[100] ;
 wire \ConfigBits[101] ;
 wire \ConfigBits[102] ;
 wire \ConfigBits[103] ;
 wire \ConfigBits[104] ;
 wire \ConfigBits[105] ;
 wire \ConfigBits[106] ;
 wire \ConfigBits[107] ;
 wire \ConfigBits[108] ;
 wire \ConfigBits[109] ;
 wire \ConfigBits[10] ;
 wire \ConfigBits[110] ;
 wire \ConfigBits[111] ;
 wire \ConfigBits[112] ;
 wire \ConfigBits[113] ;
 wire \ConfigBits[11] ;
 wire \ConfigBits[12] ;
 wire \ConfigBits[13] ;
 wire \ConfigBits[14] ;
 wire \ConfigBits[15] ;
 wire \ConfigBits[16] ;
 wire \ConfigBits[17] ;
 wire \ConfigBits[18] ;
 wire \ConfigBits[19] ;
 wire \ConfigBits[1] ;
 wire \ConfigBits[20] ;
 wire \ConfigBits[21] ;
 wire \ConfigBits[22] ;
 wire \ConfigBits[23] ;
 wire \ConfigBits[24] ;
 wire \ConfigBits[25] ;
 wire \ConfigBits[26] ;
 wire \ConfigBits[27] ;
 wire \ConfigBits[28] ;
 wire \ConfigBits[29] ;
 wire \ConfigBits[2] ;
 wire \ConfigBits[30] ;
 wire \ConfigBits[31] ;
 wire \ConfigBits[32] ;
 wire \ConfigBits[33] ;
 wire \ConfigBits[34] ;
 wire \ConfigBits[35] ;
 wire \ConfigBits[36] ;
 wire \ConfigBits[37] ;
 wire \ConfigBits[38] ;
 wire \ConfigBits[39] ;
 wire \ConfigBits[3] ;
 wire \ConfigBits[40] ;
 wire \ConfigBits[41] ;
 wire \ConfigBits[42] ;
 wire \ConfigBits[43] ;
 wire \ConfigBits[44] ;
 wire \ConfigBits[45] ;
 wire \ConfigBits[46] ;
 wire \ConfigBits[47] ;
 wire \ConfigBits[48] ;
 wire \ConfigBits[49] ;
 wire \ConfigBits[4] ;
 wire \ConfigBits[50] ;
 wire \ConfigBits[51] ;
 wire \ConfigBits[52] ;
 wire \ConfigBits[53] ;
 wire \ConfigBits[54] ;
 wire \ConfigBits[55] ;
 wire \ConfigBits[56] ;
 wire \ConfigBits[57] ;
 wire \ConfigBits[58] ;
 wire \ConfigBits[59] ;
 wire \ConfigBits[5] ;
 wire \ConfigBits[60] ;
 wire \ConfigBits[61] ;
 wire \ConfigBits[62] ;
 wire \ConfigBits[63] ;
 wire \ConfigBits[64] ;
 wire \ConfigBits[65] ;
 wire \ConfigBits[66] ;
 wire \ConfigBits[67] ;
 wire \ConfigBits[68] ;
 wire \ConfigBits[69] ;
 wire \ConfigBits[6] ;
 wire \ConfigBits[70] ;
 wire \ConfigBits[71] ;
 wire \ConfigBits[72] ;
 wire \ConfigBits[73] ;
 wire \ConfigBits[74] ;
 wire \ConfigBits[75] ;
 wire \ConfigBits[76] ;
 wire \ConfigBits[77] ;
 wire \ConfigBits[78] ;
 wire \ConfigBits[79] ;
 wire \ConfigBits[7] ;
 wire \ConfigBits[80] ;
 wire \ConfigBits[81] ;
 wire \ConfigBits[82] ;
 wire \ConfigBits[83] ;
 wire \ConfigBits[84] ;
 wire \ConfigBits[85] ;
 wire \ConfigBits[86] ;
 wire \ConfigBits[87] ;
 wire \ConfigBits[88] ;
 wire \ConfigBits[89] ;
 wire \ConfigBits[8] ;
 wire \ConfigBits[90] ;
 wire \ConfigBits[91] ;
 wire \ConfigBits[92] ;
 wire \ConfigBits[93] ;
 wire \ConfigBits[94] ;
 wire \ConfigBits[95] ;
 wire \ConfigBits[96] ;
 wire \ConfigBits[97] ;
 wire \ConfigBits[98] ;
 wire \ConfigBits[99] ;
 wire \ConfigBits[9] ;
 wire \ConfigBits_N[0] ;
 wire \ConfigBits_N[100] ;
 wire \ConfigBits_N[101] ;
 wire \ConfigBits_N[102] ;
 wire \ConfigBits_N[103] ;
 wire \ConfigBits_N[104] ;
 wire \ConfigBits_N[105] ;
 wire \ConfigBits_N[106] ;
 wire \ConfigBits_N[107] ;
 wire \ConfigBits_N[108] ;
 wire \ConfigBits_N[109] ;
 wire \ConfigBits_N[10] ;
 wire \ConfigBits_N[110] ;
 wire \ConfigBits_N[111] ;
 wire \ConfigBits_N[112] ;
 wire \ConfigBits_N[113] ;
 wire \ConfigBits_N[11] ;
 wire \ConfigBits_N[12] ;
 wire \ConfigBits_N[13] ;
 wire \ConfigBits_N[14] ;
 wire \ConfigBits_N[15] ;
 wire \ConfigBits_N[16] ;
 wire \ConfigBits_N[17] ;
 wire \ConfigBits_N[18] ;
 wire \ConfigBits_N[19] ;
 wire \ConfigBits_N[1] ;
 wire \ConfigBits_N[20] ;
 wire \ConfigBits_N[21] ;
 wire \ConfigBits_N[22] ;
 wire \ConfigBits_N[23] ;
 wire \ConfigBits_N[24] ;
 wire \ConfigBits_N[25] ;
 wire \ConfigBits_N[26] ;
 wire \ConfigBits_N[27] ;
 wire \ConfigBits_N[28] ;
 wire \ConfigBits_N[29] ;
 wire \ConfigBits_N[2] ;
 wire \ConfigBits_N[30] ;
 wire \ConfigBits_N[31] ;
 wire \ConfigBits_N[32] ;
 wire \ConfigBits_N[33] ;
 wire \ConfigBits_N[34] ;
 wire \ConfigBits_N[35] ;
 wire \ConfigBits_N[36] ;
 wire \ConfigBits_N[37] ;
 wire \ConfigBits_N[38] ;
 wire \ConfigBits_N[39] ;
 wire \ConfigBits_N[3] ;
 wire \ConfigBits_N[40] ;
 wire \ConfigBits_N[41] ;
 wire \ConfigBits_N[42] ;
 wire \ConfigBits_N[43] ;
 wire \ConfigBits_N[44] ;
 wire \ConfigBits_N[45] ;
 wire \ConfigBits_N[46] ;
 wire \ConfigBits_N[47] ;
 wire \ConfigBits_N[48] ;
 wire \ConfigBits_N[49] ;
 wire \ConfigBits_N[4] ;
 wire \ConfigBits_N[50] ;
 wire \ConfigBits_N[51] ;
 wire \ConfigBits_N[52] ;
 wire \ConfigBits_N[53] ;
 wire \ConfigBits_N[54] ;
 wire \ConfigBits_N[55] ;
 wire \ConfigBits_N[56] ;
 wire \ConfigBits_N[57] ;
 wire \ConfigBits_N[58] ;
 wire \ConfigBits_N[59] ;
 wire \ConfigBits_N[5] ;
 wire \ConfigBits_N[60] ;
 wire \ConfigBits_N[61] ;
 wire \ConfigBits_N[62] ;
 wire \ConfigBits_N[63] ;
 wire \ConfigBits_N[64] ;
 wire \ConfigBits_N[65] ;
 wire \ConfigBits_N[66] ;
 wire \ConfigBits_N[67] ;
 wire \ConfigBits_N[68] ;
 wire \ConfigBits_N[69] ;
 wire \ConfigBits_N[6] ;
 wire \ConfigBits_N[70] ;
 wire \ConfigBits_N[71] ;
 wire \ConfigBits_N[72] ;
 wire \ConfigBits_N[73] ;
 wire \ConfigBits_N[74] ;
 wire \ConfigBits_N[75] ;
 wire \ConfigBits_N[76] ;
 wire \ConfigBits_N[77] ;
 wire \ConfigBits_N[78] ;
 wire \ConfigBits_N[79] ;
 wire \ConfigBits_N[7] ;
 wire \ConfigBits_N[80] ;
 wire \ConfigBits_N[81] ;
 wire \ConfigBits_N[82] ;
 wire \ConfigBits_N[83] ;
 wire \ConfigBits_N[84] ;
 wire \ConfigBits_N[85] ;
 wire \ConfigBits_N[86] ;
 wire \ConfigBits_N[87] ;
 wire \ConfigBits_N[88] ;
 wire \ConfigBits_N[89] ;
 wire \ConfigBits_N[8] ;
 wire \ConfigBits_N[90] ;
 wire \ConfigBits_N[91] ;
 wire \ConfigBits_N[92] ;
 wire \ConfigBits_N[93] ;
 wire \ConfigBits_N[94] ;
 wire \ConfigBits_N[95] ;
 wire \ConfigBits_N[96] ;
 wire \ConfigBits_N[97] ;
 wire \ConfigBits_N[98] ;
 wire \ConfigBits_N[99] ;
 wire \ConfigBits_N[9] ;
 wire \FrameData_O_i[0] ;
 wire \FrameData_O_i[10] ;
 wire \FrameData_O_i[11] ;
 wire \FrameData_O_i[12] ;
 wire \FrameData_O_i[13] ;
 wire \FrameData_O_i[14] ;
 wire \FrameData_O_i[15] ;
 wire \FrameData_O_i[16] ;
 wire \FrameData_O_i[17] ;
 wire \FrameData_O_i[18] ;
 wire \FrameData_O_i[19] ;
 wire \FrameData_O_i[1] ;
 wire \FrameData_O_i[20] ;
 wire \FrameData_O_i[21] ;
 wire \FrameData_O_i[22] ;
 wire \FrameData_O_i[23] ;
 wire \FrameData_O_i[24] ;
 wire \FrameData_O_i[25] ;
 wire \FrameData_O_i[26] ;
 wire \FrameData_O_i[27] ;
 wire \FrameData_O_i[28] ;
 wire \FrameData_O_i[29] ;
 wire \FrameData_O_i[2] ;
 wire \FrameData_O_i[30] ;
 wire \FrameData_O_i[31] ;
 wire \FrameData_O_i[3] ;
 wire \FrameData_O_i[4] ;
 wire \FrameData_O_i[5] ;
 wire \FrameData_O_i[6] ;
 wire \FrameData_O_i[7] ;
 wire \FrameData_O_i[8] ;
 wire \FrameData_O_i[9] ;
 wire \FrameStrobe_O_i[0] ;
 wire \FrameStrobe_O_i[10] ;
 wire \FrameStrobe_O_i[11] ;
 wire \FrameStrobe_O_i[12] ;
 wire \FrameStrobe_O_i[13] ;
 wire \FrameStrobe_O_i[14] ;
 wire \FrameStrobe_O_i[15] ;
 wire \FrameStrobe_O_i[16] ;
 wire \FrameStrobe_O_i[17] ;
 wire \FrameStrobe_O_i[18] ;
 wire \FrameStrobe_O_i[19] ;
 wire \FrameStrobe_O_i[1] ;
 wire \FrameStrobe_O_i[2] ;
 wire \FrameStrobe_O_i[3] ;
 wire \FrameStrobe_O_i[4] ;
 wire \FrameStrobe_O_i[5] ;
 wire \FrameStrobe_O_i[6] ;
 wire \FrameStrobe_O_i[7] ;
 wire \FrameStrobe_O_i[8] ;
 wire \FrameStrobe_O_i[9] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out1 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out2 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out3 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out1 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out2 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out3 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out1 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[0] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[1] ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_0_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_1_ ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out1 ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net95));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_73 ();
 sky130_fd_sc_hd__inv_2 \Inst_A_IO_1_bidirectional_frame_config_pass/_0_  (.A(A_T),
    .Y(net104));
 sky130_fd_sc_hd__dfxtp_1 \Inst_A_IO_1_bidirectional_frame_config_pass/_1_  (.CLK(UserCLK),
    .D(net1),
    .Q(A_Q));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_IO_1_bidirectional_frame_config_pass/_2_  (.A(A_I),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 \Inst_A_IO_1_bidirectional_frame_config_pass/_3_  (.A(net1),
    .X(A_O));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access/_0_  (.A(\ConfigBits[0] ),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access/_1_  (.A(\ConfigBits[1] ),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access/_2_  (.A(\ConfigBits[2] ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access/_3_  (.A(\ConfigBits[3] ),
    .X(net108));
 sky130_fd_sc_hd__inv_2 \Inst_B_IO_1_bidirectional_frame_config_pass/_0_  (.A(B_T),
    .Y(net110));
 sky130_fd_sc_hd__dfxtp_1 \Inst_B_IO_1_bidirectional_frame_config_pass/_1_  (.CLK(UserCLK),
    .D(net2),
    .Q(B_Q));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_IO_1_bidirectional_frame_config_pass/_2_  (.A(B_I),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 \Inst_B_IO_1_bidirectional_frame_config_pass/_3_  (.A(net2),
    .X(B_O));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access/_0_  (.A(\ConfigBits[4] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access/_1_  (.A(\ConfigBits[5] ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access/_2_  (.A(\ConfigBits[6] ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access/_3_  (.A(\ConfigBits[7] ),
    .X(net114));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit0  (.D(net3),
    .GATE(net35),
    .Q(\ConfigBits[82] ),
    .Q_N(\ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit1  (.D(net14),
    .GATE(net35),
    .Q(\ConfigBits[83] ),
    .Q_N(\ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit10  (.D(net4),
    .GATE(net35),
    .Q(\ConfigBits[92] ),
    .Q_N(\ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit11  (.D(net5),
    .GATE(net35),
    .Q(\ConfigBits[93] ),
    .Q_N(\ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit12  (.D(net6),
    .GATE(net35),
    .Q(\ConfigBits[94] ),
    .Q_N(\ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit13  (.D(net7),
    .GATE(net35),
    .Q(\ConfigBits[95] ),
    .Q_N(\ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit14  (.D(net8),
    .GATE(net35),
    .Q(\ConfigBits[96] ),
    .Q_N(\ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit15  (.D(net9),
    .GATE(net35),
    .Q(\ConfigBits[97] ),
    .Q_N(\ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit16  (.D(net10),
    .GATE(net35),
    .Q(\ConfigBits[98] ),
    .Q_N(\ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit17  (.D(net11),
    .GATE(net35),
    .Q(\ConfigBits[99] ),
    .Q_N(\ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit18  (.D(net12),
    .GATE(net35),
    .Q(\ConfigBits[100] ),
    .Q_N(\ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit19  (.D(net13),
    .GATE(net35),
    .Q(\ConfigBits[101] ),
    .Q_N(\ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit2  (.D(net25),
    .GATE(net35),
    .Q(\ConfigBits[84] ),
    .Q_N(\ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit20  (.D(net15),
    .GATE(net35),
    .Q(\ConfigBits[102] ),
    .Q_N(\ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit21  (.D(net16),
    .GATE(net35),
    .Q(\ConfigBits[103] ),
    .Q_N(\ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit22  (.D(net17),
    .GATE(net35),
    .Q(\ConfigBits[104] ),
    .Q_N(\ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit23  (.D(net18),
    .GATE(net35),
    .Q(\ConfigBits[105] ),
    .Q_N(\ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit24  (.D(net19),
    .GATE(net35),
    .Q(\ConfigBits[106] ),
    .Q_N(\ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit25  (.D(net20),
    .GATE(net35),
    .Q(\ConfigBits[107] ),
    .Q_N(\ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit26  (.D(net21),
    .GATE(net35),
    .Q(\ConfigBits[108] ),
    .Q_N(\ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit27  (.D(net22),
    .GATE(net35),
    .Q(\ConfigBits[109] ),
    .Q_N(\ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit28  (.D(net23),
    .GATE(net35),
    .Q(\ConfigBits[110] ),
    .Q_N(\ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit29  (.D(net24),
    .GATE(net35),
    .Q(\ConfigBits[111] ),
    .Q_N(\ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit3  (.D(net28),
    .GATE(net35),
    .Q(\ConfigBits[85] ),
    .Q_N(\ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit30  (.D(net26),
    .GATE(net35),
    .Q(\ConfigBits[112] ),
    .Q_N(\ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit31  (.D(net27),
    .GATE(net35),
    .Q(\ConfigBits[113] ),
    .Q_N(\ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit4  (.D(net29),
    .GATE(net35),
    .Q(\ConfigBits[86] ),
    .Q_N(\ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit5  (.D(net30),
    .GATE(net35),
    .Q(\ConfigBits[87] ),
    .Q_N(\ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit6  (.D(net31),
    .GATE(net35),
    .Q(\ConfigBits[88] ),
    .Q_N(\ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit7  (.D(net32),
    .GATE(net35),
    .Q(\ConfigBits[89] ),
    .Q_N(\ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit8  (.D(net33),
    .GATE(net35),
    .Q(\ConfigBits[90] ),
    .Q_N(\ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame0_bit9  (.D(net34),
    .GATE(net35),
    .Q(\ConfigBits[91] ),
    .Q_N(\ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit0  (.D(net3),
    .GATE(net46),
    .Q(\ConfigBits[50] ),
    .Q_N(\ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit1  (.D(net14),
    .GATE(net46),
    .Q(\ConfigBits[51] ),
    .Q_N(\ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit10  (.D(net4),
    .GATE(net46),
    .Q(\ConfigBits[60] ),
    .Q_N(\ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit11  (.D(net5),
    .GATE(net46),
    .Q(\ConfigBits[61] ),
    .Q_N(\ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit12  (.D(net6),
    .GATE(net46),
    .Q(\ConfigBits[62] ),
    .Q_N(\ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit13  (.D(net7),
    .GATE(net46),
    .Q(\ConfigBits[63] ),
    .Q_N(\ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit14  (.D(net8),
    .GATE(net46),
    .Q(\ConfigBits[64] ),
    .Q_N(\ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit15  (.D(net9),
    .GATE(net46),
    .Q(\ConfigBits[65] ),
    .Q_N(\ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit16  (.D(net10),
    .GATE(net46),
    .Q(\ConfigBits[66] ),
    .Q_N(\ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit17  (.D(net11),
    .GATE(net46),
    .Q(\ConfigBits[67] ),
    .Q_N(\ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit18  (.D(net12),
    .GATE(net46),
    .Q(\ConfigBits[68] ),
    .Q_N(\ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit19  (.D(net13),
    .GATE(net46),
    .Q(\ConfigBits[69] ),
    .Q_N(\ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit2  (.D(net25),
    .GATE(net46),
    .Q(\ConfigBits[52] ),
    .Q_N(\ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit20  (.D(net15),
    .GATE(net46),
    .Q(\ConfigBits[70] ),
    .Q_N(\ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit21  (.D(net16),
    .GATE(net46),
    .Q(\ConfigBits[71] ),
    .Q_N(\ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit22  (.D(net17),
    .GATE(net46),
    .Q(\ConfigBits[72] ),
    .Q_N(\ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit23  (.D(net18),
    .GATE(net46),
    .Q(\ConfigBits[73] ),
    .Q_N(\ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit24  (.D(net19),
    .GATE(net46),
    .Q(\ConfigBits[74] ),
    .Q_N(\ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit25  (.D(net20),
    .GATE(net46),
    .Q(\ConfigBits[75] ),
    .Q_N(\ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit26  (.D(net21),
    .GATE(net46),
    .Q(\ConfigBits[76] ),
    .Q_N(\ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit27  (.D(net22),
    .GATE(net46),
    .Q(\ConfigBits[77] ),
    .Q_N(\ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit28  (.D(net23),
    .GATE(net46),
    .Q(\ConfigBits[78] ),
    .Q_N(\ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit29  (.D(net24),
    .GATE(net46),
    .Q(\ConfigBits[79] ),
    .Q_N(\ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit3  (.D(net28),
    .GATE(net46),
    .Q(\ConfigBits[53] ),
    .Q_N(\ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit30  (.D(net26),
    .GATE(net46),
    .Q(\ConfigBits[80] ),
    .Q_N(\ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit31  (.D(net27),
    .GATE(net46),
    .Q(\ConfigBits[81] ),
    .Q_N(\ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit4  (.D(net29),
    .GATE(net46),
    .Q(\ConfigBits[54] ),
    .Q_N(\ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit5  (.D(net30),
    .GATE(net46),
    .Q(\ConfigBits[55] ),
    .Q_N(\ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit6  (.D(net31),
    .GATE(net46),
    .Q(\ConfigBits[56] ),
    .Q_N(\ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit7  (.D(net32),
    .GATE(net46),
    .Q(\ConfigBits[57] ),
    .Q_N(\ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit8  (.D(net33),
    .GATE(net46),
    .Q(\ConfigBits[58] ),
    .Q_N(\ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame1_bit9  (.D(net34),
    .GATE(net46),
    .Q(\ConfigBits[59] ),
    .Q_N(\ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit0  (.D(net3),
    .GATE(net47),
    .Q(\ConfigBits[18] ),
    .Q_N(\ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit1  (.D(net14),
    .GATE(net47),
    .Q(\ConfigBits[19] ),
    .Q_N(\ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit10  (.D(net4),
    .GATE(net47),
    .Q(\ConfigBits[28] ),
    .Q_N(\ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit11  (.D(net5),
    .GATE(net47),
    .Q(\ConfigBits[29] ),
    .Q_N(\ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit12  (.D(net6),
    .GATE(net47),
    .Q(\ConfigBits[30] ),
    .Q_N(\ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit13  (.D(net7),
    .GATE(net47),
    .Q(\ConfigBits[31] ),
    .Q_N(\ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit14  (.D(net8),
    .GATE(net47),
    .Q(\ConfigBits[32] ),
    .Q_N(\ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit15  (.D(net9),
    .GATE(net47),
    .Q(\ConfigBits[33] ),
    .Q_N(\ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit16  (.D(net10),
    .GATE(net47),
    .Q(\ConfigBits[34] ),
    .Q_N(\ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit17  (.D(net11),
    .GATE(net47),
    .Q(\ConfigBits[35] ),
    .Q_N(\ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit18  (.D(net12),
    .GATE(net47),
    .Q(\ConfigBits[36] ),
    .Q_N(\ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit19  (.D(net13),
    .GATE(net47),
    .Q(\ConfigBits[37] ),
    .Q_N(\ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit2  (.D(net25),
    .GATE(net47),
    .Q(\ConfigBits[20] ),
    .Q_N(\ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit20  (.D(net15),
    .GATE(net47),
    .Q(\ConfigBits[38] ),
    .Q_N(\ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit21  (.D(net16),
    .GATE(net47),
    .Q(\ConfigBits[39] ),
    .Q_N(\ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit22  (.D(net17),
    .GATE(net47),
    .Q(\ConfigBits[40] ),
    .Q_N(\ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit23  (.D(net18),
    .GATE(net47),
    .Q(\ConfigBits[41] ),
    .Q_N(\ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit24  (.D(net19),
    .GATE(net47),
    .Q(\ConfigBits[42] ),
    .Q_N(\ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit25  (.D(net20),
    .GATE(net47),
    .Q(\ConfigBits[43] ),
    .Q_N(\ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit26  (.D(net21),
    .GATE(net47),
    .Q(\ConfigBits[44] ),
    .Q_N(\ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit27  (.D(net22),
    .GATE(net47),
    .Q(\ConfigBits[45] ),
    .Q_N(\ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit28  (.D(net23),
    .GATE(net47),
    .Q(\ConfigBits[46] ),
    .Q_N(\ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit29  (.D(net24),
    .GATE(net47),
    .Q(\ConfigBits[47] ),
    .Q_N(\ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit3  (.D(net28),
    .GATE(net47),
    .Q(\ConfigBits[21] ),
    .Q_N(\ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit30  (.D(net26),
    .GATE(net47),
    .Q(\ConfigBits[48] ),
    .Q_N(\ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit31  (.D(net27),
    .GATE(net47),
    .Q(\ConfigBits[49] ),
    .Q_N(\ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit4  (.D(net29),
    .GATE(net47),
    .Q(\ConfigBits[22] ),
    .Q_N(\ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit5  (.D(net30),
    .GATE(net47),
    .Q(\ConfigBits[23] ),
    .Q_N(\ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit6  (.D(net31),
    .GATE(net47),
    .Q(\ConfigBits[24] ),
    .Q_N(\ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit7  (.D(net32),
    .GATE(net47),
    .Q(\ConfigBits[25] ),
    .Q_N(\ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit8  (.D(net33),
    .GATE(net47),
    .Q(\ConfigBits[26] ),
    .Q_N(\ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame2_bit9  (.D(net34),
    .GATE(net47),
    .Q(\ConfigBits[27] ),
    .Q_N(\ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit14  (.D(net8),
    .GATE(net48),
    .Q(\ConfigBits[0] ),
    .Q_N(\ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit15  (.D(net9),
    .GATE(net48),
    .Q(\ConfigBits[1] ),
    .Q_N(\ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit16  (.D(net10),
    .GATE(net48),
    .Q(\ConfigBits[2] ),
    .Q_N(\ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit17  (.D(net11),
    .GATE(net48),
    .Q(\ConfigBits[3] ),
    .Q_N(\ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit18  (.D(net12),
    .GATE(net48),
    .Q(\ConfigBits[4] ),
    .Q_N(\ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit19  (.D(net13),
    .GATE(net48),
    .Q(\ConfigBits[5] ),
    .Q_N(\ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit20  (.D(net15),
    .GATE(net48),
    .Q(\ConfigBits[6] ),
    .Q_N(\ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit21  (.D(net16),
    .GATE(net48),
    .Q(\ConfigBits[7] ),
    .Q_N(\ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit22  (.D(net17),
    .GATE(net48),
    .Q(\ConfigBits[8] ),
    .Q_N(\ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit23  (.D(net18),
    .GATE(net48),
    .Q(\ConfigBits[9] ),
    .Q_N(\ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit24  (.D(net19),
    .GATE(net48),
    .Q(\ConfigBits[10] ),
    .Q_N(\ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit25  (.D(net20),
    .GATE(net48),
    .Q(\ConfigBits[11] ),
    .Q_N(\ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit26  (.D(net21),
    .GATE(net48),
    .Q(\ConfigBits[12] ),
    .Q_N(\ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit27  (.D(net22),
    .GATE(net48),
    .Q(\ConfigBits[13] ),
    .Q_N(\ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit28  (.D(net23),
    .GATE(net48),
    .Q(\ConfigBits[14] ),
    .Q_N(\ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit29  (.D(net24),
    .GATE(net48),
    .Q(\ConfigBits[15] ),
    .Q_N(\ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit30  (.D(net26),
    .GATE(net48),
    .Q(\ConfigBits[16] ),
    .Q_N(\ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem/Inst_frame3_bit31  (.D(net27),
    .GATE(net48),
    .Q(\ConfigBits[17] ),
    .Q_N(\ConfigBits_N[17] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_inst0  (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_inst1  (.A0(net71),
    .A1(net72),
    .A2(net73),
    .A3(net74),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_inst2  (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_inst3  (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_inst4  (.A0(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out0 ),
    .A1(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out1 ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out2 ),
    .A3(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[102] ),
    .S1(\ConfigBits[103] ),
    .X(A_I));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_inst0  (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\ConfigBits[107] ),
    .S1(\ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_inst1  (.A0(net71),
    .A1(net72),
    .A2(net73),
    .A3(net74),
    .S0(\ConfigBits[107] ),
    .S1(\ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_inst2  (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\ConfigBits[107] ),
    .S1(\ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_inst3  (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\ConfigBits[107] ),
    .S1(\ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_inst4  (.A0(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out0 ),
    .A1(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out1 ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out2 ),
    .A3(\Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[109] ),
    .S1(\ConfigBits[110] ),
    .X(B_I));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[1] ),
    .B(\ConfigBits[8] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_4_  (.A1(\ConfigBits[8] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_1_ ),
    .Y(net115));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/break_comb_loop_inst0/_0_  (.A(net58),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/break_comb_loop_inst1/_0_  (.A(A_O),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[1] ),
    .B(\ConfigBits[9] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_4_  (.A1(\ConfigBits[9] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_1_ ),
    .Y(net116));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/break_comb_loop_inst0/_0_  (.A(net57),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/break_comb_loop_inst1/_0_  (.A(A_Q),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[1] ),
    .B(\ConfigBits[10] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_4_  (.A1(\ConfigBits[10] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_1_ ),
    .Y(net117));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/break_comb_loop_inst0/_0_  (.A(net56),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/break_comb_loop_inst1/_0_  (.A(B_O),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[1] ),
    .B(\ConfigBits[11] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_4_  (.A1(\ConfigBits[11] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_1_ ),
    .Y(net118));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/break_comb_loop_inst0/_0_  (.A(net55),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/break_comb_loop_inst1/_0_  (.A(B_Q),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG0  (.A0(net74),
    .A1(net100),
    .A2(net93),
    .A3(net84),
    .S0(\ConfigBits[12] ),
    .S1(\ConfigBits[13] ),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG1  (.A0(net73),
    .A1(net99),
    .A2(net92),
    .A3(net83),
    .S0(\ConfigBits[14] ),
    .S1(\ConfigBits[15] ),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG2  (.A0(net72),
    .A1(net98),
    .A2(net91),
    .A3(net82),
    .S0(\ConfigBits[16] ),
    .S1(\ConfigBits[17] ),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG3  (.A0(net71),
    .A1(net97),
    .A2(net90),
    .A3(net81),
    .S0(\ConfigBits[18] ),
    .S1(\ConfigBits[19] ),
    .X(net122));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG4  (.A0(net70),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\ConfigBits[20] ),
    .S1(\ConfigBits[21] ),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG5  (.A0(net69),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\ConfigBits[22] ),
    .S1(\ConfigBits[23] ),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG6  (.A0(net68),
    .A1(net94),
    .A2(net102),
    .A3(net78),
    .S0(\ConfigBits[24] ),
    .S1(\ConfigBits[25] ),
    .X(net125));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEG7  (.A0(net67),
    .A1(net87),
    .A2(net101),
    .A3(net75),
    .S0(\ConfigBits[26] ),
    .S1(\ConfigBits[27] ),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb0  (.A0(net66),
    .A1(net100),
    .A2(net93),
    .A3(net84),
    .S0(\ConfigBits[28] ),
    .S1(\ConfigBits[29] ),
    .X(net127));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb1  (.A0(net65),
    .A1(net99),
    .A2(net92),
    .A3(net83),
    .S0(\ConfigBits[30] ),
    .S1(\ConfigBits[31] ),
    .X(net128));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb2  (.A0(net64),
    .A1(net98),
    .A2(net91),
    .A3(net82),
    .S0(\ConfigBits[32] ),
    .S1(\ConfigBits[33] ),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb3  (.A0(net63),
    .A1(net97),
    .A2(net90),
    .A3(net81),
    .S0(\ConfigBits[34] ),
    .S1(\ConfigBits[35] ),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb4  (.A0(net62),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\ConfigBits[36] ),
    .S1(\ConfigBits[37] ),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb5  (.A0(net61),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\ConfigBits[38] ),
    .S1(\ConfigBits[39] ),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb6  (.A0(net60),
    .A1(net94),
    .A2(net102),
    .A3(net78),
    .S0(\ConfigBits[40] ),
    .S1(\ConfigBits[41] ),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E2BEGb7  (.A0(net59),
    .A1(net87),
    .A2(net101),
    .A3(net75),
    .S0(\ConfigBits[42] ),
    .S1(\ConfigBits[43] ),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG0  (.A0(net57),
    .A1(net89),
    .A2(net77),
    .A3(A_O),
    .S0(\ConfigBits[76] ),
    .S1(\ConfigBits[77] ),
    .X(net135));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG1  (.A0(net58),
    .A1(net88),
    .A2(net76),
    .A3(B_O),
    .S0(\ConfigBits[78] ),
    .S1(\ConfigBits[79] ),
    .X(net138));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG10  (.A0(net56),
    .A1(net94),
    .A2(net78),
    .A3(A_Q),
    .S0(\ConfigBits[96] ),
    .S1(\ConfigBits[97] ),
    .X(net136));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG11  (.A0(net55),
    .A1(net87),
    .A2(net75),
    .A3(B_Q),
    .S0(\ConfigBits[98] ),
    .S1(\ConfigBits[99] ),
    .X(net137));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG2  (.A0(net100),
    .A1(net93),
    .A2(net84),
    .A3(A_O),
    .S0(\ConfigBits[80] ),
    .S1(\ConfigBits[81] ),
    .X(net139));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG3  (.A0(net99),
    .A1(net92),
    .A2(net83),
    .A3(B_O),
    .S0(\ConfigBits[82] ),
    .S1(\ConfigBits[83] ),
    .X(net140));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG4  (.A0(net57),
    .A1(net96),
    .A2(net80),
    .A3(A_O),
    .S0(\ConfigBits[84] ),
    .S1(\ConfigBits[85] ),
    .X(net141));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG5  (.A0(net58),
    .A1(net95),
    .A2(net79),
    .A3(B_O),
    .S0(\ConfigBits[86] ),
    .S1(\ConfigBits[87] ),
    .X(net142));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG6  (.A0(net56),
    .A1(net102),
    .A2(net86),
    .A3(A_Q),
    .S0(\ConfigBits[88] ),
    .S1(\ConfigBits[89] ),
    .X(net143));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG7  (.A0(net55),
    .A1(net101),
    .A2(net85),
    .A3(B_Q),
    .S0(\ConfigBits[90] ),
    .S1(\ConfigBits[91] ),
    .X(net144));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG8  (.A0(net98),
    .A1(net91),
    .A2(net82),
    .A3(A_Q),
    .S0(\ConfigBits[92] ),
    .S1(\ConfigBits[93] ),
    .X(net145));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_E6BEG9  (.A0(net97),
    .A1(net90),
    .A2(net81),
    .A3(B_Q),
    .S0(\ConfigBits[94] ),
    .S1(\ConfigBits[95] ),
    .X(net146));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG0  (.A0(net75),
    .A1(net79),
    .A2(net81),
    .A3(A_O),
    .S0(\ConfigBits[44] ),
    .S1(\ConfigBits[45] ),
    .X(net147));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG1  (.A0(net83),
    .A1(net85),
    .A2(net76),
    .A3(B_O),
    .S0(\ConfigBits[46] ),
    .S1(\ConfigBits[47] ),
    .X(net154));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG10  (.A0(net75),
    .A1(net79),
    .A2(net81),
    .A3(A_O),
    .S0(\ConfigBits[64] ),
    .S1(\ConfigBits[65] ),
    .X(net148));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG11  (.A0(net83),
    .A1(net85),
    .A2(net76),
    .A3(B_O),
    .S0(\ConfigBits[66] ),
    .S1(\ConfigBits[67] ),
    .X(net149));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG12  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(A_Q),
    .S0(\ConfigBits[68] ),
    .S1(\ConfigBits[69] ),
    .X(net150));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG13  (.A0(net84),
    .A1(net86),
    .A2(net77),
    .A3(B_Q),
    .S0(\ConfigBits[70] ),
    .S1(\ConfigBits[71] ),
    .X(net151));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG14  (.A0(net67),
    .A1(net69),
    .A2(net71),
    .A3(net73),
    .S0(\ConfigBits[72] ),
    .S1(\ConfigBits[73] ),
    .X(net152));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG15  (.A0(net68),
    .A1(net70),
    .A2(net72),
    .A3(net74),
    .S0(\ConfigBits[74] ),
    .S1(\ConfigBits[75] ),
    .X(net153));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG2  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(A_Q),
    .S0(\ConfigBits[48] ),
    .S1(\ConfigBits[49] ),
    .X(net155));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG3  (.A0(net84),
    .A1(net86),
    .A2(net77),
    .A3(B_Q),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(net156));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG4  (.A0(net59),
    .A1(net61),
    .A2(net63),
    .A3(net65),
    .S0(\ConfigBits[52] ),
    .S1(\ConfigBits[53] ),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG5  (.A0(net60),
    .A1(net62),
    .A2(net64),
    .A3(net66),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(net158));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG6  (.A0(net67),
    .A1(net69),
    .A2(net71),
    .A3(net73),
    .S0(\ConfigBits[56] ),
    .S1(\ConfigBits[57] ),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG7  (.A0(net68),
    .A1(net70),
    .A2(net72),
    .A3(net74),
    .S0(\ConfigBits[58] ),
    .S1(\ConfigBits[59] ),
    .X(net160));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG8  (.A0(net81),
    .A1(net83),
    .A2(net85),
    .A3(net76),
    .S0(\ConfigBits[60] ),
    .S1(\ConfigBits[61] ),
    .X(net161));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux41_buf_EE4BEG9  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(net84),
    .S0(\ConfigBits[62] ),
    .S1(\ConfigBits[63] ),
    .X(net162));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[106] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_4_  (.A1(\ConfigBits[106] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_1_ ),
    .Y(A_T));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out0 ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out1 ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_inst0  (.A0(net74),
    .A1(net59),
    .A2(net60),
    .A3(net61),
    .S0(\ConfigBits[104] ),
    .S1(\ConfigBits[105] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_inst1  (.A0(net62),
    .A1(net63),
    .A2(net216),
    .A3(net218),
    .S0(\ConfigBits[104] ),
    .S1(\ConfigBits[105] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_inst1_216  (.LO(net216));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_inst1_218  (.HI(net218));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_2_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_3_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[113] ),
    .Y(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_4_  (.A1(\ConfigBits[113] ),
    .A2(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_0_ ),
    .B1(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_1_ ),
    .Y(B_T));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out0 ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out1 ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_inst0  (.A0(net73),
    .A1(net74),
    .A2(net59),
    .A3(net63),
    .S0(\ConfigBits[111] ),
    .S1(\ConfigBits[112] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_inst1  (.A0(net64),
    .A1(net65),
    .A2(net217),
    .A3(net219),
    .S0(\ConfigBits[111] ),
    .S1(\ConfigBits[112] ),
    .X(\Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_inst1_217  (.LO(net217));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_inst1_219  (.HI(net219));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0/_0_  (.A(net3),
    .X(\FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1/_0_  (.A(net14),
    .X(\FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10/_0_  (.A(net4),
    .X(\FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11/_0_  (.A(net5),
    .X(\FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12/_0_  (.A(net6),
    .X(\FrameData_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13/_0_  (.A(net7),
    .X(\FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14/_0_  (.A(net8),
    .X(\FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15/_0_  (.A(net9),
    .X(\FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16/_0_  (.A(net10),
    .X(\FrameData_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17/_0_  (.A(net11),
    .X(\FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18/_0_  (.A(net12),
    .X(\FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19/_0_  (.A(net13),
    .X(\FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2/_0_  (.A(net25),
    .X(\FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20/_0_  (.A(net15),
    .X(\FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21/_0_  (.A(net16),
    .X(\FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22/_0_  (.A(net17),
    .X(\FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23/_0_  (.A(net18),
    .X(\FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24/_0_  (.A(net19),
    .X(\FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25/_0_  (.A(net20),
    .X(\FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26/_0_  (.A(net21),
    .X(\FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27/_0_  (.A(net22),
    .X(\FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28/_0_  (.A(net23),
    .X(\FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29/_0_  (.A(net24),
    .X(\FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3/_0_  (.A(net28),
    .X(\FrameData_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30/_0_  (.A(net26),
    .X(\FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31/_0_  (.A(net27),
    .X(\FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4/_0_  (.A(net29),
    .X(\FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5/_0_  (.A(net30),
    .X(\FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6/_0_  (.A(net31),
    .X(\FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7/_0_  (.A(net32),
    .X(\FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8/_0_  (.A(net33),
    .X(\FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9/_0_  (.A(net34),
    .X(\FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0/_0_  (.A(\FrameData_O_i[0] ),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1/_0_  (.A(\FrameData_O_i[1] ),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10/_0_  (.A(\FrameData_O_i[10] ),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11/_0_  (.A(\FrameData_O_i[11] ),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12/_0_  (.A(\FrameData_O_i[12] ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13/_0_  (.A(\FrameData_O_i[13] ),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14/_0_  (.A(\FrameData_O_i[14] ),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15/_0_  (.A(\FrameData_O_i[15] ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16/_0_  (.A(\FrameData_O_i[16] ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17/_0_  (.A(\FrameData_O_i[17] ),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18/_0_  (.A(\FrameData_O_i[18] ),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19/_0_  (.A(\FrameData_O_i[19] ),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2/_0_  (.A(\FrameData_O_i[2] ),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20/_0_  (.A(\FrameData_O_i[20] ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21/_0_  (.A(\FrameData_O_i[21] ),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22/_0_  (.A(\FrameData_O_i[22] ),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23/_0_  (.A(\FrameData_O_i[23] ),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24/_0_  (.A(\FrameData_O_i[24] ),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25/_0_  (.A(\FrameData_O_i[25] ),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26/_0_  (.A(\FrameData_O_i[26] ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27/_0_  (.A(\FrameData_O_i[27] ),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28/_0_  (.A(\FrameData_O_i[28] ),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29/_0_  (.A(\FrameData_O_i[29] ),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3/_0_  (.A(\FrameData_O_i[3] ),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30/_0_  (.A(\FrameData_O_i[30] ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31/_0_  (.A(\FrameData_O_i[31] ),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4/_0_  (.A(\FrameData_O_i[4] ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5/_0_  (.A(\FrameData_O_i[5] ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6/_0_  (.A(\FrameData_O_i[6] ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7/_0_  (.A(\FrameData_O_i[7] ),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8/_0_  (.A(\FrameData_O_i[8] ),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9/_0_  (.A(\FrameData_O_i[9] ),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input1 (.A(A_O_top),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(FrameData[16]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input100 (.A(WW4END[7]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(WW4END[8]),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 input102 (.A(WW4END[9]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input11 (.A(FrameData[17]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(FrameData[18]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(FrameData[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(FrameData[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(FrameData[20]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(FrameData[21]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(FrameData[22]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(FrameData[23]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(FrameData[24]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(B_O_top),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(FrameData[25]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(FrameData[26]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(FrameData[27]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(FrameData[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(FrameData[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(FrameData[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(FrameData[30]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(FrameData[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(FrameData[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(FrameData[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(FrameData[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(FrameData[5]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(FrameData[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(FrameData[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(FrameData[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(FrameData[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_8 input35 (.A(FrameStrobe[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(FrameStrobe[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(FrameStrobe[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(FrameStrobe[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(FrameStrobe[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(FrameData[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(FrameStrobe[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(FrameStrobe[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(FrameStrobe[16]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(FrameStrobe[17]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(FrameStrobe[18]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(FrameStrobe[19]),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(FrameStrobe[1]),
    .X(net46));
 sky130_fd_sc_hd__buf_8 input47 (.A(FrameStrobe[2]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(FrameStrobe[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(FrameStrobe[4]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(FrameData[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(FrameStrobe[5]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(FrameStrobe[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(FrameStrobe[7]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(FrameStrobe[8]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(FrameStrobe[9]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(W1END[0]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(W1END[1]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(W1END[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(W1END[3]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(W2END[0]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(FrameData[12]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(W2END[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(W2END[2]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(W2END[3]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(W2END[4]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(W2END[5]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(W2END[6]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(W2END[7]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(W2MID[0]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(W2MID[1]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(W2MID[2]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(FrameData[13]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(W2MID[3]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(W2MID[4]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(W2MID[5]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(W2MID[6]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(W2MID[7]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(W6END[0]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(W6END[10]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(W6END[11]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(W6END[1]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(W6END[2]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(FrameData[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(W6END[3]),
    .X(net80));
 sky130_fd_sc_hd__dlymetal6s2s_1 input81 (.A(W6END[4]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(W6END[5]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(W6END[6]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(W6END[7]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(W6END[8]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(W6END[9]),
    .X(net86));
 sky130_fd_sc_hd__dlymetal6s2s_1 input87 (.A(WW4END[0]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(WW4END[10]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(WW4END[11]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(FrameData[15]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input90 (.A(WW4END[12]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(WW4END[13]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(WW4END[14]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(WW4END[15]),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(WW4END[1]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(WW4END[2]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(WW4END[3]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(WW4END[4]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(WW4END[5]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(WW4END[6]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(A_I_top));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(A_T_top));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(A_config_C_bit0));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(A_config_C_bit1));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(A_config_C_bit2));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(A_config_C_bit3));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(B_I_top));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(B_T_top));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(B_config_C_bit0));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(B_config_C_bit1));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(B_config_C_bit2));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(B_config_C_bit3));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net134),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net146),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net159),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output167 (.A(net167),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net170),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net172),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net175),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net176),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net177),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__clkbuf_4 output183 (.A(net183),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output185 (.A(net185),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output186 (.A(net186),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output188 (.A(net188),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output189 (.A(net189),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output190 (.A(net190),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output191 (.A(net191),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output192 (.A(net192),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output193 (.A(net193),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output194 (.A(net194),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net199),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output201 (.A(net201),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output203 (.A(net203),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output204 (.A(net204),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output205 (.A(net205),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output207 (.A(net207),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output209 (.A(net209),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_1 output215 (.A(net215),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0/_0_  (.A(net35),
    .X(\FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__buf_1 \strobe_inbuf_1/_0_  (.A(net46),
    .X(\FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_10/_0_  (.A(net36),
    .X(\FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_11/_0_  (.A(net37),
    .X(\FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_12/_0_  (.A(net38),
    .X(\FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_13/_0_  (.A(net39),
    .X(\FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_14/_0_  (.A(net40),
    .X(\FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_15/_0_  (.A(net41),
    .X(\FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_16/_0_  (.A(net42),
    .X(\FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_17/_0_  (.A(net43),
    .X(\FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_18/_0_  (.A(net44),
    .X(\FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_19/_0_  (.A(net45),
    .X(\FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2/_0_  (.A(net47),
    .X(\FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__buf_1 \strobe_inbuf_3/_0_  (.A(net48),
    .X(\FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4/_0_  (.A(net49),
    .X(\FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_5/_0_  (.A(net50),
    .X(\FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6/_0_  (.A(net51),
    .X(\FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_7/_0_  (.A(net52),
    .X(\FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_8/_0_  (.A(net53),
    .X(\FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_9/_0_  (.A(net54),
    .X(\FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0/_0_  (.A(\FrameStrobe_O_i[0] ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1/_0_  (.A(\FrameStrobe_O_i[1] ),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10/_0_  (.A(\FrameStrobe_O_i[10] ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11/_0_  (.A(\FrameStrobe_O_i[11] ),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12/_0_  (.A(\FrameStrobe_O_i[12] ),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13/_0_  (.A(\FrameStrobe_O_i[13] ),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14/_0_  (.A(\FrameStrobe_O_i[14] ),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15/_0_  (.A(\FrameStrobe_O_i[15] ),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16/_0_  (.A(\FrameStrobe_O_i[16] ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17/_0_  (.A(\FrameStrobe_O_i[17] ),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18/_0_  (.A(\FrameStrobe_O_i[18] ),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19/_0_  (.A(\FrameStrobe_O_i[19] ),
    .X(net205));
 sky130_fd_sc_hd__buf_1 \strobe_outbuf_2/_0_  (.A(\FrameStrobe_O_i[2] ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3/_0_  (.A(\FrameStrobe_O_i[3] ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4/_0_  (.A(\FrameStrobe_O_i[4] ),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5/_0_  (.A(\FrameStrobe_O_i[5] ),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6/_0_  (.A(\FrameStrobe_O_i[6] ),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7/_0_  (.A(\FrameStrobe_O_i[7] ),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8/_0_  (.A(\FrameStrobe_O_i[8] ),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9/_0_  (.A(\FrameStrobe_O_i[9] ),
    .X(net214));
endmodule

