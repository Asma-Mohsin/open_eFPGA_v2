magic
tech sky130A
magscale 1 2
timestamp 1733618559
<< viali >>
rect 1593 8585 1627 8619
rect 3525 8585 3559 8619
rect 5457 8585 5491 8619
rect 7757 8585 7791 8619
rect 9689 8585 9723 8619
rect 11989 8585 12023 8619
rect 14289 8585 14323 8619
rect 16221 8585 16255 8619
rect 18153 8585 18187 8619
rect 20453 8585 20487 8619
rect 22569 8585 22603 8619
rect 24685 8585 24719 8619
rect 27169 8585 27203 8619
rect 28917 8585 28951 8619
rect 31033 8585 31067 8619
rect 32965 8585 32999 8619
rect 35265 8585 35299 8619
rect 37473 8585 37507 8619
rect 39497 8585 39531 8619
rect 41613 8585 41647 8619
rect 43085 8585 43119 8619
rect 1501 8449 1535 8483
rect 3341 8449 3375 8483
rect 5365 8449 5399 8483
rect 7573 8449 7607 8483
rect 9229 8449 9263 8483
rect 9597 8449 9631 8483
rect 11805 8449 11839 8483
rect 14197 8449 14231 8483
rect 16037 8449 16071 8483
rect 18061 8449 18095 8483
rect 20269 8449 20303 8483
rect 22385 8449 22419 8483
rect 24501 8449 24535 8483
rect 26985 8449 27019 8483
rect 28733 8449 28767 8483
rect 30849 8449 30883 8483
rect 32873 8449 32907 8483
rect 35081 8449 35115 8483
rect 37381 8449 37415 8483
rect 39313 8449 39347 8483
rect 41521 8449 41555 8483
rect 42901 8449 42935 8483
rect 2237 8313 2271 8347
rect 28181 3145 28215 3179
rect 29193 3145 29227 3179
rect 21465 3009 21499 3043
rect 22017 3009 22051 3043
rect 25605 3009 25639 3043
rect 27537 3009 27571 3043
rect 27813 3009 27847 3043
rect 28089 3009 28123 3043
rect 28365 3009 28399 3043
rect 29377 3009 29411 3043
rect 29745 3009 29779 3043
rect 27905 2873 27939 2907
rect 29561 2873 29595 2907
rect 21281 2805 21315 2839
rect 21833 2805 21867 2839
rect 25421 2805 25455 2839
rect 27353 2805 27387 2839
rect 27629 2805 27663 2839
rect 15301 2601 15335 2635
rect 15853 2601 15887 2635
rect 17233 2601 17267 2635
rect 18429 2601 18463 2635
rect 22385 2601 22419 2635
rect 22753 2601 22787 2635
rect 25973 2601 26007 2635
rect 27353 2601 27387 2635
rect 27813 2601 27847 2635
rect 28181 2601 28215 2635
rect 30205 2601 30239 2635
rect 31125 2601 31159 2635
rect 33241 2601 33275 2635
rect 35817 2601 35851 2635
rect 37565 2601 37599 2635
rect 39221 2601 39255 2635
rect 40509 2601 40543 2635
rect 42441 2601 42475 2635
rect 15577 2533 15611 2567
rect 16681 2533 16715 2567
rect 18337 2533 18371 2567
rect 19533 2533 19567 2567
rect 20453 2533 20487 2567
rect 20729 2533 20763 2567
rect 23213 2533 23247 2567
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 17049 2397 17083 2431
rect 17601 2397 17635 2431
rect 18153 2397 18187 2431
rect 18613 2397 18647 2431
rect 18981 2397 19015 2431
rect 19349 2397 19383 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 20361 2397 20395 2431
rect 20637 2397 20671 2431
rect 20913 2397 20947 2431
rect 21005 2397 21039 2431
rect 21741 2397 21775 2431
rect 22109 2397 22143 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 22937 2397 22971 2431
rect 23029 2397 23063 2431
rect 23489 2397 23523 2431
rect 25053 2397 25087 2431
rect 25145 2397 25179 2431
rect 25605 2397 25639 2431
rect 25881 2397 25915 2431
rect 26157 2397 26191 2431
rect 26433 2397 26467 2431
rect 26709 2397 26743 2431
rect 26985 2397 27019 2431
rect 27261 2397 27295 2431
rect 27537 2397 27571 2431
rect 27629 2397 27663 2431
rect 28549 2397 28583 2431
rect 28825 2397 28859 2431
rect 29101 2397 29135 2431
rect 29377 2397 29411 2431
rect 29745 2397 29779 2431
rect 30113 2397 30147 2431
rect 30389 2397 30423 2431
rect 31309 2397 31343 2431
rect 31401 2397 31435 2431
rect 33425 2397 33459 2431
rect 34805 2397 34839 2431
rect 36001 2397 36035 2431
rect 37749 2397 37783 2431
rect 39405 2397 39439 2431
rect 40693 2397 40727 2431
rect 42625 2397 42659 2431
rect 28089 2329 28123 2363
rect 16405 2261 16439 2295
rect 17417 2261 17451 2295
rect 18797 2261 18831 2295
rect 19809 2261 19843 2295
rect 19901 2261 19935 2295
rect 20177 2261 20211 2295
rect 21189 2261 21223 2295
rect 21557 2261 21591 2295
rect 21925 2261 21959 2295
rect 22477 2261 22511 2295
rect 23305 2261 23339 2295
rect 24869 2261 24903 2295
rect 25329 2261 25363 2295
rect 25421 2261 25455 2295
rect 25697 2261 25731 2295
rect 26249 2261 26283 2295
rect 26525 2261 26559 2295
rect 26801 2261 26835 2295
rect 27077 2261 27111 2295
rect 28365 2261 28399 2295
rect 28641 2261 28675 2295
rect 28917 2261 28951 2295
rect 29193 2261 29227 2295
rect 29561 2261 29595 2295
rect 30573 2261 30607 2295
rect 31585 2261 31619 2295
rect 34897 2261 34931 2295
rect 9321 2057 9355 2091
rect 14289 2057 14323 2091
rect 14841 2057 14875 2091
rect 15669 2057 15703 2091
rect 15945 2057 15979 2091
rect 17325 2057 17359 2091
rect 17601 2057 17635 2091
rect 19993 2057 20027 2091
rect 23213 2057 23247 2091
rect 23765 2057 23799 2091
rect 24041 2057 24075 2091
rect 27997 2057 28031 2091
rect 30757 2057 30791 2091
rect 31769 2057 31803 2091
rect 34529 2057 34563 2091
rect 35449 2057 35483 2091
rect 36461 2057 36495 2091
rect 37473 2057 37507 2091
rect 37933 2057 37967 2091
rect 38577 2057 38611 2091
rect 39773 2057 39807 2091
rect 20545 1989 20579 2023
rect 21281 1989 21315 2023
rect 22201 1989 22235 2023
rect 25789 1989 25823 2023
rect 26341 1989 26375 2023
rect 27905 1989 27939 2023
rect 28457 1989 28491 2023
rect 29009 1989 29043 2023
rect 29561 1989 29595 2023
rect 30113 1989 30147 2023
rect 30665 1989 30699 2023
rect 32229 1989 32263 2023
rect 9137 1921 9171 1955
rect 14105 1921 14139 1955
rect 14565 1921 14599 1955
rect 14657 1921 14691 1955
rect 14933 1921 14967 1955
rect 15209 1921 15243 1955
rect 15485 1921 15519 1955
rect 15761 1921 15795 1955
rect 16037 1921 16071 1955
rect 16313 1921 16347 1955
rect 16865 1921 16899 1955
rect 17141 1921 17175 1955
rect 17417 1921 17451 1955
rect 17877 1921 17911 1955
rect 18153 1945 18187 1979
rect 18245 1921 18279 1955
rect 18705 1921 18739 1955
rect 18981 1921 19015 1955
rect 19257 1921 19291 1955
rect 19533 1921 19567 1955
rect 19717 1921 19751 1955
rect 20361 1921 20395 1955
rect 22017 1921 22051 1955
rect 22661 1921 22695 1955
rect 23397 1921 23431 1955
rect 23673 1921 23707 1955
rect 23949 1921 23983 1955
rect 24225 1921 24259 1955
rect 24409 1921 24443 1955
rect 24961 1921 24995 1955
rect 25237 1921 25271 1955
rect 25513 1921 25547 1955
rect 27169 1921 27203 1955
rect 27721 1921 27755 1955
rect 31217 1921 31251 1955
rect 31953 1921 31987 1955
rect 32781 1921 32815 1955
rect 33333 1921 33367 1955
rect 33885 1921 33919 1955
rect 34989 1921 35023 1955
rect 35633 1921 35667 1955
rect 36645 1921 36679 1955
rect 36737 1921 36771 1955
rect 37657 1921 37691 1955
rect 38117 1921 38151 1955
rect 38761 1921 38795 1955
rect 39957 1921 39991 1955
rect 40233 1921 40267 1955
rect 30389 1853 30423 1887
rect 14381 1785 14415 1819
rect 15117 1785 15151 1819
rect 15393 1785 15427 1819
rect 16221 1785 16255 1819
rect 18429 1785 18463 1819
rect 18797 1785 18831 1819
rect 20177 1785 20211 1819
rect 20729 1785 20763 1819
rect 23489 1785 23523 1819
rect 25329 1785 25363 1819
rect 36921 1785 36955 1819
rect 40049 1785 40083 1819
rect 16497 1717 16531 1751
rect 17049 1717 17083 1751
rect 17693 1717 17727 1751
rect 17969 1717 18003 1751
rect 18521 1717 18555 1751
rect 19073 1717 19107 1751
rect 19349 1717 19383 1751
rect 21373 1717 21407 1751
rect 21833 1717 21867 1751
rect 22293 1717 22327 1751
rect 22845 1717 22879 1751
rect 24593 1717 24627 1751
rect 24777 1717 24811 1751
rect 25053 1717 25087 1751
rect 25881 1717 25915 1751
rect 26433 1717 26467 1751
rect 27537 1717 27571 1751
rect 28549 1717 28583 1751
rect 29101 1717 29135 1751
rect 29653 1717 29687 1751
rect 31309 1717 31343 1751
rect 32321 1717 32355 1751
rect 32873 1717 32907 1751
rect 33425 1717 33459 1751
rect 33977 1717 34011 1751
rect 35081 1717 35115 1751
rect 5917 1513 5951 1547
rect 9689 1513 9723 1547
rect 11069 1513 11103 1547
rect 11345 1513 11379 1547
rect 12817 1513 12851 1547
rect 14105 1513 14139 1547
rect 15485 1513 15519 1547
rect 17049 1513 17083 1547
rect 17509 1513 17543 1547
rect 23673 1513 23707 1547
rect 24961 1513 24995 1547
rect 25513 1513 25547 1547
rect 27721 1513 27755 1547
rect 28825 1513 28859 1547
rect 29193 1513 29227 1547
rect 31401 1513 31435 1547
rect 32873 1513 32907 1547
rect 33977 1513 34011 1547
rect 35817 1513 35851 1547
rect 36369 1513 36403 1547
rect 37473 1513 37507 1547
rect 39865 1513 39899 1547
rect 41521 1513 41555 1547
rect 41797 1513 41831 1547
rect 5365 1445 5399 1479
rect 6837 1445 6871 1479
rect 14657 1445 14691 1479
rect 16037 1445 16071 1479
rect 20913 1445 20947 1479
rect 27261 1445 27295 1479
rect 30941 1445 30975 1479
rect 31769 1445 31803 1479
rect 32505 1445 32539 1479
rect 34345 1445 34379 1479
rect 37749 1445 37783 1479
rect 40969 1445 41003 1479
rect 41245 1445 41279 1479
rect 20453 1377 20487 1411
rect 22385 1377 22419 1411
rect 29929 1377 29963 1411
rect 4629 1309 4663 1343
rect 4905 1309 4939 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 6929 1309 6963 1343
rect 7205 1309 7239 1343
rect 7481 1309 7515 1343
rect 7757 1309 7791 1343
rect 8033 1309 8067 1343
rect 8309 1309 8343 1343
rect 8585 1309 8619 1343
rect 8953 1309 8987 1343
rect 9229 1309 9263 1343
rect 9505 1309 9539 1343
rect 9965 1309 9999 1343
rect 10057 1309 10091 1343
rect 10333 1309 10367 1343
rect 10609 1309 10643 1343
rect 10885 1309 10919 1343
rect 11161 1309 11195 1343
rect 11529 1309 11563 1343
rect 11805 1309 11839 1343
rect 12081 1309 12115 1343
rect 12357 1309 12391 1343
rect 12633 1309 12667 1343
rect 12909 1309 12943 1343
rect 13185 1309 13219 1343
rect 13461 1309 13495 1343
rect 13921 1309 13955 1343
rect 14289 1309 14323 1343
rect 14565 1309 14599 1343
rect 14841 1309 14875 1343
rect 15117 1309 15151 1343
rect 15393 1309 15427 1343
rect 15669 1309 15703 1343
rect 15945 1309 15979 1343
rect 16221 1309 16255 1343
rect 16497 1309 16531 1343
rect 16865 1309 16899 1343
rect 17417 1309 17451 1343
rect 17693 1309 17727 1343
rect 17969 1309 18003 1343
rect 18061 1309 18095 1343
rect 18521 1309 18555 1343
rect 18613 1309 18647 1343
rect 19073 1309 19107 1343
rect 19349 1309 19383 1343
rect 19717 1309 19751 1343
rect 20177 1309 20211 1343
rect 21373 1309 21407 1343
rect 22109 1309 22143 1343
rect 22753 1309 22787 1343
rect 23121 1309 23155 1343
rect 23581 1309 23615 1343
rect 24409 1309 24443 1343
rect 25421 1309 25455 1343
rect 26433 1309 26467 1343
rect 27629 1309 27663 1343
rect 28733 1309 28767 1343
rect 29377 1309 29411 1343
rect 30205 1309 30239 1343
rect 31953 1309 31987 1343
rect 34529 1309 34563 1343
rect 35725 1309 35759 1343
rect 36737 1309 36771 1343
rect 37289 1309 37323 1343
rect 37565 1309 37599 1343
rect 37841 1309 37875 1343
rect 38117 1309 38151 1343
rect 38393 1309 38427 1343
rect 38669 1309 38703 1343
rect 38945 1309 38979 1343
rect 39221 1309 39255 1343
rect 39497 1309 39531 1343
rect 40049 1309 40083 1343
rect 40325 1309 40359 1343
rect 40601 1309 40635 1343
rect 40877 1309 40911 1343
rect 41153 1309 41187 1343
rect 41429 1309 41463 1343
rect 41705 1309 41739 1343
rect 41981 1309 42015 1343
rect 20729 1241 20763 1275
rect 24869 1241 24903 1275
rect 25973 1241 26007 1275
rect 27077 1241 27111 1275
rect 28181 1241 28215 1275
rect 29653 1241 29687 1275
rect 30757 1241 30791 1275
rect 31309 1241 31343 1275
rect 32229 1241 32263 1275
rect 32781 1241 32815 1275
rect 33885 1241 33919 1275
rect 34805 1241 34839 1275
rect 35449 1241 35483 1275
rect 36277 1241 36311 1275
rect 4813 1173 4847 1207
rect 5089 1173 5123 1207
rect 5641 1173 5675 1207
rect 6193 1173 6227 1207
rect 6561 1173 6595 1207
rect 7113 1173 7147 1207
rect 7389 1173 7423 1207
rect 7665 1173 7699 1207
rect 7941 1173 7975 1207
rect 8217 1173 8251 1207
rect 8493 1173 8527 1207
rect 8769 1173 8803 1207
rect 9137 1173 9171 1207
rect 9413 1173 9447 1207
rect 9781 1173 9815 1207
rect 10241 1173 10275 1207
rect 10517 1173 10551 1207
rect 10793 1173 10827 1207
rect 11713 1173 11747 1207
rect 11989 1173 12023 1207
rect 12265 1173 12299 1207
rect 12541 1173 12575 1207
rect 13093 1173 13127 1207
rect 13369 1173 13403 1207
rect 13645 1173 13679 1207
rect 13737 1173 13771 1207
rect 14381 1173 14415 1207
rect 14933 1173 14967 1207
rect 15209 1173 15243 1207
rect 15761 1173 15795 1207
rect 16313 1173 16347 1207
rect 17233 1173 17267 1207
rect 17785 1173 17819 1207
rect 18245 1173 18279 1207
rect 18337 1173 18371 1207
rect 18797 1173 18831 1207
rect 18889 1173 18923 1207
rect 19533 1173 19567 1207
rect 19901 1173 19935 1207
rect 21557 1173 21591 1207
rect 22937 1173 22971 1207
rect 23305 1173 23339 1207
rect 24593 1173 24627 1207
rect 26065 1173 26099 1207
rect 26617 1173 26651 1207
rect 28273 1173 28307 1207
rect 30297 1173 30331 1207
rect 33425 1173 33459 1207
rect 34897 1173 34931 1207
rect 36921 1173 36955 1207
rect 38025 1173 38059 1207
rect 38301 1173 38335 1207
rect 38577 1173 38611 1207
rect 38853 1173 38887 1207
rect 39129 1173 39163 1207
rect 39405 1173 39439 1207
rect 39681 1173 39715 1207
rect 40141 1173 40175 1207
rect 40417 1173 40451 1207
rect 40693 1173 40727 1207
<< metal1 >>
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 25314 8820 25320 8832
rect 7616 8792 25320 8820
rect 7616 8780 7622 8792
rect 25314 8780 25320 8792
rect 25372 8780 25378 8832
rect 1104 8730 43675 8752
rect 1104 8678 11552 8730
rect 11604 8678 11616 8730
rect 11668 8678 11680 8730
rect 11732 8678 11744 8730
rect 11796 8678 11808 8730
rect 11860 8678 22155 8730
rect 22207 8678 22219 8730
rect 22271 8678 22283 8730
rect 22335 8678 22347 8730
rect 22399 8678 22411 8730
rect 22463 8678 32758 8730
rect 32810 8678 32822 8730
rect 32874 8678 32886 8730
rect 32938 8678 32950 8730
rect 33002 8678 33014 8730
rect 33066 8678 43361 8730
rect 43413 8678 43425 8730
rect 43477 8678 43489 8730
rect 43541 8678 43553 8730
rect 43605 8678 43617 8730
rect 43669 8678 43675 8730
rect 1104 8656 43675 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1268 8588 1593 8616
rect 1268 8576 1274 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3292 8588 3525 8616
rect 3292 8576 3298 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7524 8588 7757 8616
rect 7524 8576 7530 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 9640 8588 9689 8616
rect 9640 8576 9646 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11940 8588 11989 8616
rect 11940 8576 11946 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 11977 8579 12035 8585
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13872 8588 14289 8616
rect 13872 8576 13878 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15988 8588 16221 8616
rect 15988 8576 15994 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 18138 8576 18144 8628
rect 18196 8576 18202 8628
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20220 8588 20453 8616
rect 20220 8576 20226 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 20441 8579 20499 8585
rect 22554 8576 22560 8628
rect 22612 8576 22618 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24673 8619 24731 8625
rect 24673 8616 24685 8619
rect 24452 8588 24685 8616
rect 24452 8576 24458 8588
rect 24673 8585 24685 8588
rect 24719 8585 24731 8619
rect 24673 8579 24731 8585
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 26568 8588 27169 8616
rect 26568 8576 26574 8588
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 27157 8579 27215 8585
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 28905 8619 28963 8625
rect 28905 8616 28917 8619
rect 28684 8588 28917 8616
rect 28684 8576 28690 8588
rect 28905 8585 28917 8588
rect 28951 8585 28963 8619
rect 28905 8579 28963 8585
rect 30742 8576 30748 8628
rect 30800 8616 30806 8628
rect 31021 8619 31079 8625
rect 31021 8616 31033 8619
rect 30800 8588 31033 8616
rect 30800 8576 30806 8588
rect 31021 8585 31033 8588
rect 31067 8585 31079 8619
rect 31021 8579 31079 8585
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 32953 8619 33011 8625
rect 32953 8616 32965 8619
rect 32732 8588 32965 8616
rect 32732 8576 32738 8588
rect 32953 8585 32965 8588
rect 32999 8585 33011 8619
rect 32953 8579 33011 8585
rect 34974 8576 34980 8628
rect 35032 8616 35038 8628
rect 35253 8619 35311 8625
rect 35253 8616 35265 8619
rect 35032 8588 35265 8616
rect 35032 8576 35038 8588
rect 35253 8585 35265 8588
rect 35299 8585 35311 8619
rect 35253 8579 35311 8585
rect 37090 8576 37096 8628
rect 37148 8616 37154 8628
rect 37461 8619 37519 8625
rect 37461 8616 37473 8619
rect 37148 8588 37473 8616
rect 37148 8576 37154 8588
rect 37461 8585 37473 8588
rect 37507 8585 37519 8619
rect 37461 8579 37519 8585
rect 39206 8576 39212 8628
rect 39264 8616 39270 8628
rect 39485 8619 39543 8625
rect 39485 8616 39497 8619
rect 39264 8588 39497 8616
rect 39264 8576 39270 8588
rect 39485 8585 39497 8588
rect 39531 8585 39543 8619
rect 39485 8579 39543 8585
rect 41322 8576 41328 8628
rect 41380 8616 41386 8628
rect 41601 8619 41659 8625
rect 41601 8616 41613 8619
rect 41380 8588 41613 8616
rect 41380 8576 41386 8588
rect 41601 8585 41613 8588
rect 41647 8585 41659 8619
rect 41601 8579 41659 8585
rect 43073 8619 43131 8625
rect 43073 8585 43085 8619
rect 43119 8616 43131 8619
rect 43254 8616 43260 8628
rect 43119 8588 43260 8616
rect 43119 8585 43131 8588
rect 43073 8579 43131 8585
rect 43254 8576 43260 8588
rect 43312 8576 43318 8628
rect 28166 8548 28172 8560
rect 3344 8520 28172 8548
rect 3344 8489 3372 8520
rect 28166 8508 28172 8520
rect 28224 8508 28230 8560
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 3329 8483 3387 8489
rect 1535 8452 2268 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 2240 8356 2268 8452
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5399 8452 6914 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 2222 8304 2228 8356
rect 2280 8304 2286 8356
rect 6886 8344 6914 8452
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9582 8480 9588 8492
rect 9263 8452 9588 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8480 11851 8483
rect 14090 8480 14096 8492
rect 11839 8452 14096 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 15286 8480 15292 8492
rect 14231 8452 15292 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 18046 8440 18052 8492
rect 18104 8440 18110 8492
rect 20254 8440 20260 8492
rect 20312 8440 20318 8492
rect 22373 8483 22431 8489
rect 22373 8449 22385 8483
rect 22419 8480 22431 8483
rect 22738 8480 22744 8492
rect 22419 8452 22744 8480
rect 22419 8449 22431 8452
rect 22373 8443 22431 8449
rect 22738 8440 22744 8452
rect 22796 8440 22802 8492
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8480 24547 8483
rect 24854 8480 24860 8492
rect 24535 8452 24860 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 26970 8440 26976 8492
rect 27028 8440 27034 8492
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 30834 8440 30840 8492
rect 30892 8440 30898 8492
rect 32861 8483 32919 8489
rect 32861 8449 32873 8483
rect 32907 8480 32919 8483
rect 33226 8480 33232 8492
rect 32907 8452 33232 8480
rect 32907 8449 32919 8452
rect 32861 8443 32919 8449
rect 33226 8440 33232 8452
rect 33284 8440 33290 8492
rect 35066 8440 35072 8492
rect 35124 8440 35130 8492
rect 37366 8440 37372 8492
rect 37424 8440 37430 8492
rect 39298 8440 39304 8492
rect 39356 8440 39362 8492
rect 40494 8440 40500 8492
rect 40552 8480 40558 8492
rect 41509 8483 41567 8489
rect 41509 8480 41521 8483
rect 40552 8452 41521 8480
rect 40552 8440 40558 8452
rect 41509 8449 41521 8452
rect 41555 8449 41567 8483
rect 41509 8443 41567 8449
rect 42886 8440 42892 8492
rect 42944 8440 42950 8492
rect 23198 8412 23204 8424
rect 14200 8384 23204 8412
rect 14200 8344 14228 8384
rect 23198 8372 23204 8384
rect 23256 8372 23262 8424
rect 6886 8316 14228 8344
rect 14274 8304 14280 8356
rect 14332 8344 14338 8356
rect 22554 8344 22560 8356
rect 14332 8316 22560 8344
rect 14332 8304 14338 8316
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 1104 8186 43516 8208
rect 1104 8134 6251 8186
rect 6303 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 16854 8186
rect 16906 8134 16918 8186
rect 16970 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 27457 8186
rect 27509 8134 27521 8186
rect 27573 8134 27585 8186
rect 27637 8134 27649 8186
rect 27701 8134 27713 8186
rect 27765 8134 38060 8186
rect 38112 8134 38124 8186
rect 38176 8134 38188 8186
rect 38240 8134 38252 8186
rect 38304 8134 38316 8186
rect 38368 8134 43516 8186
rect 1104 8112 43516 8134
rect 1104 7642 43675 7664
rect 1104 7590 11552 7642
rect 11604 7590 11616 7642
rect 11668 7590 11680 7642
rect 11732 7590 11744 7642
rect 11796 7590 11808 7642
rect 11860 7590 22155 7642
rect 22207 7590 22219 7642
rect 22271 7590 22283 7642
rect 22335 7590 22347 7642
rect 22399 7590 22411 7642
rect 22463 7590 32758 7642
rect 32810 7590 32822 7642
rect 32874 7590 32886 7642
rect 32938 7590 32950 7642
rect 33002 7590 33014 7642
rect 33066 7590 43361 7642
rect 43413 7590 43425 7642
rect 43477 7590 43489 7642
rect 43541 7590 43553 7642
rect 43605 7590 43617 7642
rect 43669 7590 43675 7642
rect 1104 7568 43675 7590
rect 1104 7098 43516 7120
rect 1104 7046 6251 7098
rect 6303 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 16854 7098
rect 16906 7046 16918 7098
rect 16970 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 27457 7098
rect 27509 7046 27521 7098
rect 27573 7046 27585 7098
rect 27637 7046 27649 7098
rect 27701 7046 27713 7098
rect 27765 7046 38060 7098
rect 38112 7046 38124 7098
rect 38176 7046 38188 7098
rect 38240 7046 38252 7098
rect 38304 7046 38316 7098
rect 38368 7046 43516 7098
rect 1104 7024 43516 7046
rect 1104 6554 43675 6576
rect 1104 6502 11552 6554
rect 11604 6502 11616 6554
rect 11668 6502 11680 6554
rect 11732 6502 11744 6554
rect 11796 6502 11808 6554
rect 11860 6502 22155 6554
rect 22207 6502 22219 6554
rect 22271 6502 22283 6554
rect 22335 6502 22347 6554
rect 22399 6502 22411 6554
rect 22463 6502 32758 6554
rect 32810 6502 32822 6554
rect 32874 6502 32886 6554
rect 32938 6502 32950 6554
rect 33002 6502 33014 6554
rect 33066 6502 43361 6554
rect 43413 6502 43425 6554
rect 43477 6502 43489 6554
rect 43541 6502 43553 6554
rect 43605 6502 43617 6554
rect 43669 6502 43675 6554
rect 1104 6480 43675 6502
rect 1104 6010 43516 6032
rect 1104 5958 6251 6010
rect 6303 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 16854 6010
rect 16906 5958 16918 6010
rect 16970 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 27457 6010
rect 27509 5958 27521 6010
rect 27573 5958 27585 6010
rect 27637 5958 27649 6010
rect 27701 5958 27713 6010
rect 27765 5958 38060 6010
rect 38112 5958 38124 6010
rect 38176 5958 38188 6010
rect 38240 5958 38252 6010
rect 38304 5958 38316 6010
rect 38368 5958 43516 6010
rect 1104 5936 43516 5958
rect 1104 5466 43675 5488
rect 1104 5414 11552 5466
rect 11604 5414 11616 5466
rect 11668 5414 11680 5466
rect 11732 5414 11744 5466
rect 11796 5414 11808 5466
rect 11860 5414 22155 5466
rect 22207 5414 22219 5466
rect 22271 5414 22283 5466
rect 22335 5414 22347 5466
rect 22399 5414 22411 5466
rect 22463 5414 32758 5466
rect 32810 5414 32822 5466
rect 32874 5414 32886 5466
rect 32938 5414 32950 5466
rect 33002 5414 33014 5466
rect 33066 5414 43361 5466
rect 43413 5414 43425 5466
rect 43477 5414 43489 5466
rect 43541 5414 43553 5466
rect 43605 5414 43617 5466
rect 43669 5414 43675 5466
rect 1104 5392 43675 5414
rect 1104 4922 43516 4944
rect 1104 4870 6251 4922
rect 6303 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 16854 4922
rect 16906 4870 16918 4922
rect 16970 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 27457 4922
rect 27509 4870 27521 4922
rect 27573 4870 27585 4922
rect 27637 4870 27649 4922
rect 27701 4870 27713 4922
rect 27765 4870 38060 4922
rect 38112 4870 38124 4922
rect 38176 4870 38188 4922
rect 38240 4870 38252 4922
rect 38304 4870 38316 4922
rect 38368 4870 43516 4922
rect 1104 4848 43516 4870
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 23382 4536 23388 4548
rect 8628 4508 23388 4536
rect 8628 4496 8634 4508
rect 23382 4496 23388 4508
rect 23440 4496 23446 4548
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 23658 4468 23664 4480
rect 9272 4440 23664 4468
rect 9272 4428 9278 4440
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 1104 4378 43675 4400
rect 1104 4326 11552 4378
rect 11604 4326 11616 4378
rect 11668 4326 11680 4378
rect 11732 4326 11744 4378
rect 11796 4326 11808 4378
rect 11860 4326 22155 4378
rect 22207 4326 22219 4378
rect 22271 4326 22283 4378
rect 22335 4326 22347 4378
rect 22399 4326 22411 4378
rect 22463 4326 32758 4378
rect 32810 4326 32822 4378
rect 32874 4326 32886 4378
rect 32938 4326 32950 4378
rect 33002 4326 33014 4378
rect 33066 4326 43361 4378
rect 43413 4326 43425 4378
rect 43477 4326 43489 4378
rect 43541 4326 43553 4378
rect 43605 4326 43617 4378
rect 43669 4326 43675 4378
rect 1104 4304 43675 4326
rect 11330 4224 11336 4276
rect 11388 4264 11394 4276
rect 28074 4264 28080 4276
rect 11388 4236 28080 4264
rect 11388 4224 11394 4236
rect 28074 4224 28080 4236
rect 28132 4224 28138 4276
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 25130 4196 25136 4208
rect 7248 4168 25136 4196
rect 7248 4156 7254 4168
rect 25130 4156 25136 4168
rect 25188 4156 25194 4208
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 28350 3924 28356 3936
rect 12032 3896 28356 3924
rect 12032 3884 12038 3896
rect 28350 3884 28356 3896
rect 28408 3884 28414 3936
rect 1104 3834 43516 3856
rect 1104 3782 6251 3834
rect 6303 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 16854 3834
rect 16906 3782 16918 3834
rect 16970 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 27457 3834
rect 27509 3782 27521 3834
rect 27573 3782 27585 3834
rect 27637 3782 27649 3834
rect 27701 3782 27713 3834
rect 27765 3782 38060 3834
rect 38112 3782 38124 3834
rect 38176 3782 38188 3834
rect 38240 3782 38252 3834
rect 38304 3782 38316 3834
rect 38368 3782 43516 3834
rect 1104 3760 43516 3782
rect 17954 3544 17960 3596
rect 18012 3584 18018 3596
rect 18012 3556 26188 3584
rect 18012 3544 18018 3556
rect 26160 3528 26188 3556
rect 36814 3544 36820 3596
rect 36872 3584 36878 3596
rect 38930 3584 38936 3596
rect 36872 3556 38936 3584
rect 36872 3544 36878 3556
rect 38930 3544 38936 3556
rect 38988 3544 38994 3596
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 25590 3516 25596 3528
rect 13688 3488 25596 3516
rect 13688 3476 13694 3488
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 26142 3476 26148 3528
rect 26200 3476 26206 3528
rect 38470 3476 38476 3528
rect 38528 3516 38534 3528
rect 40862 3516 40868 3528
rect 38528 3488 40868 3516
rect 38528 3476 38534 3488
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 16206 3408 16212 3460
rect 16264 3448 16270 3460
rect 30190 3448 30196 3460
rect 16264 3420 30196 3448
rect 16264 3408 16270 3420
rect 30190 3408 30196 3420
rect 30248 3408 30254 3460
rect 37826 3408 37832 3460
rect 37884 3448 37890 3460
rect 40310 3448 40316 3460
rect 37884 3420 40316 3448
rect 37884 3408 37890 3420
rect 40310 3408 40316 3420
rect 40368 3408 40374 3460
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 20438 3380 20444 3392
rect 8352 3352 20444 3380
rect 8352 3340 8358 3352
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 37182 3340 37188 3392
rect 37240 3380 37246 3392
rect 39482 3380 39488 3392
rect 37240 3352 39488 3380
rect 37240 3340 37246 3352
rect 39482 3340 39488 3352
rect 39540 3340 39546 3392
rect 1104 3290 43675 3312
rect 1104 3238 11552 3290
rect 11604 3238 11616 3290
rect 11668 3238 11680 3290
rect 11732 3238 11744 3290
rect 11796 3238 11808 3290
rect 11860 3238 22155 3290
rect 22207 3238 22219 3290
rect 22271 3238 22283 3290
rect 22335 3238 22347 3290
rect 22399 3238 22411 3290
rect 22463 3238 32758 3290
rect 32810 3238 32822 3290
rect 32874 3238 32886 3290
rect 32938 3238 32950 3290
rect 33002 3238 33014 3290
rect 33066 3238 43361 3290
rect 43413 3238 43425 3290
rect 43477 3238 43489 3290
rect 43541 3238 43553 3290
rect 43605 3238 43617 3290
rect 43669 3238 43675 3290
rect 1104 3216 43675 3238
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 23566 3176 23572 3188
rect 19024 3148 23572 3176
rect 19024 3136 19030 3148
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 28169 3179 28227 3185
rect 28169 3145 28181 3179
rect 28215 3145 28227 3179
rect 28169 3139 28227 3145
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 25682 3108 25688 3120
rect 17736 3080 25688 3108
rect 17736 3068 17742 3080
rect 25682 3068 25688 3080
rect 25740 3068 25746 3120
rect 28184 3108 28212 3139
rect 28718 3136 28724 3188
rect 28776 3176 28782 3188
rect 29181 3179 29239 3185
rect 29181 3176 29193 3179
rect 28776 3148 29193 3176
rect 28776 3136 28782 3148
rect 29181 3145 29193 3148
rect 29227 3145 29239 3179
rect 29181 3139 29239 3145
rect 37550 3136 37556 3188
rect 37608 3176 37614 3188
rect 40034 3176 40040 3188
rect 37608 3148 40040 3176
rect 37608 3136 37614 3148
rect 40034 3136 40040 3148
rect 40092 3136 40098 3188
rect 30098 3108 30104 3120
rect 28184 3080 30104 3108
rect 30098 3068 30104 3080
rect 30156 3068 30162 3120
rect 38010 3068 38016 3120
rect 38068 3108 38074 3120
rect 40586 3108 40592 3120
rect 38068 3080 40592 3108
rect 38068 3068 38074 3080
rect 40586 3068 40592 3080
rect 40644 3068 40650 3120
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 21453 3043 21511 3049
rect 21453 3040 21465 3043
rect 11020 3012 21465 3040
rect 11020 3000 11026 3012
rect 21453 3009 21465 3012
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22005 3043 22063 3049
rect 22005 3009 22017 3043
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 22020 2972 22048 3003
rect 25590 3000 25596 3052
rect 25648 3000 25654 3052
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 27798 3000 27804 3052
rect 27856 3000 27862 3052
rect 28074 3000 28080 3052
rect 28132 3000 28138 3052
rect 28350 3000 28356 3052
rect 28408 3000 28414 3052
rect 29365 3043 29423 3049
rect 29365 3009 29377 3043
rect 29411 3040 29423 3043
rect 29733 3043 29791 3049
rect 29411 3012 29592 3040
rect 29411 3009 29423 3012
rect 29365 3003 29423 3009
rect 26510 2972 26516 2984
rect 7892 2944 22048 2972
rect 22112 2944 26516 2972
rect 7892 2932 7898 2944
rect 15746 2864 15752 2916
rect 15804 2904 15810 2916
rect 17494 2904 17500 2916
rect 15804 2876 17500 2904
rect 15804 2864 15810 2876
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 18196 2876 19196 2904
rect 18196 2864 18202 2876
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 19058 2836 19064 2848
rect 15528 2808 19064 2836
rect 15528 2796 15534 2808
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 19168 2836 19196 2876
rect 20346 2864 20352 2916
rect 20404 2904 20410 2916
rect 22112 2904 22140 2944
rect 26510 2932 26516 2944
rect 26568 2932 26574 2984
rect 20404 2876 22140 2904
rect 27893 2907 27951 2913
rect 20404 2864 20410 2876
rect 27893 2873 27905 2907
rect 27939 2904 27951 2907
rect 29454 2904 29460 2916
rect 27939 2876 29460 2904
rect 27939 2873 27951 2876
rect 27893 2867 27951 2873
rect 29454 2864 29460 2876
rect 29512 2864 29518 2916
rect 29564 2913 29592 3012
rect 29733 3009 29745 3043
rect 29779 3040 29791 3043
rect 29779 3012 35894 3040
rect 29779 3009 29791 3012
rect 29733 3003 29791 3009
rect 29549 2907 29607 2913
rect 29549 2873 29561 2907
rect 29595 2873 29607 2907
rect 35866 2904 35894 3012
rect 38562 3000 38568 3052
rect 38620 3040 38626 3052
rect 41138 3040 41144 3052
rect 38620 3012 41144 3040
rect 38620 3000 38626 3012
rect 41138 3000 41144 3012
rect 41196 3000 41202 3052
rect 38378 2972 38384 2984
rect 37108 2944 38384 2972
rect 37108 2904 37136 2944
rect 38378 2932 38384 2944
rect 38436 2932 38442 2984
rect 35866 2876 37136 2904
rect 29549 2867 29607 2873
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 39206 2904 39212 2916
rect 37240 2876 39212 2904
rect 37240 2864 37246 2876
rect 39206 2864 39212 2876
rect 39264 2864 39270 2916
rect 21174 2836 21180 2848
rect 19168 2808 21180 2836
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21269 2839 21327 2845
rect 21269 2805 21281 2839
rect 21315 2836 21327 2839
rect 21726 2836 21732 2848
rect 21315 2808 21732 2836
rect 21315 2805 21327 2808
rect 21269 2799 21327 2805
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 21821 2839 21879 2845
rect 21821 2805 21833 2839
rect 21867 2836 21879 2839
rect 23474 2836 23480 2848
rect 21867 2808 23480 2836
rect 21867 2805 21879 2808
rect 21821 2799 21879 2805
rect 23474 2796 23480 2808
rect 23532 2796 23538 2848
rect 25409 2839 25467 2845
rect 25409 2805 25421 2839
rect 25455 2836 25467 2839
rect 26234 2836 26240 2848
rect 25455 2808 26240 2836
rect 25455 2805 25467 2808
rect 25409 2799 25467 2805
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 27338 2796 27344 2848
rect 27396 2796 27402 2848
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27798 2836 27804 2848
rect 27663 2808 27804 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28718 2796 28724 2848
rect 28776 2836 28782 2848
rect 30742 2836 30748 2848
rect 28776 2808 30748 2836
rect 28776 2796 28782 2808
rect 30742 2796 30748 2808
rect 30800 2796 30806 2848
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 38654 2836 38660 2848
rect 36412 2808 38660 2836
rect 36412 2796 36418 2808
rect 38654 2796 38660 2808
rect 38712 2836 38718 2848
rect 38712 2808 38759 2836
rect 38712 2796 38718 2808
rect 1104 2746 43516 2768
rect 1104 2694 6251 2746
rect 6303 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 16854 2746
rect 16906 2694 16918 2746
rect 16970 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 27457 2746
rect 27509 2694 27521 2746
rect 27573 2694 27585 2746
rect 27637 2694 27649 2746
rect 27701 2694 27713 2746
rect 27765 2694 38060 2746
rect 38112 2694 38124 2746
rect 38176 2694 38188 2746
rect 38240 2694 38252 2746
rect 38304 2694 38316 2746
rect 38368 2694 43516 2746
rect 1104 2672 43516 2694
rect 15286 2592 15292 2644
rect 15344 2592 15350 2644
rect 15746 2632 15752 2644
rect 15396 2604 15752 2632
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 15396 2564 15424 2604
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 16022 2632 16028 2644
rect 15887 2604 16028 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 17862 2632 17868 2644
rect 17267 2604 17868 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18046 2592 18052 2644
rect 18104 2632 18110 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 18104 2604 18429 2632
rect 18104 2592 18110 2604
rect 18417 2601 18429 2604
rect 18463 2601 18475 2635
rect 18417 2595 18475 2601
rect 22373 2635 22431 2641
rect 22373 2601 22385 2635
rect 22419 2632 22431 2635
rect 22554 2632 22560 2644
rect 22419 2604 22560 2632
rect 22419 2601 22431 2604
rect 22373 2595 22431 2601
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 22738 2592 22744 2644
rect 22796 2592 22802 2644
rect 25590 2632 25596 2644
rect 22848 2604 25596 2632
rect 11112 2536 15424 2564
rect 11112 2524 11118 2536
rect 15562 2524 15568 2576
rect 15620 2524 15626 2576
rect 16669 2567 16727 2573
rect 16669 2533 16681 2567
rect 16715 2533 16727 2567
rect 16669 2527 16727 2533
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 15286 2496 15292 2508
rect 13780 2468 15292 2496
rect 13780 2456 13786 2468
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 16482 2496 16488 2508
rect 15764 2468 16488 2496
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2428 15531 2431
rect 15562 2428 15568 2440
rect 15519 2400 15568 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15764 2437 15792 2468
rect 16482 2456 16488 2468
rect 16540 2456 16546 2508
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16684 2428 16712 2527
rect 16850 2524 16856 2576
rect 16908 2564 16914 2576
rect 17954 2564 17960 2576
rect 16908 2536 17960 2564
rect 16908 2524 16914 2536
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 18325 2567 18383 2573
rect 18325 2533 18337 2567
rect 18371 2533 18383 2567
rect 18325 2527 18383 2533
rect 19521 2567 19579 2573
rect 19521 2533 19533 2567
rect 19567 2564 19579 2567
rect 20070 2564 20076 2576
rect 19567 2536 20076 2564
rect 19567 2533 19579 2536
rect 19521 2527 19579 2533
rect 17218 2496 17224 2508
rect 16868 2468 17224 2496
rect 16071 2400 16712 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16868 2437 16896 2468
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18340 2496 18368 2527
rect 20070 2524 20076 2536
rect 20128 2524 20134 2576
rect 20254 2524 20260 2576
rect 20312 2564 20318 2576
rect 20441 2567 20499 2573
rect 20441 2564 20453 2567
rect 20312 2536 20453 2564
rect 20312 2524 20318 2536
rect 20441 2533 20453 2536
rect 20487 2533 20499 2567
rect 20441 2527 20499 2533
rect 20717 2567 20775 2573
rect 20717 2533 20729 2567
rect 20763 2533 20775 2567
rect 22848 2564 22876 2604
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 25884 2604 25973 2632
rect 25884 2576 25912 2604
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 25961 2595 26019 2601
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27341 2635 27399 2641
rect 27341 2632 27353 2635
rect 27212 2604 27353 2632
rect 27212 2592 27218 2604
rect 27341 2601 27353 2604
rect 27387 2601 27399 2635
rect 27341 2595 27399 2601
rect 27801 2635 27859 2641
rect 27801 2601 27813 2635
rect 27847 2632 27859 2635
rect 27890 2632 27896 2644
rect 27847 2604 27896 2632
rect 27847 2601 27859 2604
rect 27801 2595 27859 2601
rect 27890 2592 27896 2604
rect 27948 2592 27954 2644
rect 28166 2592 28172 2644
rect 28224 2592 28230 2644
rect 30190 2592 30196 2644
rect 30248 2592 30254 2644
rect 30834 2592 30840 2644
rect 30892 2632 30898 2644
rect 31113 2635 31171 2641
rect 31113 2632 31125 2635
rect 30892 2604 31125 2632
rect 30892 2592 30898 2604
rect 31113 2601 31125 2604
rect 31159 2601 31171 2635
rect 31113 2595 31171 2601
rect 33226 2592 33232 2644
rect 33284 2592 33290 2644
rect 35066 2592 35072 2644
rect 35124 2632 35130 2644
rect 35805 2635 35863 2641
rect 35805 2632 35817 2635
rect 35124 2604 35817 2632
rect 35124 2592 35130 2604
rect 35805 2601 35817 2604
rect 35851 2601 35863 2635
rect 35805 2595 35863 2601
rect 37366 2592 37372 2644
rect 37424 2632 37430 2644
rect 37553 2635 37611 2641
rect 37553 2632 37565 2635
rect 37424 2604 37565 2632
rect 37424 2592 37430 2604
rect 37553 2601 37565 2604
rect 37599 2601 37611 2635
rect 37553 2595 37611 2601
rect 39209 2635 39267 2641
rect 39209 2601 39221 2635
rect 39255 2632 39267 2635
rect 39298 2632 39304 2644
rect 39255 2604 39304 2632
rect 39255 2601 39267 2604
rect 39209 2595 39267 2601
rect 39298 2592 39304 2604
rect 39356 2592 39362 2644
rect 40494 2592 40500 2644
rect 40552 2592 40558 2644
rect 42429 2635 42487 2641
rect 42429 2601 42441 2635
rect 42475 2632 42487 2635
rect 42886 2632 42892 2644
rect 42475 2604 42892 2632
rect 42475 2601 42487 2604
rect 42429 2595 42487 2601
rect 42886 2592 42892 2604
rect 42944 2592 42950 2644
rect 20717 2527 20775 2533
rect 20824 2536 22876 2564
rect 18104 2468 18368 2496
rect 18524 2468 20576 2496
rect 18104 2456 18110 2468
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 17052 2360 17080 2391
rect 17310 2388 17316 2440
rect 17368 2428 17374 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17368 2400 17601 2428
rect 17368 2388 17374 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18414 2428 18420 2440
rect 18187 2400 18420 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18524 2360 18552 2468
rect 18601 2431 18659 2437
rect 18601 2397 18613 2431
rect 18647 2428 18659 2431
rect 18647 2400 18828 2428
rect 18647 2397 18659 2400
rect 18601 2391 18659 2397
rect 15252 2332 17080 2360
rect 17144 2332 18552 2360
rect 15252 2320 15258 2332
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 16298 2292 16304 2304
rect 14884 2264 16304 2292
rect 14884 2252 14890 2264
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 16393 2295 16451 2301
rect 16393 2261 16405 2295
rect 16439 2292 16451 2295
rect 16758 2292 16764 2304
rect 16439 2264 16764 2292
rect 16439 2261 16451 2264
rect 16393 2255 16451 2261
rect 16758 2252 16764 2264
rect 16816 2252 16822 2304
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 17144 2292 17172 2332
rect 16908 2264 17172 2292
rect 16908 2252 16914 2264
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 18800 2301 18828 2400
rect 18966 2388 18972 2440
rect 19024 2388 19030 2440
rect 19337 2431 19395 2437
rect 19337 2397 19349 2431
rect 19383 2428 19395 2431
rect 19383 2400 19564 2428
rect 19383 2397 19395 2400
rect 19337 2391 19395 2397
rect 19536 2360 19564 2400
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20162 2388 20168 2440
rect 20220 2428 20226 2440
rect 20349 2431 20407 2437
rect 20349 2428 20361 2431
rect 20220 2400 20361 2428
rect 20220 2388 20226 2400
rect 20349 2397 20361 2400
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 19702 2360 19708 2372
rect 19536 2332 19708 2360
rect 19702 2320 19708 2332
rect 19760 2320 19766 2372
rect 20254 2360 20260 2372
rect 19812 2332 20260 2360
rect 19812 2301 19840 2332
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 20548 2360 20576 2468
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20732 2428 20760 2527
rect 20671 2400 20760 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20824 2360 20852 2536
rect 23198 2524 23204 2576
rect 23256 2524 23262 2576
rect 25866 2524 25872 2576
rect 25924 2524 25930 2576
rect 26694 2564 26700 2576
rect 26436 2536 26700 2564
rect 23750 2496 23756 2508
rect 22940 2468 23756 2496
rect 20898 2388 20904 2440
rect 20956 2388 20962 2440
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 20548 2332 20852 2360
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 17276 2264 17417 2292
rect 17276 2252 17282 2264
rect 17405 2261 17417 2264
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 19886 2252 19892 2304
rect 19944 2252 19950 2304
rect 20165 2295 20223 2301
rect 20165 2261 20177 2295
rect 20211 2292 20223 2295
rect 21008 2292 21036 2391
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21729 2431 21787 2437
rect 21729 2428 21741 2431
rect 21324 2400 21741 2428
rect 21324 2388 21330 2400
rect 21729 2397 21741 2400
rect 21775 2397 21787 2431
rect 21729 2391 21787 2397
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 21876 2400 22109 2428
rect 21876 2388 21882 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22204 2360 22232 2391
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22940 2437 22968 2468
rect 23750 2456 23756 2468
rect 23808 2456 23814 2508
rect 25148 2468 25820 2496
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22336 2400 22661 2428
rect 22336 2388 22342 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2428 23075 2431
rect 23477 2431 23535 2437
rect 23063 2400 23428 2428
rect 23063 2397 23075 2400
rect 23017 2391 23075 2397
rect 23400 2360 23428 2400
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 24578 2428 24584 2440
rect 23523 2400 24584 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 25148 2437 25176 2468
rect 25041 2431 25099 2437
rect 25041 2397 25053 2431
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 24026 2360 24032 2372
rect 22204 2332 23336 2360
rect 23400 2332 24032 2360
rect 20211 2264 21036 2292
rect 21177 2295 21235 2301
rect 20211 2261 20223 2264
rect 20165 2255 20223 2261
rect 21177 2261 21189 2295
rect 21223 2292 21235 2295
rect 21450 2292 21456 2304
rect 21223 2264 21456 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21450 2252 21456 2264
rect 21508 2252 21514 2304
rect 21542 2252 21548 2304
rect 21600 2252 21606 2304
rect 21910 2252 21916 2304
rect 21968 2252 21974 2304
rect 22465 2295 22523 2301
rect 22465 2261 22477 2295
rect 22511 2292 22523 2295
rect 22922 2292 22928 2304
rect 22511 2264 22928 2292
rect 22511 2261 22523 2264
rect 22465 2255 22523 2261
rect 22922 2252 22928 2264
rect 22980 2252 22986 2304
rect 23308 2301 23336 2332
rect 24026 2320 24032 2332
rect 24084 2320 24090 2372
rect 25056 2360 25084 2391
rect 25590 2388 25596 2440
rect 25648 2388 25654 2440
rect 25056 2332 25728 2360
rect 23293 2295 23351 2301
rect 23293 2261 23305 2295
rect 23339 2261 23351 2295
rect 23293 2255 23351 2261
rect 24854 2252 24860 2304
rect 24912 2252 24918 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 25188 2264 25329 2292
rect 25188 2252 25194 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 25409 2295 25467 2301
rect 25409 2261 25421 2295
rect 25455 2292 25467 2295
rect 25590 2292 25596 2304
rect 25455 2264 25596 2292
rect 25455 2261 25467 2264
rect 25409 2255 25467 2261
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 25700 2301 25728 2332
rect 25685 2295 25743 2301
rect 25685 2261 25697 2295
rect 25731 2261 25743 2295
rect 25792 2292 25820 2468
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 25884 2360 25912 2391
rect 26142 2388 26148 2440
rect 26200 2388 26206 2440
rect 26436 2437 26464 2536
rect 26694 2524 26700 2536
rect 26752 2524 26758 2576
rect 26878 2524 26884 2576
rect 26936 2564 26942 2576
rect 36446 2564 36452 2576
rect 26936 2536 36452 2564
rect 26936 2524 26942 2536
rect 36446 2524 36452 2536
rect 36504 2524 36510 2576
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 26568 2468 29132 2496
rect 26568 2456 26574 2468
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2397 26479 2431
rect 26421 2391 26479 2397
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 26697 2431 26755 2437
rect 26697 2428 26709 2431
rect 26660 2400 26709 2428
rect 26660 2388 26666 2400
rect 26697 2397 26709 2400
rect 26743 2397 26755 2431
rect 26697 2391 26755 2397
rect 26970 2388 26976 2440
rect 27028 2388 27034 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27249 2431 27307 2437
rect 27249 2428 27261 2431
rect 27120 2400 27261 2428
rect 27120 2388 27126 2400
rect 27249 2397 27261 2400
rect 27295 2397 27307 2431
rect 27249 2391 27307 2397
rect 27522 2388 27528 2440
rect 27580 2388 27586 2440
rect 27614 2388 27620 2440
rect 27672 2388 27678 2440
rect 28534 2388 28540 2440
rect 28592 2388 28598 2440
rect 28626 2388 28632 2440
rect 28684 2428 28690 2440
rect 29104 2437 29132 2468
rect 30116 2468 31754 2496
rect 28813 2431 28871 2437
rect 28813 2428 28825 2431
rect 28684 2400 28825 2428
rect 28684 2388 28690 2400
rect 28813 2397 28825 2400
rect 28859 2397 28871 2431
rect 28813 2391 28871 2397
rect 29089 2431 29147 2437
rect 29089 2397 29101 2431
rect 29135 2397 29147 2431
rect 29089 2391 29147 2397
rect 29362 2388 29368 2440
rect 29420 2388 29426 2440
rect 30116 2437 30144 2468
rect 29733 2431 29791 2437
rect 29733 2397 29745 2431
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30101 2431 30159 2437
rect 30101 2397 30113 2431
rect 30147 2397 30159 2431
rect 30101 2391 30159 2397
rect 30377 2431 30435 2437
rect 30377 2397 30389 2431
rect 30423 2428 30435 2431
rect 31018 2428 31024 2440
rect 30423 2400 31024 2428
rect 30423 2397 30435 2400
rect 30377 2391 30435 2397
rect 27154 2360 27160 2372
rect 25884 2332 27160 2360
rect 27154 2320 27160 2332
rect 27212 2320 27218 2372
rect 28077 2363 28135 2369
rect 28077 2329 28089 2363
rect 28123 2360 28135 2363
rect 29748 2360 29776 2391
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 31294 2388 31300 2440
rect 31352 2388 31358 2440
rect 31386 2388 31392 2440
rect 31444 2388 31450 2440
rect 31726 2428 31754 2468
rect 33336 2468 34836 2496
rect 33336 2440 33364 2468
rect 33134 2428 33140 2440
rect 31726 2400 33140 2428
rect 33134 2388 33140 2400
rect 33192 2388 33198 2440
rect 33318 2388 33324 2440
rect 33376 2388 33382 2440
rect 33413 2431 33471 2437
rect 33413 2397 33425 2431
rect 33459 2428 33471 2431
rect 34698 2428 34704 2440
rect 33459 2400 34704 2428
rect 33459 2397 33471 2400
rect 33413 2391 33471 2397
rect 34698 2388 34704 2400
rect 34756 2388 34762 2440
rect 34808 2437 34836 2468
rect 34793 2431 34851 2437
rect 34793 2397 34805 2431
rect 34839 2397 34851 2431
rect 34793 2391 34851 2397
rect 35986 2388 35992 2440
rect 36044 2388 36050 2440
rect 37734 2388 37740 2440
rect 37792 2388 37798 2440
rect 39390 2388 39396 2440
rect 39448 2388 39454 2440
rect 40678 2388 40684 2440
rect 40736 2388 40742 2440
rect 42610 2388 42616 2440
rect 42668 2388 42674 2440
rect 35434 2360 35440 2372
rect 28123 2332 29592 2360
rect 29748 2332 35440 2360
rect 28123 2329 28135 2332
rect 28077 2323 28135 2329
rect 26237 2295 26295 2301
rect 26237 2292 26249 2295
rect 25792 2264 26249 2292
rect 25685 2255 25743 2261
rect 26237 2261 26249 2264
rect 26283 2261 26295 2295
rect 26237 2255 26295 2261
rect 26510 2252 26516 2304
rect 26568 2252 26574 2304
rect 26786 2252 26792 2304
rect 26844 2252 26850 2304
rect 27065 2295 27123 2301
rect 27065 2261 27077 2295
rect 27111 2292 27123 2295
rect 27890 2292 27896 2304
rect 27111 2264 27896 2292
rect 27111 2261 27123 2264
rect 27065 2255 27123 2261
rect 27890 2252 27896 2264
rect 27948 2252 27954 2304
rect 28350 2252 28356 2304
rect 28408 2252 28414 2304
rect 28629 2295 28687 2301
rect 28629 2261 28641 2295
rect 28675 2292 28687 2295
rect 28810 2292 28816 2304
rect 28675 2264 28816 2292
rect 28675 2261 28687 2264
rect 28629 2255 28687 2261
rect 28810 2252 28816 2264
rect 28868 2252 28874 2304
rect 28902 2252 28908 2304
rect 28960 2252 28966 2304
rect 29178 2252 29184 2304
rect 29236 2252 29242 2304
rect 29564 2301 29592 2332
rect 35434 2320 35440 2332
rect 35492 2320 35498 2372
rect 29549 2295 29607 2301
rect 29549 2261 29561 2295
rect 29595 2261 29607 2295
rect 29549 2255 29607 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 30561 2295 30619 2301
rect 30561 2292 30573 2295
rect 29696 2264 30573 2292
rect 29696 2252 29702 2264
rect 30561 2261 30573 2264
rect 30607 2261 30619 2295
rect 30561 2255 30619 2261
rect 30650 2252 30656 2304
rect 30708 2292 30714 2304
rect 31573 2295 31631 2301
rect 31573 2292 31585 2295
rect 30708 2264 31585 2292
rect 30708 2252 30714 2264
rect 31573 2261 31585 2264
rect 31619 2261 31631 2295
rect 31573 2255 31631 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 33560 2264 34897 2292
rect 33560 2252 33566 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 1104 2202 43675 2224
rect 1104 2150 11552 2202
rect 11604 2150 11616 2202
rect 11668 2150 11680 2202
rect 11732 2150 11744 2202
rect 11796 2150 11808 2202
rect 11860 2150 22155 2202
rect 22207 2150 22219 2202
rect 22271 2150 22283 2202
rect 22335 2150 22347 2202
rect 22399 2150 22411 2202
rect 22463 2150 32758 2202
rect 32810 2150 32822 2202
rect 32874 2150 32886 2202
rect 32938 2150 32950 2202
rect 33002 2150 33014 2202
rect 33066 2150 43361 2202
rect 43413 2150 43425 2202
rect 43477 2150 43489 2202
rect 43541 2150 43553 2202
rect 43605 2150 43617 2202
rect 43669 2150 43675 2202
rect 1104 2128 43675 2150
rect 9309 2091 9367 2097
rect 9309 2057 9321 2091
rect 9355 2088 9367 2091
rect 10962 2088 10968 2100
rect 9355 2060 10968 2088
rect 9355 2057 9367 2060
rect 9309 2051 9367 2057
rect 10962 2048 10968 2060
rect 11020 2048 11026 2100
rect 14274 2048 14280 2100
rect 14332 2048 14338 2100
rect 14829 2091 14887 2097
rect 14829 2057 14841 2091
rect 14875 2088 14887 2091
rect 15286 2088 15292 2100
rect 14875 2060 15292 2088
rect 14875 2057 14887 2060
rect 14829 2051 14887 2057
rect 15286 2048 15292 2060
rect 15344 2048 15350 2100
rect 15470 2048 15476 2100
rect 15528 2088 15534 2100
rect 15528 2060 15608 2088
rect 15528 2048 15534 2060
rect 15102 2020 15108 2032
rect 14568 1992 15108 2020
rect 9122 1912 9128 1964
rect 9180 1912 9186 1964
rect 14090 1912 14096 1964
rect 14148 1912 14154 1964
rect 14568 1961 14596 1992
rect 15102 1980 15108 1992
rect 15160 1980 15166 2032
rect 15580 2020 15608 2060
rect 15654 2048 15660 2100
rect 15712 2048 15718 2100
rect 15933 2091 15991 2097
rect 15933 2057 15945 2091
rect 15979 2088 15991 2091
rect 16206 2088 16212 2100
rect 15979 2060 16212 2088
rect 15979 2057 15991 2060
rect 15933 2051 15991 2057
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 16850 2048 16856 2100
rect 16908 2048 16914 2100
rect 17034 2048 17040 2100
rect 17092 2048 17098 2100
rect 17126 2048 17132 2100
rect 17184 2088 17190 2100
rect 17313 2091 17371 2097
rect 17313 2088 17325 2091
rect 17184 2060 17325 2088
rect 17184 2048 17190 2060
rect 17313 2057 17325 2060
rect 17359 2057 17371 2091
rect 17313 2051 17371 2057
rect 17589 2091 17647 2097
rect 17589 2057 17601 2091
rect 17635 2088 17647 2091
rect 18414 2088 18420 2100
rect 17635 2060 18420 2088
rect 17635 2057 17647 2060
rect 17589 2051 17647 2057
rect 18414 2048 18420 2060
rect 18472 2048 18478 2100
rect 19981 2091 20039 2097
rect 19981 2057 19993 2091
rect 20027 2088 20039 2091
rect 20990 2088 20996 2100
rect 20027 2060 20996 2088
rect 20027 2057 20039 2060
rect 19981 2051 20039 2057
rect 20990 2048 20996 2060
rect 21048 2048 21054 2100
rect 23201 2091 23259 2097
rect 23201 2057 23213 2091
rect 23247 2057 23259 2091
rect 23201 2051 23259 2057
rect 16868 2020 16896 2048
rect 15580 1992 16896 2020
rect 14553 1955 14611 1961
rect 14553 1921 14565 1955
rect 14599 1921 14611 1955
rect 14553 1915 14611 1921
rect 14642 1912 14648 1964
rect 14700 1912 14706 1964
rect 14918 1912 14924 1964
rect 14976 1912 14982 1964
rect 15197 1955 15255 1961
rect 15197 1921 15209 1955
rect 15243 1921 15255 1955
rect 15197 1915 15255 1921
rect 15212 1884 15240 1915
rect 15286 1912 15292 1964
rect 15344 1952 15350 1964
rect 15473 1955 15531 1961
rect 15473 1952 15485 1955
rect 15344 1924 15485 1952
rect 15344 1912 15350 1924
rect 15473 1921 15485 1924
rect 15519 1921 15531 1955
rect 15473 1915 15531 1921
rect 15749 1955 15807 1961
rect 15749 1921 15761 1955
rect 15795 1921 15807 1955
rect 15749 1915 15807 1921
rect 15764 1884 15792 1915
rect 15838 1912 15844 1964
rect 15896 1952 15902 1964
rect 16025 1955 16083 1961
rect 16025 1952 16037 1955
rect 15896 1924 16037 1952
rect 15896 1912 15902 1924
rect 16025 1921 16037 1924
rect 16071 1921 16083 1955
rect 16025 1915 16083 1921
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 16390 1912 16396 1964
rect 16448 1952 16454 1964
rect 16853 1955 16911 1961
rect 16853 1952 16865 1955
rect 16448 1924 16865 1952
rect 16448 1912 16454 1924
rect 16853 1921 16865 1924
rect 16899 1921 16911 1955
rect 17052 1952 17080 2048
rect 17218 1980 17224 2032
rect 17276 2020 17282 2032
rect 20533 2023 20591 2029
rect 20533 2020 20545 2023
rect 17276 1992 17356 2020
rect 17276 1980 17282 1992
rect 17328 1976 17356 1992
rect 17604 1992 18092 2020
rect 17328 1961 17448 1976
rect 17129 1955 17187 1961
rect 17129 1952 17141 1955
rect 17052 1924 17141 1952
rect 16853 1915 16911 1921
rect 17129 1921 17141 1924
rect 17175 1921 17187 1955
rect 17328 1955 17463 1961
rect 17328 1948 17417 1955
rect 17129 1915 17187 1921
rect 17405 1921 17417 1948
rect 17451 1921 17463 1955
rect 17405 1915 17463 1921
rect 14384 1856 15240 1884
rect 15304 1856 15792 1884
rect 14384 1825 14412 1856
rect 14369 1819 14427 1825
rect 14369 1785 14381 1819
rect 14415 1785 14427 1819
rect 14369 1779 14427 1785
rect 15105 1819 15163 1825
rect 15105 1785 15117 1819
rect 15151 1816 15163 1819
rect 15194 1816 15200 1828
rect 15151 1788 15200 1816
rect 15151 1785 15163 1788
rect 15105 1779 15163 1785
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
rect 14458 1708 14464 1760
rect 14516 1748 14522 1760
rect 15304 1748 15332 1856
rect 16574 1844 16580 1896
rect 16632 1884 16638 1896
rect 16632 1856 17448 1884
rect 16632 1844 16638 1856
rect 15378 1776 15384 1828
rect 15436 1776 15442 1828
rect 16209 1819 16267 1825
rect 16209 1785 16221 1819
rect 16255 1816 16267 1819
rect 16666 1816 16672 1828
rect 16255 1788 16672 1816
rect 16255 1785 16267 1788
rect 16209 1779 16267 1785
rect 16666 1776 16672 1788
rect 16724 1776 16730 1828
rect 14516 1720 15332 1748
rect 14516 1708 14522 1720
rect 16482 1708 16488 1760
rect 16540 1708 16546 1760
rect 16850 1708 16856 1760
rect 16908 1748 16914 1760
rect 17037 1751 17095 1757
rect 17037 1748 17049 1751
rect 16908 1720 17049 1748
rect 16908 1708 16914 1720
rect 17037 1717 17049 1720
rect 17083 1717 17095 1751
rect 17420 1748 17448 1856
rect 17604 1748 17632 1992
rect 18064 1964 18092 1992
rect 18616 1992 19840 2020
rect 17865 1955 17923 1961
rect 17865 1936 17877 1955
rect 17788 1921 17877 1936
rect 17911 1921 17923 1955
rect 17788 1915 17923 1921
rect 17788 1908 17908 1915
rect 18046 1912 18052 1964
rect 18104 1912 18110 1964
rect 18138 1936 18144 1988
rect 18196 1936 18202 1988
rect 18233 1955 18291 1961
rect 18233 1921 18245 1955
rect 18279 1921 18291 1955
rect 18233 1915 18291 1921
rect 17678 1844 17684 1896
rect 17736 1884 17742 1896
rect 17788 1884 17816 1908
rect 18248 1884 18276 1915
rect 17736 1856 17816 1884
rect 17926 1856 18276 1884
rect 17736 1844 17742 1856
rect 17926 1816 17954 1856
rect 17880 1788 17954 1816
rect 18417 1819 18475 1825
rect 17880 1760 17908 1788
rect 18417 1785 18429 1819
rect 18463 1816 18475 1819
rect 18616 1816 18644 1992
rect 18690 1912 18696 1964
rect 18748 1912 18754 1964
rect 18782 1912 18788 1964
rect 18840 1952 18846 1964
rect 18969 1955 19027 1961
rect 18969 1952 18981 1955
rect 18840 1924 18981 1952
rect 18840 1912 18846 1924
rect 18969 1921 18981 1924
rect 19015 1921 19027 1955
rect 18969 1915 19027 1921
rect 19058 1912 19064 1964
rect 19116 1952 19122 1964
rect 19245 1955 19303 1961
rect 19245 1952 19257 1955
rect 19116 1924 19257 1952
rect 19116 1912 19122 1924
rect 19245 1921 19257 1924
rect 19291 1921 19303 1955
rect 19245 1915 19303 1921
rect 19426 1912 19432 1964
rect 19484 1952 19490 1964
rect 19521 1955 19579 1961
rect 19521 1952 19533 1955
rect 19484 1924 19533 1952
rect 19484 1912 19490 1924
rect 19521 1921 19533 1924
rect 19567 1921 19579 1955
rect 19521 1915 19579 1921
rect 19705 1955 19763 1961
rect 19705 1921 19717 1955
rect 19751 1921 19763 1955
rect 19705 1915 19763 1921
rect 19720 1884 19748 1915
rect 18708 1856 19748 1884
rect 18708 1828 18736 1856
rect 18463 1788 18644 1816
rect 18463 1785 18475 1788
rect 18417 1779 18475 1785
rect 18690 1776 18696 1828
rect 18748 1776 18754 1828
rect 18785 1819 18843 1825
rect 18785 1785 18797 1819
rect 18831 1816 18843 1819
rect 19518 1816 19524 1828
rect 18831 1788 19524 1816
rect 18831 1785 18843 1788
rect 18785 1779 18843 1785
rect 19518 1776 19524 1788
rect 19576 1776 19582 1828
rect 17420 1720 17632 1748
rect 17037 1711 17095 1717
rect 17678 1708 17684 1760
rect 17736 1708 17742 1760
rect 17862 1708 17868 1760
rect 17920 1708 17926 1760
rect 17954 1708 17960 1760
rect 18012 1708 18018 1760
rect 18509 1751 18567 1757
rect 18509 1717 18521 1751
rect 18555 1748 18567 1751
rect 18966 1748 18972 1760
rect 18555 1720 18972 1748
rect 18555 1717 18567 1720
rect 18509 1711 18567 1717
rect 18966 1708 18972 1720
rect 19024 1708 19030 1760
rect 19061 1751 19119 1757
rect 19061 1717 19073 1751
rect 19107 1748 19119 1751
rect 19242 1748 19248 1760
rect 19107 1720 19248 1748
rect 19107 1717 19119 1720
rect 19061 1711 19119 1717
rect 19242 1708 19248 1720
rect 19300 1708 19306 1760
rect 19334 1708 19340 1760
rect 19392 1708 19398 1760
rect 19812 1748 19840 1992
rect 19904 1992 20545 2020
rect 19904 1964 19932 1992
rect 20533 1989 20545 1992
rect 20579 1989 20591 2023
rect 20533 1983 20591 1989
rect 20714 1980 20720 2032
rect 20772 2020 20778 2032
rect 21269 2023 21327 2029
rect 21269 2020 21281 2023
rect 20772 1992 21281 2020
rect 20772 1980 20778 1992
rect 21269 1989 21281 1992
rect 21315 1989 21327 2023
rect 21269 1983 21327 1989
rect 21726 1980 21732 2032
rect 21784 2020 21790 2032
rect 22189 2023 22247 2029
rect 22189 2020 22201 2023
rect 21784 1992 22201 2020
rect 21784 1980 21790 1992
rect 22189 1989 22201 1992
rect 22235 1989 22247 2023
rect 23216 2020 23244 2051
rect 23750 2048 23756 2100
rect 23808 2048 23814 2100
rect 24026 2048 24032 2100
rect 24084 2048 24090 2100
rect 24136 2060 24440 2088
rect 24136 2020 24164 2060
rect 23216 1992 24164 2020
rect 22189 1983 22247 1989
rect 19886 1912 19892 1964
rect 19944 1912 19950 1964
rect 20349 1955 20407 1961
rect 20349 1921 20361 1955
rect 20395 1952 20407 1955
rect 20622 1952 20628 1964
rect 20395 1924 20628 1952
rect 20395 1921 20407 1924
rect 20349 1915 20407 1921
rect 20622 1912 20628 1924
rect 20680 1912 20686 1964
rect 20806 1912 20812 1964
rect 20864 1952 20870 1964
rect 22005 1955 22063 1961
rect 22005 1952 22017 1955
rect 20864 1924 22017 1952
rect 20864 1912 20870 1924
rect 22005 1921 22017 1924
rect 22051 1921 22063 1955
rect 22005 1915 22063 1921
rect 22649 1955 22707 1961
rect 22649 1921 22661 1955
rect 22695 1921 22707 1955
rect 22649 1915 22707 1921
rect 22664 1884 22692 1915
rect 23382 1912 23388 1964
rect 23440 1912 23446 1964
rect 23658 1912 23664 1964
rect 23716 1912 23722 1964
rect 23842 1912 23848 1964
rect 23900 1952 23906 1964
rect 23937 1955 23995 1961
rect 23937 1952 23949 1955
rect 23900 1924 23949 1952
rect 23900 1912 23906 1924
rect 23937 1921 23949 1924
rect 23983 1921 23995 1955
rect 23937 1915 23995 1921
rect 24118 1912 24124 1964
rect 24176 1952 24182 1964
rect 24412 1961 24440 2060
rect 25866 2048 25872 2100
rect 25924 2048 25930 2100
rect 26786 2048 26792 2100
rect 26844 2048 26850 2100
rect 26970 2048 26976 2100
rect 27028 2088 27034 2100
rect 27985 2091 28043 2097
rect 27985 2088 27997 2091
rect 27028 2060 27997 2088
rect 27028 2048 27034 2060
rect 27985 2057 27997 2060
rect 28031 2057 28043 2091
rect 27985 2051 28043 2057
rect 28350 2048 28356 2100
rect 28408 2048 28414 2100
rect 28902 2048 28908 2100
rect 28960 2048 28966 2100
rect 29178 2048 29184 2100
rect 29236 2088 29242 2100
rect 29236 2060 30696 2088
rect 29236 2048 29242 2060
rect 25777 2023 25835 2029
rect 25777 1989 25789 2023
rect 25823 2020 25835 2023
rect 25884 2020 25912 2048
rect 25823 1992 25912 2020
rect 25823 1989 25835 1992
rect 25777 1983 25835 1989
rect 26234 1980 26240 2032
rect 26292 2020 26298 2032
rect 26329 2023 26387 2029
rect 26329 2020 26341 2023
rect 26292 1992 26341 2020
rect 26292 1980 26298 1992
rect 26329 1989 26341 1992
rect 26375 1989 26387 2023
rect 26804 2020 26832 2048
rect 27893 2023 27951 2029
rect 27893 2020 27905 2023
rect 26804 1992 27905 2020
rect 26329 1983 26387 1989
rect 27893 1989 27905 1992
rect 27939 1989 27951 2023
rect 28368 2020 28396 2048
rect 28445 2023 28503 2029
rect 28445 2020 28457 2023
rect 28368 1992 28457 2020
rect 27893 1983 27951 1989
rect 28445 1989 28457 1992
rect 28491 1989 28503 2023
rect 28920 2020 28948 2048
rect 28997 2023 29055 2029
rect 28997 2020 29009 2023
rect 28920 1992 29009 2020
rect 28445 1983 28503 1989
rect 28997 1989 29009 1992
rect 29043 1989 29055 2023
rect 29549 2023 29607 2029
rect 29549 2020 29561 2023
rect 28997 1983 29055 1989
rect 29472 1992 29561 2020
rect 29472 1964 29500 1992
rect 29549 1989 29561 1992
rect 29595 1989 29607 2023
rect 29549 1983 29607 1989
rect 29730 1980 29736 2032
rect 29788 2020 29794 2032
rect 30101 2023 30159 2029
rect 30101 2020 30113 2023
rect 29788 1992 30113 2020
rect 29788 1980 29794 1992
rect 30101 1989 30113 1992
rect 30147 1989 30159 2023
rect 30101 1983 30159 1989
rect 30190 1980 30196 2032
rect 30248 2020 30254 2032
rect 30668 2029 30696 2060
rect 30742 2048 30748 2100
rect 30800 2048 30806 2100
rect 31294 2048 31300 2100
rect 31352 2088 31358 2100
rect 31757 2091 31815 2097
rect 31757 2088 31769 2091
rect 31352 2060 31769 2088
rect 31352 2048 31358 2060
rect 31757 2057 31769 2060
rect 31803 2057 31815 2091
rect 31757 2051 31815 2057
rect 32582 2048 32588 2100
rect 32640 2088 32646 2100
rect 34517 2091 34575 2097
rect 34517 2088 34529 2091
rect 32640 2060 34529 2088
rect 32640 2048 32646 2060
rect 34517 2057 34529 2060
rect 34563 2057 34575 2091
rect 34517 2051 34575 2057
rect 30653 2023 30711 2029
rect 30248 1992 30604 2020
rect 30248 1980 30254 1992
rect 24213 1955 24271 1961
rect 24213 1952 24225 1955
rect 24176 1924 24225 1952
rect 24176 1912 24182 1924
rect 24213 1921 24225 1924
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 24397 1955 24455 1961
rect 24397 1921 24409 1955
rect 24443 1921 24455 1955
rect 24397 1915 24455 1921
rect 24946 1912 24952 1964
rect 25004 1912 25010 1964
rect 25222 1912 25228 1964
rect 25280 1912 25286 1964
rect 25498 1912 25504 1964
rect 25556 1912 25562 1964
rect 25866 1912 25872 1964
rect 25924 1952 25930 1964
rect 27157 1955 27215 1961
rect 27157 1952 27169 1955
rect 25924 1924 27169 1952
rect 25924 1912 25930 1924
rect 27157 1921 27169 1924
rect 27203 1952 27215 1955
rect 27709 1955 27767 1961
rect 27709 1952 27721 1955
rect 27203 1924 27721 1952
rect 27203 1921 27215 1924
rect 27157 1915 27215 1921
rect 27709 1921 27721 1924
rect 27755 1921 27767 1955
rect 27709 1915 27767 1921
rect 28166 1912 28172 1964
rect 28224 1952 28230 1964
rect 28224 1924 29408 1952
rect 28224 1912 28230 1924
rect 29270 1884 29276 1896
rect 20180 1856 22692 1884
rect 23032 1856 29276 1884
rect 20180 1825 20208 1856
rect 20165 1819 20223 1825
rect 20165 1785 20177 1819
rect 20211 1785 20223 1819
rect 20165 1779 20223 1785
rect 20438 1776 20444 1828
rect 20496 1816 20502 1828
rect 20717 1819 20775 1825
rect 20717 1816 20729 1819
rect 20496 1788 20729 1816
rect 20496 1776 20502 1788
rect 20717 1785 20729 1788
rect 20763 1785 20775 1819
rect 23032 1816 23060 1856
rect 29270 1844 29276 1856
rect 29328 1844 29334 1896
rect 20717 1779 20775 1785
rect 21284 1788 23060 1816
rect 23477 1819 23535 1825
rect 21284 1748 21312 1788
rect 23477 1785 23489 1819
rect 23523 1816 23535 1819
rect 24854 1816 24860 1828
rect 23523 1788 24860 1816
rect 23523 1785 23535 1788
rect 23477 1779 23535 1785
rect 24854 1776 24860 1788
rect 24912 1776 24918 1828
rect 25317 1819 25375 1825
rect 25317 1785 25329 1819
rect 25363 1816 25375 1819
rect 26234 1816 26240 1828
rect 25363 1788 26240 1816
rect 25363 1785 25375 1788
rect 25317 1779 25375 1785
rect 26234 1776 26240 1788
rect 26292 1776 26298 1828
rect 27798 1776 27804 1828
rect 27856 1816 27862 1828
rect 29380 1816 29408 1924
rect 29454 1912 29460 1964
rect 29512 1912 29518 1964
rect 30576 1952 30604 1992
rect 30653 1989 30665 2023
rect 30699 1989 30711 2023
rect 32217 2023 32275 2029
rect 32217 2020 32229 2023
rect 30653 1983 30711 1989
rect 30760 1992 32229 2020
rect 30760 1952 30788 1992
rect 32217 1989 32229 1992
rect 32263 1989 32275 2023
rect 32217 1983 32275 1989
rect 32306 1980 32312 2032
rect 32364 2020 32370 2032
rect 32364 1992 33272 2020
rect 32364 1980 32370 1992
rect 30576 1924 30788 1952
rect 31202 1912 31208 1964
rect 31260 1912 31266 1964
rect 31938 1912 31944 1964
rect 31996 1912 32002 1964
rect 32769 1955 32827 1961
rect 32769 1921 32781 1955
rect 32815 1921 32827 1955
rect 32769 1915 32827 1921
rect 30377 1887 30435 1893
rect 30377 1884 30389 1887
rect 29546 1856 30389 1884
rect 29546 1816 29574 1856
rect 30377 1853 30389 1856
rect 30423 1853 30435 1887
rect 30377 1847 30435 1853
rect 31478 1844 31484 1896
rect 31536 1884 31542 1896
rect 32784 1884 32812 1915
rect 31536 1856 32812 1884
rect 33244 1884 33272 1992
rect 33318 1912 33324 1964
rect 33376 1912 33382 1964
rect 33870 1912 33876 1964
rect 33928 1912 33934 1964
rect 34532 1952 34560 2051
rect 34698 2048 34704 2100
rect 34756 2048 34762 2100
rect 35434 2048 35440 2100
rect 35492 2048 35498 2100
rect 35986 2048 35992 2100
rect 36044 2088 36050 2100
rect 36449 2091 36507 2097
rect 36449 2088 36461 2091
rect 36044 2060 36461 2088
rect 36044 2048 36050 2060
rect 36449 2057 36461 2060
rect 36495 2057 36507 2091
rect 36449 2051 36507 2057
rect 37461 2091 37519 2097
rect 37461 2057 37473 2091
rect 37507 2057 37519 2091
rect 37461 2051 37519 2057
rect 34716 2020 34744 2048
rect 37476 2020 37504 2051
rect 37734 2048 37740 2100
rect 37792 2088 37798 2100
rect 37921 2091 37979 2097
rect 37921 2088 37933 2091
rect 37792 2060 37933 2088
rect 37792 2048 37798 2060
rect 37921 2057 37933 2060
rect 37967 2057 37979 2091
rect 37921 2051 37979 2057
rect 38565 2091 38623 2097
rect 38565 2057 38577 2091
rect 38611 2088 38623 2091
rect 39390 2088 39396 2100
rect 38611 2060 39396 2088
rect 38611 2057 38623 2060
rect 38565 2051 38623 2057
rect 39390 2048 39396 2060
rect 39448 2048 39454 2100
rect 39761 2091 39819 2097
rect 39761 2057 39773 2091
rect 39807 2088 39819 2091
rect 40678 2088 40684 2100
rect 39807 2060 40684 2088
rect 39807 2057 39819 2060
rect 39761 2051 39819 2057
rect 40678 2048 40684 2060
rect 40736 2048 40742 2100
rect 42610 2048 42616 2100
rect 42668 2048 42674 2100
rect 40954 2020 40960 2032
rect 34716 1992 37504 2020
rect 38120 1992 40960 2020
rect 34977 1955 35035 1961
rect 34977 1952 34989 1955
rect 34532 1924 34989 1952
rect 34977 1921 34989 1924
rect 35023 1921 35035 1955
rect 34977 1915 35035 1921
rect 35621 1955 35679 1961
rect 35621 1921 35633 1955
rect 35667 1921 35679 1955
rect 35621 1915 35679 1921
rect 33244 1856 33548 1884
rect 31536 1844 31542 1856
rect 27856 1788 28580 1816
rect 29380 1788 29574 1816
rect 27856 1776 27862 1788
rect 19812 1720 21312 1748
rect 21358 1708 21364 1760
rect 21416 1708 21422 1760
rect 21818 1708 21824 1760
rect 21876 1708 21882 1760
rect 22002 1708 22008 1760
rect 22060 1748 22066 1760
rect 22281 1751 22339 1757
rect 22281 1748 22293 1751
rect 22060 1720 22293 1748
rect 22060 1708 22066 1720
rect 22281 1717 22293 1720
rect 22327 1717 22339 1751
rect 22281 1711 22339 1717
rect 22830 1708 22836 1760
rect 22888 1708 22894 1760
rect 24210 1708 24216 1760
rect 24268 1748 24274 1760
rect 24581 1751 24639 1757
rect 24581 1748 24593 1751
rect 24268 1720 24593 1748
rect 24268 1708 24274 1720
rect 24581 1717 24593 1720
rect 24627 1717 24639 1751
rect 24581 1711 24639 1717
rect 24762 1708 24768 1760
rect 24820 1708 24826 1760
rect 25038 1708 25044 1760
rect 25096 1708 25102 1760
rect 25590 1708 25596 1760
rect 25648 1748 25654 1760
rect 25869 1751 25927 1757
rect 25869 1748 25881 1751
rect 25648 1720 25881 1748
rect 25648 1708 25654 1720
rect 25869 1717 25881 1720
rect 25915 1717 25927 1751
rect 25869 1711 25927 1717
rect 26142 1708 26148 1760
rect 26200 1748 26206 1760
rect 26421 1751 26479 1757
rect 26421 1748 26433 1751
rect 26200 1720 26433 1748
rect 26200 1708 26206 1720
rect 26421 1717 26433 1720
rect 26467 1717 26479 1751
rect 26421 1711 26479 1717
rect 27338 1708 27344 1760
rect 27396 1748 27402 1760
rect 28552 1757 28580 1788
rect 31662 1776 31668 1828
rect 31720 1816 31726 1828
rect 31720 1788 33456 1816
rect 31720 1776 31726 1788
rect 27525 1751 27583 1757
rect 27525 1748 27537 1751
rect 27396 1720 27537 1748
rect 27396 1708 27402 1720
rect 27525 1717 27537 1720
rect 27571 1717 27583 1751
rect 27525 1711 27583 1717
rect 28537 1751 28595 1757
rect 28537 1717 28549 1751
rect 28583 1717 28595 1751
rect 28537 1711 28595 1717
rect 28626 1708 28632 1760
rect 28684 1748 28690 1760
rect 29089 1751 29147 1757
rect 29089 1748 29101 1751
rect 28684 1720 29101 1748
rect 28684 1708 28690 1720
rect 29089 1717 29101 1720
rect 29135 1717 29147 1751
rect 29089 1711 29147 1717
rect 29638 1708 29644 1760
rect 29696 1708 29702 1760
rect 30466 1708 30472 1760
rect 30524 1748 30530 1760
rect 31297 1751 31355 1757
rect 31297 1748 31309 1751
rect 30524 1720 31309 1748
rect 30524 1708 30530 1720
rect 31297 1717 31309 1720
rect 31343 1717 31355 1751
rect 31297 1711 31355 1717
rect 31570 1708 31576 1760
rect 31628 1748 31634 1760
rect 32309 1751 32367 1757
rect 32309 1748 32321 1751
rect 31628 1720 32321 1748
rect 31628 1708 31634 1720
rect 32309 1717 32321 1720
rect 32355 1717 32367 1751
rect 32309 1711 32367 1717
rect 32490 1708 32496 1760
rect 32548 1748 32554 1760
rect 33428 1757 33456 1788
rect 32861 1751 32919 1757
rect 32861 1748 32873 1751
rect 32548 1720 32873 1748
rect 32548 1708 32554 1720
rect 32861 1717 32873 1720
rect 32907 1717 32919 1751
rect 32861 1711 32919 1717
rect 33413 1751 33471 1757
rect 33413 1717 33425 1751
rect 33459 1717 33471 1751
rect 33520 1748 33548 1856
rect 34238 1844 34244 1896
rect 34296 1884 34302 1896
rect 35636 1884 35664 1915
rect 36538 1912 36544 1964
rect 36596 1952 36602 1964
rect 36633 1955 36691 1961
rect 36633 1952 36645 1955
rect 36596 1924 36645 1952
rect 36596 1912 36602 1924
rect 36633 1921 36645 1924
rect 36679 1921 36691 1955
rect 36633 1915 36691 1921
rect 36725 1955 36783 1961
rect 36725 1921 36737 1955
rect 36771 1921 36783 1955
rect 36725 1915 36783 1921
rect 34296 1856 35664 1884
rect 34296 1844 34302 1856
rect 35802 1844 35808 1896
rect 35860 1884 35866 1896
rect 36740 1884 36768 1915
rect 37642 1912 37648 1964
rect 37700 1912 37706 1964
rect 38120 1961 38148 1992
rect 40954 1980 40960 1992
rect 41012 1980 41018 2032
rect 38105 1955 38163 1961
rect 38105 1921 38117 1955
rect 38151 1921 38163 1955
rect 38105 1915 38163 1921
rect 38749 1955 38807 1961
rect 38749 1921 38761 1955
rect 38795 1921 38807 1955
rect 38749 1915 38807 1921
rect 39945 1955 40003 1961
rect 39945 1921 39957 1955
rect 39991 1952 40003 1955
rect 40126 1952 40132 1964
rect 39991 1924 40132 1952
rect 39991 1921 40003 1924
rect 39945 1915 40003 1921
rect 35860 1856 36768 1884
rect 38764 1884 38792 1915
rect 40126 1912 40132 1924
rect 40184 1912 40190 1964
rect 40221 1955 40279 1961
rect 40221 1921 40233 1955
rect 40267 1952 40279 1955
rect 41782 1952 41788 1964
rect 40267 1924 41788 1952
rect 40267 1921 40279 1924
rect 40221 1915 40279 1921
rect 41782 1912 41788 1924
rect 41840 1912 41846 1964
rect 41230 1884 41236 1896
rect 38764 1856 41236 1884
rect 35860 1844 35866 1856
rect 41230 1844 41236 1856
rect 41288 1844 41294 1896
rect 33594 1776 33600 1828
rect 33652 1816 33658 1828
rect 33652 1788 35112 1816
rect 33652 1776 33658 1788
rect 35084 1757 35112 1788
rect 35158 1776 35164 1828
rect 35216 1816 35222 1828
rect 36909 1819 36967 1825
rect 36909 1816 36921 1819
rect 35216 1788 36921 1816
rect 35216 1776 35222 1788
rect 36909 1785 36921 1788
rect 36955 1785 36967 1819
rect 36909 1779 36967 1785
rect 40037 1819 40095 1825
rect 40037 1785 40049 1819
rect 40083 1816 40095 1819
rect 42628 1816 42656 2048
rect 40083 1788 42656 1816
rect 40083 1785 40095 1788
rect 40037 1779 40095 1785
rect 33965 1751 34023 1757
rect 33965 1748 33977 1751
rect 33520 1720 33977 1748
rect 33413 1711 33471 1717
rect 33965 1717 33977 1720
rect 34011 1717 34023 1751
rect 33965 1711 34023 1717
rect 35069 1751 35127 1757
rect 35069 1717 35081 1751
rect 35115 1717 35127 1751
rect 35069 1711 35127 1717
rect 1104 1658 43516 1680
rect 1104 1606 6251 1658
rect 6303 1606 6315 1658
rect 6367 1606 6379 1658
rect 6431 1606 6443 1658
rect 6495 1606 6507 1658
rect 6559 1606 16854 1658
rect 16906 1606 16918 1658
rect 16970 1606 16982 1658
rect 17034 1606 17046 1658
rect 17098 1606 17110 1658
rect 17162 1606 27457 1658
rect 27509 1606 27521 1658
rect 27573 1606 27585 1658
rect 27637 1606 27649 1658
rect 27701 1606 27713 1658
rect 27765 1606 38060 1658
rect 38112 1606 38124 1658
rect 38176 1606 38188 1658
rect 38240 1606 38252 1658
rect 38304 1606 38316 1658
rect 38368 1606 43516 1658
rect 1104 1584 43516 1606
rect 5905 1547 5963 1553
rect 5905 1513 5917 1547
rect 5951 1544 5963 1547
rect 7190 1544 7196 1556
rect 5951 1516 7196 1544
rect 5951 1513 5963 1516
rect 5905 1507 5963 1513
rect 7190 1504 7196 1516
rect 7248 1504 7254 1556
rect 9677 1547 9735 1553
rect 9677 1513 9689 1547
rect 9723 1513 9735 1547
rect 9677 1507 9735 1513
rect 5353 1479 5411 1485
rect 5353 1445 5365 1479
rect 5399 1476 5411 1479
rect 5810 1476 5816 1488
rect 5399 1448 5816 1476
rect 5399 1445 5411 1448
rect 5353 1439 5411 1445
rect 5810 1436 5816 1448
rect 5868 1436 5874 1488
rect 6825 1479 6883 1485
rect 6825 1445 6837 1479
rect 6871 1476 6883 1479
rect 8570 1476 8576 1488
rect 6871 1448 8576 1476
rect 6871 1445 6883 1448
rect 6825 1439 6883 1445
rect 8570 1436 8576 1448
rect 8628 1436 8634 1488
rect 9692 1476 9720 1507
rect 11054 1504 11060 1556
rect 11112 1504 11118 1556
rect 11330 1504 11336 1556
rect 11388 1504 11394 1556
rect 12802 1504 12808 1556
rect 12860 1504 12866 1556
rect 14093 1547 14151 1553
rect 14093 1513 14105 1547
rect 14139 1544 14151 1547
rect 14458 1544 14464 1556
rect 14139 1516 14464 1544
rect 14139 1513 14151 1516
rect 14093 1507 14151 1513
rect 14458 1504 14464 1516
rect 14516 1504 14522 1556
rect 15286 1544 15292 1556
rect 14568 1516 15292 1544
rect 13722 1476 13728 1488
rect 9692 1448 13728 1476
rect 13722 1436 13728 1448
rect 13780 1436 13786 1488
rect 5902 1408 5908 1420
rect 5552 1380 5908 1408
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1309 4675 1343
rect 4617 1303 4675 1309
rect 4893 1343 4951 1349
rect 4893 1309 4905 1343
rect 4939 1340 4951 1343
rect 5169 1343 5227 1349
rect 4939 1312 5120 1340
rect 4939 1309 4951 1312
rect 4893 1303 4951 1309
rect 4632 1272 4660 1303
rect 4982 1272 4988 1284
rect 4632 1244 4988 1272
rect 4982 1232 4988 1244
rect 5040 1232 5046 1284
rect 5092 1272 5120 1312
rect 5169 1309 5181 1343
rect 5215 1340 5227 1343
rect 5445 1343 5503 1349
rect 5215 1312 5396 1340
rect 5215 1309 5227 1312
rect 5169 1303 5227 1309
rect 5258 1272 5264 1284
rect 5092 1244 5264 1272
rect 5258 1232 5264 1244
rect 5316 1232 5322 1284
rect 5368 1272 5396 1312
rect 5445 1309 5457 1343
rect 5491 1340 5503 1343
rect 5552 1340 5580 1380
rect 5902 1368 5908 1380
rect 5960 1368 5966 1420
rect 9674 1408 9680 1420
rect 9416 1380 9680 1408
rect 5491 1312 5580 1340
rect 5721 1343 5779 1349
rect 5491 1309 5503 1312
rect 5445 1303 5503 1309
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5534 1272 5540 1284
rect 5368 1244 5540 1272
rect 5534 1232 5540 1244
rect 5592 1232 5598 1284
rect 5736 1272 5764 1303
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 6730 1300 6736 1352
rect 6788 1300 6794 1352
rect 6917 1343 6975 1349
rect 6917 1309 6929 1343
rect 6963 1309 6975 1343
rect 6917 1303 6975 1309
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1340 7251 1343
rect 7374 1340 7380 1352
rect 7239 1312 7380 1340
rect 7239 1309 7251 1312
rect 7193 1303 7251 1309
rect 6270 1272 6276 1284
rect 5736 1244 6276 1272
rect 6270 1232 6276 1244
rect 6328 1232 6334 1284
rect 6748 1272 6776 1300
rect 6472 1244 6776 1272
rect 6932 1272 6960 1303
rect 7374 1300 7380 1312
rect 7432 1300 7438 1352
rect 7469 1343 7527 1349
rect 7469 1309 7481 1343
rect 7515 1340 7527 1343
rect 7650 1340 7656 1352
rect 7515 1312 7656 1340
rect 7515 1309 7527 1312
rect 7469 1303 7527 1309
rect 7650 1300 7656 1312
rect 7708 1300 7714 1352
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1340 7803 1343
rect 7926 1340 7932 1352
rect 7791 1312 7932 1340
rect 7791 1309 7803 1312
rect 7745 1303 7803 1309
rect 7926 1300 7932 1312
rect 7984 1300 7990 1352
rect 8021 1343 8079 1349
rect 8021 1309 8033 1343
rect 8067 1309 8079 1343
rect 8021 1303 8079 1309
rect 8297 1343 8355 1349
rect 8297 1309 8309 1343
rect 8343 1340 8355 1343
rect 8478 1340 8484 1352
rect 8343 1312 8484 1340
rect 8343 1309 8355 1312
rect 8297 1303 8355 1309
rect 7282 1272 7288 1284
rect 6932 1244 7288 1272
rect 4798 1164 4804 1216
rect 4856 1164 4862 1216
rect 4890 1164 4896 1216
rect 4948 1204 4954 1216
rect 5077 1207 5135 1213
rect 5077 1204 5089 1207
rect 4948 1176 5089 1204
rect 4948 1164 4954 1176
rect 5077 1173 5089 1176
rect 5123 1173 5135 1207
rect 5077 1167 5135 1173
rect 5629 1207 5687 1213
rect 5629 1173 5641 1207
rect 5675 1204 5687 1207
rect 6086 1204 6092 1216
rect 5675 1176 6092 1204
rect 5675 1173 5687 1176
rect 5629 1167 5687 1173
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 6181 1207 6239 1213
rect 6181 1173 6193 1207
rect 6227 1204 6239 1207
rect 6472 1204 6500 1244
rect 7282 1232 7288 1244
rect 7340 1232 7346 1284
rect 7834 1272 7840 1284
rect 7392 1244 7840 1272
rect 6227 1176 6500 1204
rect 6227 1173 6239 1176
rect 6181 1167 6239 1173
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 7101 1207 7159 1213
rect 7101 1173 7113 1207
rect 7147 1204 7159 1207
rect 7190 1204 7196 1216
rect 7147 1176 7196 1204
rect 7147 1173 7159 1176
rect 7101 1167 7159 1173
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
rect 7392 1213 7420 1244
rect 7834 1232 7840 1244
rect 7892 1232 7898 1284
rect 8036 1272 8064 1303
rect 8478 1300 8484 1312
rect 8536 1300 8542 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8846 1340 8852 1352
rect 8619 1312 8852 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8846 1300 8852 1312
rect 8904 1300 8910 1352
rect 8941 1343 8999 1349
rect 8941 1309 8953 1343
rect 8987 1309 8999 1343
rect 8941 1303 8999 1309
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1340 9275 1343
rect 9416 1340 9444 1380
rect 9674 1368 9680 1380
rect 9732 1368 9738 1420
rect 12434 1408 12440 1420
rect 10244 1380 10456 1408
rect 9263 1312 9444 1340
rect 9493 1343 9551 1349
rect 9263 1309 9275 1312
rect 9217 1303 9275 1309
rect 9493 1309 9505 1343
rect 9539 1340 9551 1343
rect 9858 1340 9864 1352
rect 9539 1312 9864 1340
rect 9539 1309 9551 1312
rect 9493 1303 9551 1309
rect 8386 1272 8392 1284
rect 8036 1244 8392 1272
rect 8386 1232 8392 1244
rect 8444 1232 8450 1284
rect 8956 1272 8984 1303
rect 9858 1300 9864 1312
rect 9916 1300 9922 1352
rect 9953 1343 10011 1349
rect 9953 1309 9965 1343
rect 9999 1309 10011 1343
rect 9953 1303 10011 1309
rect 10045 1343 10103 1349
rect 10045 1309 10057 1343
rect 10091 1340 10103 1343
rect 10244 1340 10272 1380
rect 10091 1312 10272 1340
rect 10091 1309 10103 1312
rect 10045 1303 10103 1309
rect 9582 1272 9588 1284
rect 8956 1244 9588 1272
rect 9582 1232 9588 1244
rect 9640 1232 9646 1284
rect 9968 1272 9996 1303
rect 10318 1300 10324 1352
rect 10376 1300 10382 1352
rect 10428 1340 10456 1380
rect 10980 1380 11468 1408
rect 10502 1340 10508 1352
rect 10428 1312 10508 1340
rect 10502 1300 10508 1312
rect 10560 1300 10566 1352
rect 10597 1343 10655 1349
rect 10597 1309 10609 1343
rect 10643 1309 10655 1343
rect 10597 1303 10655 1309
rect 10873 1343 10931 1349
rect 10873 1309 10885 1343
rect 10919 1340 10931 1343
rect 10980 1340 11008 1380
rect 11440 1352 11468 1380
rect 12268 1380 12440 1408
rect 10919 1312 11008 1340
rect 11149 1343 11207 1349
rect 10919 1309 10931 1312
rect 10873 1303 10931 1309
rect 11149 1309 11161 1343
rect 11195 1309 11207 1343
rect 11149 1303 11207 1309
rect 10410 1272 10416 1284
rect 9968 1244 10416 1272
rect 10410 1232 10416 1244
rect 10468 1232 10474 1284
rect 10612 1272 10640 1303
rect 10962 1272 10968 1284
rect 10612 1244 10968 1272
rect 10962 1232 10968 1244
rect 11020 1232 11026 1284
rect 11164 1216 11192 1303
rect 11422 1300 11428 1352
rect 11480 1300 11486 1352
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1309 11575 1343
rect 11517 1303 11575 1309
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1340 11851 1343
rect 12069 1343 12127 1349
rect 11839 1312 12020 1340
rect 11839 1309 11851 1312
rect 11793 1303 11851 1309
rect 11532 1272 11560 1303
rect 11882 1272 11888 1284
rect 11532 1244 11888 1272
rect 11882 1232 11888 1244
rect 11940 1232 11946 1284
rect 11992 1272 12020 1312
rect 12069 1309 12081 1343
rect 12115 1340 12127 1343
rect 12268 1340 12296 1380
rect 12434 1368 12440 1380
rect 12492 1368 12498 1420
rect 14568 1408 14596 1516
rect 15286 1504 15292 1516
rect 15344 1504 15350 1556
rect 15473 1547 15531 1553
rect 15473 1513 15485 1547
rect 15519 1544 15531 1547
rect 16390 1544 16396 1556
rect 15519 1516 16396 1544
rect 15519 1513 15531 1516
rect 15473 1507 15531 1513
rect 16390 1504 16396 1516
rect 16448 1504 16454 1556
rect 17037 1547 17095 1553
rect 17037 1513 17049 1547
rect 17083 1544 17095 1547
rect 17402 1544 17408 1556
rect 17083 1516 17408 1544
rect 17083 1513 17095 1516
rect 17037 1507 17095 1513
rect 17402 1504 17408 1516
rect 17460 1504 17466 1556
rect 17497 1547 17555 1553
rect 17497 1513 17509 1547
rect 17543 1544 17555 1547
rect 17862 1544 17868 1556
rect 17543 1516 17868 1544
rect 17543 1513 17555 1516
rect 17497 1507 17555 1513
rect 17862 1504 17868 1516
rect 17920 1504 17926 1556
rect 18506 1504 18512 1556
rect 18564 1544 18570 1556
rect 22646 1544 22652 1556
rect 18564 1516 22652 1544
rect 18564 1504 18570 1516
rect 22646 1504 22652 1516
rect 22704 1504 22710 1556
rect 23382 1504 23388 1556
rect 23440 1544 23446 1556
rect 23661 1547 23719 1553
rect 23661 1544 23673 1547
rect 23440 1516 23673 1544
rect 23440 1504 23446 1516
rect 23661 1513 23673 1516
rect 23707 1513 23719 1547
rect 23661 1507 23719 1513
rect 24302 1504 24308 1556
rect 24360 1544 24366 1556
rect 24949 1547 25007 1553
rect 24949 1544 24961 1547
rect 24360 1516 24961 1544
rect 24360 1504 24366 1516
rect 24949 1513 24961 1516
rect 24995 1513 25007 1547
rect 24949 1507 25007 1513
rect 25501 1547 25559 1553
rect 25501 1513 25513 1547
rect 25547 1513 25559 1547
rect 25501 1507 25559 1513
rect 14645 1479 14703 1485
rect 14645 1445 14657 1479
rect 14691 1476 14703 1479
rect 14826 1476 14832 1488
rect 14691 1448 14832 1476
rect 14691 1445 14703 1448
rect 14645 1439 14703 1445
rect 14826 1436 14832 1448
rect 14884 1436 14890 1488
rect 15654 1476 15660 1488
rect 14936 1448 15660 1476
rect 14200 1380 14596 1408
rect 12115 1312 12296 1340
rect 12345 1343 12403 1349
rect 12115 1309 12127 1312
rect 12069 1303 12127 1309
rect 12345 1309 12357 1343
rect 12391 1340 12403 1343
rect 12526 1340 12532 1352
rect 12391 1312 12532 1340
rect 12391 1309 12403 1312
rect 12345 1303 12403 1309
rect 12526 1300 12532 1312
rect 12584 1300 12590 1352
rect 12618 1300 12624 1352
rect 12676 1300 12682 1352
rect 12897 1343 12955 1349
rect 12897 1309 12909 1343
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 12912 1272 12940 1303
rect 13170 1300 13176 1352
rect 13228 1300 13234 1352
rect 13354 1300 13360 1352
rect 13412 1300 13418 1352
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1340 13507 1343
rect 13722 1340 13728 1352
rect 13495 1312 13728 1340
rect 13495 1309 13507 1312
rect 13449 1303 13507 1309
rect 13722 1300 13728 1312
rect 13780 1300 13786 1352
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 13262 1272 13268 1284
rect 11992 1244 12388 1272
rect 12912 1244 13268 1272
rect 12360 1216 12388 1244
rect 13262 1232 13268 1244
rect 13320 1232 13326 1284
rect 7377 1207 7435 1213
rect 7377 1173 7389 1207
rect 7423 1173 7435 1207
rect 7377 1167 7435 1173
rect 7650 1164 7656 1216
rect 7708 1164 7714 1216
rect 7929 1207 7987 1213
rect 7929 1173 7941 1207
rect 7975 1204 7987 1207
rect 8110 1204 8116 1216
rect 7975 1176 8116 1204
rect 7975 1173 7987 1176
rect 7929 1167 7987 1173
rect 8110 1164 8116 1176
rect 8168 1164 8174 1216
rect 8205 1207 8263 1213
rect 8205 1173 8217 1207
rect 8251 1204 8263 1207
rect 8294 1204 8300 1216
rect 8251 1176 8300 1204
rect 8251 1173 8263 1176
rect 8205 1167 8263 1173
rect 8294 1164 8300 1176
rect 8352 1164 8358 1216
rect 8481 1207 8539 1213
rect 8481 1173 8493 1207
rect 8527 1204 8539 1207
rect 8662 1204 8668 1216
rect 8527 1176 8668 1204
rect 8527 1173 8539 1176
rect 8481 1167 8539 1173
rect 8662 1164 8668 1176
rect 8720 1164 8726 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9125 1207 9183 1213
rect 9125 1173 9137 1207
rect 9171 1204 9183 1207
rect 9306 1204 9312 1216
rect 9171 1176 9312 1204
rect 9171 1173 9183 1176
rect 9125 1167 9183 1173
rect 9306 1164 9312 1176
rect 9364 1164 9370 1216
rect 9398 1164 9404 1216
rect 9456 1164 9462 1216
rect 9769 1207 9827 1213
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10134 1204 10140 1216
rect 9815 1176 10140 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10134 1164 10140 1176
rect 10192 1164 10198 1216
rect 10226 1164 10232 1216
rect 10284 1164 10290 1216
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 10686 1204 10692 1216
rect 10551 1176 10692 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 10686 1164 10692 1176
rect 10744 1164 10750 1216
rect 10778 1164 10784 1216
rect 10836 1164 10842 1216
rect 11146 1164 11152 1216
rect 11204 1164 11210 1216
rect 11238 1164 11244 1216
rect 11296 1204 11302 1216
rect 11701 1207 11759 1213
rect 11701 1204 11713 1207
rect 11296 1176 11713 1204
rect 11296 1164 11302 1176
rect 11701 1173 11713 1176
rect 11747 1173 11759 1207
rect 11701 1167 11759 1173
rect 11974 1164 11980 1216
rect 12032 1164 12038 1216
rect 12250 1164 12256 1216
rect 12308 1164 12314 1216
rect 12342 1164 12348 1216
rect 12400 1164 12406 1216
rect 12529 1207 12587 1213
rect 12529 1173 12541 1207
rect 12575 1204 12587 1207
rect 12894 1204 12900 1216
rect 12575 1176 12900 1204
rect 12575 1173 12587 1176
rect 12529 1167 12587 1173
rect 12894 1164 12900 1176
rect 12952 1164 12958 1216
rect 12986 1164 12992 1216
rect 13044 1204 13050 1216
rect 13372 1213 13400 1300
rect 13081 1207 13139 1213
rect 13081 1204 13093 1207
rect 13044 1176 13093 1204
rect 13044 1164 13050 1176
rect 13081 1173 13093 1176
rect 13127 1173 13139 1207
rect 13081 1167 13139 1173
rect 13357 1207 13415 1213
rect 13357 1173 13369 1207
rect 13403 1173 13415 1207
rect 13357 1167 13415 1173
rect 13630 1164 13636 1216
rect 13688 1164 13694 1216
rect 13725 1207 13783 1213
rect 13725 1173 13737 1207
rect 13771 1204 13783 1207
rect 14200 1204 14228 1380
rect 14277 1343 14335 1349
rect 14277 1309 14289 1343
rect 14323 1309 14335 1343
rect 14277 1303 14335 1309
rect 14553 1343 14611 1349
rect 14553 1309 14565 1343
rect 14599 1340 14611 1343
rect 14734 1340 14740 1352
rect 14599 1312 14740 1340
rect 14599 1309 14611 1312
rect 14553 1303 14611 1309
rect 14292 1272 14320 1303
rect 14734 1300 14740 1312
rect 14792 1300 14798 1352
rect 14829 1343 14887 1349
rect 14829 1309 14841 1343
rect 14875 1340 14887 1343
rect 14936 1340 14964 1448
rect 15654 1436 15660 1448
rect 15712 1436 15718 1488
rect 16025 1479 16083 1485
rect 16025 1445 16037 1479
rect 16071 1476 16083 1479
rect 17126 1476 17132 1488
rect 16071 1448 17132 1476
rect 16071 1445 16083 1448
rect 16025 1439 16083 1445
rect 17126 1436 17132 1448
rect 17184 1436 17190 1488
rect 17770 1476 17776 1488
rect 17236 1448 17776 1476
rect 15562 1408 15568 1420
rect 14875 1312 14964 1340
rect 15028 1380 15568 1408
rect 14875 1309 14887 1312
rect 14829 1303 14887 1309
rect 15028 1272 15056 1380
rect 15562 1368 15568 1380
rect 15620 1368 15626 1420
rect 16758 1368 16764 1420
rect 16816 1408 16822 1420
rect 17236 1408 17264 1448
rect 17770 1436 17776 1448
rect 17828 1436 17834 1488
rect 18046 1436 18052 1488
rect 18104 1476 18110 1488
rect 18598 1476 18604 1488
rect 18104 1448 18604 1476
rect 18104 1436 18110 1448
rect 18598 1436 18604 1448
rect 18656 1436 18662 1488
rect 18690 1436 18696 1488
rect 18748 1476 18754 1488
rect 18748 1448 19380 1476
rect 18748 1436 18754 1448
rect 16816 1380 17264 1408
rect 17328 1380 18092 1408
rect 16816 1368 16822 1380
rect 15105 1343 15163 1349
rect 15105 1309 15117 1343
rect 15151 1340 15163 1343
rect 15194 1340 15200 1352
rect 15151 1312 15200 1340
rect 15151 1309 15163 1312
rect 15105 1303 15163 1309
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
rect 15378 1300 15384 1352
rect 15436 1300 15442 1352
rect 15654 1300 15660 1352
rect 15712 1300 15718 1352
rect 15930 1300 15936 1352
rect 15988 1300 15994 1352
rect 16209 1343 16267 1349
rect 16209 1309 16221 1343
rect 16255 1340 16267 1343
rect 16390 1340 16396 1352
rect 16255 1312 16396 1340
rect 16255 1309 16267 1312
rect 16209 1303 16267 1309
rect 16390 1300 16396 1312
rect 16448 1300 16454 1352
rect 16482 1300 16488 1352
rect 16540 1300 16546 1352
rect 16853 1343 16911 1349
rect 16853 1309 16865 1343
rect 16899 1309 16911 1343
rect 17328 1340 17356 1380
rect 16853 1303 16911 1309
rect 16960 1312 17356 1340
rect 16868 1272 16896 1303
rect 14292 1244 15056 1272
rect 15212 1244 16896 1272
rect 13771 1176 14228 1204
rect 13771 1173 13783 1176
rect 13725 1167 13783 1173
rect 14366 1164 14372 1216
rect 14424 1164 14430 1216
rect 14921 1207 14979 1213
rect 14921 1173 14933 1207
rect 14967 1204 14979 1207
rect 15010 1204 15016 1216
rect 14967 1176 15016 1204
rect 14967 1173 14979 1176
rect 14921 1167 14979 1173
rect 15010 1164 15016 1176
rect 15068 1164 15074 1216
rect 15212 1213 15240 1244
rect 15197 1207 15255 1213
rect 15197 1173 15209 1207
rect 15243 1173 15255 1207
rect 15197 1167 15255 1173
rect 15746 1164 15752 1216
rect 15804 1164 15810 1216
rect 16301 1207 16359 1213
rect 16301 1173 16313 1207
rect 16347 1204 16359 1207
rect 16960 1204 16988 1312
rect 17402 1300 17408 1352
rect 17460 1300 17466 1352
rect 17678 1300 17684 1352
rect 17736 1300 17742 1352
rect 17954 1300 17960 1352
rect 18012 1300 18018 1352
rect 18064 1349 18092 1380
rect 18432 1380 18644 1408
rect 18049 1343 18107 1349
rect 18049 1309 18061 1343
rect 18095 1309 18107 1343
rect 18049 1303 18107 1309
rect 18432 1272 18460 1380
rect 18616 1349 18644 1380
rect 18874 1368 18880 1420
rect 18932 1408 18938 1420
rect 18932 1380 19104 1408
rect 18932 1368 18938 1380
rect 18509 1343 18567 1349
rect 18509 1309 18521 1343
rect 18555 1309 18567 1343
rect 18509 1303 18567 1309
rect 18601 1343 18659 1349
rect 18601 1309 18613 1343
rect 18647 1309 18659 1343
rect 18966 1340 18972 1352
rect 18601 1303 18659 1309
rect 18800 1312 18972 1340
rect 17236 1244 18460 1272
rect 18524 1272 18552 1303
rect 18800 1272 18828 1312
rect 18966 1300 18972 1312
rect 19024 1300 19030 1352
rect 19076 1349 19104 1380
rect 19352 1349 19380 1448
rect 20162 1436 20168 1488
rect 20220 1476 20226 1488
rect 20220 1448 20392 1476
rect 20220 1436 20226 1448
rect 19536 1380 20208 1408
rect 19536 1352 19564 1380
rect 19061 1343 19119 1349
rect 19061 1309 19073 1343
rect 19107 1309 19119 1343
rect 19061 1303 19119 1309
rect 19337 1343 19395 1349
rect 19337 1309 19349 1343
rect 19383 1309 19395 1343
rect 19337 1303 19395 1309
rect 19518 1300 19524 1352
rect 19576 1300 19582 1352
rect 20180 1349 20208 1380
rect 19705 1343 19763 1349
rect 19705 1340 19717 1343
rect 19702 1309 19717 1340
rect 19751 1309 19763 1343
rect 19702 1303 19763 1309
rect 20165 1343 20223 1349
rect 20165 1309 20177 1343
rect 20211 1309 20223 1343
rect 20364 1340 20392 1448
rect 20898 1436 20904 1488
rect 20956 1436 20962 1488
rect 24670 1436 24676 1488
rect 24728 1476 24734 1488
rect 25516 1476 25544 1507
rect 26142 1504 26148 1556
rect 26200 1544 26206 1556
rect 27709 1547 27767 1553
rect 27709 1544 27721 1547
rect 26200 1516 27721 1544
rect 26200 1504 26206 1516
rect 27709 1513 27721 1516
rect 27755 1513 27767 1547
rect 27709 1507 27767 1513
rect 28813 1547 28871 1553
rect 28813 1513 28825 1547
rect 28859 1513 28871 1547
rect 28813 1507 28871 1513
rect 29181 1547 29239 1553
rect 29181 1513 29193 1547
rect 29227 1544 29239 1547
rect 29454 1544 29460 1556
rect 29227 1516 29460 1544
rect 29227 1513 29239 1516
rect 29181 1507 29239 1513
rect 24728 1448 25544 1476
rect 27249 1479 27307 1485
rect 24728 1436 24734 1448
rect 27249 1445 27261 1479
rect 27295 1445 27307 1479
rect 27249 1439 27307 1445
rect 20438 1368 20444 1420
rect 20496 1368 20502 1420
rect 22373 1411 22431 1417
rect 22373 1377 22385 1411
rect 22419 1408 22431 1411
rect 22554 1408 22560 1420
rect 22419 1380 22560 1408
rect 22419 1377 22431 1380
rect 22373 1371 22431 1377
rect 22554 1368 22560 1380
rect 22612 1368 22618 1420
rect 25498 1368 25504 1420
rect 25556 1408 25562 1420
rect 27264 1408 27292 1439
rect 27614 1436 27620 1488
rect 27672 1476 27678 1488
rect 28828 1476 28856 1507
rect 29454 1504 29460 1516
rect 29512 1504 29518 1556
rect 30834 1504 30840 1556
rect 30892 1544 30898 1556
rect 31389 1547 31447 1553
rect 31389 1544 31401 1547
rect 30892 1516 31401 1544
rect 30892 1504 30898 1516
rect 31389 1513 31401 1516
rect 31435 1513 31447 1547
rect 32861 1547 32919 1553
rect 32861 1544 32873 1547
rect 31389 1507 31447 1513
rect 31864 1516 32873 1544
rect 27672 1448 28856 1476
rect 27672 1436 27678 1448
rect 29086 1436 29092 1488
rect 29144 1476 29150 1488
rect 29546 1476 29552 1488
rect 29144 1448 29552 1476
rect 29144 1436 29150 1448
rect 29546 1436 29552 1448
rect 29604 1436 29610 1488
rect 29638 1436 29644 1488
rect 29696 1476 29702 1488
rect 30929 1479 30987 1485
rect 30929 1476 30941 1479
rect 29696 1448 30941 1476
rect 29696 1436 29702 1448
rect 30929 1445 30941 1448
rect 30975 1445 30987 1479
rect 30929 1439 30987 1445
rect 31018 1436 31024 1488
rect 31076 1476 31082 1488
rect 31757 1479 31815 1485
rect 31757 1476 31769 1479
rect 31076 1448 31769 1476
rect 31076 1436 31082 1448
rect 31757 1445 31769 1448
rect 31803 1445 31815 1479
rect 31757 1439 31815 1445
rect 25556 1380 27292 1408
rect 25556 1368 25562 1380
rect 27706 1368 27712 1420
rect 27764 1408 27770 1420
rect 29917 1411 29975 1417
rect 29917 1408 29929 1411
rect 27764 1380 29929 1408
rect 27764 1368 27770 1380
rect 29917 1377 29929 1380
rect 29963 1377 29975 1411
rect 29917 1371 29975 1377
rect 30466 1368 30472 1420
rect 30524 1408 30530 1420
rect 31864 1408 31892 1516
rect 32861 1513 32873 1516
rect 32907 1513 32919 1547
rect 32861 1507 32919 1513
rect 32950 1504 32956 1556
rect 33008 1544 33014 1556
rect 33965 1547 34023 1553
rect 33965 1544 33977 1547
rect 33008 1516 33977 1544
rect 33008 1504 33014 1516
rect 33965 1513 33977 1516
rect 34011 1513 34023 1547
rect 33965 1507 34023 1513
rect 34974 1504 34980 1556
rect 35032 1544 35038 1556
rect 35805 1547 35863 1553
rect 35805 1544 35817 1547
rect 35032 1516 35817 1544
rect 35032 1504 35038 1516
rect 35805 1513 35817 1516
rect 35851 1513 35863 1547
rect 35805 1507 35863 1513
rect 35894 1504 35900 1556
rect 35952 1544 35958 1556
rect 36357 1547 36415 1553
rect 36357 1544 36369 1547
rect 35952 1516 36369 1544
rect 35952 1504 35958 1516
rect 36357 1513 36369 1516
rect 36403 1513 36415 1547
rect 36357 1507 36415 1513
rect 36446 1504 36452 1556
rect 36504 1544 36510 1556
rect 37461 1547 37519 1553
rect 37461 1544 37473 1547
rect 36504 1516 37473 1544
rect 36504 1504 36510 1516
rect 37461 1513 37473 1516
rect 37507 1513 37519 1547
rect 37461 1507 37519 1513
rect 37642 1504 37648 1556
rect 37700 1544 37706 1556
rect 37700 1516 38332 1544
rect 37700 1504 37706 1516
rect 32490 1436 32496 1488
rect 32548 1436 32554 1488
rect 33134 1436 33140 1488
rect 33192 1476 33198 1488
rect 34333 1479 34391 1485
rect 34333 1476 34345 1479
rect 33192 1448 34345 1476
rect 33192 1436 33198 1448
rect 34333 1445 34345 1448
rect 34379 1445 34391 1479
rect 34333 1439 34391 1445
rect 35710 1436 35716 1488
rect 35768 1476 35774 1488
rect 37737 1479 37795 1485
rect 37737 1476 37749 1479
rect 35768 1448 37749 1476
rect 35768 1436 35774 1448
rect 37737 1445 37749 1448
rect 37783 1445 37795 1479
rect 37737 1439 37795 1445
rect 38304 1408 38332 1516
rect 38378 1504 38384 1556
rect 38436 1544 38442 1556
rect 39853 1547 39911 1553
rect 39853 1544 39865 1547
rect 38436 1516 39865 1544
rect 38436 1504 38442 1516
rect 39853 1513 39865 1516
rect 39899 1513 39911 1547
rect 39853 1507 39911 1513
rect 40126 1504 40132 1556
rect 40184 1544 40190 1556
rect 41509 1547 41567 1553
rect 41509 1544 41521 1547
rect 40184 1516 41521 1544
rect 40184 1504 40190 1516
rect 41509 1513 41521 1516
rect 41555 1513 41567 1547
rect 41509 1507 41567 1513
rect 41782 1504 41788 1556
rect 41840 1504 41846 1556
rect 40954 1436 40960 1488
rect 41012 1436 41018 1488
rect 41230 1436 41236 1488
rect 41288 1436 41294 1488
rect 30524 1380 31892 1408
rect 35084 1380 35848 1408
rect 30524 1368 30530 1380
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 20364 1312 21373 1340
rect 20165 1303 20223 1309
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 21361 1303 21419 1309
rect 19702 1272 19730 1303
rect 21542 1300 21548 1352
rect 21600 1340 21606 1352
rect 22097 1343 22155 1349
rect 22097 1340 22109 1343
rect 21600 1312 22109 1340
rect 21600 1300 21606 1312
rect 22097 1309 22109 1312
rect 22143 1309 22155 1343
rect 22097 1303 22155 1309
rect 22741 1343 22799 1349
rect 22741 1309 22753 1343
rect 22787 1309 22799 1343
rect 22741 1303 22799 1309
rect 18524 1244 18828 1272
rect 18892 1244 19730 1272
rect 17236 1213 17264 1244
rect 16347 1176 16988 1204
rect 17221 1207 17279 1213
rect 16347 1173 16359 1176
rect 16301 1167 16359 1173
rect 17221 1173 17233 1207
rect 17267 1173 17279 1207
rect 17221 1167 17279 1173
rect 17770 1164 17776 1216
rect 17828 1164 17834 1216
rect 18230 1164 18236 1216
rect 18288 1164 18294 1216
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1204 18383 1207
rect 18690 1204 18696 1216
rect 18371 1176 18696 1204
rect 18371 1173 18383 1176
rect 18325 1167 18383 1173
rect 18690 1164 18696 1176
rect 18748 1164 18754 1216
rect 18782 1164 18788 1216
rect 18840 1164 18846 1216
rect 18892 1213 18920 1244
rect 20530 1232 20536 1284
rect 20588 1272 20594 1284
rect 20717 1275 20775 1281
rect 20717 1272 20729 1275
rect 20588 1244 20729 1272
rect 20588 1232 20594 1244
rect 20717 1241 20729 1244
rect 20763 1241 20775 1275
rect 20717 1235 20775 1241
rect 21910 1232 21916 1284
rect 21968 1272 21974 1284
rect 22756 1272 22784 1303
rect 22922 1300 22928 1352
rect 22980 1340 22986 1352
rect 23109 1343 23167 1349
rect 23109 1340 23121 1343
rect 22980 1312 23121 1340
rect 22980 1300 22986 1312
rect 23109 1309 23121 1312
rect 23155 1309 23167 1343
rect 23109 1303 23167 1309
rect 23474 1300 23480 1352
rect 23532 1340 23538 1352
rect 23569 1343 23627 1349
rect 23569 1340 23581 1343
rect 23532 1312 23581 1340
rect 23532 1300 23538 1312
rect 23569 1309 23581 1312
rect 23615 1309 23627 1343
rect 23569 1303 23627 1309
rect 24397 1343 24455 1349
rect 24397 1309 24409 1343
rect 24443 1309 24455 1343
rect 24397 1303 24455 1309
rect 24412 1272 24440 1303
rect 24762 1300 24768 1352
rect 24820 1340 24826 1352
rect 25409 1343 25467 1349
rect 25409 1340 25421 1343
rect 24820 1312 25421 1340
rect 24820 1300 24826 1312
rect 25409 1309 25421 1312
rect 25455 1309 25467 1343
rect 25409 1303 25467 1309
rect 25682 1300 25688 1352
rect 25740 1340 25746 1352
rect 25740 1312 26188 1340
rect 25740 1300 25746 1312
rect 21968 1244 22784 1272
rect 22848 1244 24440 1272
rect 21968 1232 21974 1244
rect 18877 1207 18935 1213
rect 18877 1173 18889 1207
rect 18923 1173 18935 1207
rect 18877 1167 18935 1173
rect 19521 1207 19579 1213
rect 19521 1173 19533 1207
rect 19567 1204 19579 1207
rect 19794 1204 19800 1216
rect 19567 1176 19800 1204
rect 19567 1173 19579 1176
rect 19521 1167 19579 1173
rect 19794 1164 19800 1176
rect 19852 1164 19858 1216
rect 19886 1164 19892 1216
rect 19944 1164 19950 1216
rect 21542 1164 21548 1216
rect 21600 1164 21606 1216
rect 21818 1164 21824 1216
rect 21876 1204 21882 1216
rect 22848 1204 22876 1244
rect 24854 1232 24860 1284
rect 24912 1232 24918 1284
rect 25038 1232 25044 1284
rect 25096 1272 25102 1284
rect 25961 1275 26019 1281
rect 25961 1272 25973 1275
rect 25096 1244 25973 1272
rect 25096 1232 25102 1244
rect 25961 1241 25973 1244
rect 26007 1241 26019 1275
rect 26160 1272 26188 1312
rect 26234 1300 26240 1352
rect 26292 1340 26298 1352
rect 26421 1343 26479 1349
rect 26421 1340 26433 1343
rect 26292 1312 26433 1340
rect 26292 1300 26298 1312
rect 26421 1309 26433 1312
rect 26467 1309 26479 1343
rect 26421 1303 26479 1309
rect 26510 1300 26516 1352
rect 26568 1340 26574 1352
rect 26568 1312 27292 1340
rect 26568 1300 26574 1312
rect 27065 1275 27123 1281
rect 27065 1272 27077 1275
rect 26160 1244 27077 1272
rect 25961 1235 26019 1241
rect 27065 1241 27077 1244
rect 27111 1241 27123 1275
rect 27264 1272 27292 1312
rect 27338 1300 27344 1352
rect 27396 1340 27402 1352
rect 27617 1343 27675 1349
rect 27617 1340 27629 1343
rect 27396 1312 27629 1340
rect 27396 1300 27402 1312
rect 27617 1309 27629 1312
rect 27663 1309 27675 1343
rect 27617 1303 27675 1309
rect 27890 1300 27896 1352
rect 27948 1340 27954 1352
rect 28721 1343 28779 1349
rect 28721 1340 28733 1343
rect 27948 1312 28733 1340
rect 27948 1300 27954 1312
rect 28721 1309 28733 1312
rect 28767 1309 28779 1343
rect 28721 1303 28779 1309
rect 28810 1300 28816 1352
rect 28868 1300 28874 1352
rect 28994 1300 29000 1352
rect 29052 1340 29058 1352
rect 29365 1343 29423 1349
rect 29365 1340 29377 1343
rect 29052 1312 29377 1340
rect 29052 1300 29058 1312
rect 29365 1309 29377 1312
rect 29411 1309 29423 1343
rect 29365 1303 29423 1309
rect 30098 1300 30104 1352
rect 30156 1340 30162 1352
rect 30193 1343 30251 1349
rect 30193 1340 30205 1343
rect 30156 1312 30205 1340
rect 30156 1300 30162 1312
rect 30193 1309 30205 1312
rect 30239 1309 30251 1343
rect 30193 1303 30251 1309
rect 31938 1300 31944 1352
rect 31996 1300 32002 1352
rect 33962 1300 33968 1352
rect 34020 1340 34026 1352
rect 34517 1343 34575 1349
rect 34517 1340 34529 1343
rect 34020 1312 34529 1340
rect 34020 1300 34026 1312
rect 34517 1309 34529 1312
rect 34563 1309 34575 1343
rect 35084 1340 35112 1380
rect 34517 1303 34575 1309
rect 34624 1312 35112 1340
rect 28169 1275 28227 1281
rect 28169 1272 28181 1275
rect 27264 1244 28181 1272
rect 27065 1235 27123 1241
rect 28169 1241 28181 1244
rect 28215 1241 28227 1275
rect 28828 1272 28856 1300
rect 29641 1275 29699 1281
rect 29641 1272 29653 1275
rect 28828 1244 29653 1272
rect 28169 1235 28227 1241
rect 29641 1241 29653 1244
rect 29687 1241 29699 1275
rect 29641 1235 29699 1241
rect 30742 1232 30748 1284
rect 30800 1232 30806 1284
rect 30926 1232 30932 1284
rect 30984 1272 30990 1284
rect 31297 1275 31355 1281
rect 31297 1272 31309 1275
rect 30984 1244 31309 1272
rect 30984 1232 30990 1244
rect 31297 1241 31309 1244
rect 31343 1241 31355 1275
rect 31297 1235 31355 1241
rect 32214 1232 32220 1284
rect 32272 1232 32278 1284
rect 32306 1232 32312 1284
rect 32364 1272 32370 1284
rect 32769 1275 32827 1281
rect 32769 1272 32781 1275
rect 32364 1244 32781 1272
rect 32364 1232 32370 1244
rect 32769 1241 32781 1244
rect 32815 1241 32827 1275
rect 32769 1235 32827 1241
rect 33873 1275 33931 1281
rect 33873 1241 33885 1275
rect 33919 1241 33931 1275
rect 33873 1235 33931 1241
rect 21876 1176 22876 1204
rect 21876 1164 21882 1176
rect 22922 1164 22928 1216
rect 22980 1164 22986 1216
rect 23290 1164 23296 1216
rect 23348 1164 23354 1216
rect 23658 1164 23664 1216
rect 23716 1204 23722 1216
rect 24581 1207 24639 1213
rect 24581 1204 24593 1207
rect 23716 1176 24593 1204
rect 23716 1164 23722 1176
rect 24581 1173 24593 1176
rect 24627 1173 24639 1207
rect 24581 1167 24639 1173
rect 24762 1164 24768 1216
rect 24820 1204 24826 1216
rect 26053 1207 26111 1213
rect 26053 1204 26065 1207
rect 24820 1176 26065 1204
rect 24820 1164 24826 1176
rect 26053 1173 26065 1176
rect 26099 1173 26111 1207
rect 26053 1167 26111 1173
rect 26142 1164 26148 1216
rect 26200 1204 26206 1216
rect 26605 1207 26663 1213
rect 26605 1204 26617 1207
rect 26200 1176 26617 1204
rect 26200 1164 26206 1176
rect 26605 1173 26617 1176
rect 26651 1173 26663 1207
rect 26605 1167 26663 1173
rect 26878 1164 26884 1216
rect 26936 1204 26942 1216
rect 28261 1207 28319 1213
rect 28261 1204 28273 1207
rect 26936 1176 28273 1204
rect 26936 1164 26942 1176
rect 28261 1173 28273 1176
rect 28307 1173 28319 1207
rect 28261 1167 28319 1173
rect 30282 1164 30288 1216
rect 30340 1164 30346 1216
rect 32122 1164 32128 1216
rect 32180 1204 32186 1216
rect 33413 1207 33471 1213
rect 33413 1204 33425 1207
rect 32180 1176 33425 1204
rect 32180 1164 32186 1176
rect 33413 1173 33425 1176
rect 33459 1204 33471 1207
rect 33888 1204 33916 1235
rect 34422 1232 34428 1284
rect 34480 1272 34486 1284
rect 34624 1272 34652 1312
rect 35158 1300 35164 1352
rect 35216 1340 35222 1352
rect 35713 1343 35771 1349
rect 35713 1340 35725 1343
rect 35216 1312 35725 1340
rect 35216 1300 35222 1312
rect 35713 1309 35725 1312
rect 35759 1309 35771 1343
rect 35820 1340 35848 1380
rect 37384 1380 37780 1408
rect 38304 1380 38608 1408
rect 36725 1343 36783 1349
rect 36725 1340 36737 1343
rect 35820 1312 36737 1340
rect 35713 1303 35771 1309
rect 36725 1309 36737 1312
rect 36771 1309 36783 1343
rect 36725 1303 36783 1309
rect 36814 1300 36820 1352
rect 36872 1340 36878 1352
rect 37277 1343 37335 1349
rect 37277 1340 37289 1343
rect 36872 1312 37289 1340
rect 36872 1300 36878 1312
rect 37277 1309 37289 1312
rect 37323 1309 37335 1343
rect 37277 1303 37335 1309
rect 34480 1244 34652 1272
rect 34793 1275 34851 1281
rect 34480 1232 34486 1244
rect 34793 1241 34805 1275
rect 34839 1272 34851 1275
rect 35437 1275 35495 1281
rect 35437 1272 35449 1275
rect 34839 1244 35449 1272
rect 34839 1241 34851 1244
rect 34793 1235 34851 1241
rect 35437 1241 35449 1244
rect 35483 1241 35495 1275
rect 35437 1235 35495 1241
rect 33459 1176 33916 1204
rect 33459 1173 33471 1176
rect 33413 1167 33471 1173
rect 34514 1164 34520 1216
rect 34572 1204 34578 1216
rect 34808 1204 34836 1235
rect 36262 1232 36268 1284
rect 36320 1232 36326 1284
rect 37384 1272 37412 1380
rect 37458 1300 37464 1352
rect 37516 1300 37522 1352
rect 37553 1343 37611 1349
rect 37553 1309 37565 1343
rect 37599 1340 37611 1343
rect 37642 1340 37648 1352
rect 37599 1312 37648 1340
rect 37599 1309 37611 1312
rect 37553 1303 37611 1309
rect 37642 1300 37648 1312
rect 37700 1300 37706 1352
rect 37752 1340 37780 1380
rect 37829 1343 37887 1349
rect 37829 1340 37841 1343
rect 37752 1312 37841 1340
rect 37829 1309 37841 1312
rect 37875 1309 37887 1343
rect 37829 1303 37887 1309
rect 38102 1300 38108 1352
rect 38160 1300 38166 1352
rect 38378 1300 38384 1352
rect 38436 1300 38442 1352
rect 36372 1244 37412 1272
rect 37476 1272 37504 1300
rect 38580 1272 38608 1380
rect 39574 1368 39580 1420
rect 39632 1408 39638 1420
rect 39632 1380 41828 1408
rect 39632 1368 39638 1380
rect 38654 1300 38660 1352
rect 38712 1300 38718 1352
rect 38930 1300 38936 1352
rect 38988 1300 38994 1352
rect 39206 1300 39212 1352
rect 39264 1300 39270 1352
rect 39482 1300 39488 1352
rect 39540 1300 39546 1352
rect 40034 1300 40040 1352
rect 40092 1300 40098 1352
rect 40310 1300 40316 1352
rect 40368 1300 40374 1352
rect 40586 1300 40592 1352
rect 40644 1300 40650 1352
rect 40862 1300 40868 1352
rect 40920 1300 40926 1352
rect 41138 1300 41144 1352
rect 41196 1300 41202 1352
rect 41414 1300 41420 1352
rect 41472 1300 41478 1352
rect 41690 1300 41696 1352
rect 41748 1300 41754 1352
rect 41800 1340 41828 1380
rect 41969 1343 42027 1349
rect 41969 1340 41981 1343
rect 41800 1312 41981 1340
rect 41969 1309 41981 1312
rect 42015 1309 42027 1343
rect 41969 1303 42027 1309
rect 37476 1244 38332 1272
rect 38580 1244 40448 1272
rect 34572 1176 34836 1204
rect 34572 1164 34578 1176
rect 34882 1164 34888 1216
rect 34940 1164 34946 1216
rect 35710 1164 35716 1216
rect 35768 1204 35774 1216
rect 36372 1204 36400 1244
rect 35768 1176 36400 1204
rect 35768 1164 35774 1176
rect 36906 1164 36912 1216
rect 36964 1164 36970 1216
rect 37826 1164 37832 1216
rect 37884 1204 37890 1216
rect 38304 1213 38332 1244
rect 38013 1207 38071 1213
rect 38013 1204 38025 1207
rect 37884 1176 38025 1204
rect 37884 1164 37890 1176
rect 38013 1173 38025 1176
rect 38059 1173 38071 1207
rect 38013 1167 38071 1173
rect 38289 1207 38347 1213
rect 38289 1173 38301 1207
rect 38335 1173 38347 1207
rect 38289 1167 38347 1173
rect 38565 1207 38623 1213
rect 38565 1173 38577 1207
rect 38611 1204 38623 1207
rect 38654 1204 38660 1216
rect 38611 1176 38660 1204
rect 38611 1173 38623 1176
rect 38565 1167 38623 1173
rect 38654 1164 38660 1176
rect 38712 1164 38718 1216
rect 38838 1164 38844 1216
rect 38896 1164 38902 1216
rect 39114 1164 39120 1216
rect 39172 1164 39178 1216
rect 39298 1164 39304 1216
rect 39356 1204 39362 1216
rect 39393 1207 39451 1213
rect 39393 1204 39405 1207
rect 39356 1176 39405 1204
rect 39356 1164 39362 1176
rect 39393 1173 39405 1176
rect 39439 1173 39451 1207
rect 39393 1167 39451 1173
rect 39666 1164 39672 1216
rect 39724 1164 39730 1216
rect 40126 1164 40132 1216
rect 40184 1164 40190 1216
rect 40420 1213 40448 1244
rect 40405 1207 40463 1213
rect 40405 1173 40417 1207
rect 40451 1173 40463 1207
rect 40405 1167 40463 1173
rect 40678 1164 40684 1216
rect 40736 1164 40742 1216
rect 1104 1114 43675 1136
rect 1104 1062 11552 1114
rect 11604 1062 11616 1114
rect 11668 1062 11680 1114
rect 11732 1062 11744 1114
rect 11796 1062 11808 1114
rect 11860 1062 22155 1114
rect 22207 1062 22219 1114
rect 22271 1062 22283 1114
rect 22335 1062 22347 1114
rect 22399 1062 22411 1114
rect 22463 1062 32758 1114
rect 32810 1062 32822 1114
rect 32874 1062 32886 1114
rect 32938 1062 32950 1114
rect 33002 1062 33014 1114
rect 33066 1062 43361 1114
rect 43413 1062 43425 1114
rect 43477 1062 43489 1114
rect 43541 1062 43553 1114
rect 43605 1062 43617 1114
rect 43669 1062 43675 1114
rect 1104 1040 43675 1062
rect 4798 960 4804 1012
rect 4856 960 4862 1012
rect 6546 960 6552 1012
rect 6604 1000 6610 1012
rect 9214 1000 9220 1012
rect 6604 972 9220 1000
rect 6604 960 6610 972
rect 9214 960 9220 972
rect 9272 960 9278 1012
rect 12894 960 12900 1012
rect 12952 1000 12958 1012
rect 13630 1000 13636 1012
rect 12952 972 13636 1000
rect 12952 960 12958 972
rect 13630 960 13636 972
rect 13688 960 13694 1012
rect 14366 960 14372 1012
rect 14424 1000 14430 1012
rect 15470 1000 15476 1012
rect 14424 972 15476 1000
rect 14424 960 14430 972
rect 15470 960 15476 972
rect 15528 960 15534 1012
rect 15930 960 15936 1012
rect 15988 1000 15994 1012
rect 17494 1000 17500 1012
rect 15988 972 17500 1000
rect 15988 960 15994 972
rect 17494 960 17500 972
rect 17552 960 17558 1012
rect 18230 960 18236 1012
rect 18288 960 18294 1012
rect 18782 960 18788 1012
rect 18840 1000 18846 1012
rect 32306 1000 32312 1012
rect 18840 972 32312 1000
rect 18840 960 18846 972
rect 32306 960 32312 972
rect 32364 960 32370 1012
rect 32766 960 32772 1012
rect 32824 1000 32830 1012
rect 34974 1000 34980 1012
rect 32824 972 34980 1000
rect 32824 960 32830 972
rect 34974 960 34980 972
rect 35032 960 35038 1012
rect 36078 960 36084 1012
rect 36136 1000 36142 1012
rect 38378 1000 38384 1012
rect 36136 972 38384 1000
rect 36136 960 36142 972
rect 38378 960 38384 972
rect 38436 960 38442 1012
rect 40126 1000 40132 1012
rect 38626 972 40132 1000
rect 4816 932 4844 960
rect 9030 932 9036 944
rect 4816 904 9036 932
rect 9030 892 9036 904
rect 9088 892 9094 944
rect 10226 892 10232 944
rect 10284 932 10290 944
rect 16482 932 16488 944
rect 10284 904 12572 932
rect 10284 892 10290 904
rect 5810 824 5816 876
rect 5868 864 5874 876
rect 5868 836 6914 864
rect 5868 824 5874 836
rect 4890 416 4896 468
rect 4948 416 4954 468
rect 6086 416 6092 468
rect 6144 416 6150 468
rect 6886 456 6914 836
rect 9306 824 9312 876
rect 9364 864 9370 876
rect 12544 864 12572 904
rect 15672 904 16488 932
rect 15672 864 15700 904
rect 16482 892 16488 904
rect 16540 892 16546 944
rect 18046 932 18052 944
rect 16592 904 18052 932
rect 9364 836 12434 864
rect 12544 836 15700 864
rect 9364 824 9370 836
rect 7650 756 7656 808
rect 7708 796 7714 808
rect 12158 796 12164 808
rect 7708 768 12164 796
rect 7708 756 7714 768
rect 12158 756 12164 768
rect 12216 756 12222 808
rect 12406 796 12434 836
rect 15746 824 15752 876
rect 15804 864 15810 876
rect 16592 864 16620 904
rect 18046 892 18052 904
rect 18104 892 18110 944
rect 18248 932 18276 960
rect 23750 932 23756 944
rect 18248 904 23756 932
rect 23750 892 23756 904
rect 23808 892 23814 944
rect 23842 892 23848 944
rect 23900 932 23906 944
rect 23900 904 31754 932
rect 23900 892 23906 904
rect 15804 836 16620 864
rect 15804 824 15810 836
rect 17402 824 17408 876
rect 17460 864 17466 876
rect 18414 864 18420 876
rect 17460 836 18420 864
rect 17460 824 17466 836
rect 18414 824 18420 836
rect 18472 824 18478 876
rect 18690 824 18696 876
rect 18748 864 18754 876
rect 19610 864 19616 876
rect 18748 836 19616 864
rect 18748 824 18754 836
rect 19610 824 19616 836
rect 19668 824 19674 876
rect 20162 824 20168 876
rect 20220 824 20226 876
rect 27154 824 27160 876
rect 27212 864 27218 876
rect 31202 864 31208 876
rect 27212 836 31208 864
rect 27212 824 27218 836
rect 31202 824 31208 836
rect 31260 824 31266 876
rect 13538 796 13544 808
rect 12406 768 13544 796
rect 13538 756 13544 768
rect 13596 756 13602 808
rect 15378 756 15384 808
rect 15436 796 15442 808
rect 16482 796 16488 808
rect 15436 768 16488 796
rect 15436 756 15442 768
rect 16482 756 16488 768
rect 16540 756 16546 808
rect 17770 756 17776 808
rect 17828 796 17834 808
rect 19702 796 19708 808
rect 17828 768 19708 796
rect 17828 756 17834 768
rect 19702 756 19708 768
rect 19760 756 19766 808
rect 8662 688 8668 740
rect 8720 688 8726 740
rect 8846 688 8852 740
rect 8904 728 8910 740
rect 9306 728 9312 740
rect 8904 700 9312 728
rect 8904 688 8910 700
rect 9306 688 9312 700
rect 9364 688 9370 740
rect 10318 688 10324 740
rect 10376 728 10382 740
rect 10962 728 10968 740
rect 10376 700 10968 728
rect 10376 688 10382 700
rect 10962 688 10968 700
rect 11020 688 11026 740
rect 11146 688 11152 740
rect 11204 728 11210 740
rect 11790 728 11796 740
rect 11204 700 11796 728
rect 11204 688 11210 700
rect 11790 688 11796 700
rect 11848 688 11854 740
rect 13170 688 13176 740
rect 13228 728 13234 740
rect 13722 728 13728 740
rect 13228 700 13728 728
rect 13228 688 13234 700
rect 13722 688 13728 700
rect 13780 688 13786 740
rect 15654 688 15660 740
rect 15712 728 15718 740
rect 17034 728 17040 740
rect 15712 700 17040 728
rect 15712 688 15718 700
rect 17034 688 17040 700
rect 17092 688 17098 740
rect 17678 688 17684 740
rect 17736 728 17742 740
rect 18598 728 18604 740
rect 17736 700 18604 728
rect 17736 688 17742 700
rect 18598 688 18604 700
rect 18656 688 18662 740
rect 20180 728 20208 824
rect 31726 796 31754 904
rect 31846 892 31852 944
rect 31904 892 31910 944
rect 33042 892 33048 944
rect 33100 932 33106 944
rect 35894 932 35900 944
rect 33100 904 35900 932
rect 33100 892 33106 904
rect 35894 892 35900 904
rect 35952 892 35958 944
rect 31864 864 31892 892
rect 38626 864 38654 972
rect 40126 960 40132 972
rect 40184 960 40190 1012
rect 31864 836 38654 864
rect 39114 796 39120 808
rect 31726 768 34744 796
rect 20180 700 26372 728
rect 8680 660 8708 688
rect 8680 632 14688 660
rect 8754 552 8760 604
rect 8812 592 8818 604
rect 13998 592 14004 604
rect 8812 564 14004 592
rect 8812 552 8818 564
rect 13998 552 14004 564
rect 14056 552 14062 604
rect 14660 592 14688 632
rect 14734 620 14740 672
rect 14792 660 14798 672
rect 15746 660 15752 672
rect 14792 632 15752 660
rect 14792 620 14798 632
rect 15746 620 15752 632
rect 15804 620 15810 672
rect 16390 620 16396 672
rect 16448 660 16454 672
rect 17770 660 17776 672
rect 16448 632 17776 660
rect 16448 620 16454 632
rect 17770 620 17776 632
rect 17828 620 17834 672
rect 17954 620 17960 672
rect 18012 660 18018 672
rect 18966 660 18972 672
rect 18012 632 18972 660
rect 18012 620 18018 632
rect 18966 620 18972 632
rect 19024 620 19030 672
rect 19518 620 19524 672
rect 19576 660 19582 672
rect 20990 660 20996 672
rect 19576 632 20996 660
rect 19576 620 19582 632
rect 20990 620 20996 632
rect 21048 620 21054 672
rect 25038 620 25044 672
rect 25096 660 25102 672
rect 26142 660 26148 672
rect 25096 632 26148 660
rect 25096 620 25102 632
rect 26142 620 26148 632
rect 26200 620 26206 672
rect 15010 592 15016 604
rect 14660 564 15016 592
rect 15010 552 15016 564
rect 15068 552 15074 604
rect 15194 552 15200 604
rect 15252 592 15258 604
rect 16298 592 16304 604
rect 15252 564 16304 592
rect 15252 552 15258 564
rect 16298 552 16304 564
rect 16356 552 16362 604
rect 18322 552 18328 604
rect 18380 592 18386 604
rect 21910 592 21916 604
rect 18380 564 21916 592
rect 18380 552 18386 564
rect 21910 552 21916 564
rect 21968 552 21974 604
rect 26344 592 26372 700
rect 26786 688 26792 740
rect 26844 728 26850 740
rect 26844 700 31754 728
rect 26844 688 26850 700
rect 27614 620 27620 672
rect 27672 660 27678 672
rect 30926 660 30932 672
rect 27672 632 30932 660
rect 27672 620 27678 632
rect 30926 620 30932 632
rect 30984 620 30990 672
rect 31726 660 31754 700
rect 32214 688 32220 740
rect 32272 688 32278 740
rect 34716 728 34744 768
rect 34992 768 39120 796
rect 34992 728 35020 768
rect 39114 756 39120 768
rect 39172 756 39178 808
rect 34716 700 35020 728
rect 36538 688 36544 740
rect 36596 728 36602 740
rect 40678 728 40684 740
rect 36596 700 40684 728
rect 36596 688 36602 700
rect 40678 688 40684 700
rect 40736 688 40742 740
rect 32122 660 32128 672
rect 31726 632 32128 660
rect 32122 620 32128 632
rect 32180 620 32186 672
rect 32232 592 32260 688
rect 35342 620 35348 672
rect 35400 660 35406 672
rect 37642 660 37648 672
rect 35400 632 37648 660
rect 35400 620 35406 632
rect 37642 620 37648 632
rect 37700 620 37706 672
rect 26344 564 32260 592
rect 34882 552 34888 604
rect 34940 592 34946 604
rect 36814 592 36820 604
rect 34940 564 36820 592
rect 34940 552 34946 564
rect 36814 552 36820 564
rect 36872 552 36878 604
rect 18874 524 18880 536
rect 12912 496 13124 524
rect 11330 456 11336 468
rect 6886 428 11336 456
rect 11330 416 11336 428
rect 11388 416 11394 468
rect 4908 320 4936 416
rect 6104 388 6132 416
rect 8938 388 8944 400
rect 6104 360 8944 388
rect 8938 348 8944 360
rect 8996 348 9002 400
rect 12912 320 12940 496
rect 12986 416 12992 468
rect 13044 416 13050 468
rect 13096 456 13124 496
rect 13832 496 18880 524
rect 13832 456 13860 496
rect 18874 484 18880 496
rect 18932 484 18938 536
rect 23566 484 23572 536
rect 23624 524 23630 536
rect 38654 524 38660 536
rect 23624 496 38660 524
rect 23624 484 23630 496
rect 38654 484 38660 496
rect 38712 484 38718 536
rect 39206 484 39212 536
rect 39264 524 39270 536
rect 41690 524 41696 536
rect 39264 496 41696 524
rect 39264 484 39270 496
rect 41690 484 41696 496
rect 41748 484 41754 536
rect 13096 428 13860 456
rect 13906 416 13912 468
rect 13964 456 13970 468
rect 15194 456 15200 468
rect 13964 428 15200 456
rect 13964 416 13970 428
rect 15194 416 15200 428
rect 15252 416 15258 468
rect 30742 456 30748 468
rect 26436 428 30748 456
rect 4908 292 12940 320
rect 7190 212 7196 264
rect 7248 212 7254 264
rect 13004 252 13032 416
rect 13998 348 14004 400
rect 14056 388 14062 400
rect 19426 388 19432 400
rect 14056 360 19432 388
rect 14056 348 14062 360
rect 19426 348 19432 360
rect 19484 348 19490 400
rect 20254 348 20260 400
rect 20312 388 20318 400
rect 26436 388 26464 428
rect 30742 416 30748 428
rect 30800 416 30806 468
rect 31662 416 31668 468
rect 31720 456 31726 468
rect 34790 456 34796 468
rect 31720 428 34796 456
rect 31720 416 31726 428
rect 34790 416 34796 428
rect 34848 416 34854 468
rect 20312 360 26464 388
rect 20312 348 20318 360
rect 27522 348 27528 400
rect 27580 388 27586 400
rect 30282 388 30288 400
rect 27580 360 30288 388
rect 27580 348 27586 360
rect 30282 348 30288 360
rect 30340 348 30346 400
rect 36906 388 36912 400
rect 31726 360 36912 388
rect 13630 280 13636 332
rect 13688 320 13694 332
rect 26878 320 26884 332
rect 13688 292 26884 320
rect 13688 280 13694 292
rect 26878 280 26884 292
rect 26936 280 26942 332
rect 31726 320 31754 360
rect 36906 348 36912 360
rect 36964 348 36970 400
rect 38838 348 38844 400
rect 38896 388 38902 400
rect 41414 388 41420 400
rect 38896 360 41420 388
rect 38896 348 38902 360
rect 41414 348 41420 360
rect 41472 348 41478 400
rect 28966 292 31754 320
rect 23014 252 23020 264
rect 13004 224 23020 252
rect 23014 212 23020 224
rect 23072 212 23078 264
rect 24394 212 24400 264
rect 24452 252 24458 264
rect 28966 252 28994 292
rect 37826 280 37832 332
rect 37884 280 37890 332
rect 24452 224 28994 252
rect 24452 212 24458 224
rect 29730 212 29736 264
rect 29788 252 29794 264
rect 32490 252 32496 264
rect 29788 224 32496 252
rect 29788 212 29794 224
rect 32490 212 32496 224
rect 32548 212 32554 264
rect 7208 184 7236 212
rect 20806 184 20812 196
rect 7208 156 20812 184
rect 20806 144 20812 156
rect 20864 144 20870 196
rect 21266 144 21272 196
rect 21324 144 21330 196
rect 24578 144 24584 196
rect 24636 184 24642 196
rect 37844 184 37872 280
rect 24636 156 37872 184
rect 24636 144 24642 156
rect 6086 76 6092 128
rect 6144 116 6150 128
rect 6362 116 6368 128
rect 6144 88 6368 116
rect 6144 76 6150 88
rect 6362 76 6368 88
rect 6420 76 6426 128
rect 10226 76 10232 128
rect 10284 116 10290 128
rect 18506 116 18512 128
rect 10284 88 18512 116
rect 10284 76 10290 88
rect 18506 76 18512 88
rect 18564 76 18570 128
rect 15010 8 15016 60
rect 15068 48 15074 60
rect 21284 48 21312 144
rect 21910 76 21916 128
rect 21968 116 21974 128
rect 26786 116 26792 128
rect 21968 88 26792 116
rect 21968 76 21974 88
rect 26786 76 26792 88
rect 26844 76 26850 128
rect 35710 76 35716 128
rect 35768 116 35774 128
rect 38102 116 38108 128
rect 35768 88 38108 116
rect 35768 76 35774 88
rect 38102 76 38108 88
rect 38160 76 38166 128
rect 15068 20 21312 48
rect 15068 8 15074 20
<< via1 >>
rect 7564 8780 7616 8832
rect 25320 8780 25372 8832
rect 11552 8678 11604 8730
rect 11616 8678 11668 8730
rect 11680 8678 11732 8730
rect 11744 8678 11796 8730
rect 11808 8678 11860 8730
rect 22155 8678 22207 8730
rect 22219 8678 22271 8730
rect 22283 8678 22335 8730
rect 22347 8678 22399 8730
rect 22411 8678 22463 8730
rect 32758 8678 32810 8730
rect 32822 8678 32874 8730
rect 32886 8678 32938 8730
rect 32950 8678 33002 8730
rect 33014 8678 33066 8730
rect 43361 8678 43413 8730
rect 43425 8678 43477 8730
rect 43489 8678 43541 8730
rect 43553 8678 43605 8730
rect 43617 8678 43669 8730
rect 1216 8576 1268 8628
rect 3240 8576 3292 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 7472 8576 7524 8628
rect 9588 8576 9640 8628
rect 11888 8576 11940 8628
rect 13820 8576 13872 8628
rect 15936 8576 15988 8628
rect 18144 8619 18196 8628
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 20168 8576 20220 8628
rect 22560 8619 22612 8628
rect 22560 8585 22569 8619
rect 22569 8585 22603 8619
rect 22603 8585 22612 8619
rect 22560 8576 22612 8585
rect 24400 8576 24452 8628
rect 26516 8576 26568 8628
rect 28632 8576 28684 8628
rect 30748 8576 30800 8628
rect 32680 8576 32732 8628
rect 34980 8576 35032 8628
rect 37096 8576 37148 8628
rect 39212 8576 39264 8628
rect 41328 8576 41380 8628
rect 43260 8576 43312 8628
rect 28172 8508 28224 8560
rect 2228 8347 2280 8356
rect 2228 8313 2237 8347
rect 2237 8313 2271 8347
rect 2271 8313 2280 8347
rect 2228 8304 2280 8313
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 14096 8440 14148 8492
rect 15292 8440 15344 8492
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 22744 8440 22796 8492
rect 24860 8440 24912 8492
rect 26976 8483 27028 8492
rect 26976 8449 26985 8483
rect 26985 8449 27019 8483
rect 27019 8449 27028 8483
rect 26976 8440 27028 8449
rect 28724 8483 28776 8492
rect 28724 8449 28733 8483
rect 28733 8449 28767 8483
rect 28767 8449 28776 8483
rect 28724 8440 28776 8449
rect 30840 8483 30892 8492
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 33232 8440 33284 8492
rect 35072 8483 35124 8492
rect 35072 8449 35081 8483
rect 35081 8449 35115 8483
rect 35115 8449 35124 8483
rect 35072 8440 35124 8449
rect 37372 8483 37424 8492
rect 37372 8449 37381 8483
rect 37381 8449 37415 8483
rect 37415 8449 37424 8483
rect 37372 8440 37424 8449
rect 39304 8483 39356 8492
rect 39304 8449 39313 8483
rect 39313 8449 39347 8483
rect 39347 8449 39356 8483
rect 39304 8440 39356 8449
rect 40500 8440 40552 8492
rect 42892 8483 42944 8492
rect 42892 8449 42901 8483
rect 42901 8449 42935 8483
rect 42935 8449 42944 8483
rect 42892 8440 42944 8449
rect 23204 8372 23256 8424
rect 14280 8304 14332 8356
rect 22560 8304 22612 8356
rect 6251 8134 6303 8186
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 16854 8134 16906 8186
rect 16918 8134 16970 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 27457 8134 27509 8186
rect 27521 8134 27573 8186
rect 27585 8134 27637 8186
rect 27649 8134 27701 8186
rect 27713 8134 27765 8186
rect 38060 8134 38112 8186
rect 38124 8134 38176 8186
rect 38188 8134 38240 8186
rect 38252 8134 38304 8186
rect 38316 8134 38368 8186
rect 11552 7590 11604 7642
rect 11616 7590 11668 7642
rect 11680 7590 11732 7642
rect 11744 7590 11796 7642
rect 11808 7590 11860 7642
rect 22155 7590 22207 7642
rect 22219 7590 22271 7642
rect 22283 7590 22335 7642
rect 22347 7590 22399 7642
rect 22411 7590 22463 7642
rect 32758 7590 32810 7642
rect 32822 7590 32874 7642
rect 32886 7590 32938 7642
rect 32950 7590 33002 7642
rect 33014 7590 33066 7642
rect 43361 7590 43413 7642
rect 43425 7590 43477 7642
rect 43489 7590 43541 7642
rect 43553 7590 43605 7642
rect 43617 7590 43669 7642
rect 6251 7046 6303 7098
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 16854 7046 16906 7098
rect 16918 7046 16970 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 27457 7046 27509 7098
rect 27521 7046 27573 7098
rect 27585 7046 27637 7098
rect 27649 7046 27701 7098
rect 27713 7046 27765 7098
rect 38060 7046 38112 7098
rect 38124 7046 38176 7098
rect 38188 7046 38240 7098
rect 38252 7046 38304 7098
rect 38316 7046 38368 7098
rect 11552 6502 11604 6554
rect 11616 6502 11668 6554
rect 11680 6502 11732 6554
rect 11744 6502 11796 6554
rect 11808 6502 11860 6554
rect 22155 6502 22207 6554
rect 22219 6502 22271 6554
rect 22283 6502 22335 6554
rect 22347 6502 22399 6554
rect 22411 6502 22463 6554
rect 32758 6502 32810 6554
rect 32822 6502 32874 6554
rect 32886 6502 32938 6554
rect 32950 6502 33002 6554
rect 33014 6502 33066 6554
rect 43361 6502 43413 6554
rect 43425 6502 43477 6554
rect 43489 6502 43541 6554
rect 43553 6502 43605 6554
rect 43617 6502 43669 6554
rect 6251 5958 6303 6010
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 16854 5958 16906 6010
rect 16918 5958 16970 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 27457 5958 27509 6010
rect 27521 5958 27573 6010
rect 27585 5958 27637 6010
rect 27649 5958 27701 6010
rect 27713 5958 27765 6010
rect 38060 5958 38112 6010
rect 38124 5958 38176 6010
rect 38188 5958 38240 6010
rect 38252 5958 38304 6010
rect 38316 5958 38368 6010
rect 11552 5414 11604 5466
rect 11616 5414 11668 5466
rect 11680 5414 11732 5466
rect 11744 5414 11796 5466
rect 11808 5414 11860 5466
rect 22155 5414 22207 5466
rect 22219 5414 22271 5466
rect 22283 5414 22335 5466
rect 22347 5414 22399 5466
rect 22411 5414 22463 5466
rect 32758 5414 32810 5466
rect 32822 5414 32874 5466
rect 32886 5414 32938 5466
rect 32950 5414 33002 5466
rect 33014 5414 33066 5466
rect 43361 5414 43413 5466
rect 43425 5414 43477 5466
rect 43489 5414 43541 5466
rect 43553 5414 43605 5466
rect 43617 5414 43669 5466
rect 6251 4870 6303 4922
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 16854 4870 16906 4922
rect 16918 4870 16970 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 27457 4870 27509 4922
rect 27521 4870 27573 4922
rect 27585 4870 27637 4922
rect 27649 4870 27701 4922
rect 27713 4870 27765 4922
rect 38060 4870 38112 4922
rect 38124 4870 38176 4922
rect 38188 4870 38240 4922
rect 38252 4870 38304 4922
rect 38316 4870 38368 4922
rect 8576 4496 8628 4548
rect 23388 4496 23440 4548
rect 9220 4428 9272 4480
rect 23664 4428 23716 4480
rect 11552 4326 11604 4378
rect 11616 4326 11668 4378
rect 11680 4326 11732 4378
rect 11744 4326 11796 4378
rect 11808 4326 11860 4378
rect 22155 4326 22207 4378
rect 22219 4326 22271 4378
rect 22283 4326 22335 4378
rect 22347 4326 22399 4378
rect 22411 4326 22463 4378
rect 32758 4326 32810 4378
rect 32822 4326 32874 4378
rect 32886 4326 32938 4378
rect 32950 4326 33002 4378
rect 33014 4326 33066 4378
rect 43361 4326 43413 4378
rect 43425 4326 43477 4378
rect 43489 4326 43541 4378
rect 43553 4326 43605 4378
rect 43617 4326 43669 4378
rect 11336 4224 11388 4276
rect 28080 4224 28132 4276
rect 7196 4156 7248 4208
rect 25136 4156 25188 4208
rect 11980 3884 12032 3936
rect 28356 3884 28408 3936
rect 6251 3782 6303 3834
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 16854 3782 16906 3834
rect 16918 3782 16970 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 27457 3782 27509 3834
rect 27521 3782 27573 3834
rect 27585 3782 27637 3834
rect 27649 3782 27701 3834
rect 27713 3782 27765 3834
rect 38060 3782 38112 3834
rect 38124 3782 38176 3834
rect 38188 3782 38240 3834
rect 38252 3782 38304 3834
rect 38316 3782 38368 3834
rect 17960 3544 18012 3596
rect 36820 3544 36872 3596
rect 38936 3544 38988 3596
rect 13636 3476 13688 3528
rect 25596 3476 25648 3528
rect 26148 3476 26200 3528
rect 38476 3476 38528 3528
rect 40868 3476 40920 3528
rect 16212 3408 16264 3460
rect 30196 3408 30248 3460
rect 37832 3408 37884 3460
rect 40316 3408 40368 3460
rect 8300 3340 8352 3392
rect 20444 3340 20496 3392
rect 37188 3340 37240 3392
rect 39488 3340 39540 3392
rect 11552 3238 11604 3290
rect 11616 3238 11668 3290
rect 11680 3238 11732 3290
rect 11744 3238 11796 3290
rect 11808 3238 11860 3290
rect 22155 3238 22207 3290
rect 22219 3238 22271 3290
rect 22283 3238 22335 3290
rect 22347 3238 22399 3290
rect 22411 3238 22463 3290
rect 32758 3238 32810 3290
rect 32822 3238 32874 3290
rect 32886 3238 32938 3290
rect 32950 3238 33002 3290
rect 33014 3238 33066 3290
rect 43361 3238 43413 3290
rect 43425 3238 43477 3290
rect 43489 3238 43541 3290
rect 43553 3238 43605 3290
rect 43617 3238 43669 3290
rect 18972 3136 19024 3188
rect 23572 3136 23624 3188
rect 17684 3068 17736 3120
rect 25688 3068 25740 3120
rect 28724 3136 28776 3188
rect 37556 3136 37608 3188
rect 40040 3136 40092 3188
rect 30104 3068 30156 3120
rect 38016 3068 38068 3120
rect 40592 3068 40644 3120
rect 10968 3000 11020 3052
rect 7840 2932 7892 2984
rect 25596 3043 25648 3052
rect 25596 3009 25605 3043
rect 25605 3009 25639 3043
rect 25639 3009 25648 3043
rect 25596 3000 25648 3009
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 27804 3043 27856 3052
rect 27804 3009 27813 3043
rect 27813 3009 27847 3043
rect 27847 3009 27856 3043
rect 27804 3000 27856 3009
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 15752 2864 15804 2916
rect 17500 2864 17552 2916
rect 18144 2864 18196 2916
rect 15476 2796 15528 2848
rect 19064 2796 19116 2848
rect 20352 2864 20404 2916
rect 26516 2932 26568 2984
rect 29460 2864 29512 2916
rect 38568 3000 38620 3052
rect 41144 3000 41196 3052
rect 38384 2932 38436 2984
rect 37188 2864 37240 2916
rect 39212 2864 39264 2916
rect 21180 2796 21232 2848
rect 21732 2796 21784 2848
rect 23480 2796 23532 2848
rect 26240 2796 26292 2848
rect 27344 2839 27396 2848
rect 27344 2805 27353 2839
rect 27353 2805 27387 2839
rect 27387 2805 27396 2839
rect 27344 2796 27396 2805
rect 27804 2796 27856 2848
rect 28724 2796 28776 2848
rect 30748 2796 30800 2848
rect 36360 2796 36412 2848
rect 38660 2796 38712 2848
rect 6251 2694 6303 2746
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 16854 2694 16906 2746
rect 16918 2694 16970 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 27457 2694 27509 2746
rect 27521 2694 27573 2746
rect 27585 2694 27637 2746
rect 27649 2694 27701 2746
rect 27713 2694 27765 2746
rect 38060 2694 38112 2746
rect 38124 2694 38176 2746
rect 38188 2694 38240 2746
rect 38252 2694 38304 2746
rect 38316 2694 38368 2746
rect 15292 2635 15344 2644
rect 15292 2601 15301 2635
rect 15301 2601 15335 2635
rect 15335 2601 15344 2635
rect 15292 2592 15344 2601
rect 11060 2524 11112 2576
rect 15752 2592 15804 2644
rect 16028 2592 16080 2644
rect 17868 2592 17920 2644
rect 18052 2592 18104 2644
rect 22560 2592 22612 2644
rect 22744 2635 22796 2644
rect 22744 2601 22753 2635
rect 22753 2601 22787 2635
rect 22787 2601 22796 2635
rect 22744 2592 22796 2601
rect 15568 2567 15620 2576
rect 15568 2533 15577 2567
rect 15577 2533 15611 2567
rect 15611 2533 15620 2567
rect 15568 2524 15620 2533
rect 13728 2456 13780 2508
rect 15292 2456 15344 2508
rect 15568 2388 15620 2440
rect 16488 2456 16540 2508
rect 16856 2524 16908 2576
rect 17960 2524 18012 2576
rect 16764 2388 16816 2440
rect 17224 2456 17276 2508
rect 18052 2456 18104 2508
rect 20076 2524 20128 2576
rect 20260 2524 20312 2576
rect 25596 2592 25648 2644
rect 27160 2592 27212 2644
rect 27896 2592 27948 2644
rect 28172 2635 28224 2644
rect 28172 2601 28181 2635
rect 28181 2601 28215 2635
rect 28215 2601 28224 2635
rect 28172 2592 28224 2601
rect 30196 2635 30248 2644
rect 30196 2601 30205 2635
rect 30205 2601 30239 2635
rect 30239 2601 30248 2635
rect 30196 2592 30248 2601
rect 30840 2592 30892 2644
rect 33232 2635 33284 2644
rect 33232 2601 33241 2635
rect 33241 2601 33275 2635
rect 33275 2601 33284 2635
rect 33232 2592 33284 2601
rect 35072 2592 35124 2644
rect 37372 2592 37424 2644
rect 39304 2592 39356 2644
rect 40500 2635 40552 2644
rect 40500 2601 40509 2635
rect 40509 2601 40543 2635
rect 40543 2601 40552 2635
rect 40500 2592 40552 2601
rect 42892 2592 42944 2644
rect 15200 2320 15252 2372
rect 17316 2388 17368 2440
rect 18420 2388 18472 2440
rect 14832 2252 14884 2304
rect 16304 2252 16356 2304
rect 16764 2252 16816 2304
rect 16856 2252 16908 2304
rect 17224 2252 17276 2304
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19984 2388 20036 2440
rect 20168 2388 20220 2440
rect 19708 2320 19760 2372
rect 20260 2320 20312 2372
rect 23204 2567 23256 2576
rect 23204 2533 23213 2567
rect 23213 2533 23247 2567
rect 23247 2533 23256 2567
rect 23204 2524 23256 2533
rect 25872 2524 25924 2576
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 19892 2295 19944 2304
rect 19892 2261 19901 2295
rect 19901 2261 19935 2295
rect 19935 2261 19944 2295
rect 19892 2252 19944 2261
rect 21272 2388 21324 2440
rect 21824 2388 21876 2440
rect 22284 2388 22336 2440
rect 23756 2456 23808 2508
rect 24584 2388 24636 2440
rect 21456 2252 21508 2304
rect 21548 2295 21600 2304
rect 21548 2261 21557 2295
rect 21557 2261 21591 2295
rect 21591 2261 21600 2295
rect 21548 2252 21600 2261
rect 21916 2295 21968 2304
rect 21916 2261 21925 2295
rect 21925 2261 21959 2295
rect 21959 2261 21968 2295
rect 21916 2252 21968 2261
rect 22928 2252 22980 2304
rect 24032 2320 24084 2372
rect 25596 2431 25648 2440
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 24860 2295 24912 2304
rect 24860 2261 24869 2295
rect 24869 2261 24903 2295
rect 24903 2261 24912 2295
rect 24860 2252 24912 2261
rect 25136 2252 25188 2304
rect 25596 2252 25648 2304
rect 26148 2431 26200 2440
rect 26148 2397 26157 2431
rect 26157 2397 26191 2431
rect 26191 2397 26200 2431
rect 26148 2388 26200 2397
rect 26700 2524 26752 2576
rect 26884 2524 26936 2576
rect 36452 2524 36504 2576
rect 26516 2456 26568 2508
rect 26608 2388 26660 2440
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 27068 2388 27120 2440
rect 27528 2431 27580 2440
rect 27528 2397 27537 2431
rect 27537 2397 27571 2431
rect 27571 2397 27580 2431
rect 27528 2388 27580 2397
rect 27620 2431 27672 2440
rect 27620 2397 27629 2431
rect 27629 2397 27663 2431
rect 27663 2397 27672 2431
rect 27620 2388 27672 2397
rect 28540 2431 28592 2440
rect 28540 2397 28549 2431
rect 28549 2397 28583 2431
rect 28583 2397 28592 2431
rect 28540 2388 28592 2397
rect 28632 2388 28684 2440
rect 29368 2431 29420 2440
rect 29368 2397 29377 2431
rect 29377 2397 29411 2431
rect 29411 2397 29420 2431
rect 29368 2388 29420 2397
rect 27160 2320 27212 2372
rect 31024 2388 31076 2440
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 31392 2431 31444 2440
rect 31392 2397 31401 2431
rect 31401 2397 31435 2431
rect 31435 2397 31444 2431
rect 31392 2388 31444 2397
rect 33140 2388 33192 2440
rect 33324 2388 33376 2440
rect 34704 2388 34756 2440
rect 35992 2431 36044 2440
rect 35992 2397 36001 2431
rect 36001 2397 36035 2431
rect 36035 2397 36044 2431
rect 35992 2388 36044 2397
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 39396 2431 39448 2440
rect 39396 2397 39405 2431
rect 39405 2397 39439 2431
rect 39439 2397 39448 2431
rect 39396 2388 39448 2397
rect 40684 2431 40736 2440
rect 40684 2397 40693 2431
rect 40693 2397 40727 2431
rect 40727 2397 40736 2431
rect 40684 2388 40736 2397
rect 42616 2431 42668 2440
rect 42616 2397 42625 2431
rect 42625 2397 42659 2431
rect 42659 2397 42668 2431
rect 42616 2388 42668 2397
rect 26516 2295 26568 2304
rect 26516 2261 26525 2295
rect 26525 2261 26559 2295
rect 26559 2261 26568 2295
rect 26516 2252 26568 2261
rect 26792 2295 26844 2304
rect 26792 2261 26801 2295
rect 26801 2261 26835 2295
rect 26835 2261 26844 2295
rect 26792 2252 26844 2261
rect 27896 2252 27948 2304
rect 28356 2295 28408 2304
rect 28356 2261 28365 2295
rect 28365 2261 28399 2295
rect 28399 2261 28408 2295
rect 28356 2252 28408 2261
rect 28816 2252 28868 2304
rect 28908 2295 28960 2304
rect 28908 2261 28917 2295
rect 28917 2261 28951 2295
rect 28951 2261 28960 2295
rect 28908 2252 28960 2261
rect 29184 2295 29236 2304
rect 29184 2261 29193 2295
rect 29193 2261 29227 2295
rect 29227 2261 29236 2295
rect 29184 2252 29236 2261
rect 35440 2320 35492 2372
rect 29644 2252 29696 2304
rect 30656 2252 30708 2304
rect 33508 2252 33560 2304
rect 11552 2150 11604 2202
rect 11616 2150 11668 2202
rect 11680 2150 11732 2202
rect 11744 2150 11796 2202
rect 11808 2150 11860 2202
rect 22155 2150 22207 2202
rect 22219 2150 22271 2202
rect 22283 2150 22335 2202
rect 22347 2150 22399 2202
rect 22411 2150 22463 2202
rect 32758 2150 32810 2202
rect 32822 2150 32874 2202
rect 32886 2150 32938 2202
rect 32950 2150 33002 2202
rect 33014 2150 33066 2202
rect 43361 2150 43413 2202
rect 43425 2150 43477 2202
rect 43489 2150 43541 2202
rect 43553 2150 43605 2202
rect 43617 2150 43669 2202
rect 10968 2048 11020 2100
rect 14280 2091 14332 2100
rect 14280 2057 14289 2091
rect 14289 2057 14323 2091
rect 14323 2057 14332 2091
rect 14280 2048 14332 2057
rect 15292 2048 15344 2100
rect 15476 2048 15528 2100
rect 9128 1955 9180 1964
rect 9128 1921 9137 1955
rect 9137 1921 9171 1955
rect 9171 1921 9180 1955
rect 9128 1912 9180 1921
rect 14096 1955 14148 1964
rect 14096 1921 14105 1955
rect 14105 1921 14139 1955
rect 14139 1921 14148 1955
rect 14096 1912 14148 1921
rect 15108 1980 15160 2032
rect 15660 2091 15712 2100
rect 15660 2057 15669 2091
rect 15669 2057 15703 2091
rect 15703 2057 15712 2091
rect 15660 2048 15712 2057
rect 16212 2048 16264 2100
rect 16856 2048 16908 2100
rect 17040 2048 17092 2100
rect 17132 2048 17184 2100
rect 18420 2048 18472 2100
rect 20996 2048 21048 2100
rect 14648 1955 14700 1964
rect 14648 1921 14657 1955
rect 14657 1921 14691 1955
rect 14691 1921 14700 1955
rect 14648 1912 14700 1921
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 14924 1912 14976 1921
rect 15292 1912 15344 1964
rect 15844 1912 15896 1964
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 16396 1912 16448 1964
rect 17224 1980 17276 2032
rect 15200 1776 15252 1828
rect 14464 1708 14516 1760
rect 16580 1844 16632 1896
rect 15384 1819 15436 1828
rect 15384 1785 15393 1819
rect 15393 1785 15427 1819
rect 15427 1785 15436 1819
rect 15384 1776 15436 1785
rect 16672 1776 16724 1828
rect 16488 1751 16540 1760
rect 16488 1717 16497 1751
rect 16497 1717 16531 1751
rect 16531 1717 16540 1751
rect 16488 1708 16540 1717
rect 16856 1708 16908 1760
rect 18052 1912 18104 1964
rect 18144 1979 18196 1988
rect 18144 1945 18153 1979
rect 18153 1945 18187 1979
rect 18187 1945 18196 1979
rect 18144 1936 18196 1945
rect 17684 1844 17736 1896
rect 18696 1955 18748 1964
rect 18696 1921 18705 1955
rect 18705 1921 18739 1955
rect 18739 1921 18748 1955
rect 18696 1912 18748 1921
rect 18788 1912 18840 1964
rect 19064 1912 19116 1964
rect 19432 1912 19484 1964
rect 18696 1776 18748 1828
rect 19524 1776 19576 1828
rect 17684 1751 17736 1760
rect 17684 1717 17693 1751
rect 17693 1717 17727 1751
rect 17727 1717 17736 1751
rect 17684 1708 17736 1717
rect 17868 1708 17920 1760
rect 17960 1751 18012 1760
rect 17960 1717 17969 1751
rect 17969 1717 18003 1751
rect 18003 1717 18012 1751
rect 17960 1708 18012 1717
rect 18972 1708 19024 1760
rect 19248 1708 19300 1760
rect 19340 1751 19392 1760
rect 19340 1717 19349 1751
rect 19349 1717 19383 1751
rect 19383 1717 19392 1751
rect 19340 1708 19392 1717
rect 20720 1980 20772 2032
rect 21732 1980 21784 2032
rect 23756 2091 23808 2100
rect 23756 2057 23765 2091
rect 23765 2057 23799 2091
rect 23799 2057 23808 2091
rect 23756 2048 23808 2057
rect 24032 2091 24084 2100
rect 24032 2057 24041 2091
rect 24041 2057 24075 2091
rect 24075 2057 24084 2091
rect 24032 2048 24084 2057
rect 19892 1912 19944 1964
rect 20628 1912 20680 1964
rect 20812 1912 20864 1964
rect 23388 1955 23440 1964
rect 23388 1921 23397 1955
rect 23397 1921 23431 1955
rect 23431 1921 23440 1955
rect 23388 1912 23440 1921
rect 23664 1955 23716 1964
rect 23664 1921 23673 1955
rect 23673 1921 23707 1955
rect 23707 1921 23716 1955
rect 23664 1912 23716 1921
rect 23848 1912 23900 1964
rect 24124 1912 24176 1964
rect 25872 2048 25924 2100
rect 26792 2048 26844 2100
rect 26976 2048 27028 2100
rect 28356 2048 28408 2100
rect 28908 2048 28960 2100
rect 29184 2048 29236 2100
rect 26240 1980 26292 2032
rect 29736 1980 29788 2032
rect 30196 1980 30248 2032
rect 30748 2091 30800 2100
rect 30748 2057 30757 2091
rect 30757 2057 30791 2091
rect 30791 2057 30800 2091
rect 30748 2048 30800 2057
rect 31300 2048 31352 2100
rect 32588 2048 32640 2100
rect 24952 1955 25004 1964
rect 24952 1921 24961 1955
rect 24961 1921 24995 1955
rect 24995 1921 25004 1955
rect 24952 1912 25004 1921
rect 25228 1955 25280 1964
rect 25228 1921 25237 1955
rect 25237 1921 25271 1955
rect 25271 1921 25280 1955
rect 25228 1912 25280 1921
rect 25504 1955 25556 1964
rect 25504 1921 25513 1955
rect 25513 1921 25547 1955
rect 25547 1921 25556 1955
rect 25504 1912 25556 1921
rect 25872 1912 25924 1964
rect 28172 1912 28224 1964
rect 20444 1776 20496 1828
rect 29276 1844 29328 1896
rect 24860 1776 24912 1828
rect 26240 1776 26292 1828
rect 27804 1776 27856 1828
rect 29460 1912 29512 1964
rect 32312 1980 32364 2032
rect 31208 1955 31260 1964
rect 31208 1921 31217 1955
rect 31217 1921 31251 1955
rect 31251 1921 31260 1955
rect 31208 1912 31260 1921
rect 31944 1955 31996 1964
rect 31944 1921 31953 1955
rect 31953 1921 31987 1955
rect 31987 1921 31996 1955
rect 31944 1912 31996 1921
rect 31484 1844 31536 1896
rect 33324 1955 33376 1964
rect 33324 1921 33333 1955
rect 33333 1921 33367 1955
rect 33367 1921 33376 1955
rect 33324 1912 33376 1921
rect 33876 1955 33928 1964
rect 33876 1921 33885 1955
rect 33885 1921 33919 1955
rect 33919 1921 33928 1955
rect 33876 1912 33928 1921
rect 34704 2048 34756 2100
rect 35440 2091 35492 2100
rect 35440 2057 35449 2091
rect 35449 2057 35483 2091
rect 35483 2057 35492 2091
rect 35440 2048 35492 2057
rect 35992 2048 36044 2100
rect 37740 2048 37792 2100
rect 39396 2048 39448 2100
rect 40684 2048 40736 2100
rect 42616 2048 42668 2100
rect 21364 1751 21416 1760
rect 21364 1717 21373 1751
rect 21373 1717 21407 1751
rect 21407 1717 21416 1751
rect 21364 1708 21416 1717
rect 21824 1751 21876 1760
rect 21824 1717 21833 1751
rect 21833 1717 21867 1751
rect 21867 1717 21876 1751
rect 21824 1708 21876 1717
rect 22008 1708 22060 1760
rect 22836 1751 22888 1760
rect 22836 1717 22845 1751
rect 22845 1717 22879 1751
rect 22879 1717 22888 1751
rect 22836 1708 22888 1717
rect 24216 1708 24268 1760
rect 24768 1751 24820 1760
rect 24768 1717 24777 1751
rect 24777 1717 24811 1751
rect 24811 1717 24820 1751
rect 24768 1708 24820 1717
rect 25044 1751 25096 1760
rect 25044 1717 25053 1751
rect 25053 1717 25087 1751
rect 25087 1717 25096 1751
rect 25044 1708 25096 1717
rect 25596 1708 25648 1760
rect 26148 1708 26200 1760
rect 27344 1708 27396 1760
rect 31668 1776 31720 1828
rect 28632 1708 28684 1760
rect 29644 1751 29696 1760
rect 29644 1717 29653 1751
rect 29653 1717 29687 1751
rect 29687 1717 29696 1751
rect 29644 1708 29696 1717
rect 30472 1708 30524 1760
rect 31576 1708 31628 1760
rect 32496 1708 32548 1760
rect 34244 1844 34296 1896
rect 36544 1912 36596 1964
rect 35808 1844 35860 1896
rect 37648 1955 37700 1964
rect 37648 1921 37657 1955
rect 37657 1921 37691 1955
rect 37691 1921 37700 1955
rect 37648 1912 37700 1921
rect 40960 1980 41012 2032
rect 40132 1912 40184 1964
rect 41788 1912 41840 1964
rect 41236 1844 41288 1896
rect 33600 1776 33652 1828
rect 35164 1776 35216 1828
rect 6251 1606 6303 1658
rect 6315 1606 6367 1658
rect 6379 1606 6431 1658
rect 6443 1606 6495 1658
rect 6507 1606 6559 1658
rect 16854 1606 16906 1658
rect 16918 1606 16970 1658
rect 16982 1606 17034 1658
rect 17046 1606 17098 1658
rect 17110 1606 17162 1658
rect 27457 1606 27509 1658
rect 27521 1606 27573 1658
rect 27585 1606 27637 1658
rect 27649 1606 27701 1658
rect 27713 1606 27765 1658
rect 38060 1606 38112 1658
rect 38124 1606 38176 1658
rect 38188 1606 38240 1658
rect 38252 1606 38304 1658
rect 38316 1606 38368 1658
rect 7196 1504 7248 1556
rect 5816 1436 5868 1488
rect 8576 1436 8628 1488
rect 11060 1547 11112 1556
rect 11060 1513 11069 1547
rect 11069 1513 11103 1547
rect 11103 1513 11112 1547
rect 11060 1504 11112 1513
rect 11336 1547 11388 1556
rect 11336 1513 11345 1547
rect 11345 1513 11379 1547
rect 11379 1513 11388 1547
rect 11336 1504 11388 1513
rect 12808 1547 12860 1556
rect 12808 1513 12817 1547
rect 12817 1513 12851 1547
rect 12851 1513 12860 1547
rect 12808 1504 12860 1513
rect 14464 1504 14516 1556
rect 13728 1436 13780 1488
rect 4988 1232 5040 1284
rect 5264 1232 5316 1284
rect 5908 1368 5960 1420
rect 5540 1232 5592 1284
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 6736 1300 6788 1352
rect 6276 1232 6328 1284
rect 7380 1300 7432 1352
rect 7656 1300 7708 1352
rect 7932 1300 7984 1352
rect 4804 1207 4856 1216
rect 4804 1173 4813 1207
rect 4813 1173 4847 1207
rect 4847 1173 4856 1207
rect 4804 1164 4856 1173
rect 4896 1164 4948 1216
rect 6092 1164 6144 1216
rect 7288 1232 7340 1284
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 7196 1164 7248 1216
rect 7840 1232 7892 1284
rect 8484 1300 8536 1352
rect 8852 1300 8904 1352
rect 9680 1368 9732 1420
rect 8392 1232 8444 1284
rect 9864 1300 9916 1352
rect 9588 1232 9640 1284
rect 10324 1343 10376 1352
rect 10324 1309 10333 1343
rect 10333 1309 10367 1343
rect 10367 1309 10376 1343
rect 10324 1300 10376 1309
rect 10508 1300 10560 1352
rect 10416 1232 10468 1284
rect 10968 1232 11020 1284
rect 11428 1300 11480 1352
rect 11888 1232 11940 1284
rect 12440 1368 12492 1420
rect 15292 1504 15344 1556
rect 16396 1504 16448 1556
rect 17408 1504 17460 1556
rect 17868 1504 17920 1556
rect 18512 1504 18564 1556
rect 22652 1504 22704 1556
rect 23388 1504 23440 1556
rect 24308 1504 24360 1556
rect 14832 1436 14884 1488
rect 12532 1300 12584 1352
rect 12624 1343 12676 1352
rect 12624 1309 12633 1343
rect 12633 1309 12667 1343
rect 12667 1309 12676 1343
rect 12624 1300 12676 1309
rect 13176 1343 13228 1352
rect 13176 1309 13185 1343
rect 13185 1309 13219 1343
rect 13219 1309 13228 1343
rect 13176 1300 13228 1309
rect 13360 1300 13412 1352
rect 13728 1300 13780 1352
rect 13912 1343 13964 1352
rect 13912 1309 13921 1343
rect 13921 1309 13955 1343
rect 13955 1309 13964 1343
rect 13912 1300 13964 1309
rect 13268 1232 13320 1284
rect 7656 1207 7708 1216
rect 7656 1173 7665 1207
rect 7665 1173 7699 1207
rect 7699 1173 7708 1207
rect 7656 1164 7708 1173
rect 8116 1164 8168 1216
rect 8300 1164 8352 1216
rect 8668 1164 8720 1216
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9312 1164 9364 1216
rect 9404 1207 9456 1216
rect 9404 1173 9413 1207
rect 9413 1173 9447 1207
rect 9447 1173 9456 1207
rect 9404 1164 9456 1173
rect 10140 1164 10192 1216
rect 10232 1207 10284 1216
rect 10232 1173 10241 1207
rect 10241 1173 10275 1207
rect 10275 1173 10284 1207
rect 10232 1164 10284 1173
rect 10692 1164 10744 1216
rect 10784 1207 10836 1216
rect 10784 1173 10793 1207
rect 10793 1173 10827 1207
rect 10827 1173 10836 1207
rect 10784 1164 10836 1173
rect 11152 1164 11204 1216
rect 11244 1164 11296 1216
rect 11980 1207 12032 1216
rect 11980 1173 11989 1207
rect 11989 1173 12023 1207
rect 12023 1173 12032 1207
rect 11980 1164 12032 1173
rect 12256 1207 12308 1216
rect 12256 1173 12265 1207
rect 12265 1173 12299 1207
rect 12299 1173 12308 1207
rect 12256 1164 12308 1173
rect 12348 1164 12400 1216
rect 12900 1164 12952 1216
rect 12992 1164 13044 1216
rect 13636 1207 13688 1216
rect 13636 1173 13645 1207
rect 13645 1173 13679 1207
rect 13679 1173 13688 1207
rect 13636 1164 13688 1173
rect 14740 1300 14792 1352
rect 15660 1436 15712 1488
rect 17132 1436 17184 1488
rect 15568 1368 15620 1420
rect 16764 1368 16816 1420
rect 17776 1436 17828 1488
rect 18052 1436 18104 1488
rect 18604 1436 18656 1488
rect 18696 1436 18748 1488
rect 15200 1300 15252 1352
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 15660 1343 15712 1352
rect 15660 1309 15669 1343
rect 15669 1309 15703 1343
rect 15703 1309 15712 1343
rect 15660 1300 15712 1309
rect 15936 1343 15988 1352
rect 15936 1309 15945 1343
rect 15945 1309 15979 1343
rect 15979 1309 15988 1343
rect 15936 1300 15988 1309
rect 16396 1300 16448 1352
rect 16488 1343 16540 1352
rect 16488 1309 16497 1343
rect 16497 1309 16531 1343
rect 16531 1309 16540 1343
rect 16488 1300 16540 1309
rect 14372 1207 14424 1216
rect 14372 1173 14381 1207
rect 14381 1173 14415 1207
rect 14415 1173 14424 1207
rect 14372 1164 14424 1173
rect 15016 1164 15068 1216
rect 15752 1207 15804 1216
rect 15752 1173 15761 1207
rect 15761 1173 15795 1207
rect 15795 1173 15804 1207
rect 15752 1164 15804 1173
rect 17408 1343 17460 1352
rect 17408 1309 17417 1343
rect 17417 1309 17451 1343
rect 17451 1309 17460 1343
rect 17408 1300 17460 1309
rect 17684 1343 17736 1352
rect 17684 1309 17693 1343
rect 17693 1309 17727 1343
rect 17727 1309 17736 1343
rect 17684 1300 17736 1309
rect 17960 1343 18012 1352
rect 17960 1309 17969 1343
rect 17969 1309 18003 1343
rect 18003 1309 18012 1343
rect 17960 1300 18012 1309
rect 18880 1368 18932 1420
rect 18972 1300 19024 1352
rect 20168 1436 20220 1488
rect 19524 1300 19576 1352
rect 20904 1479 20956 1488
rect 20904 1445 20913 1479
rect 20913 1445 20947 1479
rect 20947 1445 20956 1479
rect 20904 1436 20956 1445
rect 24676 1436 24728 1488
rect 26148 1504 26200 1556
rect 20444 1411 20496 1420
rect 20444 1377 20453 1411
rect 20453 1377 20487 1411
rect 20487 1377 20496 1411
rect 20444 1368 20496 1377
rect 22560 1368 22612 1420
rect 25504 1368 25556 1420
rect 27620 1436 27672 1488
rect 29460 1504 29512 1556
rect 30840 1504 30892 1556
rect 29092 1436 29144 1488
rect 29552 1436 29604 1488
rect 29644 1436 29696 1488
rect 31024 1436 31076 1488
rect 27712 1368 27764 1420
rect 30472 1368 30524 1420
rect 32956 1504 33008 1556
rect 34980 1504 35032 1556
rect 35900 1504 35952 1556
rect 36452 1504 36504 1556
rect 37648 1504 37700 1556
rect 32496 1479 32548 1488
rect 32496 1445 32505 1479
rect 32505 1445 32539 1479
rect 32539 1445 32548 1479
rect 32496 1436 32548 1445
rect 33140 1436 33192 1488
rect 35716 1436 35768 1488
rect 38384 1504 38436 1556
rect 40132 1504 40184 1556
rect 41788 1547 41840 1556
rect 41788 1513 41797 1547
rect 41797 1513 41831 1547
rect 41831 1513 41840 1547
rect 41788 1504 41840 1513
rect 40960 1479 41012 1488
rect 40960 1445 40969 1479
rect 40969 1445 41003 1479
rect 41003 1445 41012 1479
rect 40960 1436 41012 1445
rect 41236 1479 41288 1488
rect 41236 1445 41245 1479
rect 41245 1445 41279 1479
rect 41279 1445 41288 1479
rect 41236 1436 41288 1445
rect 21548 1300 21600 1352
rect 17776 1207 17828 1216
rect 17776 1173 17785 1207
rect 17785 1173 17819 1207
rect 17819 1173 17828 1207
rect 17776 1164 17828 1173
rect 18236 1207 18288 1216
rect 18236 1173 18245 1207
rect 18245 1173 18279 1207
rect 18279 1173 18288 1207
rect 18236 1164 18288 1173
rect 18696 1164 18748 1216
rect 18788 1207 18840 1216
rect 18788 1173 18797 1207
rect 18797 1173 18831 1207
rect 18831 1173 18840 1207
rect 18788 1164 18840 1173
rect 20536 1232 20588 1284
rect 21916 1232 21968 1284
rect 22928 1300 22980 1352
rect 23480 1300 23532 1352
rect 24768 1300 24820 1352
rect 25688 1300 25740 1352
rect 19800 1164 19852 1216
rect 19892 1207 19944 1216
rect 19892 1173 19901 1207
rect 19901 1173 19935 1207
rect 19935 1173 19944 1207
rect 19892 1164 19944 1173
rect 21548 1207 21600 1216
rect 21548 1173 21557 1207
rect 21557 1173 21591 1207
rect 21591 1173 21600 1207
rect 21548 1164 21600 1173
rect 21824 1164 21876 1216
rect 24860 1275 24912 1284
rect 24860 1241 24869 1275
rect 24869 1241 24903 1275
rect 24903 1241 24912 1275
rect 24860 1232 24912 1241
rect 25044 1232 25096 1284
rect 26240 1300 26292 1352
rect 26516 1300 26568 1352
rect 27344 1300 27396 1352
rect 27896 1300 27948 1352
rect 28816 1300 28868 1352
rect 29000 1300 29052 1352
rect 30104 1300 30156 1352
rect 31944 1343 31996 1352
rect 31944 1309 31953 1343
rect 31953 1309 31987 1343
rect 31987 1309 31996 1343
rect 31944 1300 31996 1309
rect 33968 1300 34020 1352
rect 30748 1275 30800 1284
rect 30748 1241 30757 1275
rect 30757 1241 30791 1275
rect 30791 1241 30800 1275
rect 30748 1232 30800 1241
rect 30932 1232 30984 1284
rect 32220 1275 32272 1284
rect 32220 1241 32229 1275
rect 32229 1241 32263 1275
rect 32263 1241 32272 1275
rect 32220 1232 32272 1241
rect 32312 1232 32364 1284
rect 22928 1207 22980 1216
rect 22928 1173 22937 1207
rect 22937 1173 22971 1207
rect 22971 1173 22980 1207
rect 22928 1164 22980 1173
rect 23296 1207 23348 1216
rect 23296 1173 23305 1207
rect 23305 1173 23339 1207
rect 23339 1173 23348 1207
rect 23296 1164 23348 1173
rect 23664 1164 23716 1216
rect 24768 1164 24820 1216
rect 26148 1164 26200 1216
rect 26884 1164 26936 1216
rect 30288 1207 30340 1216
rect 30288 1173 30297 1207
rect 30297 1173 30331 1207
rect 30331 1173 30340 1207
rect 30288 1164 30340 1173
rect 32128 1164 32180 1216
rect 34428 1232 34480 1284
rect 35164 1300 35216 1352
rect 36820 1300 36872 1352
rect 34520 1164 34572 1216
rect 36268 1275 36320 1284
rect 36268 1241 36277 1275
rect 36277 1241 36311 1275
rect 36311 1241 36320 1275
rect 36268 1232 36320 1241
rect 37464 1300 37516 1352
rect 37648 1300 37700 1352
rect 38108 1343 38160 1352
rect 38108 1309 38117 1343
rect 38117 1309 38151 1343
rect 38151 1309 38160 1343
rect 38108 1300 38160 1309
rect 38384 1343 38436 1352
rect 38384 1309 38393 1343
rect 38393 1309 38427 1343
rect 38427 1309 38436 1343
rect 38384 1300 38436 1309
rect 39580 1368 39632 1420
rect 38660 1343 38712 1352
rect 38660 1309 38669 1343
rect 38669 1309 38703 1343
rect 38703 1309 38712 1343
rect 38660 1300 38712 1309
rect 38936 1343 38988 1352
rect 38936 1309 38945 1343
rect 38945 1309 38979 1343
rect 38979 1309 38988 1343
rect 38936 1300 38988 1309
rect 39212 1343 39264 1352
rect 39212 1309 39221 1343
rect 39221 1309 39255 1343
rect 39255 1309 39264 1343
rect 39212 1300 39264 1309
rect 39488 1343 39540 1352
rect 39488 1309 39497 1343
rect 39497 1309 39531 1343
rect 39531 1309 39540 1343
rect 39488 1300 39540 1309
rect 40040 1343 40092 1352
rect 40040 1309 40049 1343
rect 40049 1309 40083 1343
rect 40083 1309 40092 1343
rect 40040 1300 40092 1309
rect 40316 1343 40368 1352
rect 40316 1309 40325 1343
rect 40325 1309 40359 1343
rect 40359 1309 40368 1343
rect 40316 1300 40368 1309
rect 40592 1343 40644 1352
rect 40592 1309 40601 1343
rect 40601 1309 40635 1343
rect 40635 1309 40644 1343
rect 40592 1300 40644 1309
rect 40868 1343 40920 1352
rect 40868 1309 40877 1343
rect 40877 1309 40911 1343
rect 40911 1309 40920 1343
rect 40868 1300 40920 1309
rect 41144 1343 41196 1352
rect 41144 1309 41153 1343
rect 41153 1309 41187 1343
rect 41187 1309 41196 1343
rect 41144 1300 41196 1309
rect 41420 1343 41472 1352
rect 41420 1309 41429 1343
rect 41429 1309 41463 1343
rect 41463 1309 41472 1343
rect 41420 1300 41472 1309
rect 41696 1343 41748 1352
rect 41696 1309 41705 1343
rect 41705 1309 41739 1343
rect 41739 1309 41748 1343
rect 41696 1300 41748 1309
rect 34888 1207 34940 1216
rect 34888 1173 34897 1207
rect 34897 1173 34931 1207
rect 34931 1173 34940 1207
rect 34888 1164 34940 1173
rect 35716 1164 35768 1216
rect 36912 1207 36964 1216
rect 36912 1173 36921 1207
rect 36921 1173 36955 1207
rect 36955 1173 36964 1207
rect 36912 1164 36964 1173
rect 37832 1164 37884 1216
rect 38660 1164 38712 1216
rect 38844 1207 38896 1216
rect 38844 1173 38853 1207
rect 38853 1173 38887 1207
rect 38887 1173 38896 1207
rect 38844 1164 38896 1173
rect 39120 1207 39172 1216
rect 39120 1173 39129 1207
rect 39129 1173 39163 1207
rect 39163 1173 39172 1207
rect 39120 1164 39172 1173
rect 39304 1164 39356 1216
rect 39672 1207 39724 1216
rect 39672 1173 39681 1207
rect 39681 1173 39715 1207
rect 39715 1173 39724 1207
rect 39672 1164 39724 1173
rect 40132 1207 40184 1216
rect 40132 1173 40141 1207
rect 40141 1173 40175 1207
rect 40175 1173 40184 1207
rect 40132 1164 40184 1173
rect 40684 1207 40736 1216
rect 40684 1173 40693 1207
rect 40693 1173 40727 1207
rect 40727 1173 40736 1207
rect 40684 1164 40736 1173
rect 11552 1062 11604 1114
rect 11616 1062 11668 1114
rect 11680 1062 11732 1114
rect 11744 1062 11796 1114
rect 11808 1062 11860 1114
rect 22155 1062 22207 1114
rect 22219 1062 22271 1114
rect 22283 1062 22335 1114
rect 22347 1062 22399 1114
rect 22411 1062 22463 1114
rect 32758 1062 32810 1114
rect 32822 1062 32874 1114
rect 32886 1062 32938 1114
rect 32950 1062 33002 1114
rect 33014 1062 33066 1114
rect 43361 1062 43413 1114
rect 43425 1062 43477 1114
rect 43489 1062 43541 1114
rect 43553 1062 43605 1114
rect 43617 1062 43669 1114
rect 4804 960 4856 1012
rect 6552 960 6604 1012
rect 9220 960 9272 1012
rect 12900 960 12952 1012
rect 13636 960 13688 1012
rect 14372 960 14424 1012
rect 15476 960 15528 1012
rect 15936 960 15988 1012
rect 17500 960 17552 1012
rect 18236 960 18288 1012
rect 18788 960 18840 1012
rect 32312 960 32364 1012
rect 32772 960 32824 1012
rect 34980 960 35032 1012
rect 36084 960 36136 1012
rect 38384 960 38436 1012
rect 9036 892 9088 944
rect 10232 892 10284 944
rect 5816 824 5868 876
rect 4896 416 4948 468
rect 6092 416 6144 468
rect 9312 824 9364 876
rect 16488 892 16540 944
rect 7656 756 7708 808
rect 12164 756 12216 808
rect 15752 824 15804 876
rect 18052 892 18104 944
rect 23756 892 23808 944
rect 23848 892 23900 944
rect 17408 824 17460 876
rect 18420 824 18472 876
rect 18696 824 18748 876
rect 19616 824 19668 876
rect 20168 824 20220 876
rect 27160 824 27212 876
rect 31208 824 31260 876
rect 13544 756 13596 808
rect 15384 756 15436 808
rect 16488 756 16540 808
rect 17776 756 17828 808
rect 19708 756 19760 808
rect 8668 688 8720 740
rect 8852 688 8904 740
rect 9312 688 9364 740
rect 10324 688 10376 740
rect 10968 688 11020 740
rect 11152 688 11204 740
rect 11796 688 11848 740
rect 13176 688 13228 740
rect 13728 688 13780 740
rect 15660 688 15712 740
rect 17040 688 17092 740
rect 17684 688 17736 740
rect 18604 688 18656 740
rect 31852 892 31904 944
rect 33048 892 33100 944
rect 35900 892 35952 944
rect 40132 960 40184 1012
rect 8760 552 8812 604
rect 14004 552 14056 604
rect 14740 620 14792 672
rect 15752 620 15804 672
rect 16396 620 16448 672
rect 17776 620 17828 672
rect 17960 620 18012 672
rect 18972 620 19024 672
rect 19524 620 19576 672
rect 20996 620 21048 672
rect 25044 620 25096 672
rect 26148 620 26200 672
rect 15016 552 15068 604
rect 15200 552 15252 604
rect 16304 552 16356 604
rect 18328 552 18380 604
rect 21916 552 21968 604
rect 26792 688 26844 740
rect 27620 620 27672 672
rect 30932 620 30984 672
rect 32220 688 32272 740
rect 39120 756 39172 808
rect 36544 688 36596 740
rect 40684 688 40736 740
rect 32128 620 32180 672
rect 35348 620 35400 672
rect 37648 620 37700 672
rect 34888 552 34940 604
rect 36820 552 36872 604
rect 11336 416 11388 468
rect 8944 348 8996 400
rect 12992 416 13044 468
rect 18880 484 18932 536
rect 23572 484 23624 536
rect 38660 484 38712 536
rect 39212 484 39264 536
rect 41696 484 41748 536
rect 13912 416 13964 468
rect 15200 416 15252 468
rect 7196 212 7248 264
rect 14004 348 14056 400
rect 19432 348 19484 400
rect 20260 348 20312 400
rect 30748 416 30800 468
rect 31668 416 31720 468
rect 34796 416 34848 468
rect 27528 348 27580 400
rect 30288 348 30340 400
rect 13636 280 13688 332
rect 26884 280 26936 332
rect 36912 348 36964 400
rect 38844 348 38896 400
rect 41420 348 41472 400
rect 23020 212 23072 264
rect 24400 212 24452 264
rect 37832 280 37884 332
rect 29736 212 29788 264
rect 32496 212 32548 264
rect 20812 144 20864 196
rect 21272 144 21324 196
rect 24584 144 24636 196
rect 6092 76 6144 128
rect 6368 76 6420 128
rect 10232 76 10284 128
rect 18512 76 18564 128
rect 15016 8 15068 60
rect 21916 76 21968 128
rect 26792 76 26844 128
rect 35716 76 35768 128
rect 38108 76 38160 128
<< metal2 >>
rect 1122 9840 1178 10300
rect 3238 9840 3294 10300
rect 5354 9840 5410 10300
rect 7470 9840 7526 10300
rect 9586 9840 9642 10300
rect 11702 9840 11758 10300
rect 13818 9840 13874 10300
rect 15934 9840 15990 10300
rect 18050 9840 18106 10300
rect 20166 9840 20222 10300
rect 22282 9840 22338 10300
rect 22388 9846 22600 9874
rect 1136 9058 1164 9840
rect 1136 9030 1256 9058
rect 1228 8634 1256 9030
rect 3252 8634 3280 9840
rect 5368 9058 5396 9840
rect 5368 9030 5488 9058
rect 5460 8634 5488 9030
rect 7484 8634 7512 9840
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7576 8498 7604 8774
rect 9600 8634 9628 9840
rect 11716 8922 11744 9840
rect 11716 8894 11928 8922
rect 11552 8732 11860 8741
rect 11552 8730 11558 8732
rect 11614 8730 11638 8732
rect 11694 8730 11718 8732
rect 11774 8730 11798 8732
rect 11854 8730 11860 8732
rect 11614 8678 11616 8730
rect 11796 8678 11798 8730
rect 11552 8676 11558 8678
rect 11614 8676 11638 8678
rect 11694 8676 11718 8678
rect 11774 8676 11798 8678
rect 11854 8676 11860 8678
rect 11552 8667 11860 8676
rect 11900 8634 11928 8894
rect 13832 8634 13860 9840
rect 15948 8634 15976 9840
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 15936 8628 15988 8634
rect 18064 8616 18092 9840
rect 20180 8634 20208 9840
rect 22296 9738 22324 9840
rect 22388 9738 22416 9846
rect 22296 9710 22416 9738
rect 22155 8732 22463 8741
rect 22155 8730 22161 8732
rect 22217 8730 22241 8732
rect 22297 8730 22321 8732
rect 22377 8730 22401 8732
rect 22457 8730 22463 8732
rect 22217 8678 22219 8730
rect 22399 8678 22401 8730
rect 22155 8676 22161 8678
rect 22217 8676 22241 8678
rect 22297 8676 22321 8678
rect 22377 8676 22401 8678
rect 22457 8676 22463 8678
rect 22155 8667 22463 8676
rect 22572 8634 22600 9846
rect 24398 9840 24454 10300
rect 26514 9840 26570 10300
rect 28630 9840 28686 10300
rect 30746 9840 30802 10300
rect 32862 9840 32918 10300
rect 34978 9840 35034 10300
rect 37094 9840 37150 10300
rect 39210 9840 39266 10300
rect 41326 9840 41382 10300
rect 43442 9840 43498 10300
rect 24412 8634 24440 9840
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 18144 8628 18196 8634
rect 18064 8588 18144 8616
rect 15936 8570 15988 8576
rect 18144 8570 18196 8576
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 9586 8528 9642 8537
rect 7564 8492 7616 8498
rect 9586 8463 9588 8472
rect 7564 8434 7616 8440
rect 9640 8463 9642 8472
rect 14096 8492 14148 8498
rect 9588 8434 9640 8440
rect 14096 8434 14148 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 2226 8392 2282 8401
rect 14108 8378 14136 8434
rect 14108 8362 14320 8378
rect 14108 8356 14332 8362
rect 14108 8350 14280 8356
rect 2226 8327 2228 8336
rect 2280 8327 2282 8336
rect 2228 8298 2280 8304
rect 14280 8298 14332 8304
rect 6251 8188 6559 8197
rect 6251 8186 6257 8188
rect 6313 8186 6337 8188
rect 6393 8186 6417 8188
rect 6473 8186 6497 8188
rect 6553 8186 6559 8188
rect 6313 8134 6315 8186
rect 6495 8134 6497 8186
rect 6251 8132 6257 8134
rect 6313 8132 6337 8134
rect 6393 8132 6417 8134
rect 6473 8132 6497 8134
rect 6553 8132 6559 8134
rect 6251 8123 6559 8132
rect 11552 7644 11860 7653
rect 11552 7642 11558 7644
rect 11614 7642 11638 7644
rect 11694 7642 11718 7644
rect 11774 7642 11798 7644
rect 11854 7642 11860 7644
rect 11614 7590 11616 7642
rect 11796 7590 11798 7642
rect 11552 7588 11558 7590
rect 11614 7588 11638 7590
rect 11694 7588 11718 7590
rect 11774 7588 11798 7590
rect 11854 7588 11860 7590
rect 11552 7579 11860 7588
rect 6251 7100 6559 7109
rect 6251 7098 6257 7100
rect 6313 7098 6337 7100
rect 6393 7098 6417 7100
rect 6473 7098 6497 7100
rect 6553 7098 6559 7100
rect 6313 7046 6315 7098
rect 6495 7046 6497 7098
rect 6251 7044 6257 7046
rect 6313 7044 6337 7046
rect 6393 7044 6417 7046
rect 6473 7044 6497 7046
rect 6553 7044 6559 7046
rect 6251 7035 6559 7044
rect 11552 6556 11860 6565
rect 11552 6554 11558 6556
rect 11614 6554 11638 6556
rect 11694 6554 11718 6556
rect 11774 6554 11798 6556
rect 11854 6554 11860 6556
rect 11614 6502 11616 6554
rect 11796 6502 11798 6554
rect 11552 6500 11558 6502
rect 11614 6500 11638 6502
rect 11694 6500 11718 6502
rect 11774 6500 11798 6502
rect 11854 6500 11860 6502
rect 11552 6491 11860 6500
rect 6251 6012 6559 6021
rect 6251 6010 6257 6012
rect 6313 6010 6337 6012
rect 6393 6010 6417 6012
rect 6473 6010 6497 6012
rect 6553 6010 6559 6012
rect 6313 5958 6315 6010
rect 6495 5958 6497 6010
rect 6251 5956 6257 5958
rect 6313 5956 6337 5958
rect 6393 5956 6417 5958
rect 6473 5956 6497 5958
rect 6553 5956 6559 5958
rect 6251 5947 6559 5956
rect 11552 5468 11860 5477
rect 11552 5466 11558 5468
rect 11614 5466 11638 5468
rect 11694 5466 11718 5468
rect 11774 5466 11798 5468
rect 11854 5466 11860 5468
rect 11614 5414 11616 5466
rect 11796 5414 11798 5466
rect 11552 5412 11558 5414
rect 11614 5412 11638 5414
rect 11694 5412 11718 5414
rect 11774 5412 11798 5414
rect 11854 5412 11860 5414
rect 11552 5403 11860 5412
rect 6251 4924 6559 4933
rect 6251 4922 6257 4924
rect 6313 4922 6337 4924
rect 6393 4922 6417 4924
rect 6473 4922 6497 4924
rect 6553 4922 6559 4924
rect 6313 4870 6315 4922
rect 6495 4870 6497 4922
rect 6251 4868 6257 4870
rect 6313 4868 6337 4870
rect 6393 4868 6417 4870
rect 6473 4868 6497 4870
rect 6553 4868 6559 4870
rect 6251 4859 6559 4868
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 7196 4208 7248 4214
rect 6734 4176 6790 4185
rect 7196 4150 7248 4156
rect 6734 4111 6790 4120
rect 6251 3836 6559 3845
rect 6251 3834 6257 3836
rect 6313 3834 6337 3836
rect 6393 3834 6417 3836
rect 6473 3834 6497 3836
rect 6553 3834 6559 3836
rect 6313 3782 6315 3834
rect 6495 3782 6497 3834
rect 6251 3780 6257 3782
rect 6313 3780 6337 3782
rect 6393 3780 6417 3782
rect 6473 3780 6497 3782
rect 6553 3780 6559 3782
rect 6251 3771 6559 3780
rect 6251 2748 6559 2757
rect 6251 2746 6257 2748
rect 6313 2746 6337 2748
rect 6393 2746 6417 2748
rect 6473 2746 6497 2748
rect 6553 2746 6559 2748
rect 6313 2694 6315 2746
rect 6495 2694 6497 2746
rect 6251 2692 6257 2694
rect 6313 2692 6337 2694
rect 6393 2692 6417 2694
rect 6473 2692 6497 2694
rect 6553 2692 6559 2694
rect 6251 2683 6559 2692
rect 6251 1660 6559 1669
rect 6251 1658 6257 1660
rect 6313 1658 6337 1660
rect 6393 1658 6417 1660
rect 6473 1658 6497 1660
rect 6553 1658 6559 1660
rect 6313 1606 6315 1658
rect 6495 1606 6497 1658
rect 6251 1604 6257 1606
rect 6313 1604 6337 1606
rect 6393 1604 6417 1606
rect 6473 1604 6497 1606
rect 6553 1604 6559 1606
rect 6251 1595 6559 1604
rect 5816 1488 5868 1494
rect 5816 1430 5868 1436
rect 4988 1284 5040 1290
rect 5264 1284 5316 1290
rect 5040 1244 5212 1272
rect 4988 1226 5040 1232
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 4816 1018 4844 1158
rect 4804 1012 4856 1018
rect 4804 954 4856 960
rect 4908 474 4936 1158
rect 4896 468 4948 474
rect 4896 410 4948 416
rect 5184 160 5212 1244
rect 5540 1284 5592 1290
rect 5316 1244 5488 1272
rect 5264 1226 5316 1232
rect 5460 160 5488 1244
rect 5592 1244 5764 1272
rect 5540 1226 5592 1232
rect 5736 160 5764 1244
rect 5828 882 5856 1430
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 5816 876 5868 882
rect 5816 818 5868 824
rect 5920 218 5948 1362
rect 6748 1358 6776 4111
rect 7208 1562 7236 4150
rect 8206 4040 8262 4049
rect 8128 3998 8206 4026
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 7380 1352 7432 1358
rect 7656 1352 7708 1358
rect 7432 1312 7512 1340
rect 7380 1294 7432 1300
rect 6012 354 6040 1294
rect 6276 1284 6328 1290
rect 6276 1226 6328 1232
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 474 6132 1158
rect 6092 468 6144 474
rect 6092 410 6144 416
rect 6012 326 6132 354
rect 5920 190 6040 218
rect 6012 160 6040 190
rect 5170 -300 5226 160
rect 5446 -300 5502 160
rect 5722 -300 5778 160
rect 5998 -300 6054 160
rect 6104 134 6132 326
rect 6288 160 6316 1226
rect 6380 218 6408 1294
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6564 1018 6592 1158
rect 6552 1012 6604 1018
rect 6552 954 6604 960
rect 6656 626 6684 1294
rect 7288 1284 7340 1290
rect 7288 1226 7340 1232
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 6656 598 6776 626
rect 6748 490 6776 598
rect 6748 462 6960 490
rect 6380 190 6684 218
rect 6092 128 6144 134
rect 6092 70 6144 76
rect 6274 -300 6330 160
rect 6368 128 6420 134
rect 6550 82 6606 160
rect 6420 76 6606 82
rect 6368 70 6606 76
rect 6380 54 6606 70
rect 6656 82 6684 190
rect 6826 82 6882 160
rect 6656 54 6882 82
rect 6932 82 6960 462
rect 7208 270 7236 1158
rect 7196 264 7248 270
rect 7196 206 7248 212
rect 7102 82 7158 160
rect 6932 54 7158 82
rect 7300 82 7328 1226
rect 7378 82 7434 160
rect 7300 54 7434 82
rect 7484 82 7512 1312
rect 7708 1312 7788 1340
rect 7656 1294 7708 1300
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7668 814 7696 1158
rect 7656 808 7708 814
rect 7656 750 7708 756
rect 7654 82 7710 160
rect 7484 54 7710 82
rect 7760 82 7788 1312
rect 7852 1290 7880 2926
rect 7932 1352 7984 1358
rect 7984 1312 8064 1340
rect 7932 1294 7984 1300
rect 7840 1284 7892 1290
rect 7840 1226 7892 1232
rect 7930 82 7986 160
rect 7760 54 7986 82
rect 8036 82 8064 1312
rect 8128 1222 8156 3998
rect 8206 3975 8262 3984
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 1222 8340 3334
rect 8588 1494 8616 4490
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9034 2000 9090 2009
rect 9034 1935 9090 1944
rect 9128 1964 9180 1970
rect 8942 1864 8998 1873
rect 8942 1799 8998 1808
rect 8576 1488 8628 1494
rect 8576 1430 8628 1436
rect 8484 1352 8536 1358
rect 8852 1352 8904 1358
rect 8536 1312 8616 1340
rect 8484 1294 8536 1300
rect 8392 1284 8444 1290
rect 8392 1226 8444 1232
rect 8116 1216 8168 1222
rect 8116 1158 8168 1164
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8404 762 8432 1226
rect 8404 734 8524 762
rect 8496 160 8524 734
rect 8206 82 8262 160
rect 8036 54 8262 82
rect 6550 -300 6606 54
rect 6826 -300 6882 54
rect 7102 -300 7158 54
rect 7378 -300 7434 54
rect 7654 -300 7710 54
rect 7930 -300 7986 54
rect 8206 -300 8262 54
rect 8482 -300 8538 160
rect 8588 82 8616 1312
rect 8852 1294 8904 1300
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8680 746 8708 1158
rect 8668 740 8720 746
rect 8668 682 8720 688
rect 8772 610 8800 1158
rect 8864 746 8892 1294
rect 8852 740 8904 746
rect 8852 682 8904 688
rect 8760 604 8812 610
rect 8760 546 8812 552
rect 8956 406 8984 1799
rect 9048 950 9076 1935
rect 9128 1906 9180 1912
rect 9036 944 9088 950
rect 9036 886 9088 892
rect 8944 400 8996 406
rect 8944 342 8996 348
rect 8758 82 8814 160
rect 8588 54 8814 82
rect 8758 -300 8814 54
rect 9034 82 9090 160
rect 9140 82 9168 1906
rect 9232 1018 9260 4422
rect 11552 4380 11860 4389
rect 11552 4378 11558 4380
rect 11614 4378 11638 4380
rect 11694 4378 11718 4380
rect 11774 4378 11798 4380
rect 11854 4378 11860 4380
rect 11614 4326 11616 4378
rect 11796 4326 11798 4378
rect 11552 4324 11558 4326
rect 11614 4324 11638 4326
rect 11694 4324 11718 4326
rect 11774 4324 11798 4326
rect 11854 4324 11860 4326
rect 11552 4315 11860 4324
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10980 2106 11008 2994
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11072 1562 11100 2518
rect 11348 1562 11376 4218
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11552 3292 11860 3301
rect 11552 3290 11558 3292
rect 11614 3290 11638 3292
rect 11694 3290 11718 3292
rect 11774 3290 11798 3292
rect 11854 3290 11860 3292
rect 11614 3238 11616 3290
rect 11796 3238 11798 3290
rect 11552 3236 11558 3238
rect 11614 3236 11638 3238
rect 11694 3236 11718 3238
rect 11774 3236 11798 3238
rect 11854 3236 11860 3238
rect 11552 3227 11860 3236
rect 11426 3088 11482 3097
rect 11426 3023 11482 3032
rect 11060 1556 11112 1562
rect 11060 1498 11112 1504
rect 11336 1556 11388 1562
rect 11336 1498 11388 1504
rect 11440 1442 11468 3023
rect 11552 2204 11860 2213
rect 11552 2202 11558 2204
rect 11614 2202 11638 2204
rect 11694 2202 11718 2204
rect 11774 2202 11798 2204
rect 11854 2202 11860 2204
rect 11614 2150 11616 2202
rect 11796 2150 11798 2202
rect 11552 2148 11558 2150
rect 11614 2148 11638 2150
rect 11694 2148 11718 2150
rect 11774 2148 11798 2150
rect 11854 2148 11860 2150
rect 11552 2139 11860 2148
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 11348 1414 11468 1442
rect 9402 1320 9458 1329
rect 9402 1255 9458 1264
rect 9588 1284 9640 1290
rect 9416 1222 9444 1255
rect 9588 1226 9640 1232
rect 9312 1216 9364 1222
rect 9312 1158 9364 1164
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9220 1012 9272 1018
rect 9220 954 9272 960
rect 9324 882 9352 1158
rect 9312 876 9364 882
rect 9312 818 9364 824
rect 9312 740 9364 746
rect 9312 682 9364 688
rect 9324 160 9352 682
rect 9600 160 9628 1226
rect 9034 54 9168 82
rect 9034 -300 9090 54
rect 9310 -300 9366 160
rect 9586 -300 9642 160
rect 9692 82 9720 1362
rect 9864 1352 9916 1358
rect 10324 1352 10376 1358
rect 9916 1312 9996 1340
rect 9864 1294 9916 1300
rect 9862 82 9918 160
rect 9692 54 9918 82
rect 9968 82 9996 1312
rect 10324 1294 10376 1300
rect 10508 1352 10560 1358
rect 10508 1294 10560 1300
rect 10140 1216 10192 1222
rect 10140 1158 10192 1164
rect 10232 1216 10284 1222
rect 10232 1158 10284 1164
rect 10152 388 10180 1158
rect 10244 950 10272 1158
rect 10232 944 10284 950
rect 10232 886 10284 892
rect 10336 746 10364 1294
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10324 740 10376 746
rect 10324 682 10376 688
rect 10152 360 10272 388
rect 10138 82 10194 160
rect 10244 134 10272 360
rect 10428 160 10456 1226
rect 9968 54 10194 82
rect 10232 128 10284 134
rect 10232 70 10284 76
rect 9862 -300 9918 54
rect 10138 -300 10194 54
rect 10414 -300 10470 160
rect 10520 82 10548 1294
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10784 1216 10836 1222
rect 10784 1158 10836 1164
rect 10704 649 10732 1158
rect 10690 640 10746 649
rect 10690 575 10746 584
rect 10796 241 10824 1158
rect 10980 898 11008 1226
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 10980 870 11100 898
rect 10968 740 11020 746
rect 10968 682 11020 688
rect 10782 232 10838 241
rect 10782 167 10838 176
rect 10980 160 11008 682
rect 10690 82 10746 160
rect 10520 54 10746 82
rect 10690 -300 10746 54
rect 10966 -300 11022 160
rect 11072 82 11100 870
rect 11164 746 11192 1158
rect 11152 740 11204 746
rect 11152 682 11204 688
rect 11256 513 11284 1158
rect 11242 504 11298 513
rect 11348 474 11376 1414
rect 11428 1352 11480 1358
rect 11428 1294 11480 1300
rect 11440 762 11468 1294
rect 11888 1284 11940 1290
rect 11888 1226 11940 1232
rect 11552 1116 11860 1125
rect 11552 1114 11558 1116
rect 11614 1114 11638 1116
rect 11694 1114 11718 1116
rect 11774 1114 11798 1116
rect 11854 1114 11860 1116
rect 11614 1062 11616 1114
rect 11796 1062 11798 1114
rect 11552 1060 11558 1062
rect 11614 1060 11638 1062
rect 11694 1060 11718 1062
rect 11774 1060 11798 1062
rect 11854 1060 11860 1062
rect 11552 1051 11860 1060
rect 11900 762 11928 1226
rect 11992 1222 12020 3878
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 12254 3224 12310 3233
rect 12254 3159 12310 3168
rect 12268 1340 12296 3159
rect 13358 2952 13414 2961
rect 13358 2887 13414 2896
rect 12806 2136 12862 2145
rect 12806 2071 12862 2080
rect 12820 1562 12848 2071
rect 12808 1556 12860 1562
rect 12808 1498 12860 1504
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12176 1312 12296 1340
rect 11980 1216 12032 1222
rect 11980 1158 12032 1164
rect 12176 814 12204 1312
rect 12256 1216 12308 1222
rect 12256 1158 12308 1164
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12164 808 12216 814
rect 11440 734 11560 762
rect 11242 439 11298 448
rect 11336 468 11388 474
rect 11336 410 11388 416
rect 11532 160 11560 734
rect 11796 740 11848 746
rect 11900 734 12112 762
rect 12164 750 12216 756
rect 11796 682 11848 688
rect 11808 160 11836 682
rect 12084 160 12112 734
rect 12268 377 12296 1158
rect 12254 368 12310 377
rect 12254 303 12310 312
rect 12360 160 12388 1158
rect 12452 762 12480 1362
rect 13372 1358 13400 2887
rect 13542 2544 13598 2553
rect 13542 2479 13598 2488
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 12624 1352 12676 1358
rect 13176 1352 13228 1358
rect 12676 1312 13124 1340
rect 12624 1294 12676 1300
rect 12544 898 12572 1294
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12992 1216 13044 1222
rect 12992 1158 13044 1164
rect 12912 1018 12940 1158
rect 12900 1012 12952 1018
rect 12900 954 12952 960
rect 12544 870 12940 898
rect 12452 734 12664 762
rect 12636 160 12664 734
rect 12912 160 12940 870
rect 13004 474 13032 1158
rect 13096 626 13124 1312
rect 13176 1294 13228 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 13188 746 13216 1294
rect 13268 1284 13320 1290
rect 13268 1226 13320 1232
rect 13280 762 13308 1226
rect 13556 814 13584 2479
rect 13648 1222 13676 3470
rect 15304 2650 15332 8434
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15488 2530 15516 2790
rect 15764 2650 15792 2858
rect 16040 2650 16068 8434
rect 16854 8188 17162 8197
rect 16854 8186 16860 8188
rect 16916 8186 16940 8188
rect 16996 8186 17020 8188
rect 17076 8186 17100 8188
rect 17156 8186 17162 8188
rect 16916 8134 16918 8186
rect 17098 8134 17100 8186
rect 16854 8132 16860 8134
rect 16916 8132 16940 8134
rect 16996 8132 17020 8134
rect 17076 8132 17100 8134
rect 17156 8132 17162 8134
rect 16854 8123 17162 8132
rect 16854 7100 17162 7109
rect 16854 7098 16860 7100
rect 16916 7098 16940 7100
rect 16996 7098 17020 7100
rect 17076 7098 17100 7100
rect 17156 7098 17162 7100
rect 16916 7046 16918 7098
rect 17098 7046 17100 7098
rect 16854 7044 16860 7046
rect 16916 7044 16940 7046
rect 16996 7044 17020 7046
rect 17076 7044 17100 7046
rect 17156 7044 17162 7046
rect 16854 7035 17162 7044
rect 16854 6012 17162 6021
rect 16854 6010 16860 6012
rect 16916 6010 16940 6012
rect 16996 6010 17020 6012
rect 17076 6010 17100 6012
rect 17156 6010 17162 6012
rect 16916 5958 16918 6010
rect 17098 5958 17100 6010
rect 16854 5956 16860 5958
rect 16916 5956 16940 5958
rect 16996 5956 17020 5958
rect 17076 5956 17100 5958
rect 17156 5956 17162 5958
rect 16854 5947 17162 5956
rect 16854 4924 17162 4933
rect 16854 4922 16860 4924
rect 16916 4922 16940 4924
rect 16996 4922 17020 4924
rect 17076 4922 17100 4924
rect 17156 4922 17162 4924
rect 16916 4870 16918 4922
rect 17098 4870 17100 4922
rect 16854 4868 16860 4870
rect 16916 4868 16940 4870
rect 16996 4868 17020 4870
rect 17076 4868 17100 4870
rect 17156 4868 17162 4870
rect 16854 4859 17162 4868
rect 17314 3904 17370 3913
rect 17236 3862 17314 3890
rect 16854 3836 17162 3845
rect 16854 3834 16860 3836
rect 16916 3834 16940 3836
rect 16996 3834 17020 3836
rect 17076 3834 17100 3836
rect 17156 3834 17162 3836
rect 16916 3782 16918 3834
rect 17098 3782 17100 3834
rect 16854 3780 16860 3782
rect 16916 3780 16940 3782
rect 16996 3780 17020 3782
rect 17076 3780 17100 3782
rect 17156 3780 17162 3782
rect 16854 3771 17162 3780
rect 16578 3632 16634 3641
rect 16578 3567 16634 3576
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 15304 2514 15516 2530
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 15292 2508 15516 2514
rect 15344 2502 15516 2508
rect 15292 2450 15344 2456
rect 13740 1494 13768 2450
rect 15580 2446 15608 2518
rect 15568 2440 15620 2446
rect 14278 2408 14334 2417
rect 15568 2382 15620 2388
rect 14278 2343 14334 2352
rect 15200 2372 15252 2378
rect 14292 2106 14320 2343
rect 15200 2314 15252 2320
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 13728 1488 13780 1494
rect 13728 1430 13780 1436
rect 13728 1352 13780 1358
rect 13912 1352 13964 1358
rect 13780 1312 13860 1340
rect 13728 1294 13780 1300
rect 13636 1216 13688 1222
rect 13636 1158 13688 1164
rect 13636 1012 13688 1018
rect 13636 954 13688 960
rect 13544 808 13596 814
rect 13176 740 13228 746
rect 13280 734 13492 762
rect 13544 750 13596 756
rect 13176 682 13228 688
rect 13096 598 13216 626
rect 12992 468 13044 474
rect 12992 410 13044 416
rect 13188 160 13216 598
rect 13464 160 13492 734
rect 13648 338 13676 954
rect 13728 740 13780 746
rect 13728 682 13780 688
rect 13636 332 13688 338
rect 13636 274 13688 280
rect 13740 160 13768 682
rect 11242 82 11298 160
rect 11072 54 11298 82
rect 11242 -300 11298 54
rect 11518 -300 11574 160
rect 11794 -300 11850 160
rect 12070 -300 12126 160
rect 12346 -300 12402 160
rect 12622 -300 12678 160
rect 12898 -300 12954 160
rect 13174 -300 13230 160
rect 13450 -300 13506 160
rect 13726 -300 13782 160
rect 13832 82 13860 1312
rect 13912 1294 13964 1300
rect 13924 474 13952 1294
rect 14108 1034 14136 1906
rect 14464 1760 14516 1766
rect 14464 1702 14516 1708
rect 14476 1562 14504 1702
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 14372 1216 14424 1222
rect 14372 1158 14424 1164
rect 14108 1006 14320 1034
rect 14384 1018 14412 1158
rect 14660 1034 14688 1906
rect 14844 1494 14872 2246
rect 15212 2122 15240 2314
rect 15658 2272 15714 2281
rect 15658 2207 15714 2216
rect 15028 2094 15240 2122
rect 15672 2106 15700 2207
rect 16224 2106 16252 3402
rect 16592 2802 16620 3567
rect 16762 3496 16818 3505
rect 16500 2774 16620 2802
rect 16684 3454 16762 3482
rect 16500 2514 16528 2774
rect 16488 2508 16540 2514
rect 16488 2450 16540 2456
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 15292 2100 15344 2106
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 14832 1488 14884 1494
rect 14832 1430 14884 1436
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 14004 604 14056 610
rect 14004 546 14056 552
rect 13912 468 13964 474
rect 13912 410 13964 416
rect 14016 406 14044 546
rect 14004 400 14056 406
rect 14004 342 14056 348
rect 14292 160 14320 1006
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 14568 1006 14688 1034
rect 14568 160 14596 1006
rect 14752 678 14780 1294
rect 14936 1034 14964 1906
rect 15028 1222 15056 2094
rect 15476 2100 15528 2106
rect 15344 2060 15476 2088
rect 15292 2042 15344 2048
rect 15476 2042 15528 2048
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 15108 2032 15160 2038
rect 15108 1974 15160 1980
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 14844 1006 14964 1034
rect 14740 672 14792 678
rect 14740 614 14792 620
rect 14844 160 14872 1006
rect 15016 604 15068 610
rect 15016 546 15068 552
rect 14002 82 14058 160
rect 13832 54 14058 82
rect 14002 -300 14058 54
rect 14278 -300 14334 160
rect 14554 -300 14610 160
rect 14830 -300 14886 160
rect 15028 66 15056 546
rect 15120 160 15148 1974
rect 16316 1970 16344 2246
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16396 1964 16448 1970
rect 16396 1906 16448 1912
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 15212 1737 15240 1770
rect 15198 1728 15254 1737
rect 15198 1663 15254 1672
rect 15304 1562 15332 1906
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 15292 1556 15344 1562
rect 15292 1498 15344 1504
rect 15396 1442 15424 1770
rect 15856 1578 15884 1906
rect 15304 1414 15424 1442
rect 15488 1550 15884 1578
rect 16408 1562 16436 1906
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 16488 1760 16540 1766
rect 16592 1737 16620 1838
rect 16684 1834 16712 3454
rect 16762 3431 16818 3440
rect 16854 2748 17162 2757
rect 16854 2746 16860 2748
rect 16916 2746 16940 2748
rect 16996 2746 17020 2748
rect 17076 2746 17100 2748
rect 17156 2746 17162 2748
rect 16916 2694 16918 2746
rect 17098 2694 17100 2746
rect 16854 2692 16860 2694
rect 16916 2692 16940 2694
rect 16996 2692 17020 2694
rect 17076 2692 17100 2694
rect 17156 2692 17162 2694
rect 16854 2683 17162 2692
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16764 2440 16816 2446
rect 16868 2417 16896 2518
rect 17236 2514 17264 3862
rect 17314 3839 17370 3848
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17696 2961 17724 3062
rect 17682 2952 17738 2961
rect 17500 2916 17552 2922
rect 17682 2887 17738 2896
rect 17866 2952 17922 2961
rect 17866 2887 17922 2896
rect 17500 2858 17552 2864
rect 17512 2689 17540 2858
rect 17774 2816 17830 2825
rect 17604 2774 17774 2802
rect 17498 2680 17554 2689
rect 17498 2615 17554 2624
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17316 2440 17368 2446
rect 16764 2382 16816 2388
rect 16854 2408 16910 2417
rect 16776 2310 16804 2382
rect 17316 2382 17368 2388
rect 16854 2343 16910 2352
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16856 2304 16908 2310
rect 17224 2304 17276 2310
rect 16856 2246 16908 2252
rect 17052 2264 17224 2292
rect 16868 2106 16896 2246
rect 17052 2106 17080 2264
rect 17224 2246 17276 2252
rect 17130 2136 17186 2145
rect 16856 2100 16908 2106
rect 16856 2042 16908 2048
rect 17040 2100 17092 2106
rect 17130 2071 17132 2080
rect 17040 2042 17092 2048
rect 17184 2071 17186 2080
rect 17132 2042 17184 2048
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 16856 1760 16908 1766
rect 16488 1702 16540 1708
rect 16578 1728 16634 1737
rect 16396 1556 16448 1562
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15212 610 15240 1294
rect 15304 785 15332 1414
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15396 814 15424 1294
rect 15488 1018 15516 1550
rect 16396 1498 16448 1504
rect 15660 1488 15712 1494
rect 16500 1465 16528 1702
rect 16578 1663 16634 1672
rect 16776 1720 16856 1748
rect 16486 1456 16542 1465
rect 15712 1436 16252 1442
rect 15660 1430 16252 1436
rect 15568 1420 15620 1426
rect 15672 1414 16252 1430
rect 15568 1362 15620 1368
rect 15476 1012 15528 1018
rect 15476 954 15528 960
rect 15384 808 15436 814
rect 15290 776 15346 785
rect 15384 750 15436 756
rect 15290 711 15346 720
rect 15580 626 15608 1362
rect 15660 1352 15712 1358
rect 15660 1294 15712 1300
rect 15936 1352 15988 1358
rect 15936 1294 15988 1300
rect 15672 746 15700 1294
rect 15752 1216 15804 1222
rect 15752 1158 15804 1164
rect 15764 882 15792 1158
rect 15948 1018 15976 1294
rect 15936 1012 15988 1018
rect 15936 954 15988 960
rect 15752 876 15804 882
rect 15752 818 15804 824
rect 15660 740 15712 746
rect 15660 682 15712 688
rect 15752 672 15804 678
rect 15200 604 15252 610
rect 15580 598 15700 626
rect 15804 620 15976 626
rect 15752 614 15976 620
rect 15764 598 15976 614
rect 15200 546 15252 552
rect 15200 468 15252 474
rect 15200 410 15252 416
rect 15212 354 15240 410
rect 15212 326 15424 354
rect 15396 160 15424 326
rect 15672 160 15700 598
rect 15948 160 15976 598
rect 16224 160 16252 1414
rect 16776 1426 16804 1720
rect 16856 1702 16908 1708
rect 16854 1660 17162 1669
rect 16854 1658 16860 1660
rect 16916 1658 16940 1660
rect 16996 1658 17020 1660
rect 17076 1658 17100 1660
rect 17156 1658 17162 1660
rect 16916 1606 16918 1658
rect 17098 1606 17100 1658
rect 16854 1604 16860 1606
rect 16916 1604 16940 1606
rect 16996 1604 17020 1606
rect 17076 1604 17100 1606
rect 17156 1604 17162 1606
rect 16854 1595 17162 1604
rect 17132 1488 17184 1494
rect 17236 1476 17264 1974
rect 17184 1448 17264 1476
rect 17132 1430 17184 1436
rect 16486 1391 16542 1400
rect 16764 1420 16816 1426
rect 16764 1362 16816 1368
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 16488 1352 16540 1358
rect 16488 1294 16540 1300
rect 16408 678 16436 1294
rect 16500 1057 16528 1294
rect 16486 1048 16542 1057
rect 16486 983 16542 992
rect 16488 944 16540 950
rect 16486 912 16488 921
rect 16540 912 16542 921
rect 16486 847 16542 856
rect 16488 808 16540 814
rect 16540 768 16620 796
rect 16488 750 16540 756
rect 16396 672 16448 678
rect 16396 614 16448 620
rect 16304 604 16356 610
rect 16304 546 16356 552
rect 16316 490 16344 546
rect 16316 462 16528 490
rect 16500 160 16528 462
rect 15016 60 15068 66
rect 15016 2 15068 8
rect 15106 -300 15162 160
rect 15382 -300 15438 160
rect 15658 -300 15714 160
rect 15934 -300 15990 160
rect 16210 -300 16266 160
rect 16486 -300 16542 160
rect 16592 82 16620 768
rect 17040 740 17092 746
rect 17040 682 17092 688
rect 17052 160 17080 682
rect 17328 160 17356 2382
rect 17604 1986 17632 2774
rect 17774 2751 17830 2760
rect 17880 2650 17908 2887
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17972 2582 18000 3538
rect 18064 2650 18092 8434
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18234 3088 18290 3097
rect 18234 3023 18290 3032
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18064 2417 18092 2450
rect 18050 2408 18106 2417
rect 18050 2343 18106 2352
rect 18156 2258 18184 2858
rect 17420 1958 17632 1986
rect 18064 2230 18184 2258
rect 18064 1970 18092 2230
rect 18144 1988 18196 1994
rect 18052 1964 18104 1970
rect 17420 1562 17448 1958
rect 18248 1986 18276 3023
rect 18984 2446 19012 3130
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18420 2440 18472 2446
rect 18972 2440 19024 2446
rect 18472 2400 18644 2428
rect 18420 2382 18472 2388
rect 18420 2100 18472 2106
rect 18472 2060 18552 2088
rect 18420 2042 18472 2048
rect 18196 1958 18276 1986
rect 18144 1930 18196 1936
rect 18052 1906 18104 1912
rect 17684 1896 17736 1902
rect 17512 1873 17684 1884
rect 17498 1864 17684 1873
rect 17554 1856 17684 1864
rect 17684 1838 17736 1844
rect 17866 1864 17922 1873
rect 17498 1799 17554 1808
rect 18050 1864 18106 1873
rect 17922 1822 18050 1850
rect 17866 1799 17922 1808
rect 18050 1799 18106 1808
rect 17684 1760 17736 1766
rect 17682 1728 17684 1737
rect 17868 1760 17920 1766
rect 17736 1728 17738 1737
rect 17868 1702 17920 1708
rect 17960 1760 18012 1766
rect 18012 1737 18276 1748
rect 18012 1728 18290 1737
rect 18012 1720 18234 1728
rect 17960 1702 18012 1708
rect 17682 1663 17738 1672
rect 17774 1592 17830 1601
rect 17408 1556 17460 1562
rect 17880 1562 17908 1702
rect 18234 1663 18290 1672
rect 18524 1562 18552 2060
rect 17774 1527 17830 1536
rect 17868 1556 17920 1562
rect 17408 1498 17460 1504
rect 17788 1494 17816 1527
rect 17868 1498 17920 1504
rect 18512 1556 18564 1562
rect 18512 1498 18564 1504
rect 18616 1494 18644 2400
rect 18972 2382 19024 2388
rect 18694 2000 18750 2009
rect 19076 1970 19104 2790
rect 20272 2582 20300 8434
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22155 7644 22463 7653
rect 22155 7642 22161 7644
rect 22217 7642 22241 7644
rect 22297 7642 22321 7644
rect 22377 7642 22401 7644
rect 22457 7642 22463 7644
rect 22217 7590 22219 7642
rect 22399 7590 22401 7642
rect 22155 7588 22161 7590
rect 22217 7588 22241 7590
rect 22297 7588 22321 7590
rect 22377 7588 22401 7590
rect 22457 7588 22463 7590
rect 22155 7579 22463 7588
rect 22155 6556 22463 6565
rect 22155 6554 22161 6556
rect 22217 6554 22241 6556
rect 22297 6554 22321 6556
rect 22377 6554 22401 6556
rect 22457 6554 22463 6556
rect 22217 6502 22219 6554
rect 22399 6502 22401 6554
rect 22155 6500 22161 6502
rect 22217 6500 22241 6502
rect 22297 6500 22321 6502
rect 22377 6500 22401 6502
rect 22457 6500 22463 6502
rect 22155 6491 22463 6500
rect 22155 5468 22463 5477
rect 22155 5466 22161 5468
rect 22217 5466 22241 5468
rect 22297 5466 22321 5468
rect 22377 5466 22401 5468
rect 22457 5466 22463 5468
rect 22217 5414 22219 5466
rect 22399 5414 22401 5466
rect 22155 5412 22161 5414
rect 22217 5412 22241 5414
rect 22297 5412 22321 5414
rect 22377 5412 22401 5414
rect 22457 5412 22463 5414
rect 22155 5403 22463 5412
rect 22155 4380 22463 4389
rect 22155 4378 22161 4380
rect 22217 4378 22241 4380
rect 22297 4378 22321 4380
rect 22377 4378 22401 4380
rect 22457 4378 22463 4380
rect 22217 4326 22219 4378
rect 22399 4326 22401 4378
rect 22155 4324 22161 4326
rect 22217 4324 22241 4326
rect 22297 4324 22321 4326
rect 22377 4324 22401 4326
rect 22457 4324 22463 4326
rect 22155 4315 22463 4324
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20364 2689 20392 2858
rect 20456 2774 20484 3334
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 20456 2746 20668 2774
rect 20350 2680 20406 2689
rect 20350 2615 20406 2624
rect 20076 2576 20128 2582
rect 20260 2576 20312 2582
rect 20076 2518 20128 2524
rect 20166 2544 20222 2553
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19430 2136 19486 2145
rect 19168 2094 19430 2122
rect 18694 1935 18696 1944
rect 18748 1935 18750 1944
rect 18788 1964 18840 1970
rect 18696 1906 18748 1912
rect 18788 1906 18840 1912
rect 19064 1964 19116 1970
rect 19064 1906 19116 1912
rect 18694 1864 18750 1873
rect 18694 1799 18696 1808
rect 18748 1799 18750 1808
rect 18696 1770 18748 1776
rect 18694 1728 18750 1737
rect 18694 1663 18750 1672
rect 18708 1494 18736 1663
rect 17776 1488 17828 1494
rect 17776 1430 17828 1436
rect 18052 1488 18104 1494
rect 18604 1488 18656 1494
rect 18052 1430 18104 1436
rect 18142 1456 18198 1465
rect 17408 1352 17460 1358
rect 17408 1294 17460 1300
rect 17684 1352 17736 1358
rect 17684 1294 17736 1300
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 17420 882 17448 1294
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 17408 876 17460 882
rect 17408 818 17460 824
rect 17512 762 17540 954
rect 17512 734 17632 762
rect 17696 746 17724 1294
rect 17776 1216 17828 1222
rect 17776 1158 17828 1164
rect 17788 814 17816 1158
rect 17776 808 17828 814
rect 17776 750 17828 756
rect 17604 160 17632 734
rect 17684 740 17736 746
rect 17684 682 17736 688
rect 17972 678 18000 1294
rect 18064 950 18092 1430
rect 18604 1430 18656 1436
rect 18696 1488 18748 1494
rect 18696 1430 18748 1436
rect 18142 1391 18198 1400
rect 18156 1306 18184 1391
rect 18800 1306 18828 1906
rect 18972 1760 19024 1766
rect 19168 1748 19196 2094
rect 19430 2071 19486 2080
rect 19432 1964 19484 1970
rect 19432 1906 19484 1912
rect 19024 1720 19196 1748
rect 19248 1760 19300 1766
rect 18972 1702 19024 1708
rect 19340 1760 19392 1766
rect 19248 1702 19300 1708
rect 19338 1728 19340 1737
rect 19392 1728 19394 1737
rect 18880 1420 18932 1426
rect 18880 1362 18932 1368
rect 18156 1278 18368 1306
rect 18236 1216 18288 1222
rect 18236 1158 18288 1164
rect 18142 1048 18198 1057
rect 18248 1018 18276 1158
rect 18142 983 18198 992
rect 18236 1012 18288 1018
rect 18052 944 18104 950
rect 18052 886 18104 892
rect 17776 672 17828 678
rect 17960 672 18012 678
rect 17828 620 17908 626
rect 17776 614 17908 620
rect 17960 614 18012 620
rect 17788 598 17908 614
rect 17880 160 17908 598
rect 18156 160 18184 983
rect 18236 954 18288 960
rect 18340 610 18368 1278
rect 18524 1278 18828 1306
rect 18420 876 18472 882
rect 18420 818 18472 824
rect 18328 604 18380 610
rect 18328 546 18380 552
rect 18432 160 18460 818
rect 16762 82 16818 160
rect 16592 54 16818 82
rect 16762 -300 16818 54
rect 17038 -300 17094 160
rect 17314 -300 17370 160
rect 17590 -300 17646 160
rect 17866 -300 17922 160
rect 18142 -300 18198 160
rect 18418 -300 18474 160
rect 18524 134 18552 1278
rect 18696 1216 18748 1222
rect 18696 1158 18748 1164
rect 18788 1216 18840 1222
rect 18788 1158 18840 1164
rect 18708 882 18736 1158
rect 18800 1018 18828 1158
rect 18788 1012 18840 1018
rect 18788 954 18840 960
rect 18696 876 18748 882
rect 18696 818 18748 824
rect 18604 740 18656 746
rect 18604 682 18656 688
rect 18616 626 18644 682
rect 18616 598 18736 626
rect 18708 160 18736 598
rect 18892 542 18920 1362
rect 18972 1352 19024 1358
rect 19260 1340 19288 1702
rect 19338 1663 19394 1672
rect 19024 1312 19104 1340
rect 19260 1312 19380 1340
rect 18972 1294 19024 1300
rect 18972 672 19024 678
rect 18972 614 19024 620
rect 18880 536 18932 542
rect 18880 478 18932 484
rect 18984 160 19012 614
rect 19076 354 19104 1312
rect 19352 1193 19380 1312
rect 19338 1184 19394 1193
rect 19338 1119 19394 1128
rect 19444 406 19472 1906
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 19536 1358 19564 1770
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19628 882 19656 2382
rect 19708 2372 19760 2378
rect 19708 2314 19760 2320
rect 19720 1816 19748 2314
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19904 2145 19932 2246
rect 19890 2136 19946 2145
rect 19890 2071 19946 2080
rect 19890 2000 19946 2009
rect 19890 1935 19892 1944
rect 19944 1935 19946 1944
rect 19892 1906 19944 1912
rect 19702 1788 19748 1816
rect 19702 1578 19730 1788
rect 19702 1550 19748 1578
rect 19616 876 19668 882
rect 19616 818 19668 824
rect 19720 814 19748 1550
rect 19996 1329 20024 2382
rect 19982 1320 20038 1329
rect 19982 1255 20038 1264
rect 20088 1272 20116 2518
rect 20260 2518 20312 2524
rect 20166 2479 20222 2488
rect 20180 2446 20208 2479
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20166 1728 20222 1737
rect 20166 1663 20222 1672
rect 20180 1494 20208 1663
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 20088 1244 20208 1272
rect 19800 1216 19852 1222
rect 19800 1158 19852 1164
rect 19892 1216 19944 1222
rect 19944 1176 20116 1204
rect 19892 1158 19944 1164
rect 19708 808 19760 814
rect 19708 750 19760 756
rect 19524 672 19576 678
rect 19524 614 19576 620
rect 19432 400 19484 406
rect 19076 326 19288 354
rect 19432 342 19484 348
rect 19260 160 19288 326
rect 19536 160 19564 614
rect 19812 160 19840 1158
rect 20088 160 20116 1176
rect 20180 882 20208 1244
rect 20168 876 20220 882
rect 20168 818 20220 824
rect 20272 406 20300 2314
rect 20640 1970 20668 2746
rect 20718 2680 20774 2689
rect 20718 2615 20774 2624
rect 20732 2281 20760 2615
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20718 2272 20774 2281
rect 20718 2207 20774 2216
rect 20718 2136 20774 2145
rect 20718 2071 20774 2080
rect 20732 2038 20760 2071
rect 20720 2032 20772 2038
rect 20720 1974 20772 1980
rect 20628 1964 20680 1970
rect 20628 1906 20680 1912
rect 20812 1964 20864 1970
rect 20812 1906 20864 1912
rect 20364 1834 20484 1850
rect 20364 1828 20496 1834
rect 20364 1822 20444 1828
rect 20260 400 20312 406
rect 20260 342 20312 348
rect 20364 160 20392 1822
rect 20444 1770 20496 1776
rect 20444 1420 20496 1426
rect 20444 1362 20496 1368
rect 20456 626 20484 1362
rect 20536 1284 20588 1290
rect 20536 1226 20588 1232
rect 20548 1193 20576 1226
rect 20534 1184 20590 1193
rect 20534 1119 20590 1128
rect 20456 598 20668 626
rect 20640 160 20668 598
rect 20824 202 20852 1906
rect 20916 1601 20944 2382
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 20902 1592 20958 1601
rect 20902 1527 20958 1536
rect 20904 1488 20956 1494
rect 20904 1430 20956 1436
rect 20812 196 20864 202
rect 18512 128 18564 134
rect 18512 70 18564 76
rect 18694 -300 18750 160
rect 18970 -300 19026 160
rect 19246 -300 19302 160
rect 19522 -300 19578 160
rect 19798 -300 19854 160
rect 20074 -300 20130 160
rect 20350 -300 20406 160
rect 20626 -300 20682 160
rect 20916 160 20944 1430
rect 21008 678 21036 2042
rect 21192 2009 21220 2790
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21178 2000 21234 2009
rect 21178 1935 21234 1944
rect 20996 672 21048 678
rect 20996 614 21048 620
rect 21284 202 21312 2382
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21364 1760 21416 1766
rect 21364 1702 21416 1708
rect 21272 196 21324 202
rect 20812 138 20864 144
rect 20902 -300 20958 160
rect 21178 82 21234 160
rect 21272 138 21324 144
rect 21376 82 21404 1702
rect 21468 160 21496 2246
rect 21560 1358 21588 2246
rect 21744 2038 21772 2790
rect 21836 2446 21864 3975
rect 22155 3292 22463 3301
rect 22155 3290 22161 3292
rect 22217 3290 22241 3292
rect 22297 3290 22321 3292
rect 22377 3290 22401 3292
rect 22457 3290 22463 3292
rect 22217 3238 22219 3290
rect 22399 3238 22401 3290
rect 22155 3236 22161 3238
rect 22217 3236 22241 3238
rect 22297 3236 22321 3238
rect 22377 3236 22401 3238
rect 22457 3236 22463 3238
rect 22155 3227 22463 3236
rect 22282 3088 22338 3097
rect 22282 3023 22338 3032
rect 22296 2446 22324 3023
rect 22572 2650 22600 8298
rect 22756 2650 22784 8434
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 23216 2582 23244 8366
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22928 2304 22980 2310
rect 23294 2272 23350 2281
rect 22928 2246 22980 2252
rect 21732 2032 21784 2038
rect 21732 1974 21784 1980
rect 21824 1760 21876 1766
rect 21824 1702 21876 1708
rect 21548 1352 21600 1358
rect 21548 1294 21600 1300
rect 21836 1222 21864 1702
rect 21928 1290 21956 2246
rect 22155 2204 22463 2213
rect 22155 2202 22161 2204
rect 22217 2202 22241 2204
rect 22297 2202 22321 2204
rect 22377 2202 22401 2204
rect 22457 2202 22463 2204
rect 22217 2150 22219 2202
rect 22399 2150 22401 2202
rect 22155 2148 22161 2150
rect 22217 2148 22241 2150
rect 22297 2148 22321 2150
rect 22377 2148 22401 2150
rect 22457 2148 22463 2150
rect 22155 2139 22463 2148
rect 22008 1760 22060 1766
rect 22836 1760 22888 1766
rect 22008 1702 22060 1708
rect 22756 1720 22836 1748
rect 21916 1284 21968 1290
rect 21916 1226 21968 1232
rect 21548 1216 21600 1222
rect 21824 1216 21876 1222
rect 21600 1176 21772 1204
rect 21548 1158 21600 1164
rect 21744 160 21772 1176
rect 21824 1158 21876 1164
rect 21916 604 21968 610
rect 21916 546 21968 552
rect 21178 54 21404 82
rect 21178 -300 21234 54
rect 21454 -300 21510 160
rect 21730 -300 21786 160
rect 21928 134 21956 546
rect 22020 160 22048 1702
rect 22652 1556 22704 1562
rect 22652 1498 22704 1504
rect 22560 1420 22612 1426
rect 22560 1362 22612 1368
rect 22155 1116 22463 1125
rect 22155 1114 22161 1116
rect 22217 1114 22241 1116
rect 22297 1114 22321 1116
rect 22377 1114 22401 1116
rect 22457 1114 22463 1116
rect 22217 1062 22219 1114
rect 22399 1062 22401 1114
rect 22155 1060 22161 1062
rect 22217 1060 22241 1062
rect 22297 1060 22321 1062
rect 22377 1060 22401 1062
rect 22457 1060 22463 1062
rect 22155 1051 22463 1060
rect 22572 218 22600 1362
rect 22664 1193 22692 1498
rect 22650 1184 22706 1193
rect 22650 1119 22706 1128
rect 22480 190 22600 218
rect 21916 128 21968 134
rect 21916 70 21968 76
rect 22006 -300 22062 160
rect 22282 82 22338 160
rect 22480 82 22508 190
rect 22282 54 22508 82
rect 22558 82 22614 160
rect 22756 82 22784 1720
rect 22836 1702 22888 1708
rect 22940 1358 22968 2246
rect 23032 2230 23294 2258
rect 22928 1352 22980 1358
rect 22928 1294 22980 1300
rect 22928 1216 22980 1222
rect 22928 1158 22980 1164
rect 22558 54 22784 82
rect 22834 82 22890 160
rect 22940 82 22968 1158
rect 23032 270 23060 2230
rect 23294 2207 23350 2216
rect 23400 1970 23428 4490
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23388 1964 23440 1970
rect 23388 1906 23440 1912
rect 23388 1556 23440 1562
rect 23388 1498 23440 1504
rect 23296 1216 23348 1222
rect 23124 1176 23296 1204
rect 23020 264 23072 270
rect 23020 206 23072 212
rect 23124 160 23152 1176
rect 23296 1158 23348 1164
rect 23400 160 23428 1498
rect 23492 1358 23520 2790
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23584 542 23612 3130
rect 23676 1970 23704 4422
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23768 2106 23796 2450
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24044 2106 24072 2314
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 23848 1964 23900 1970
rect 23848 1906 23900 1912
rect 24124 1964 24176 1970
rect 24176 1924 24440 1952
rect 24124 1906 24176 1912
rect 23664 1216 23716 1222
rect 23664 1158 23716 1164
rect 23572 536 23624 542
rect 23572 478 23624 484
rect 23676 160 23704 1158
rect 23754 1048 23810 1057
rect 23754 983 23810 992
rect 23768 950 23796 983
rect 23860 950 23888 1906
rect 24216 1760 24268 1766
rect 23952 1720 24216 1748
rect 23756 944 23808 950
rect 23756 886 23808 892
rect 23848 944 23900 950
rect 23848 886 23900 892
rect 23952 160 23980 1720
rect 24216 1702 24268 1708
rect 24308 1556 24360 1562
rect 24228 1516 24308 1544
rect 24228 160 24256 1516
rect 24308 1498 24360 1504
rect 24412 270 24440 1924
rect 24400 264 24452 270
rect 24400 206 24452 212
rect 24596 202 24624 2382
rect 24872 2310 24900 8434
rect 25136 4208 25188 4214
rect 24950 4176 25006 4185
rect 25136 4150 25188 4156
rect 24950 4111 25006 4120
rect 24860 2304 24912 2310
rect 24860 2246 24912 2252
rect 24964 1970 24992 4111
rect 25148 2774 25176 4150
rect 25056 2746 25176 2774
rect 24952 1964 25004 1970
rect 25056 1952 25084 2746
rect 25332 2530 25360 8774
rect 26528 8634 26556 9840
rect 28644 8634 28672 9840
rect 30760 8634 30788 9840
rect 32876 9058 32904 9840
rect 32692 9030 32904 9058
rect 32692 8634 32720 9030
rect 32758 8732 33066 8741
rect 32758 8730 32764 8732
rect 32820 8730 32844 8732
rect 32900 8730 32924 8732
rect 32980 8730 33004 8732
rect 33060 8730 33066 8732
rect 32820 8678 32822 8730
rect 33002 8678 33004 8730
rect 32758 8676 32764 8678
rect 32820 8676 32844 8678
rect 32900 8676 32924 8678
rect 32980 8676 33004 8678
rect 33060 8676 33066 8678
rect 32758 8667 33066 8676
rect 34992 8634 35020 9840
rect 37108 8634 37136 9840
rect 39224 8634 39252 9840
rect 41340 8634 41368 9840
rect 43456 8922 43484 9840
rect 43272 8894 43484 8922
rect 43272 8634 43300 8894
rect 43361 8732 43669 8741
rect 43361 8730 43367 8732
rect 43423 8730 43447 8732
rect 43503 8730 43527 8732
rect 43583 8730 43607 8732
rect 43663 8730 43669 8732
rect 43423 8678 43425 8730
rect 43605 8678 43607 8730
rect 43361 8676 43367 8678
rect 43423 8676 43447 8678
rect 43503 8676 43527 8678
rect 43583 8676 43607 8678
rect 43663 8676 43669 8678
rect 43361 8667 43669 8676
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 37096 8628 37148 8634
rect 37096 8570 37148 8576
rect 39212 8628 39264 8634
rect 39212 8570 39264 8576
rect 41328 8628 41380 8634
rect 41328 8570 41380 8576
rect 43260 8628 43312 8634
rect 43260 8570 43312 8576
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 26988 6914 27016 8434
rect 27457 8188 27765 8197
rect 27457 8186 27463 8188
rect 27519 8186 27543 8188
rect 27599 8186 27623 8188
rect 27679 8186 27703 8188
rect 27759 8186 27765 8188
rect 27519 8134 27521 8186
rect 27701 8134 27703 8186
rect 27457 8132 27463 8134
rect 27519 8132 27543 8134
rect 27599 8132 27623 8134
rect 27679 8132 27703 8134
rect 27759 8132 27765 8134
rect 27457 8123 27765 8132
rect 27457 7100 27765 7109
rect 27457 7098 27463 7100
rect 27519 7098 27543 7100
rect 27599 7098 27623 7100
rect 27679 7098 27703 7100
rect 27759 7098 27765 7100
rect 27519 7046 27521 7098
rect 27701 7046 27703 7098
rect 27457 7044 27463 7046
rect 27519 7044 27543 7046
rect 27599 7044 27623 7046
rect 27679 7044 27703 7046
rect 27759 7044 27765 7046
rect 27457 7035 27765 7044
rect 26988 6886 27200 6914
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 25608 3058 25636 3470
rect 25688 3120 25740 3126
rect 25688 3062 25740 3068
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 25700 2774 25728 3062
rect 25700 2746 25820 2774
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25148 2502 25360 2530
rect 25148 2310 25176 2502
rect 25608 2446 25636 2586
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25596 2304 25648 2310
rect 25648 2264 25728 2292
rect 25596 2246 25648 2252
rect 25502 2000 25558 2009
rect 25228 1964 25280 1970
rect 25056 1924 25228 1952
rect 24952 1906 25004 1912
rect 25502 1935 25504 1944
rect 25228 1906 25280 1912
rect 25556 1935 25558 1944
rect 25504 1906 25556 1912
rect 24860 1828 24912 1834
rect 24860 1770 24912 1776
rect 24768 1760 24820 1766
rect 24768 1702 24820 1708
rect 24676 1488 24728 1494
rect 24676 1430 24728 1436
rect 24584 196 24636 202
rect 22834 54 22968 82
rect 22282 -300 22338 54
rect 22558 -300 22614 54
rect 22834 -300 22890 54
rect 23110 -300 23166 160
rect 23386 -300 23442 160
rect 23662 -300 23718 160
rect 23938 -300 23994 160
rect 24214 -300 24270 160
rect 24490 82 24546 160
rect 24584 138 24636 144
rect 24688 82 24716 1430
rect 24780 1358 24808 1702
rect 24768 1352 24820 1358
rect 24768 1294 24820 1300
rect 24872 1290 24900 1770
rect 25044 1760 25096 1766
rect 25044 1702 25096 1708
rect 25596 1760 25648 1766
rect 25596 1702 25648 1708
rect 25056 1290 25084 1702
rect 25504 1420 25556 1426
rect 25504 1362 25556 1368
rect 24860 1284 24912 1290
rect 24860 1226 24912 1232
rect 25044 1284 25096 1290
rect 25044 1226 25096 1232
rect 24768 1216 24820 1222
rect 24768 1158 24820 1164
rect 24780 160 24808 1158
rect 25044 672 25096 678
rect 25044 614 25096 620
rect 25056 160 25084 614
rect 24490 54 24716 82
rect 24490 -300 24546 54
rect 24766 -300 24822 160
rect 25042 -300 25098 160
rect 25318 82 25374 160
rect 25516 82 25544 1362
rect 25608 160 25636 1702
rect 25700 1358 25728 2264
rect 25792 1952 25820 2746
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25884 2106 25912 2518
rect 26160 2446 26188 3470
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 25872 2100 25924 2106
rect 25872 2042 25924 2048
rect 26252 2038 26280 2790
rect 26528 2514 26556 2926
rect 26974 2680 27030 2689
rect 27172 2650 27200 6886
rect 27457 6012 27765 6021
rect 27457 6010 27463 6012
rect 27519 6010 27543 6012
rect 27599 6010 27623 6012
rect 27679 6010 27703 6012
rect 27759 6010 27765 6012
rect 27519 5958 27521 6010
rect 27701 5958 27703 6010
rect 27457 5956 27463 5958
rect 27519 5956 27543 5958
rect 27599 5956 27623 5958
rect 27679 5956 27703 5958
rect 27759 5956 27765 5958
rect 27457 5947 27765 5956
rect 27457 4924 27765 4933
rect 27457 4922 27463 4924
rect 27519 4922 27543 4924
rect 27599 4922 27623 4924
rect 27679 4922 27703 4924
rect 27759 4922 27765 4924
rect 27519 4870 27521 4922
rect 27701 4870 27703 4922
rect 27457 4868 27463 4870
rect 27519 4868 27543 4870
rect 27599 4868 27623 4870
rect 27679 4868 27703 4870
rect 27759 4868 27765 4870
rect 27457 4859 27765 4868
rect 28080 4276 28132 4282
rect 28080 4218 28132 4224
rect 27457 3836 27765 3845
rect 27457 3834 27463 3836
rect 27519 3834 27543 3836
rect 27599 3834 27623 3836
rect 27679 3834 27703 3836
rect 27759 3834 27765 3836
rect 27519 3782 27521 3834
rect 27701 3782 27703 3834
rect 27457 3780 27463 3782
rect 27519 3780 27543 3782
rect 27599 3780 27623 3782
rect 27679 3780 27703 3782
rect 27759 3780 27765 3782
rect 27457 3771 27765 3780
rect 27526 3088 27582 3097
rect 28092 3058 28120 4218
rect 27526 3023 27528 3032
rect 27580 3023 27582 3032
rect 27804 3052 27856 3058
rect 27528 2994 27580 3000
rect 27804 2994 27856 3000
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 27816 2961 27844 2994
rect 27802 2952 27858 2961
rect 27802 2887 27858 2896
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 26974 2615 27030 2624
rect 27160 2644 27212 2650
rect 26700 2576 26752 2582
rect 26884 2576 26936 2582
rect 26752 2536 26884 2564
rect 26700 2518 26752 2524
rect 26884 2518 26936 2524
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26988 2446 27016 2615
rect 27160 2586 27212 2592
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27068 2440 27120 2446
rect 27356 2428 27384 2790
rect 27457 2748 27765 2757
rect 27457 2746 27463 2748
rect 27519 2746 27543 2748
rect 27599 2746 27623 2748
rect 27679 2746 27703 2748
rect 27759 2746 27765 2748
rect 27519 2694 27521 2746
rect 27701 2694 27703 2746
rect 27457 2692 27463 2694
rect 27519 2692 27543 2694
rect 27599 2692 27623 2694
rect 27679 2692 27703 2694
rect 27759 2692 27765 2694
rect 27457 2683 27765 2692
rect 27528 2440 27580 2446
rect 27068 2382 27120 2388
rect 27158 2408 27214 2417
rect 26516 2304 26568 2310
rect 26620 2281 26648 2382
rect 26792 2304 26844 2310
rect 26516 2246 26568 2252
rect 26606 2272 26662 2281
rect 26240 2032 26292 2038
rect 26240 1974 26292 1980
rect 25872 1964 25924 1970
rect 25792 1924 25872 1952
rect 25872 1906 25924 1912
rect 26240 1828 26292 1834
rect 26240 1770 26292 1776
rect 26148 1760 26200 1766
rect 25884 1720 26148 1748
rect 25688 1352 25740 1358
rect 25688 1294 25740 1300
rect 25884 160 25912 1720
rect 26148 1702 26200 1708
rect 26148 1556 26200 1562
rect 26068 1516 26148 1544
rect 26068 490 26096 1516
rect 26148 1498 26200 1504
rect 26252 1358 26280 1770
rect 26528 1358 26556 2246
rect 26792 2246 26844 2252
rect 26606 2207 26662 2216
rect 26804 2106 26832 2246
rect 26792 2100 26844 2106
rect 26792 2042 26844 2048
rect 26976 2100 27028 2106
rect 26976 2042 27028 2048
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 26516 1352 26568 1358
rect 26516 1294 26568 1300
rect 26148 1216 26200 1222
rect 26884 1216 26936 1222
rect 26148 1158 26200 1164
rect 26436 1176 26884 1204
rect 26160 678 26188 1158
rect 26148 672 26200 678
rect 26148 614 26200 620
rect 26068 462 26188 490
rect 26160 160 26188 462
rect 26436 160 26464 1176
rect 26884 1158 26936 1164
rect 26988 898 27016 2042
rect 26712 870 27016 898
rect 26712 160 26740 870
rect 27080 762 27108 2382
rect 27356 2400 27528 2428
rect 27528 2382 27580 2388
rect 27620 2440 27672 2446
rect 27816 2428 27844 2790
rect 27894 2680 27950 2689
rect 28184 2650 28212 8502
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 35072 8492 35124 8498
rect 35072 8434 35124 8440
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 40500 8492 40552 8498
rect 40500 8434 40552 8440
rect 42892 8492 42944 8498
rect 42892 8434 42944 8440
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28368 3058 28396 3878
rect 28736 3194 28764 8434
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 30104 3120 30156 3126
rect 30104 3062 30156 3068
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 29460 2916 29512 2922
rect 29512 2876 29776 2904
rect 29460 2858 29512 2864
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 27894 2615 27896 2624
rect 27948 2615 27950 2624
rect 28172 2644 28224 2650
rect 27896 2586 27948 2592
rect 28172 2586 28224 2592
rect 27672 2400 27844 2428
rect 28276 2502 28672 2530
rect 27620 2382 27672 2388
rect 27158 2343 27160 2352
rect 27212 2343 27214 2352
rect 27160 2314 27212 2320
rect 27896 2304 27948 2310
rect 27896 2246 27948 2252
rect 27804 1828 27856 1834
rect 27804 1770 27856 1776
rect 27344 1760 27396 1766
rect 27344 1702 27396 1708
rect 27356 1358 27384 1702
rect 27457 1660 27765 1669
rect 27457 1658 27463 1660
rect 27519 1658 27543 1660
rect 27599 1658 27623 1660
rect 27679 1658 27703 1660
rect 27759 1658 27765 1660
rect 27519 1606 27521 1658
rect 27701 1606 27703 1658
rect 27457 1604 27463 1606
rect 27519 1604 27543 1606
rect 27599 1604 27623 1606
rect 27679 1604 27703 1606
rect 27759 1604 27765 1606
rect 27457 1595 27765 1604
rect 27620 1488 27672 1494
rect 27448 1436 27620 1442
rect 27448 1430 27672 1436
rect 27448 1414 27660 1430
rect 27712 1420 27764 1426
rect 27344 1352 27396 1358
rect 27344 1294 27396 1300
rect 27158 1048 27214 1057
rect 27158 983 27214 992
rect 27172 882 27200 983
rect 27160 876 27212 882
rect 27160 818 27212 824
rect 26792 740 26844 746
rect 26792 682 26844 688
rect 26896 734 27108 762
rect 25318 54 25544 82
rect 25318 -300 25374 54
rect 25594 -300 25650 160
rect 25870 -300 25926 160
rect 26146 -300 26202 160
rect 26422 -300 26478 160
rect 26698 -300 26754 160
rect 26804 134 26832 682
rect 26896 338 26924 734
rect 27448 626 27476 1414
rect 27712 1362 27764 1368
rect 27724 1306 27752 1362
rect 26988 598 27476 626
rect 27540 1278 27752 1306
rect 26884 332 26936 338
rect 26884 274 26936 280
rect 26988 160 27016 598
rect 27540 490 27568 1278
rect 27618 1184 27674 1193
rect 27618 1119 27674 1128
rect 27632 678 27660 1119
rect 27620 672 27672 678
rect 27620 614 27672 620
rect 27264 462 27568 490
rect 27264 160 27292 462
rect 27528 400 27580 406
rect 27528 342 27580 348
rect 27540 160 27568 342
rect 27816 160 27844 1770
rect 27908 1358 27936 2246
rect 28172 1964 28224 1970
rect 28092 1924 28172 1952
rect 27986 1456 28042 1465
rect 27986 1391 28042 1400
rect 27896 1352 27948 1358
rect 27896 1294 27948 1300
rect 28000 513 28028 1391
rect 27986 504 28042 513
rect 27986 439 28042 448
rect 28092 160 28120 1924
rect 28172 1906 28224 1912
rect 28276 241 28304 2502
rect 28644 2446 28672 2502
rect 28540 2440 28592 2446
rect 28460 2400 28540 2428
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28368 2106 28396 2246
rect 28356 2100 28408 2106
rect 28356 2042 28408 2048
rect 28460 377 28488 2400
rect 28540 2382 28592 2388
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 28632 1760 28684 1766
rect 28552 1720 28632 1748
rect 28446 368 28502 377
rect 28446 303 28502 312
rect 28262 232 28318 241
rect 28262 167 28318 176
rect 26792 128 26844 134
rect 26792 70 26844 76
rect 26974 -300 27030 160
rect 27250 -300 27306 160
rect 27526 -300 27582 160
rect 27802 -300 27858 160
rect 28078 -300 28134 160
rect 28354 82 28410 160
rect 28552 82 28580 1720
rect 28632 1702 28684 1708
rect 28354 54 28580 82
rect 28630 82 28686 160
rect 28736 82 28764 2790
rect 29366 2544 29422 2553
rect 29366 2479 29422 2488
rect 29380 2446 29408 2479
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 29184 2304 29236 2310
rect 29644 2304 29696 2310
rect 29184 2246 29236 2252
rect 29380 2264 29644 2292
rect 28828 1358 28856 2246
rect 28920 2106 28948 2246
rect 29196 2106 29224 2246
rect 29274 2136 29330 2145
rect 28908 2100 28960 2106
rect 28908 2042 28960 2048
rect 29184 2100 29236 2106
rect 29274 2071 29330 2080
rect 29184 2042 29236 2048
rect 29288 1902 29316 2071
rect 29276 1896 29328 1902
rect 29276 1838 29328 1844
rect 29092 1488 29144 1494
rect 28920 1436 29092 1442
rect 28920 1430 29144 1436
rect 28920 1414 29132 1430
rect 28816 1352 28868 1358
rect 28816 1294 28868 1300
rect 28920 160 28948 1414
rect 29000 1352 29052 1358
rect 29000 1294 29052 1300
rect 29012 649 29040 1294
rect 28998 640 29054 649
rect 28998 575 29054 584
rect 28630 54 28764 82
rect 28354 -300 28410 54
rect 28630 -300 28686 54
rect 28906 -300 28962 160
rect 29182 82 29238 160
rect 29380 82 29408 2264
rect 29644 2246 29696 2252
rect 29748 2038 29776 2876
rect 29736 2032 29788 2038
rect 29736 1974 29788 1980
rect 29460 1964 29512 1970
rect 29460 1906 29512 1912
rect 29472 1562 29500 1906
rect 29644 1760 29696 1766
rect 29564 1720 29644 1748
rect 29460 1556 29512 1562
rect 29460 1498 29512 1504
rect 29564 1494 29592 1720
rect 29644 1702 29696 1708
rect 29552 1488 29604 1494
rect 29552 1430 29604 1436
rect 29644 1488 29696 1494
rect 29644 1430 29696 1436
rect 29182 54 29408 82
rect 29458 82 29514 160
rect 29656 82 29684 1430
rect 30116 1358 30144 3062
rect 30208 2825 30236 3402
rect 30748 2848 30800 2854
rect 30194 2816 30250 2825
rect 30748 2790 30800 2796
rect 30194 2751 30250 2760
rect 30194 2680 30250 2689
rect 30194 2615 30196 2624
rect 30248 2615 30250 2624
rect 30196 2586 30248 2592
rect 30656 2304 30708 2310
rect 30194 2272 30250 2281
rect 30194 2207 30250 2216
rect 30576 2264 30656 2292
rect 30208 2038 30236 2207
rect 30196 2032 30248 2038
rect 30196 1974 30248 1980
rect 30472 1760 30524 1766
rect 30208 1720 30472 1748
rect 30104 1352 30156 1358
rect 30104 1294 30156 1300
rect 29736 264 29788 270
rect 29736 206 29788 212
rect 29748 160 29776 206
rect 29458 54 29684 82
rect 29182 -300 29238 54
rect 29458 -300 29514 54
rect 29734 -300 29790 160
rect 30010 82 30066 160
rect 30208 82 30236 1720
rect 30472 1702 30524 1708
rect 30472 1420 30524 1426
rect 30472 1362 30524 1368
rect 30288 1216 30340 1222
rect 30288 1158 30340 1164
rect 30300 406 30328 1158
rect 30288 400 30340 406
rect 30288 342 30340 348
rect 30010 54 30236 82
rect 30286 82 30342 160
rect 30484 82 30512 1362
rect 30576 160 30604 2264
rect 30656 2246 30708 2252
rect 30760 2106 30788 2790
rect 30852 2650 30880 8434
rect 32758 7644 33066 7653
rect 32758 7642 32764 7644
rect 32820 7642 32844 7644
rect 32900 7642 32924 7644
rect 32980 7642 33004 7644
rect 33060 7642 33066 7644
rect 32820 7590 32822 7642
rect 33002 7590 33004 7642
rect 32758 7588 32764 7590
rect 32820 7588 32844 7590
rect 32900 7588 32924 7590
rect 32980 7588 33004 7590
rect 33060 7588 33066 7590
rect 32758 7579 33066 7588
rect 32758 6556 33066 6565
rect 32758 6554 32764 6556
rect 32820 6554 32844 6556
rect 32900 6554 32924 6556
rect 32980 6554 33004 6556
rect 33060 6554 33066 6556
rect 32820 6502 32822 6554
rect 33002 6502 33004 6554
rect 32758 6500 32764 6502
rect 32820 6500 32844 6502
rect 32900 6500 32924 6502
rect 32980 6500 33004 6502
rect 33060 6500 33066 6502
rect 32758 6491 33066 6500
rect 32758 5468 33066 5477
rect 32758 5466 32764 5468
rect 32820 5466 32844 5468
rect 32900 5466 32924 5468
rect 32980 5466 33004 5468
rect 33060 5466 33066 5468
rect 32820 5414 32822 5466
rect 33002 5414 33004 5466
rect 32758 5412 32764 5414
rect 32820 5412 32844 5414
rect 32900 5412 32924 5414
rect 32980 5412 33004 5414
rect 33060 5412 33066 5414
rect 32758 5403 33066 5412
rect 32758 4380 33066 4389
rect 32758 4378 32764 4380
rect 32820 4378 32844 4380
rect 32900 4378 32924 4380
rect 32980 4378 33004 4380
rect 33060 4378 33066 4380
rect 32820 4326 32822 4378
rect 33002 4326 33004 4378
rect 32758 4324 32764 4326
rect 32820 4324 32844 4326
rect 32900 4324 32924 4326
rect 32980 4324 33004 4326
rect 33060 4324 33066 4326
rect 32758 4315 33066 4324
rect 32758 3292 33066 3301
rect 32758 3290 32764 3292
rect 32820 3290 32844 3292
rect 32900 3290 32924 3292
rect 32980 3290 33004 3292
rect 33060 3290 33066 3292
rect 32820 3238 32822 3290
rect 33002 3238 33004 3290
rect 32758 3236 32764 3238
rect 32820 3236 32844 3238
rect 32900 3236 32924 3238
rect 32980 3236 33004 3238
rect 33060 3236 33066 3238
rect 31482 3224 31538 3233
rect 32758 3227 33066 3236
rect 31482 3159 31538 3168
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 30748 2100 30800 2106
rect 30748 2042 30800 2048
rect 30840 1556 30892 1562
rect 30840 1498 30892 1504
rect 30748 1284 30800 1290
rect 30748 1226 30800 1232
rect 30760 474 30788 1226
rect 30748 468 30800 474
rect 30748 410 30800 416
rect 30852 160 30880 1498
rect 31036 1494 31064 2382
rect 31206 2136 31262 2145
rect 31312 2106 31340 2382
rect 31206 2071 31262 2080
rect 31300 2100 31352 2106
rect 31220 1970 31248 2071
rect 31300 2042 31352 2048
rect 31208 1964 31260 1970
rect 31208 1906 31260 1912
rect 31404 1850 31432 2382
rect 31496 1902 31524 3159
rect 33244 2650 33272 8434
rect 33322 4584 33378 4593
rect 33322 4519 33378 4528
rect 33232 2644 33284 2650
rect 33232 2586 33284 2592
rect 33336 2446 33364 4519
rect 35084 2650 35112 8434
rect 36820 3596 36872 3602
rect 36740 3556 36820 3584
rect 35714 2952 35770 2961
rect 35714 2887 35770 2896
rect 35162 2680 35218 2689
rect 35072 2644 35124 2650
rect 35162 2615 35218 2624
rect 35072 2586 35124 2592
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 32758 2204 33066 2213
rect 32758 2202 32764 2204
rect 32820 2202 32844 2204
rect 32900 2202 32924 2204
rect 32980 2202 33004 2204
rect 33060 2202 33066 2204
rect 32820 2150 32822 2202
rect 33002 2150 33004 2202
rect 32758 2148 32764 2150
rect 32820 2148 32844 2150
rect 32900 2148 32924 2150
rect 32980 2148 33004 2150
rect 33060 2148 33066 2150
rect 32758 2139 33066 2148
rect 32048 2094 32352 2122
rect 31944 1964 31996 1970
rect 31944 1906 31996 1912
rect 31220 1822 31432 1850
rect 31484 1896 31536 1902
rect 31484 1838 31536 1844
rect 31668 1828 31720 1834
rect 31024 1488 31076 1494
rect 31024 1430 31076 1436
rect 30932 1284 30984 1290
rect 30932 1226 30984 1232
rect 30944 678 30972 1226
rect 31220 882 31248 1822
rect 31668 1770 31720 1776
rect 31576 1760 31628 1766
rect 31312 1720 31576 1748
rect 31208 876 31260 882
rect 31208 818 31260 824
rect 30932 672 30984 678
rect 30932 614 30984 620
rect 30286 54 30512 82
rect 30010 -300 30066 54
rect 30286 -300 30342 54
rect 30562 -300 30618 160
rect 30838 -300 30894 160
rect 31114 82 31170 160
rect 31312 82 31340 1720
rect 31576 1702 31628 1708
rect 31680 1442 31708 1770
rect 31956 1442 31984 1906
rect 31404 1414 31708 1442
rect 31864 1414 31984 1442
rect 31404 160 31432 1414
rect 31864 950 31892 1414
rect 31944 1352 31996 1358
rect 31944 1294 31996 1300
rect 31852 944 31904 950
rect 31956 921 31984 1294
rect 31852 886 31904 892
rect 31942 912 31998 921
rect 31942 847 31998 856
rect 32048 762 32076 2094
rect 32324 2038 32352 2094
rect 32588 2100 32640 2106
rect 32588 2042 32640 2048
rect 32312 2032 32364 2038
rect 32312 1974 32364 1980
rect 32496 1760 32548 1766
rect 32416 1720 32496 1748
rect 32220 1284 32272 1290
rect 32220 1226 32272 1232
rect 32312 1284 32364 1290
rect 32312 1226 32364 1232
rect 32128 1216 32180 1222
rect 32128 1158 32180 1164
rect 31956 734 32076 762
rect 31668 468 31720 474
rect 31668 410 31720 416
rect 31680 160 31708 410
rect 31956 160 31984 734
rect 32140 678 32168 1158
rect 32232 746 32260 1226
rect 32324 1018 32352 1226
rect 32312 1012 32364 1018
rect 32312 954 32364 960
rect 32220 740 32272 746
rect 32220 682 32272 688
rect 32128 672 32180 678
rect 32128 614 32180 620
rect 31114 54 31340 82
rect 31114 -300 31170 54
rect 31390 -300 31446 160
rect 31666 -300 31722 160
rect 31942 -300 31998 160
rect 32218 82 32274 160
rect 32416 82 32444 1720
rect 32496 1702 32548 1708
rect 32496 1488 32548 1494
rect 32496 1430 32548 1436
rect 32508 270 32536 1430
rect 32600 785 32628 2042
rect 32956 1556 33008 1562
rect 32692 1516 32956 1544
rect 32586 776 32642 785
rect 32586 711 32642 720
rect 32496 264 32548 270
rect 32496 206 32548 212
rect 32218 54 32444 82
rect 32494 82 32550 160
rect 32692 82 32720 1516
rect 32956 1498 33008 1504
rect 33152 1494 33180 2382
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33324 1964 33376 1970
rect 33324 1906 33376 1912
rect 33336 1873 33364 1906
rect 33322 1864 33378 1873
rect 33322 1799 33378 1808
rect 33140 1488 33192 1494
rect 33140 1430 33192 1436
rect 32758 1116 33066 1125
rect 32758 1114 32764 1116
rect 32820 1114 32844 1116
rect 32900 1114 32924 1116
rect 32980 1114 33004 1116
rect 33060 1114 33066 1116
rect 32820 1062 32822 1114
rect 33002 1062 33004 1114
rect 32758 1060 32764 1062
rect 32820 1060 32844 1062
rect 32900 1060 32924 1062
rect 32980 1060 33004 1062
rect 33060 1060 33066 1062
rect 32758 1051 33066 1060
rect 32772 1012 32824 1018
rect 32772 954 32824 960
rect 32784 160 32812 954
rect 33048 944 33100 950
rect 33048 886 33100 892
rect 33060 160 33088 886
rect 32494 54 32720 82
rect 32218 -300 32274 54
rect 32494 -300 32550 54
rect 32770 -300 32826 160
rect 33046 -300 33102 160
rect 33322 82 33378 160
rect 33520 82 33548 2246
rect 34716 2106 34744 2382
rect 34704 2100 34756 2106
rect 34704 2042 34756 2048
rect 33874 2000 33930 2009
rect 33874 1935 33876 1944
rect 33928 1935 33930 1944
rect 33876 1906 33928 1912
rect 34244 1896 34296 1902
rect 34244 1838 34296 1844
rect 33600 1828 33652 1834
rect 33600 1770 33652 1776
rect 33612 160 33640 1770
rect 33968 1352 34020 1358
rect 33888 1312 33968 1340
rect 33888 160 33916 1312
rect 33968 1294 34020 1300
rect 34256 1034 34284 1838
rect 35176 1834 35204 2615
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 35452 2106 35480 2314
rect 35440 2100 35492 2106
rect 35440 2042 35492 2048
rect 35164 1828 35216 1834
rect 35164 1770 35216 1776
rect 34980 1556 35032 1562
rect 34980 1498 35032 1504
rect 34518 1320 34574 1329
rect 34428 1284 34480 1290
rect 34518 1255 34574 1264
rect 34428 1226 34480 1232
rect 34164 1006 34284 1034
rect 34164 160 34192 1006
rect 34440 160 34468 1226
rect 34532 1222 34560 1255
rect 34520 1216 34572 1222
rect 34888 1216 34940 1222
rect 34520 1158 34572 1164
rect 34808 1176 34888 1204
rect 34808 474 34836 1176
rect 34888 1158 34940 1164
rect 34992 1018 35020 1498
rect 35728 1494 35756 2887
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 36004 2106 36032 2382
rect 35992 2100 36044 2106
rect 35992 2042 36044 2048
rect 35808 1896 35860 1902
rect 35808 1838 35860 1844
rect 35716 1488 35768 1494
rect 35716 1430 35768 1436
rect 35164 1352 35216 1358
rect 35162 1320 35164 1329
rect 35216 1320 35218 1329
rect 35162 1255 35218 1264
rect 35716 1216 35768 1222
rect 35716 1158 35768 1164
rect 34980 1012 35032 1018
rect 34980 954 35032 960
rect 35348 672 35400 678
rect 35348 614 35400 620
rect 34888 604 34940 610
rect 34888 546 34940 552
rect 34796 468 34848 474
rect 34796 410 34848 416
rect 33322 54 33548 82
rect 33322 -300 33378 54
rect 33598 -300 33654 160
rect 33874 -300 33930 160
rect 34150 -300 34206 160
rect 34426 -300 34482 160
rect 34702 82 34758 160
rect 34900 82 34928 546
rect 35360 218 35388 614
rect 35728 218 35756 1158
rect 35176 190 35388 218
rect 35452 190 35756 218
rect 34702 54 34928 82
rect 34978 82 35034 160
rect 35176 82 35204 190
rect 34978 54 35204 82
rect 35254 82 35310 160
rect 35452 82 35480 190
rect 35820 160 35848 1838
rect 35900 1556 35952 1562
rect 35900 1498 35952 1504
rect 35912 950 35940 1498
rect 36268 1284 36320 1290
rect 36268 1226 36320 1232
rect 36280 1057 36308 1226
rect 36266 1048 36322 1057
rect 36084 1012 36136 1018
rect 36266 983 36322 992
rect 36084 954 36136 960
rect 35900 944 35952 950
rect 35900 886 35952 892
rect 36096 160 36124 954
rect 36372 160 36400 2790
rect 36740 2774 36768 3556
rect 36820 3538 36872 3544
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37200 3074 37228 3334
rect 37200 3046 37320 3074
rect 37188 2916 37240 2922
rect 36648 2746 36768 2774
rect 37108 2876 37188 2904
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 36464 1562 36492 2518
rect 36544 1964 36596 1970
rect 36544 1906 36596 1912
rect 36452 1556 36504 1562
rect 36452 1498 36504 1504
rect 36556 746 36584 1906
rect 36544 740 36596 746
rect 36544 682 36596 688
rect 36648 160 36676 2746
rect 36820 1352 36872 1358
rect 36820 1294 36872 1300
rect 36832 610 36860 1294
rect 36912 1216 36964 1222
rect 36912 1158 36964 1164
rect 36820 604 36872 610
rect 36820 546 36872 552
rect 36924 406 36952 1158
rect 36912 400 36964 406
rect 36912 342 36964 348
rect 35254 54 35480 82
rect 35530 82 35586 160
rect 35716 128 35768 134
rect 35530 76 35716 82
rect 35530 70 35768 76
rect 35530 54 35756 70
rect 34702 -300 34758 54
rect 34978 -300 35034 54
rect 35254 -300 35310 54
rect 35530 -300 35586 54
rect 35806 -300 35862 160
rect 36082 -300 36138 160
rect 36358 -300 36414 160
rect 36634 -300 36690 160
rect 36910 82 36966 160
rect 37108 82 37136 2876
rect 37188 2858 37240 2864
rect 37292 2802 37320 3046
rect 37200 2774 37320 2802
rect 37200 160 37228 2774
rect 37384 2650 37412 8434
rect 38060 8188 38368 8197
rect 38060 8186 38066 8188
rect 38122 8186 38146 8188
rect 38202 8186 38226 8188
rect 38282 8186 38306 8188
rect 38362 8186 38368 8188
rect 38122 8134 38124 8186
rect 38304 8134 38306 8186
rect 38060 8132 38066 8134
rect 38122 8132 38146 8134
rect 38202 8132 38226 8134
rect 38282 8132 38306 8134
rect 38362 8132 38368 8134
rect 38060 8123 38368 8132
rect 38060 7100 38368 7109
rect 38060 7098 38066 7100
rect 38122 7098 38146 7100
rect 38202 7098 38226 7100
rect 38282 7098 38306 7100
rect 38362 7098 38368 7100
rect 38122 7046 38124 7098
rect 38304 7046 38306 7098
rect 38060 7044 38066 7046
rect 38122 7044 38146 7046
rect 38202 7044 38226 7046
rect 38282 7044 38306 7046
rect 38362 7044 38368 7046
rect 38060 7035 38368 7044
rect 38060 6012 38368 6021
rect 38060 6010 38066 6012
rect 38122 6010 38146 6012
rect 38202 6010 38226 6012
rect 38282 6010 38306 6012
rect 38362 6010 38368 6012
rect 38122 5958 38124 6010
rect 38304 5958 38306 6010
rect 38060 5956 38066 5958
rect 38122 5956 38146 5958
rect 38202 5956 38226 5958
rect 38282 5956 38306 5958
rect 38362 5956 38368 5958
rect 38060 5947 38368 5956
rect 38060 4924 38368 4933
rect 38060 4922 38066 4924
rect 38122 4922 38146 4924
rect 38202 4922 38226 4924
rect 38282 4922 38306 4924
rect 38362 4922 38368 4924
rect 38122 4870 38124 4922
rect 38304 4870 38306 4922
rect 38060 4868 38066 4870
rect 38122 4868 38146 4870
rect 38202 4868 38226 4870
rect 38282 4868 38306 4870
rect 38362 4868 38368 4870
rect 38060 4859 38368 4868
rect 38060 3836 38368 3845
rect 38060 3834 38066 3836
rect 38122 3834 38146 3836
rect 38202 3834 38226 3836
rect 38282 3834 38306 3836
rect 38362 3834 38368 3836
rect 38122 3782 38124 3834
rect 38304 3782 38306 3834
rect 38060 3780 38066 3782
rect 38122 3780 38146 3782
rect 38202 3780 38226 3782
rect 38282 3780 38306 3782
rect 38362 3780 38368 3782
rect 38060 3771 38368 3780
rect 37462 3632 37518 3641
rect 37462 3567 37518 3576
rect 38936 3596 38988 3602
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 37476 1358 37504 3567
rect 38936 3538 38988 3544
rect 38476 3528 38528 3534
rect 38476 3470 38528 3476
rect 37832 3460 37884 3466
rect 37832 3402 37884 3408
rect 37556 3188 37608 3194
rect 37556 3130 37608 3136
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 36910 54 37136 82
rect 36910 -300 36966 54
rect 37186 -300 37242 160
rect 37462 82 37518 160
rect 37568 82 37596 3130
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37752 2106 37780 2382
rect 37740 2100 37792 2106
rect 37740 2042 37792 2048
rect 37648 1964 37700 1970
rect 37648 1906 37700 1912
rect 37660 1562 37688 1906
rect 37648 1556 37700 1562
rect 37648 1498 37700 1504
rect 37844 1442 37872 3402
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38028 2836 38056 3062
rect 38384 2984 38436 2990
rect 38384 2926 38436 2932
rect 37752 1414 37872 1442
rect 37936 2808 38056 2836
rect 37648 1352 37700 1358
rect 37648 1294 37700 1300
rect 37660 678 37688 1294
rect 37648 672 37700 678
rect 37648 614 37700 620
rect 37752 160 37780 1414
rect 37832 1216 37884 1222
rect 37832 1158 37884 1164
rect 37844 338 37872 1158
rect 37832 332 37884 338
rect 37832 274 37884 280
rect 37462 54 37596 82
rect 37462 -300 37518 54
rect 37738 -300 37794 160
rect 37936 82 37964 2808
rect 38060 2748 38368 2757
rect 38060 2746 38066 2748
rect 38122 2746 38146 2748
rect 38202 2746 38226 2748
rect 38282 2746 38306 2748
rect 38362 2746 38368 2748
rect 38122 2694 38124 2746
rect 38304 2694 38306 2746
rect 38060 2692 38066 2694
rect 38122 2692 38146 2694
rect 38202 2692 38226 2694
rect 38282 2692 38306 2694
rect 38362 2692 38368 2694
rect 38060 2683 38368 2692
rect 38060 1660 38368 1669
rect 38060 1658 38066 1660
rect 38122 1658 38146 1660
rect 38202 1658 38226 1660
rect 38282 1658 38306 1660
rect 38362 1658 38368 1660
rect 38122 1606 38124 1658
rect 38304 1606 38306 1658
rect 38060 1604 38066 1606
rect 38122 1604 38146 1606
rect 38202 1604 38226 1606
rect 38282 1604 38306 1606
rect 38362 1604 38368 1606
rect 38060 1595 38368 1604
rect 38396 1562 38424 2926
rect 38384 1556 38436 1562
rect 38384 1498 38436 1504
rect 38108 1352 38160 1358
rect 38108 1294 38160 1300
rect 38384 1352 38436 1358
rect 38384 1294 38436 1300
rect 38014 82 38070 160
rect 38120 134 38148 1294
rect 38396 1018 38424 1294
rect 38384 1012 38436 1018
rect 38384 954 38436 960
rect 37936 54 38070 82
rect 38108 128 38160 134
rect 38108 70 38160 76
rect 38290 82 38346 160
rect 38488 82 38516 3470
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 38580 160 38608 2994
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 1358 38700 2790
rect 38948 1358 38976 3538
rect 39212 2916 39264 2922
rect 39212 2858 39264 2864
rect 39224 1358 39252 2858
rect 39316 2650 39344 8434
rect 40316 3460 40368 3466
rect 40316 3402 40368 3408
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39304 2644 39356 2650
rect 39304 2586 39356 2592
rect 39396 2440 39448 2446
rect 39302 2408 39358 2417
rect 39396 2382 39448 2388
rect 39302 2343 39358 2352
rect 38660 1352 38712 1358
rect 38660 1294 38712 1300
rect 38936 1352 38988 1358
rect 38936 1294 38988 1300
rect 39212 1352 39264 1358
rect 39212 1294 39264 1300
rect 39316 1222 39344 2343
rect 39408 2106 39436 2382
rect 39396 2100 39448 2106
rect 39396 2042 39448 2048
rect 39500 1358 39528 3334
rect 40040 3188 40092 3194
rect 40040 3130 40092 3136
rect 39670 3088 39726 3097
rect 39670 3023 39726 3032
rect 39580 1420 39632 1426
rect 39580 1362 39632 1368
rect 39488 1352 39540 1358
rect 39488 1294 39540 1300
rect 38660 1216 38712 1222
rect 38660 1158 38712 1164
rect 38844 1216 38896 1222
rect 38844 1158 38896 1164
rect 39120 1216 39172 1222
rect 39120 1158 39172 1164
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 38672 542 38700 1158
rect 38660 536 38712 542
rect 38856 513 38884 1158
rect 39132 814 39160 1158
rect 39120 808 39172 814
rect 39592 762 39620 1362
rect 39684 1222 39712 3023
rect 40052 1358 40080 3130
rect 40132 1964 40184 1970
rect 40132 1906 40184 1912
rect 40144 1562 40172 1906
rect 40132 1556 40184 1562
rect 40132 1498 40184 1504
rect 40328 1358 40356 3402
rect 40512 2650 40540 8434
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 40592 3120 40644 3126
rect 40592 3062 40644 3068
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 40604 1358 40632 3062
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 40696 2106 40724 2382
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 40880 1358 40908 3470
rect 41144 3052 41196 3058
rect 41144 2994 41196 3000
rect 40960 2032 41012 2038
rect 40960 1974 41012 1980
rect 40972 1494 41000 1974
rect 40960 1488 41012 1494
rect 40960 1430 41012 1436
rect 41156 1358 41184 2994
rect 42904 2650 42932 8434
rect 43361 7644 43669 7653
rect 43361 7642 43367 7644
rect 43423 7642 43447 7644
rect 43503 7642 43527 7644
rect 43583 7642 43607 7644
rect 43663 7642 43669 7644
rect 43423 7590 43425 7642
rect 43605 7590 43607 7642
rect 43361 7588 43367 7590
rect 43423 7588 43447 7590
rect 43503 7588 43527 7590
rect 43583 7588 43607 7590
rect 43663 7588 43669 7590
rect 43361 7579 43669 7588
rect 43361 6556 43669 6565
rect 43361 6554 43367 6556
rect 43423 6554 43447 6556
rect 43503 6554 43527 6556
rect 43583 6554 43607 6556
rect 43663 6554 43669 6556
rect 43423 6502 43425 6554
rect 43605 6502 43607 6554
rect 43361 6500 43367 6502
rect 43423 6500 43447 6502
rect 43503 6500 43527 6502
rect 43583 6500 43607 6502
rect 43663 6500 43669 6502
rect 43361 6491 43669 6500
rect 43361 5468 43669 5477
rect 43361 5466 43367 5468
rect 43423 5466 43447 5468
rect 43503 5466 43527 5468
rect 43583 5466 43607 5468
rect 43663 5466 43669 5468
rect 43423 5414 43425 5466
rect 43605 5414 43607 5466
rect 43361 5412 43367 5414
rect 43423 5412 43447 5414
rect 43503 5412 43527 5414
rect 43583 5412 43607 5414
rect 43663 5412 43669 5414
rect 43361 5403 43669 5412
rect 43361 4380 43669 4389
rect 43361 4378 43367 4380
rect 43423 4378 43447 4380
rect 43503 4378 43527 4380
rect 43583 4378 43607 4380
rect 43663 4378 43669 4380
rect 43423 4326 43425 4378
rect 43605 4326 43607 4378
rect 43361 4324 43367 4326
rect 43423 4324 43447 4326
rect 43503 4324 43527 4326
rect 43583 4324 43607 4326
rect 43663 4324 43669 4326
rect 43361 4315 43669 4324
rect 43361 3292 43669 3301
rect 43361 3290 43367 3292
rect 43423 3290 43447 3292
rect 43503 3290 43527 3292
rect 43583 3290 43607 3292
rect 43663 3290 43669 3292
rect 43423 3238 43425 3290
rect 43605 3238 43607 3290
rect 43361 3236 43367 3238
rect 43423 3236 43447 3238
rect 43503 3236 43527 3238
rect 43583 3236 43607 3238
rect 43663 3236 43669 3238
rect 43361 3227 43669 3236
rect 42892 2644 42944 2650
rect 42892 2586 42944 2592
rect 42616 2440 42668 2446
rect 42616 2382 42668 2388
rect 42628 2106 42656 2382
rect 43361 2204 43669 2213
rect 43361 2202 43367 2204
rect 43423 2202 43447 2204
rect 43503 2202 43527 2204
rect 43583 2202 43607 2204
rect 43663 2202 43669 2204
rect 43423 2150 43425 2202
rect 43605 2150 43607 2202
rect 43361 2148 43367 2150
rect 43423 2148 43447 2150
rect 43503 2148 43527 2150
rect 43583 2148 43607 2150
rect 43663 2148 43669 2150
rect 43361 2139 43669 2148
rect 42616 2100 42668 2106
rect 42616 2042 42668 2048
rect 41788 1964 41840 1970
rect 41788 1906 41840 1912
rect 41236 1896 41288 1902
rect 41236 1838 41288 1844
rect 41248 1494 41276 1838
rect 41800 1562 41828 1906
rect 41788 1556 41840 1562
rect 41788 1498 41840 1504
rect 41236 1488 41288 1494
rect 41236 1430 41288 1436
rect 40040 1352 40092 1358
rect 40040 1294 40092 1300
rect 40316 1352 40368 1358
rect 40316 1294 40368 1300
rect 40592 1352 40644 1358
rect 40592 1294 40644 1300
rect 40868 1352 40920 1358
rect 40868 1294 40920 1300
rect 41144 1352 41196 1358
rect 41144 1294 41196 1300
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 41696 1352 41748 1358
rect 41696 1294 41748 1300
rect 39672 1216 39724 1222
rect 39672 1158 39724 1164
rect 40132 1216 40184 1222
rect 40132 1158 40184 1164
rect 40684 1216 40736 1222
rect 40684 1158 40736 1164
rect 40144 1018 40172 1158
rect 40132 1012 40184 1018
rect 40132 954 40184 960
rect 39120 750 39172 756
rect 39408 734 39620 762
rect 40696 746 40724 1158
rect 40684 740 40736 746
rect 39212 536 39264 542
rect 38660 478 38712 484
rect 38842 504 38898 513
rect 38842 439 38898 448
rect 39132 496 39212 524
rect 38844 400 38896 406
rect 38844 342 38896 348
rect 38856 160 38884 342
rect 39132 160 39160 496
rect 39212 478 39264 484
rect 39408 160 39436 734
rect 40684 682 40736 688
rect 41432 406 41460 1294
rect 41708 542 41736 1294
rect 43361 1116 43669 1125
rect 43361 1114 43367 1116
rect 43423 1114 43447 1116
rect 43503 1114 43527 1116
rect 43583 1114 43607 1116
rect 43663 1114 43669 1116
rect 43423 1062 43425 1114
rect 43605 1062 43607 1114
rect 43361 1060 43367 1062
rect 43423 1060 43447 1062
rect 43503 1060 43527 1062
rect 43583 1060 43607 1062
rect 43663 1060 43669 1062
rect 43361 1051 43669 1060
rect 41696 536 41748 542
rect 41696 478 41748 484
rect 41420 400 41472 406
rect 41420 342 41472 348
rect 38014 -300 38070 54
rect 38290 54 38516 82
rect 38290 -300 38346 54
rect 38566 -300 38622 160
rect 38842 -300 38898 160
rect 39118 -300 39174 160
rect 39394 -300 39450 160
<< via2 >>
rect 11558 8730 11614 8732
rect 11638 8730 11694 8732
rect 11718 8730 11774 8732
rect 11798 8730 11854 8732
rect 11558 8678 11604 8730
rect 11604 8678 11614 8730
rect 11638 8678 11668 8730
rect 11668 8678 11680 8730
rect 11680 8678 11694 8730
rect 11718 8678 11732 8730
rect 11732 8678 11744 8730
rect 11744 8678 11774 8730
rect 11798 8678 11808 8730
rect 11808 8678 11854 8730
rect 11558 8676 11614 8678
rect 11638 8676 11694 8678
rect 11718 8676 11774 8678
rect 11798 8676 11854 8678
rect 22161 8730 22217 8732
rect 22241 8730 22297 8732
rect 22321 8730 22377 8732
rect 22401 8730 22457 8732
rect 22161 8678 22207 8730
rect 22207 8678 22217 8730
rect 22241 8678 22271 8730
rect 22271 8678 22283 8730
rect 22283 8678 22297 8730
rect 22321 8678 22335 8730
rect 22335 8678 22347 8730
rect 22347 8678 22377 8730
rect 22401 8678 22411 8730
rect 22411 8678 22457 8730
rect 22161 8676 22217 8678
rect 22241 8676 22297 8678
rect 22321 8676 22377 8678
rect 22401 8676 22457 8678
rect 9586 8492 9642 8528
rect 9586 8472 9588 8492
rect 9588 8472 9640 8492
rect 9640 8472 9642 8492
rect 2226 8356 2282 8392
rect 2226 8336 2228 8356
rect 2228 8336 2280 8356
rect 2280 8336 2282 8356
rect 6257 8186 6313 8188
rect 6337 8186 6393 8188
rect 6417 8186 6473 8188
rect 6497 8186 6553 8188
rect 6257 8134 6303 8186
rect 6303 8134 6313 8186
rect 6337 8134 6367 8186
rect 6367 8134 6379 8186
rect 6379 8134 6393 8186
rect 6417 8134 6431 8186
rect 6431 8134 6443 8186
rect 6443 8134 6473 8186
rect 6497 8134 6507 8186
rect 6507 8134 6553 8186
rect 6257 8132 6313 8134
rect 6337 8132 6393 8134
rect 6417 8132 6473 8134
rect 6497 8132 6553 8134
rect 11558 7642 11614 7644
rect 11638 7642 11694 7644
rect 11718 7642 11774 7644
rect 11798 7642 11854 7644
rect 11558 7590 11604 7642
rect 11604 7590 11614 7642
rect 11638 7590 11668 7642
rect 11668 7590 11680 7642
rect 11680 7590 11694 7642
rect 11718 7590 11732 7642
rect 11732 7590 11744 7642
rect 11744 7590 11774 7642
rect 11798 7590 11808 7642
rect 11808 7590 11854 7642
rect 11558 7588 11614 7590
rect 11638 7588 11694 7590
rect 11718 7588 11774 7590
rect 11798 7588 11854 7590
rect 6257 7098 6313 7100
rect 6337 7098 6393 7100
rect 6417 7098 6473 7100
rect 6497 7098 6553 7100
rect 6257 7046 6303 7098
rect 6303 7046 6313 7098
rect 6337 7046 6367 7098
rect 6367 7046 6379 7098
rect 6379 7046 6393 7098
rect 6417 7046 6431 7098
rect 6431 7046 6443 7098
rect 6443 7046 6473 7098
rect 6497 7046 6507 7098
rect 6507 7046 6553 7098
rect 6257 7044 6313 7046
rect 6337 7044 6393 7046
rect 6417 7044 6473 7046
rect 6497 7044 6553 7046
rect 11558 6554 11614 6556
rect 11638 6554 11694 6556
rect 11718 6554 11774 6556
rect 11798 6554 11854 6556
rect 11558 6502 11604 6554
rect 11604 6502 11614 6554
rect 11638 6502 11668 6554
rect 11668 6502 11680 6554
rect 11680 6502 11694 6554
rect 11718 6502 11732 6554
rect 11732 6502 11744 6554
rect 11744 6502 11774 6554
rect 11798 6502 11808 6554
rect 11808 6502 11854 6554
rect 11558 6500 11614 6502
rect 11638 6500 11694 6502
rect 11718 6500 11774 6502
rect 11798 6500 11854 6502
rect 6257 6010 6313 6012
rect 6337 6010 6393 6012
rect 6417 6010 6473 6012
rect 6497 6010 6553 6012
rect 6257 5958 6303 6010
rect 6303 5958 6313 6010
rect 6337 5958 6367 6010
rect 6367 5958 6379 6010
rect 6379 5958 6393 6010
rect 6417 5958 6431 6010
rect 6431 5958 6443 6010
rect 6443 5958 6473 6010
rect 6497 5958 6507 6010
rect 6507 5958 6553 6010
rect 6257 5956 6313 5958
rect 6337 5956 6393 5958
rect 6417 5956 6473 5958
rect 6497 5956 6553 5958
rect 11558 5466 11614 5468
rect 11638 5466 11694 5468
rect 11718 5466 11774 5468
rect 11798 5466 11854 5468
rect 11558 5414 11604 5466
rect 11604 5414 11614 5466
rect 11638 5414 11668 5466
rect 11668 5414 11680 5466
rect 11680 5414 11694 5466
rect 11718 5414 11732 5466
rect 11732 5414 11744 5466
rect 11744 5414 11774 5466
rect 11798 5414 11808 5466
rect 11808 5414 11854 5466
rect 11558 5412 11614 5414
rect 11638 5412 11694 5414
rect 11718 5412 11774 5414
rect 11798 5412 11854 5414
rect 6257 4922 6313 4924
rect 6337 4922 6393 4924
rect 6417 4922 6473 4924
rect 6497 4922 6553 4924
rect 6257 4870 6303 4922
rect 6303 4870 6313 4922
rect 6337 4870 6367 4922
rect 6367 4870 6379 4922
rect 6379 4870 6393 4922
rect 6417 4870 6431 4922
rect 6431 4870 6443 4922
rect 6443 4870 6473 4922
rect 6497 4870 6507 4922
rect 6507 4870 6553 4922
rect 6257 4868 6313 4870
rect 6337 4868 6393 4870
rect 6417 4868 6473 4870
rect 6497 4868 6553 4870
rect 6734 4120 6790 4176
rect 6257 3834 6313 3836
rect 6337 3834 6393 3836
rect 6417 3834 6473 3836
rect 6497 3834 6553 3836
rect 6257 3782 6303 3834
rect 6303 3782 6313 3834
rect 6337 3782 6367 3834
rect 6367 3782 6379 3834
rect 6379 3782 6393 3834
rect 6417 3782 6431 3834
rect 6431 3782 6443 3834
rect 6443 3782 6473 3834
rect 6497 3782 6507 3834
rect 6507 3782 6553 3834
rect 6257 3780 6313 3782
rect 6337 3780 6393 3782
rect 6417 3780 6473 3782
rect 6497 3780 6553 3782
rect 6257 2746 6313 2748
rect 6337 2746 6393 2748
rect 6417 2746 6473 2748
rect 6497 2746 6553 2748
rect 6257 2694 6303 2746
rect 6303 2694 6313 2746
rect 6337 2694 6367 2746
rect 6367 2694 6379 2746
rect 6379 2694 6393 2746
rect 6417 2694 6431 2746
rect 6431 2694 6443 2746
rect 6443 2694 6473 2746
rect 6497 2694 6507 2746
rect 6507 2694 6553 2746
rect 6257 2692 6313 2694
rect 6337 2692 6393 2694
rect 6417 2692 6473 2694
rect 6497 2692 6553 2694
rect 6257 1658 6313 1660
rect 6337 1658 6393 1660
rect 6417 1658 6473 1660
rect 6497 1658 6553 1660
rect 6257 1606 6303 1658
rect 6303 1606 6313 1658
rect 6337 1606 6367 1658
rect 6367 1606 6379 1658
rect 6379 1606 6393 1658
rect 6417 1606 6431 1658
rect 6431 1606 6443 1658
rect 6443 1606 6473 1658
rect 6497 1606 6507 1658
rect 6507 1606 6553 1658
rect 6257 1604 6313 1606
rect 6337 1604 6393 1606
rect 6417 1604 6473 1606
rect 6497 1604 6553 1606
rect 8206 3984 8262 4040
rect 9034 1944 9090 2000
rect 8942 1808 8998 1864
rect 11558 4378 11614 4380
rect 11638 4378 11694 4380
rect 11718 4378 11774 4380
rect 11798 4378 11854 4380
rect 11558 4326 11604 4378
rect 11604 4326 11614 4378
rect 11638 4326 11668 4378
rect 11668 4326 11680 4378
rect 11680 4326 11694 4378
rect 11718 4326 11732 4378
rect 11732 4326 11744 4378
rect 11744 4326 11774 4378
rect 11798 4326 11808 4378
rect 11808 4326 11854 4378
rect 11558 4324 11614 4326
rect 11638 4324 11694 4326
rect 11718 4324 11774 4326
rect 11798 4324 11854 4326
rect 11558 3290 11614 3292
rect 11638 3290 11694 3292
rect 11718 3290 11774 3292
rect 11798 3290 11854 3292
rect 11558 3238 11604 3290
rect 11604 3238 11614 3290
rect 11638 3238 11668 3290
rect 11668 3238 11680 3290
rect 11680 3238 11694 3290
rect 11718 3238 11732 3290
rect 11732 3238 11744 3290
rect 11744 3238 11774 3290
rect 11798 3238 11808 3290
rect 11808 3238 11854 3290
rect 11558 3236 11614 3238
rect 11638 3236 11694 3238
rect 11718 3236 11774 3238
rect 11798 3236 11854 3238
rect 11426 3032 11482 3088
rect 11558 2202 11614 2204
rect 11638 2202 11694 2204
rect 11718 2202 11774 2204
rect 11798 2202 11854 2204
rect 11558 2150 11604 2202
rect 11604 2150 11614 2202
rect 11638 2150 11668 2202
rect 11668 2150 11680 2202
rect 11680 2150 11694 2202
rect 11718 2150 11732 2202
rect 11732 2150 11744 2202
rect 11744 2150 11774 2202
rect 11798 2150 11808 2202
rect 11808 2150 11854 2202
rect 11558 2148 11614 2150
rect 11638 2148 11694 2150
rect 11718 2148 11774 2150
rect 11798 2148 11854 2150
rect 9402 1264 9458 1320
rect 10690 584 10746 640
rect 10782 176 10838 232
rect 11242 448 11298 504
rect 11558 1114 11614 1116
rect 11638 1114 11694 1116
rect 11718 1114 11774 1116
rect 11798 1114 11854 1116
rect 11558 1062 11604 1114
rect 11604 1062 11614 1114
rect 11638 1062 11668 1114
rect 11668 1062 11680 1114
rect 11680 1062 11694 1114
rect 11718 1062 11732 1114
rect 11732 1062 11744 1114
rect 11744 1062 11774 1114
rect 11798 1062 11808 1114
rect 11808 1062 11854 1114
rect 11558 1060 11614 1062
rect 11638 1060 11694 1062
rect 11718 1060 11774 1062
rect 11798 1060 11854 1062
rect 12254 3168 12310 3224
rect 13358 2896 13414 2952
rect 12806 2080 12862 2136
rect 12254 312 12310 368
rect 13542 2488 13598 2544
rect 16860 8186 16916 8188
rect 16940 8186 16996 8188
rect 17020 8186 17076 8188
rect 17100 8186 17156 8188
rect 16860 8134 16906 8186
rect 16906 8134 16916 8186
rect 16940 8134 16970 8186
rect 16970 8134 16982 8186
rect 16982 8134 16996 8186
rect 17020 8134 17034 8186
rect 17034 8134 17046 8186
rect 17046 8134 17076 8186
rect 17100 8134 17110 8186
rect 17110 8134 17156 8186
rect 16860 8132 16916 8134
rect 16940 8132 16996 8134
rect 17020 8132 17076 8134
rect 17100 8132 17156 8134
rect 16860 7098 16916 7100
rect 16940 7098 16996 7100
rect 17020 7098 17076 7100
rect 17100 7098 17156 7100
rect 16860 7046 16906 7098
rect 16906 7046 16916 7098
rect 16940 7046 16970 7098
rect 16970 7046 16982 7098
rect 16982 7046 16996 7098
rect 17020 7046 17034 7098
rect 17034 7046 17046 7098
rect 17046 7046 17076 7098
rect 17100 7046 17110 7098
rect 17110 7046 17156 7098
rect 16860 7044 16916 7046
rect 16940 7044 16996 7046
rect 17020 7044 17076 7046
rect 17100 7044 17156 7046
rect 16860 6010 16916 6012
rect 16940 6010 16996 6012
rect 17020 6010 17076 6012
rect 17100 6010 17156 6012
rect 16860 5958 16906 6010
rect 16906 5958 16916 6010
rect 16940 5958 16970 6010
rect 16970 5958 16982 6010
rect 16982 5958 16996 6010
rect 17020 5958 17034 6010
rect 17034 5958 17046 6010
rect 17046 5958 17076 6010
rect 17100 5958 17110 6010
rect 17110 5958 17156 6010
rect 16860 5956 16916 5958
rect 16940 5956 16996 5958
rect 17020 5956 17076 5958
rect 17100 5956 17156 5958
rect 16860 4922 16916 4924
rect 16940 4922 16996 4924
rect 17020 4922 17076 4924
rect 17100 4922 17156 4924
rect 16860 4870 16906 4922
rect 16906 4870 16916 4922
rect 16940 4870 16970 4922
rect 16970 4870 16982 4922
rect 16982 4870 16996 4922
rect 17020 4870 17034 4922
rect 17034 4870 17046 4922
rect 17046 4870 17076 4922
rect 17100 4870 17110 4922
rect 17110 4870 17156 4922
rect 16860 4868 16916 4870
rect 16940 4868 16996 4870
rect 17020 4868 17076 4870
rect 17100 4868 17156 4870
rect 16860 3834 16916 3836
rect 16940 3834 16996 3836
rect 17020 3834 17076 3836
rect 17100 3834 17156 3836
rect 16860 3782 16906 3834
rect 16906 3782 16916 3834
rect 16940 3782 16970 3834
rect 16970 3782 16982 3834
rect 16982 3782 16996 3834
rect 17020 3782 17034 3834
rect 17034 3782 17046 3834
rect 17046 3782 17076 3834
rect 17100 3782 17110 3834
rect 17110 3782 17156 3834
rect 16860 3780 16916 3782
rect 16940 3780 16996 3782
rect 17020 3780 17076 3782
rect 17100 3780 17156 3782
rect 16578 3576 16634 3632
rect 14278 2352 14334 2408
rect 15658 2216 15714 2272
rect 15198 1672 15254 1728
rect 16762 3440 16818 3496
rect 16860 2746 16916 2748
rect 16940 2746 16996 2748
rect 17020 2746 17076 2748
rect 17100 2746 17156 2748
rect 16860 2694 16906 2746
rect 16906 2694 16916 2746
rect 16940 2694 16970 2746
rect 16970 2694 16982 2746
rect 16982 2694 16996 2746
rect 17020 2694 17034 2746
rect 17034 2694 17046 2746
rect 17046 2694 17076 2746
rect 17100 2694 17110 2746
rect 17110 2694 17156 2746
rect 16860 2692 16916 2694
rect 16940 2692 16996 2694
rect 17020 2692 17076 2694
rect 17100 2692 17156 2694
rect 17314 3848 17370 3904
rect 17682 2896 17738 2952
rect 17866 2896 17922 2952
rect 17498 2624 17554 2680
rect 16854 2352 16910 2408
rect 17130 2100 17186 2136
rect 17130 2080 17132 2100
rect 17132 2080 17184 2100
rect 17184 2080 17186 2100
rect 16578 1672 16634 1728
rect 15290 720 15346 776
rect 16486 1400 16542 1456
rect 16860 1658 16916 1660
rect 16940 1658 16996 1660
rect 17020 1658 17076 1660
rect 17100 1658 17156 1660
rect 16860 1606 16906 1658
rect 16906 1606 16916 1658
rect 16940 1606 16970 1658
rect 16970 1606 16982 1658
rect 16982 1606 16996 1658
rect 17020 1606 17034 1658
rect 17034 1606 17046 1658
rect 17046 1606 17076 1658
rect 17100 1606 17110 1658
rect 17110 1606 17156 1658
rect 16860 1604 16916 1606
rect 16940 1604 16996 1606
rect 17020 1604 17076 1606
rect 17100 1604 17156 1606
rect 16486 992 16542 1048
rect 16486 892 16488 912
rect 16488 892 16540 912
rect 16540 892 16542 912
rect 16486 856 16542 892
rect 17774 2760 17830 2816
rect 18234 3032 18290 3088
rect 18050 2352 18106 2408
rect 17498 1808 17554 1864
rect 17866 1808 17922 1864
rect 18050 1808 18106 1864
rect 17682 1708 17684 1728
rect 17684 1708 17736 1728
rect 17736 1708 17738 1728
rect 17682 1672 17738 1708
rect 17774 1536 17830 1592
rect 18234 1672 18290 1728
rect 18694 1964 18750 2000
rect 22161 7642 22217 7644
rect 22241 7642 22297 7644
rect 22321 7642 22377 7644
rect 22401 7642 22457 7644
rect 22161 7590 22207 7642
rect 22207 7590 22217 7642
rect 22241 7590 22271 7642
rect 22271 7590 22283 7642
rect 22283 7590 22297 7642
rect 22321 7590 22335 7642
rect 22335 7590 22347 7642
rect 22347 7590 22377 7642
rect 22401 7590 22411 7642
rect 22411 7590 22457 7642
rect 22161 7588 22217 7590
rect 22241 7588 22297 7590
rect 22321 7588 22377 7590
rect 22401 7588 22457 7590
rect 22161 6554 22217 6556
rect 22241 6554 22297 6556
rect 22321 6554 22377 6556
rect 22401 6554 22457 6556
rect 22161 6502 22207 6554
rect 22207 6502 22217 6554
rect 22241 6502 22271 6554
rect 22271 6502 22283 6554
rect 22283 6502 22297 6554
rect 22321 6502 22335 6554
rect 22335 6502 22347 6554
rect 22347 6502 22377 6554
rect 22401 6502 22411 6554
rect 22411 6502 22457 6554
rect 22161 6500 22217 6502
rect 22241 6500 22297 6502
rect 22321 6500 22377 6502
rect 22401 6500 22457 6502
rect 22161 5466 22217 5468
rect 22241 5466 22297 5468
rect 22321 5466 22377 5468
rect 22401 5466 22457 5468
rect 22161 5414 22207 5466
rect 22207 5414 22217 5466
rect 22241 5414 22271 5466
rect 22271 5414 22283 5466
rect 22283 5414 22297 5466
rect 22321 5414 22335 5466
rect 22335 5414 22347 5466
rect 22347 5414 22377 5466
rect 22401 5414 22411 5466
rect 22411 5414 22457 5466
rect 22161 5412 22217 5414
rect 22241 5412 22297 5414
rect 22321 5412 22377 5414
rect 22401 5412 22457 5414
rect 22161 4378 22217 4380
rect 22241 4378 22297 4380
rect 22321 4378 22377 4380
rect 22401 4378 22457 4380
rect 22161 4326 22207 4378
rect 22207 4326 22217 4378
rect 22241 4326 22271 4378
rect 22271 4326 22283 4378
rect 22283 4326 22297 4378
rect 22321 4326 22335 4378
rect 22335 4326 22347 4378
rect 22347 4326 22377 4378
rect 22401 4326 22411 4378
rect 22411 4326 22457 4378
rect 22161 4324 22217 4326
rect 22241 4324 22297 4326
rect 22321 4324 22377 4326
rect 22401 4324 22457 4326
rect 21822 3984 21878 4040
rect 20350 2624 20406 2680
rect 18694 1944 18696 1964
rect 18696 1944 18748 1964
rect 18748 1944 18750 1964
rect 18694 1828 18750 1864
rect 18694 1808 18696 1828
rect 18696 1808 18748 1828
rect 18748 1808 18750 1828
rect 18694 1672 18750 1728
rect 18142 1400 18198 1456
rect 19430 2080 19486 2136
rect 19338 1708 19340 1728
rect 19340 1708 19392 1728
rect 19392 1708 19394 1728
rect 18142 992 18198 1048
rect 19338 1672 19394 1708
rect 19338 1128 19394 1184
rect 19890 2080 19946 2136
rect 19890 1964 19946 2000
rect 19890 1944 19892 1964
rect 19892 1944 19944 1964
rect 19944 1944 19946 1964
rect 19982 1264 20038 1320
rect 20166 2488 20222 2544
rect 20166 1672 20222 1728
rect 20718 2624 20774 2680
rect 20718 2216 20774 2272
rect 20718 2080 20774 2136
rect 20534 1128 20590 1184
rect 20902 1536 20958 1592
rect 21178 1944 21234 2000
rect 22161 3290 22217 3292
rect 22241 3290 22297 3292
rect 22321 3290 22377 3292
rect 22401 3290 22457 3292
rect 22161 3238 22207 3290
rect 22207 3238 22217 3290
rect 22241 3238 22271 3290
rect 22271 3238 22283 3290
rect 22283 3238 22297 3290
rect 22321 3238 22335 3290
rect 22335 3238 22347 3290
rect 22347 3238 22377 3290
rect 22401 3238 22411 3290
rect 22411 3238 22457 3290
rect 22161 3236 22217 3238
rect 22241 3236 22297 3238
rect 22321 3236 22377 3238
rect 22401 3236 22457 3238
rect 22282 3032 22338 3088
rect 22161 2202 22217 2204
rect 22241 2202 22297 2204
rect 22321 2202 22377 2204
rect 22401 2202 22457 2204
rect 22161 2150 22207 2202
rect 22207 2150 22217 2202
rect 22241 2150 22271 2202
rect 22271 2150 22283 2202
rect 22283 2150 22297 2202
rect 22321 2150 22335 2202
rect 22335 2150 22347 2202
rect 22347 2150 22377 2202
rect 22401 2150 22411 2202
rect 22411 2150 22457 2202
rect 22161 2148 22217 2150
rect 22241 2148 22297 2150
rect 22321 2148 22377 2150
rect 22401 2148 22457 2150
rect 22161 1114 22217 1116
rect 22241 1114 22297 1116
rect 22321 1114 22377 1116
rect 22401 1114 22457 1116
rect 22161 1062 22207 1114
rect 22207 1062 22217 1114
rect 22241 1062 22271 1114
rect 22271 1062 22283 1114
rect 22283 1062 22297 1114
rect 22321 1062 22335 1114
rect 22335 1062 22347 1114
rect 22347 1062 22377 1114
rect 22401 1062 22411 1114
rect 22411 1062 22457 1114
rect 22161 1060 22217 1062
rect 22241 1060 22297 1062
rect 22321 1060 22377 1062
rect 22401 1060 22457 1062
rect 22650 1128 22706 1184
rect 23294 2216 23350 2272
rect 23754 992 23810 1048
rect 24950 4120 25006 4176
rect 32764 8730 32820 8732
rect 32844 8730 32900 8732
rect 32924 8730 32980 8732
rect 33004 8730 33060 8732
rect 32764 8678 32810 8730
rect 32810 8678 32820 8730
rect 32844 8678 32874 8730
rect 32874 8678 32886 8730
rect 32886 8678 32900 8730
rect 32924 8678 32938 8730
rect 32938 8678 32950 8730
rect 32950 8678 32980 8730
rect 33004 8678 33014 8730
rect 33014 8678 33060 8730
rect 32764 8676 32820 8678
rect 32844 8676 32900 8678
rect 32924 8676 32980 8678
rect 33004 8676 33060 8678
rect 43367 8730 43423 8732
rect 43447 8730 43503 8732
rect 43527 8730 43583 8732
rect 43607 8730 43663 8732
rect 43367 8678 43413 8730
rect 43413 8678 43423 8730
rect 43447 8678 43477 8730
rect 43477 8678 43489 8730
rect 43489 8678 43503 8730
rect 43527 8678 43541 8730
rect 43541 8678 43553 8730
rect 43553 8678 43583 8730
rect 43607 8678 43617 8730
rect 43617 8678 43663 8730
rect 43367 8676 43423 8678
rect 43447 8676 43503 8678
rect 43527 8676 43583 8678
rect 43607 8676 43663 8678
rect 27463 8186 27519 8188
rect 27543 8186 27599 8188
rect 27623 8186 27679 8188
rect 27703 8186 27759 8188
rect 27463 8134 27509 8186
rect 27509 8134 27519 8186
rect 27543 8134 27573 8186
rect 27573 8134 27585 8186
rect 27585 8134 27599 8186
rect 27623 8134 27637 8186
rect 27637 8134 27649 8186
rect 27649 8134 27679 8186
rect 27703 8134 27713 8186
rect 27713 8134 27759 8186
rect 27463 8132 27519 8134
rect 27543 8132 27599 8134
rect 27623 8132 27679 8134
rect 27703 8132 27759 8134
rect 27463 7098 27519 7100
rect 27543 7098 27599 7100
rect 27623 7098 27679 7100
rect 27703 7098 27759 7100
rect 27463 7046 27509 7098
rect 27509 7046 27519 7098
rect 27543 7046 27573 7098
rect 27573 7046 27585 7098
rect 27585 7046 27599 7098
rect 27623 7046 27637 7098
rect 27637 7046 27649 7098
rect 27649 7046 27679 7098
rect 27703 7046 27713 7098
rect 27713 7046 27759 7098
rect 27463 7044 27519 7046
rect 27543 7044 27599 7046
rect 27623 7044 27679 7046
rect 27703 7044 27759 7046
rect 25502 1964 25558 2000
rect 25502 1944 25504 1964
rect 25504 1944 25556 1964
rect 25556 1944 25558 1964
rect 26974 2624 27030 2680
rect 27463 6010 27519 6012
rect 27543 6010 27599 6012
rect 27623 6010 27679 6012
rect 27703 6010 27759 6012
rect 27463 5958 27509 6010
rect 27509 5958 27519 6010
rect 27543 5958 27573 6010
rect 27573 5958 27585 6010
rect 27585 5958 27599 6010
rect 27623 5958 27637 6010
rect 27637 5958 27649 6010
rect 27649 5958 27679 6010
rect 27703 5958 27713 6010
rect 27713 5958 27759 6010
rect 27463 5956 27519 5958
rect 27543 5956 27599 5958
rect 27623 5956 27679 5958
rect 27703 5956 27759 5958
rect 27463 4922 27519 4924
rect 27543 4922 27599 4924
rect 27623 4922 27679 4924
rect 27703 4922 27759 4924
rect 27463 4870 27509 4922
rect 27509 4870 27519 4922
rect 27543 4870 27573 4922
rect 27573 4870 27585 4922
rect 27585 4870 27599 4922
rect 27623 4870 27637 4922
rect 27637 4870 27649 4922
rect 27649 4870 27679 4922
rect 27703 4870 27713 4922
rect 27713 4870 27759 4922
rect 27463 4868 27519 4870
rect 27543 4868 27599 4870
rect 27623 4868 27679 4870
rect 27703 4868 27759 4870
rect 27463 3834 27519 3836
rect 27543 3834 27599 3836
rect 27623 3834 27679 3836
rect 27703 3834 27759 3836
rect 27463 3782 27509 3834
rect 27509 3782 27519 3834
rect 27543 3782 27573 3834
rect 27573 3782 27585 3834
rect 27585 3782 27599 3834
rect 27623 3782 27637 3834
rect 27637 3782 27649 3834
rect 27649 3782 27679 3834
rect 27703 3782 27713 3834
rect 27713 3782 27759 3834
rect 27463 3780 27519 3782
rect 27543 3780 27599 3782
rect 27623 3780 27679 3782
rect 27703 3780 27759 3782
rect 27526 3052 27582 3088
rect 27526 3032 27528 3052
rect 27528 3032 27580 3052
rect 27580 3032 27582 3052
rect 27802 2896 27858 2952
rect 27463 2746 27519 2748
rect 27543 2746 27599 2748
rect 27623 2746 27679 2748
rect 27703 2746 27759 2748
rect 27463 2694 27509 2746
rect 27509 2694 27519 2746
rect 27543 2694 27573 2746
rect 27573 2694 27585 2746
rect 27585 2694 27599 2746
rect 27623 2694 27637 2746
rect 27637 2694 27649 2746
rect 27649 2694 27679 2746
rect 27703 2694 27713 2746
rect 27713 2694 27759 2746
rect 27463 2692 27519 2694
rect 27543 2692 27599 2694
rect 27623 2692 27679 2694
rect 27703 2692 27759 2694
rect 26606 2216 26662 2272
rect 27158 2372 27214 2408
rect 27894 2644 27950 2680
rect 27894 2624 27896 2644
rect 27896 2624 27948 2644
rect 27948 2624 27950 2644
rect 27158 2352 27160 2372
rect 27160 2352 27212 2372
rect 27212 2352 27214 2372
rect 27463 1658 27519 1660
rect 27543 1658 27599 1660
rect 27623 1658 27679 1660
rect 27703 1658 27759 1660
rect 27463 1606 27509 1658
rect 27509 1606 27519 1658
rect 27543 1606 27573 1658
rect 27573 1606 27585 1658
rect 27585 1606 27599 1658
rect 27623 1606 27637 1658
rect 27637 1606 27649 1658
rect 27649 1606 27679 1658
rect 27703 1606 27713 1658
rect 27713 1606 27759 1658
rect 27463 1604 27519 1606
rect 27543 1604 27599 1606
rect 27623 1604 27679 1606
rect 27703 1604 27759 1606
rect 27158 992 27214 1048
rect 27618 1128 27674 1184
rect 27986 1400 28042 1456
rect 27986 448 28042 504
rect 28446 312 28502 368
rect 28262 176 28318 232
rect 29366 2488 29422 2544
rect 29274 2080 29330 2136
rect 28998 584 29054 640
rect 30194 2760 30250 2816
rect 30194 2644 30250 2680
rect 30194 2624 30196 2644
rect 30196 2624 30248 2644
rect 30248 2624 30250 2644
rect 30194 2216 30250 2272
rect 32764 7642 32820 7644
rect 32844 7642 32900 7644
rect 32924 7642 32980 7644
rect 33004 7642 33060 7644
rect 32764 7590 32810 7642
rect 32810 7590 32820 7642
rect 32844 7590 32874 7642
rect 32874 7590 32886 7642
rect 32886 7590 32900 7642
rect 32924 7590 32938 7642
rect 32938 7590 32950 7642
rect 32950 7590 32980 7642
rect 33004 7590 33014 7642
rect 33014 7590 33060 7642
rect 32764 7588 32820 7590
rect 32844 7588 32900 7590
rect 32924 7588 32980 7590
rect 33004 7588 33060 7590
rect 32764 6554 32820 6556
rect 32844 6554 32900 6556
rect 32924 6554 32980 6556
rect 33004 6554 33060 6556
rect 32764 6502 32810 6554
rect 32810 6502 32820 6554
rect 32844 6502 32874 6554
rect 32874 6502 32886 6554
rect 32886 6502 32900 6554
rect 32924 6502 32938 6554
rect 32938 6502 32950 6554
rect 32950 6502 32980 6554
rect 33004 6502 33014 6554
rect 33014 6502 33060 6554
rect 32764 6500 32820 6502
rect 32844 6500 32900 6502
rect 32924 6500 32980 6502
rect 33004 6500 33060 6502
rect 32764 5466 32820 5468
rect 32844 5466 32900 5468
rect 32924 5466 32980 5468
rect 33004 5466 33060 5468
rect 32764 5414 32810 5466
rect 32810 5414 32820 5466
rect 32844 5414 32874 5466
rect 32874 5414 32886 5466
rect 32886 5414 32900 5466
rect 32924 5414 32938 5466
rect 32938 5414 32950 5466
rect 32950 5414 32980 5466
rect 33004 5414 33014 5466
rect 33014 5414 33060 5466
rect 32764 5412 32820 5414
rect 32844 5412 32900 5414
rect 32924 5412 32980 5414
rect 33004 5412 33060 5414
rect 32764 4378 32820 4380
rect 32844 4378 32900 4380
rect 32924 4378 32980 4380
rect 33004 4378 33060 4380
rect 32764 4326 32810 4378
rect 32810 4326 32820 4378
rect 32844 4326 32874 4378
rect 32874 4326 32886 4378
rect 32886 4326 32900 4378
rect 32924 4326 32938 4378
rect 32938 4326 32950 4378
rect 32950 4326 32980 4378
rect 33004 4326 33014 4378
rect 33014 4326 33060 4378
rect 32764 4324 32820 4326
rect 32844 4324 32900 4326
rect 32924 4324 32980 4326
rect 33004 4324 33060 4326
rect 32764 3290 32820 3292
rect 32844 3290 32900 3292
rect 32924 3290 32980 3292
rect 33004 3290 33060 3292
rect 32764 3238 32810 3290
rect 32810 3238 32820 3290
rect 32844 3238 32874 3290
rect 32874 3238 32886 3290
rect 32886 3238 32900 3290
rect 32924 3238 32938 3290
rect 32938 3238 32950 3290
rect 32950 3238 32980 3290
rect 33004 3238 33014 3290
rect 33014 3238 33060 3290
rect 32764 3236 32820 3238
rect 32844 3236 32900 3238
rect 32924 3236 32980 3238
rect 33004 3236 33060 3238
rect 31482 3168 31538 3224
rect 31206 2080 31262 2136
rect 33322 4528 33378 4584
rect 35714 2896 35770 2952
rect 35162 2624 35218 2680
rect 32764 2202 32820 2204
rect 32844 2202 32900 2204
rect 32924 2202 32980 2204
rect 33004 2202 33060 2204
rect 32764 2150 32810 2202
rect 32810 2150 32820 2202
rect 32844 2150 32874 2202
rect 32874 2150 32886 2202
rect 32886 2150 32900 2202
rect 32924 2150 32938 2202
rect 32938 2150 32950 2202
rect 32950 2150 32980 2202
rect 33004 2150 33014 2202
rect 33014 2150 33060 2202
rect 32764 2148 32820 2150
rect 32844 2148 32900 2150
rect 32924 2148 32980 2150
rect 33004 2148 33060 2150
rect 31942 856 31998 912
rect 32586 720 32642 776
rect 33322 1808 33378 1864
rect 32764 1114 32820 1116
rect 32844 1114 32900 1116
rect 32924 1114 32980 1116
rect 33004 1114 33060 1116
rect 32764 1062 32810 1114
rect 32810 1062 32820 1114
rect 32844 1062 32874 1114
rect 32874 1062 32886 1114
rect 32886 1062 32900 1114
rect 32924 1062 32938 1114
rect 32938 1062 32950 1114
rect 32950 1062 32980 1114
rect 33004 1062 33014 1114
rect 33014 1062 33060 1114
rect 32764 1060 32820 1062
rect 32844 1060 32900 1062
rect 32924 1060 32980 1062
rect 33004 1060 33060 1062
rect 33874 1964 33930 2000
rect 33874 1944 33876 1964
rect 33876 1944 33928 1964
rect 33928 1944 33930 1964
rect 34518 1264 34574 1320
rect 35162 1300 35164 1320
rect 35164 1300 35216 1320
rect 35216 1300 35218 1320
rect 35162 1264 35218 1300
rect 36266 992 36322 1048
rect 38066 8186 38122 8188
rect 38146 8186 38202 8188
rect 38226 8186 38282 8188
rect 38306 8186 38362 8188
rect 38066 8134 38112 8186
rect 38112 8134 38122 8186
rect 38146 8134 38176 8186
rect 38176 8134 38188 8186
rect 38188 8134 38202 8186
rect 38226 8134 38240 8186
rect 38240 8134 38252 8186
rect 38252 8134 38282 8186
rect 38306 8134 38316 8186
rect 38316 8134 38362 8186
rect 38066 8132 38122 8134
rect 38146 8132 38202 8134
rect 38226 8132 38282 8134
rect 38306 8132 38362 8134
rect 38066 7098 38122 7100
rect 38146 7098 38202 7100
rect 38226 7098 38282 7100
rect 38306 7098 38362 7100
rect 38066 7046 38112 7098
rect 38112 7046 38122 7098
rect 38146 7046 38176 7098
rect 38176 7046 38188 7098
rect 38188 7046 38202 7098
rect 38226 7046 38240 7098
rect 38240 7046 38252 7098
rect 38252 7046 38282 7098
rect 38306 7046 38316 7098
rect 38316 7046 38362 7098
rect 38066 7044 38122 7046
rect 38146 7044 38202 7046
rect 38226 7044 38282 7046
rect 38306 7044 38362 7046
rect 38066 6010 38122 6012
rect 38146 6010 38202 6012
rect 38226 6010 38282 6012
rect 38306 6010 38362 6012
rect 38066 5958 38112 6010
rect 38112 5958 38122 6010
rect 38146 5958 38176 6010
rect 38176 5958 38188 6010
rect 38188 5958 38202 6010
rect 38226 5958 38240 6010
rect 38240 5958 38252 6010
rect 38252 5958 38282 6010
rect 38306 5958 38316 6010
rect 38316 5958 38362 6010
rect 38066 5956 38122 5958
rect 38146 5956 38202 5958
rect 38226 5956 38282 5958
rect 38306 5956 38362 5958
rect 38066 4922 38122 4924
rect 38146 4922 38202 4924
rect 38226 4922 38282 4924
rect 38306 4922 38362 4924
rect 38066 4870 38112 4922
rect 38112 4870 38122 4922
rect 38146 4870 38176 4922
rect 38176 4870 38188 4922
rect 38188 4870 38202 4922
rect 38226 4870 38240 4922
rect 38240 4870 38252 4922
rect 38252 4870 38282 4922
rect 38306 4870 38316 4922
rect 38316 4870 38362 4922
rect 38066 4868 38122 4870
rect 38146 4868 38202 4870
rect 38226 4868 38282 4870
rect 38306 4868 38362 4870
rect 38066 3834 38122 3836
rect 38146 3834 38202 3836
rect 38226 3834 38282 3836
rect 38306 3834 38362 3836
rect 38066 3782 38112 3834
rect 38112 3782 38122 3834
rect 38146 3782 38176 3834
rect 38176 3782 38188 3834
rect 38188 3782 38202 3834
rect 38226 3782 38240 3834
rect 38240 3782 38252 3834
rect 38252 3782 38282 3834
rect 38306 3782 38316 3834
rect 38316 3782 38362 3834
rect 38066 3780 38122 3782
rect 38146 3780 38202 3782
rect 38226 3780 38282 3782
rect 38306 3780 38362 3782
rect 37462 3576 37518 3632
rect 38066 2746 38122 2748
rect 38146 2746 38202 2748
rect 38226 2746 38282 2748
rect 38306 2746 38362 2748
rect 38066 2694 38112 2746
rect 38112 2694 38122 2746
rect 38146 2694 38176 2746
rect 38176 2694 38188 2746
rect 38188 2694 38202 2746
rect 38226 2694 38240 2746
rect 38240 2694 38252 2746
rect 38252 2694 38282 2746
rect 38306 2694 38316 2746
rect 38316 2694 38362 2746
rect 38066 2692 38122 2694
rect 38146 2692 38202 2694
rect 38226 2692 38282 2694
rect 38306 2692 38362 2694
rect 38066 1658 38122 1660
rect 38146 1658 38202 1660
rect 38226 1658 38282 1660
rect 38306 1658 38362 1660
rect 38066 1606 38112 1658
rect 38112 1606 38122 1658
rect 38146 1606 38176 1658
rect 38176 1606 38188 1658
rect 38188 1606 38202 1658
rect 38226 1606 38240 1658
rect 38240 1606 38252 1658
rect 38252 1606 38282 1658
rect 38306 1606 38316 1658
rect 38316 1606 38362 1658
rect 38066 1604 38122 1606
rect 38146 1604 38202 1606
rect 38226 1604 38282 1606
rect 38306 1604 38362 1606
rect 39302 2352 39358 2408
rect 39670 3032 39726 3088
rect 43367 7642 43423 7644
rect 43447 7642 43503 7644
rect 43527 7642 43583 7644
rect 43607 7642 43663 7644
rect 43367 7590 43413 7642
rect 43413 7590 43423 7642
rect 43447 7590 43477 7642
rect 43477 7590 43489 7642
rect 43489 7590 43503 7642
rect 43527 7590 43541 7642
rect 43541 7590 43553 7642
rect 43553 7590 43583 7642
rect 43607 7590 43617 7642
rect 43617 7590 43663 7642
rect 43367 7588 43423 7590
rect 43447 7588 43503 7590
rect 43527 7588 43583 7590
rect 43607 7588 43663 7590
rect 43367 6554 43423 6556
rect 43447 6554 43503 6556
rect 43527 6554 43583 6556
rect 43607 6554 43663 6556
rect 43367 6502 43413 6554
rect 43413 6502 43423 6554
rect 43447 6502 43477 6554
rect 43477 6502 43489 6554
rect 43489 6502 43503 6554
rect 43527 6502 43541 6554
rect 43541 6502 43553 6554
rect 43553 6502 43583 6554
rect 43607 6502 43617 6554
rect 43617 6502 43663 6554
rect 43367 6500 43423 6502
rect 43447 6500 43503 6502
rect 43527 6500 43583 6502
rect 43607 6500 43663 6502
rect 43367 5466 43423 5468
rect 43447 5466 43503 5468
rect 43527 5466 43583 5468
rect 43607 5466 43663 5468
rect 43367 5414 43413 5466
rect 43413 5414 43423 5466
rect 43447 5414 43477 5466
rect 43477 5414 43489 5466
rect 43489 5414 43503 5466
rect 43527 5414 43541 5466
rect 43541 5414 43553 5466
rect 43553 5414 43583 5466
rect 43607 5414 43617 5466
rect 43617 5414 43663 5466
rect 43367 5412 43423 5414
rect 43447 5412 43503 5414
rect 43527 5412 43583 5414
rect 43607 5412 43663 5414
rect 43367 4378 43423 4380
rect 43447 4378 43503 4380
rect 43527 4378 43583 4380
rect 43607 4378 43663 4380
rect 43367 4326 43413 4378
rect 43413 4326 43423 4378
rect 43447 4326 43477 4378
rect 43477 4326 43489 4378
rect 43489 4326 43503 4378
rect 43527 4326 43541 4378
rect 43541 4326 43553 4378
rect 43553 4326 43583 4378
rect 43607 4326 43617 4378
rect 43617 4326 43663 4378
rect 43367 4324 43423 4326
rect 43447 4324 43503 4326
rect 43527 4324 43583 4326
rect 43607 4324 43663 4326
rect 43367 3290 43423 3292
rect 43447 3290 43503 3292
rect 43527 3290 43583 3292
rect 43607 3290 43663 3292
rect 43367 3238 43413 3290
rect 43413 3238 43423 3290
rect 43447 3238 43477 3290
rect 43477 3238 43489 3290
rect 43489 3238 43503 3290
rect 43527 3238 43541 3290
rect 43541 3238 43553 3290
rect 43553 3238 43583 3290
rect 43607 3238 43617 3290
rect 43617 3238 43663 3290
rect 43367 3236 43423 3238
rect 43447 3236 43503 3238
rect 43527 3236 43583 3238
rect 43607 3236 43663 3238
rect 43367 2202 43423 2204
rect 43447 2202 43503 2204
rect 43527 2202 43583 2204
rect 43607 2202 43663 2204
rect 43367 2150 43413 2202
rect 43413 2150 43423 2202
rect 43447 2150 43477 2202
rect 43477 2150 43489 2202
rect 43489 2150 43503 2202
rect 43527 2150 43541 2202
rect 43541 2150 43553 2202
rect 43553 2150 43583 2202
rect 43607 2150 43617 2202
rect 43617 2150 43663 2202
rect 43367 2148 43423 2150
rect 43447 2148 43503 2150
rect 43527 2148 43583 2150
rect 43607 2148 43663 2150
rect 38842 448 38898 504
rect 43367 1114 43423 1116
rect 43447 1114 43503 1116
rect 43527 1114 43583 1116
rect 43607 1114 43663 1116
rect 43367 1062 43413 1114
rect 43413 1062 43423 1114
rect 43447 1062 43477 1114
rect 43477 1062 43489 1114
rect 43489 1062 43503 1114
rect 43527 1062 43541 1114
rect 43541 1062 43553 1114
rect 43553 1062 43583 1114
rect 43607 1062 43617 1114
rect 43617 1062 43663 1114
rect 43367 1060 43423 1062
rect 43447 1060 43503 1062
rect 43527 1060 43583 1062
rect 43607 1060 43663 1062
<< metal3 >>
rect 11548 8736 11864 8737
rect 11548 8672 11554 8736
rect 11618 8672 11634 8736
rect 11698 8672 11714 8736
rect 11778 8672 11794 8736
rect 11858 8672 11864 8736
rect 11548 8671 11864 8672
rect 22151 8736 22467 8737
rect 22151 8672 22157 8736
rect 22221 8672 22237 8736
rect 22301 8672 22317 8736
rect 22381 8672 22397 8736
rect 22461 8672 22467 8736
rect 22151 8671 22467 8672
rect 32754 8736 33070 8737
rect 32754 8672 32760 8736
rect 32824 8672 32840 8736
rect 32904 8672 32920 8736
rect 32984 8672 33000 8736
rect 33064 8672 33070 8736
rect 32754 8671 33070 8672
rect 43357 8736 43673 8737
rect 43357 8672 43363 8736
rect 43427 8672 43443 8736
rect 43507 8672 43523 8736
rect 43587 8672 43603 8736
rect 43667 8672 43673 8736
rect 43357 8671 43673 8672
rect 9581 8530 9647 8533
rect 27838 8530 27844 8532
rect 9581 8528 27844 8530
rect 9581 8472 9586 8528
rect 9642 8472 27844 8528
rect 9581 8470 27844 8472
rect 9581 8467 9647 8470
rect 27838 8468 27844 8470
rect 27908 8468 27914 8532
rect 2221 8394 2287 8397
rect 29494 8394 29500 8396
rect 2221 8392 29500 8394
rect 2221 8336 2226 8392
rect 2282 8336 29500 8392
rect 2221 8334 29500 8336
rect 2221 8331 2287 8334
rect 29494 8332 29500 8334
rect 29564 8332 29570 8396
rect 6247 8192 6563 8193
rect 6247 8128 6253 8192
rect 6317 8128 6333 8192
rect 6397 8128 6413 8192
rect 6477 8128 6493 8192
rect 6557 8128 6563 8192
rect 6247 8127 6563 8128
rect 16850 8192 17166 8193
rect 16850 8128 16856 8192
rect 16920 8128 16936 8192
rect 17000 8128 17016 8192
rect 17080 8128 17096 8192
rect 17160 8128 17166 8192
rect 16850 8127 17166 8128
rect 27453 8192 27769 8193
rect 27453 8128 27459 8192
rect 27523 8128 27539 8192
rect 27603 8128 27619 8192
rect 27683 8128 27699 8192
rect 27763 8128 27769 8192
rect 27453 8127 27769 8128
rect 38056 8192 38372 8193
rect 38056 8128 38062 8192
rect 38126 8128 38142 8192
rect 38206 8128 38222 8192
rect 38286 8128 38302 8192
rect 38366 8128 38372 8192
rect 38056 8127 38372 8128
rect 11548 7648 11864 7649
rect 11548 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11864 7648
rect 11548 7583 11864 7584
rect 22151 7648 22467 7649
rect 22151 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22467 7648
rect 22151 7583 22467 7584
rect 32754 7648 33070 7649
rect 32754 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33070 7648
rect 32754 7583 33070 7584
rect 43357 7648 43673 7649
rect 43357 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43673 7648
rect 43357 7583 43673 7584
rect 6247 7104 6563 7105
rect 6247 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6563 7104
rect 6247 7039 6563 7040
rect 16850 7104 17166 7105
rect 16850 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17166 7104
rect 16850 7039 17166 7040
rect 27453 7104 27769 7105
rect 27453 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27769 7104
rect 27453 7039 27769 7040
rect 38056 7104 38372 7105
rect 38056 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38372 7104
rect 38056 7039 38372 7040
rect 11548 6560 11864 6561
rect 11548 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11864 6560
rect 11548 6495 11864 6496
rect 22151 6560 22467 6561
rect 22151 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22467 6560
rect 22151 6495 22467 6496
rect 32754 6560 33070 6561
rect 32754 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33070 6560
rect 32754 6495 33070 6496
rect 43357 6560 43673 6561
rect 43357 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43673 6560
rect 43357 6495 43673 6496
rect 6247 6016 6563 6017
rect 6247 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6563 6016
rect 6247 5951 6563 5952
rect 16850 6016 17166 6017
rect 16850 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17166 6016
rect 16850 5951 17166 5952
rect 27453 6016 27769 6017
rect 27453 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27769 6016
rect 27453 5951 27769 5952
rect 38056 6016 38372 6017
rect 38056 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38372 6016
rect 38056 5951 38372 5952
rect 11548 5472 11864 5473
rect 11548 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11864 5472
rect 11548 5407 11864 5408
rect 22151 5472 22467 5473
rect 22151 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22467 5472
rect 22151 5407 22467 5408
rect 32754 5472 33070 5473
rect 32754 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33070 5472
rect 32754 5407 33070 5408
rect 43357 5472 43673 5473
rect 43357 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43673 5472
rect 43357 5407 43673 5408
rect 6247 4928 6563 4929
rect 6247 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6563 4928
rect 6247 4863 6563 4864
rect 16850 4928 17166 4929
rect 16850 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17166 4928
rect 16850 4863 17166 4864
rect 27453 4928 27769 4929
rect 27453 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27769 4928
rect 27453 4863 27769 4864
rect 38056 4928 38372 4929
rect 38056 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38372 4928
rect 38056 4863 38372 4864
rect 16062 4524 16068 4588
rect 16132 4586 16138 4588
rect 33317 4586 33383 4589
rect 16132 4584 33383 4586
rect 16132 4528 33322 4584
rect 33378 4528 33383 4584
rect 16132 4526 33383 4528
rect 16132 4524 16138 4526
rect 33317 4523 33383 4526
rect 11548 4384 11864 4385
rect 11548 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11864 4384
rect 11548 4319 11864 4320
rect 22151 4384 22467 4385
rect 22151 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22467 4384
rect 22151 4319 22467 4320
rect 32754 4384 33070 4385
rect 32754 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33070 4384
rect 32754 4319 33070 4320
rect 43357 4384 43673 4385
rect 43357 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43673 4384
rect 43357 4319 43673 4320
rect 6729 4178 6795 4181
rect 24945 4178 25011 4181
rect 6729 4176 25011 4178
rect 6729 4120 6734 4176
rect 6790 4120 24950 4176
rect 25006 4120 25011 4176
rect 6729 4118 25011 4120
rect 6729 4115 6795 4118
rect 24945 4115 25011 4118
rect 8201 4042 8267 4045
rect 21817 4042 21883 4045
rect 8201 4040 21883 4042
rect 8201 3984 8206 4040
rect 8262 3984 21822 4040
rect 21878 3984 21883 4040
rect 8201 3982 21883 3984
rect 8201 3979 8267 3982
rect 21817 3979 21883 3982
rect 26190 3982 31770 4042
rect 17309 3906 17375 3909
rect 26190 3906 26250 3982
rect 31710 3908 31770 3982
rect 17309 3904 26250 3906
rect 17309 3848 17314 3904
rect 17370 3848 26250 3904
rect 17309 3846 26250 3848
rect 17309 3843 17375 3846
rect 31702 3844 31708 3908
rect 31772 3844 31778 3908
rect 6247 3840 6563 3841
rect 6247 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6563 3840
rect 6247 3775 6563 3776
rect 16850 3840 17166 3841
rect 16850 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17166 3840
rect 16850 3775 17166 3776
rect 27453 3840 27769 3841
rect 27453 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27769 3840
rect 27453 3775 27769 3776
rect 38056 3840 38372 3841
rect 38056 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38372 3840
rect 38056 3775 38372 3776
rect 16573 3634 16639 3637
rect 37457 3634 37523 3637
rect 16573 3632 37523 3634
rect 16573 3576 16578 3632
rect 16634 3576 37462 3632
rect 37518 3576 37523 3632
rect 16573 3574 37523 3576
rect 16573 3571 16639 3574
rect 37457 3571 37523 3574
rect 16757 3498 16823 3501
rect 34646 3498 34652 3500
rect 16757 3496 34652 3498
rect 16757 3440 16762 3496
rect 16818 3440 34652 3496
rect 16757 3438 34652 3440
rect 16757 3435 16823 3438
rect 34646 3436 34652 3438
rect 34716 3436 34722 3500
rect 11548 3296 11864 3297
rect 11548 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11864 3296
rect 11548 3231 11864 3232
rect 22151 3296 22467 3297
rect 22151 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22467 3296
rect 22151 3231 22467 3232
rect 32754 3296 33070 3297
rect 32754 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33070 3296
rect 32754 3231 33070 3232
rect 43357 3296 43673 3297
rect 43357 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43673 3296
rect 43357 3231 43673 3232
rect 12249 3226 12315 3229
rect 31477 3226 31543 3229
rect 12249 3224 19350 3226
rect 12249 3168 12254 3224
rect 12310 3168 19350 3224
rect 12249 3166 19350 3168
rect 12249 3163 12315 3166
rect 11421 3090 11487 3093
rect 18229 3090 18295 3093
rect 11421 3088 18295 3090
rect 11421 3032 11426 3088
rect 11482 3032 18234 3088
rect 18290 3032 18295 3088
rect 11421 3030 18295 3032
rect 19290 3090 19350 3166
rect 26190 3224 31543 3226
rect 26190 3168 31482 3224
rect 31538 3168 31543 3224
rect 26190 3166 31543 3168
rect 22277 3090 22343 3093
rect 19290 3088 22343 3090
rect 19290 3032 22282 3088
rect 22338 3032 22343 3088
rect 19290 3030 22343 3032
rect 11421 3027 11487 3030
rect 18229 3027 18295 3030
rect 22277 3027 22343 3030
rect 13353 2954 13419 2957
rect 17677 2954 17743 2957
rect 13353 2952 17743 2954
rect 13353 2896 13358 2952
rect 13414 2896 17682 2952
rect 17738 2896 17743 2952
rect 13353 2894 17743 2896
rect 13353 2891 13419 2894
rect 17677 2891 17743 2894
rect 17861 2954 17927 2957
rect 26190 2954 26250 3166
rect 31477 3163 31543 3166
rect 27521 3090 27587 3093
rect 39665 3090 39731 3093
rect 27521 3088 39731 3090
rect 27521 3032 27526 3088
rect 27582 3032 39670 3088
rect 39726 3032 39731 3088
rect 27521 3030 39731 3032
rect 27521 3027 27587 3030
rect 39665 3027 39731 3030
rect 17861 2952 26250 2954
rect 17861 2896 17866 2952
rect 17922 2896 26250 2952
rect 17861 2894 26250 2896
rect 27797 2954 27863 2957
rect 35709 2954 35775 2957
rect 27797 2952 35775 2954
rect 27797 2896 27802 2952
rect 27858 2896 35714 2952
rect 35770 2896 35775 2952
rect 27797 2894 35775 2896
rect 17861 2891 17927 2894
rect 27797 2891 27863 2894
rect 35709 2891 35775 2894
rect 17769 2818 17835 2821
rect 30189 2820 30255 2821
rect 27286 2818 27292 2820
rect 17769 2816 27292 2818
rect 17769 2760 17774 2816
rect 17830 2760 27292 2816
rect 17769 2758 27292 2760
rect 17769 2755 17835 2758
rect 27286 2756 27292 2758
rect 27356 2756 27362 2820
rect 30189 2818 30236 2820
rect 30144 2816 30236 2818
rect 30144 2760 30194 2816
rect 30144 2758 30236 2760
rect 30189 2756 30236 2758
rect 30300 2756 30306 2820
rect 30189 2755 30255 2756
rect 6247 2752 6563 2753
rect 6247 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6563 2752
rect 6247 2687 6563 2688
rect 16850 2752 17166 2753
rect 16850 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17166 2752
rect 16850 2687 17166 2688
rect 27453 2752 27769 2753
rect 27453 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27769 2752
rect 27453 2687 27769 2688
rect 38056 2752 38372 2753
rect 38056 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38372 2752
rect 38056 2687 38372 2688
rect 17493 2682 17559 2685
rect 20345 2682 20411 2685
rect 17493 2680 20411 2682
rect 17493 2624 17498 2680
rect 17554 2624 20350 2680
rect 20406 2624 20411 2680
rect 17493 2622 20411 2624
rect 17493 2619 17559 2622
rect 20345 2619 20411 2622
rect 20713 2682 20779 2685
rect 26969 2682 27035 2685
rect 27889 2684 27955 2685
rect 20713 2680 27035 2682
rect 20713 2624 20718 2680
rect 20774 2624 26974 2680
rect 27030 2624 27035 2680
rect 20713 2622 27035 2624
rect 20713 2619 20779 2622
rect 26969 2619 27035 2622
rect 27838 2620 27844 2684
rect 27908 2682 27955 2684
rect 27908 2680 28000 2682
rect 27950 2624 28000 2680
rect 27908 2622 28000 2624
rect 27908 2620 27955 2622
rect 29494 2620 29500 2684
rect 29564 2682 29570 2684
rect 30189 2682 30255 2685
rect 29564 2680 30255 2682
rect 29564 2624 30194 2680
rect 30250 2624 30255 2680
rect 29564 2622 30255 2624
rect 29564 2620 29570 2622
rect 27889 2619 27955 2620
rect 30189 2619 30255 2622
rect 31702 2620 31708 2684
rect 31772 2682 31778 2684
rect 35157 2682 35223 2685
rect 31772 2680 35223 2682
rect 31772 2624 35162 2680
rect 35218 2624 35223 2680
rect 31772 2622 35223 2624
rect 31772 2620 31778 2622
rect 35157 2619 35223 2622
rect 13537 2546 13603 2549
rect 20161 2546 20227 2549
rect 13537 2544 20227 2546
rect 13537 2488 13542 2544
rect 13598 2488 20166 2544
rect 20222 2488 20227 2544
rect 13537 2486 20227 2488
rect 13537 2483 13603 2486
rect 20161 2483 20227 2486
rect 24894 2484 24900 2548
rect 24964 2546 24970 2548
rect 29361 2546 29427 2549
rect 24964 2544 29427 2546
rect 24964 2488 29366 2544
rect 29422 2488 29427 2544
rect 24964 2486 29427 2488
rect 24964 2484 24970 2486
rect 29361 2483 29427 2486
rect 14273 2410 14339 2413
rect 16849 2410 16915 2413
rect 14273 2408 16915 2410
rect 14273 2352 14278 2408
rect 14334 2352 16854 2408
rect 16910 2352 16915 2408
rect 14273 2350 16915 2352
rect 14273 2347 14339 2350
rect 16849 2347 16915 2350
rect 18045 2410 18111 2413
rect 27153 2410 27219 2413
rect 39297 2410 39363 2413
rect 18045 2408 26802 2410
rect 18045 2352 18050 2408
rect 18106 2352 26802 2408
rect 18045 2350 26802 2352
rect 18045 2347 18111 2350
rect 15653 2274 15719 2277
rect 16062 2274 16068 2276
rect 15653 2272 16068 2274
rect 15653 2216 15658 2272
rect 15714 2216 16068 2272
rect 15653 2214 16068 2216
rect 15653 2211 15719 2214
rect 16062 2212 16068 2214
rect 16132 2212 16138 2276
rect 20713 2274 20779 2277
rect 16254 2272 20779 2274
rect 16254 2216 20718 2272
rect 20774 2216 20779 2272
rect 16254 2214 20779 2216
rect 11548 2208 11864 2209
rect 11548 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11864 2208
rect 11548 2143 11864 2144
rect 12801 2138 12867 2141
rect 16254 2138 16314 2214
rect 20713 2211 20779 2214
rect 23289 2274 23355 2277
rect 26601 2274 26667 2277
rect 23289 2272 26667 2274
rect 23289 2216 23294 2272
rect 23350 2216 26606 2272
rect 26662 2216 26667 2272
rect 23289 2214 26667 2216
rect 26742 2274 26802 2350
rect 27153 2408 39363 2410
rect 27153 2352 27158 2408
rect 27214 2352 39302 2408
rect 39358 2352 39363 2408
rect 27153 2350 39363 2352
rect 27153 2347 27219 2350
rect 39297 2347 39363 2350
rect 30189 2274 30255 2277
rect 26742 2272 30255 2274
rect 26742 2216 30194 2272
rect 30250 2216 30255 2272
rect 26742 2214 30255 2216
rect 23289 2211 23355 2214
rect 26601 2211 26667 2214
rect 30189 2211 30255 2214
rect 22151 2208 22467 2209
rect 22151 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22467 2208
rect 22151 2143 22467 2144
rect 32754 2208 33070 2209
rect 32754 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33070 2208
rect 32754 2143 33070 2144
rect 43357 2208 43673 2209
rect 43357 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43673 2208
rect 43357 2143 43673 2144
rect 12801 2136 16314 2138
rect 12801 2080 12806 2136
rect 12862 2080 16314 2136
rect 12801 2078 16314 2080
rect 17125 2138 17191 2141
rect 17125 2136 19350 2138
rect 17125 2080 17130 2136
rect 17186 2080 19350 2136
rect 17125 2078 19350 2080
rect 12801 2075 12867 2078
rect 17125 2075 17191 2078
rect 9029 2002 9095 2005
rect 18689 2002 18755 2005
rect 9029 2000 18755 2002
rect 9029 1944 9034 2000
rect 9090 1944 18694 2000
rect 18750 1944 18755 2000
rect 9029 1942 18755 1944
rect 9029 1939 9095 1942
rect 18689 1939 18755 1942
rect 8937 1866 9003 1869
rect 17493 1866 17559 1869
rect 17861 1866 17927 1869
rect 8937 1864 17559 1866
rect 8937 1808 8942 1864
rect 8998 1808 17498 1864
rect 17554 1808 17559 1864
rect 8937 1806 17559 1808
rect 8937 1803 9003 1806
rect 17493 1803 17559 1806
rect 17680 1864 17927 1866
rect 17680 1808 17866 1864
rect 17922 1808 17927 1864
rect 17680 1806 17927 1808
rect 17680 1733 17740 1806
rect 17861 1803 17927 1806
rect 18045 1866 18111 1869
rect 18689 1866 18755 1869
rect 18045 1864 18755 1866
rect 18045 1808 18050 1864
rect 18106 1808 18694 1864
rect 18750 1808 18755 1864
rect 18045 1806 18755 1808
rect 19290 1866 19350 2078
rect 19425 2136 19491 2141
rect 19425 2080 19430 2136
rect 19486 2080 19491 2136
rect 19425 2075 19491 2080
rect 19885 2138 19951 2141
rect 20713 2138 20779 2141
rect 19885 2136 20779 2138
rect 19885 2080 19890 2136
rect 19946 2080 20718 2136
rect 20774 2080 20779 2136
rect 19885 2078 20779 2080
rect 19885 2075 19951 2078
rect 20713 2075 20779 2078
rect 29269 2138 29335 2141
rect 31201 2138 31267 2141
rect 29269 2136 31267 2138
rect 29269 2080 29274 2136
rect 29330 2080 31206 2136
rect 31262 2080 31267 2136
rect 29269 2078 31267 2080
rect 29269 2075 29335 2078
rect 31201 2075 31267 2078
rect 19428 2002 19488 2075
rect 19885 2002 19951 2005
rect 19428 2000 19951 2002
rect 19428 1944 19890 2000
rect 19946 1944 19951 2000
rect 19428 1942 19951 1944
rect 19885 1939 19951 1942
rect 21173 2002 21239 2005
rect 25497 2002 25563 2005
rect 21173 2000 25563 2002
rect 21173 1944 21178 2000
rect 21234 1944 25502 2000
rect 25558 1944 25563 2000
rect 21173 1942 25563 1944
rect 21173 1939 21239 1942
rect 25497 1939 25563 1942
rect 27286 1940 27292 2004
rect 27356 2002 27362 2004
rect 33869 2002 33935 2005
rect 27356 2000 33935 2002
rect 27356 1944 33874 2000
rect 33930 1944 33935 2000
rect 27356 1942 33935 1944
rect 27356 1940 27362 1942
rect 33869 1939 33935 1942
rect 33317 1866 33383 1869
rect 19290 1864 33383 1866
rect 19290 1808 33322 1864
rect 33378 1808 33383 1864
rect 19290 1806 33383 1808
rect 18045 1803 18111 1806
rect 18689 1803 18755 1806
rect 33317 1803 33383 1806
rect 15193 1730 15259 1733
rect 16573 1730 16639 1733
rect 15193 1728 16639 1730
rect 15193 1672 15198 1728
rect 15254 1672 16578 1728
rect 16634 1672 16639 1728
rect 15193 1670 16639 1672
rect 15193 1667 15259 1670
rect 16573 1667 16639 1670
rect 17677 1728 17743 1733
rect 17677 1672 17682 1728
rect 17738 1672 17743 1728
rect 17677 1667 17743 1672
rect 18229 1730 18295 1733
rect 18689 1730 18755 1733
rect 18229 1728 18755 1730
rect 18229 1672 18234 1728
rect 18290 1672 18694 1728
rect 18750 1672 18755 1728
rect 18229 1670 18755 1672
rect 18229 1667 18295 1670
rect 18689 1667 18755 1670
rect 19333 1730 19399 1733
rect 20161 1730 20227 1733
rect 19333 1728 20227 1730
rect 19333 1672 19338 1728
rect 19394 1672 20166 1728
rect 20222 1672 20227 1728
rect 19333 1670 20227 1672
rect 19333 1667 19399 1670
rect 20161 1667 20227 1670
rect 6247 1664 6563 1665
rect 6247 1600 6253 1664
rect 6317 1600 6333 1664
rect 6397 1600 6413 1664
rect 6477 1600 6493 1664
rect 6557 1600 6563 1664
rect 6247 1599 6563 1600
rect 16850 1664 17166 1665
rect 16850 1600 16856 1664
rect 16920 1600 16936 1664
rect 17000 1600 17016 1664
rect 17080 1600 17096 1664
rect 17160 1600 17166 1664
rect 16850 1599 17166 1600
rect 27453 1664 27769 1665
rect 27453 1600 27459 1664
rect 27523 1600 27539 1664
rect 27603 1600 27619 1664
rect 27683 1600 27699 1664
rect 27763 1600 27769 1664
rect 27453 1599 27769 1600
rect 38056 1664 38372 1665
rect 38056 1600 38062 1664
rect 38126 1600 38142 1664
rect 38206 1600 38222 1664
rect 38286 1600 38302 1664
rect 38366 1600 38372 1664
rect 38056 1599 38372 1600
rect 17769 1594 17835 1597
rect 20897 1594 20963 1597
rect 17769 1592 20178 1594
rect 17769 1536 17774 1592
rect 17830 1536 20178 1592
rect 17769 1534 20178 1536
rect 17769 1531 17835 1534
rect 16481 1458 16547 1461
rect 18137 1458 18203 1461
rect 16481 1456 18203 1458
rect 16481 1400 16486 1456
rect 16542 1400 18142 1456
rect 18198 1400 18203 1456
rect 16481 1398 18203 1400
rect 16481 1395 16547 1398
rect 18137 1395 18203 1398
rect 9397 1322 9463 1325
rect 19977 1322 20043 1325
rect 9397 1320 20043 1322
rect 9397 1264 9402 1320
rect 9458 1264 19982 1320
rect 20038 1264 20043 1320
rect 9397 1262 20043 1264
rect 20118 1322 20178 1534
rect 20897 1592 27170 1594
rect 20897 1536 20902 1592
rect 20958 1536 27170 1592
rect 20897 1534 27170 1536
rect 20897 1531 20963 1534
rect 27110 1458 27170 1534
rect 27981 1458 28047 1461
rect 27110 1456 28047 1458
rect 27110 1400 27986 1456
rect 28042 1400 28047 1456
rect 27110 1398 28047 1400
rect 27981 1395 28047 1398
rect 34513 1322 34579 1325
rect 20118 1320 34579 1322
rect 20118 1264 34518 1320
rect 34574 1264 34579 1320
rect 20118 1262 34579 1264
rect 9397 1259 9463 1262
rect 19977 1259 20043 1262
rect 34513 1259 34579 1262
rect 34646 1260 34652 1324
rect 34716 1322 34722 1324
rect 35157 1322 35223 1325
rect 34716 1320 35223 1322
rect 34716 1264 35162 1320
rect 35218 1264 35223 1320
rect 34716 1262 35223 1264
rect 34716 1260 34722 1262
rect 35157 1259 35223 1262
rect 19333 1186 19399 1189
rect 20529 1186 20595 1189
rect 19333 1184 20595 1186
rect 19333 1128 19338 1184
rect 19394 1128 20534 1184
rect 20590 1128 20595 1184
rect 19333 1126 20595 1128
rect 19333 1123 19399 1126
rect 20529 1123 20595 1126
rect 22645 1186 22711 1189
rect 27613 1186 27679 1189
rect 22645 1184 27679 1186
rect 22645 1128 22650 1184
rect 22706 1128 27618 1184
rect 27674 1128 27679 1184
rect 22645 1126 27679 1128
rect 22645 1123 22711 1126
rect 27613 1123 27679 1126
rect 11548 1120 11864 1121
rect 11548 1056 11554 1120
rect 11618 1056 11634 1120
rect 11698 1056 11714 1120
rect 11778 1056 11794 1120
rect 11858 1056 11864 1120
rect 11548 1055 11864 1056
rect 22151 1120 22467 1121
rect 22151 1056 22157 1120
rect 22221 1056 22237 1120
rect 22301 1056 22317 1120
rect 22381 1056 22397 1120
rect 22461 1056 22467 1120
rect 22151 1055 22467 1056
rect 32754 1120 33070 1121
rect 32754 1056 32760 1120
rect 32824 1056 32840 1120
rect 32904 1056 32920 1120
rect 32984 1056 33000 1120
rect 33064 1056 33070 1120
rect 32754 1055 33070 1056
rect 43357 1120 43673 1121
rect 43357 1056 43363 1120
rect 43427 1056 43443 1120
rect 43507 1056 43523 1120
rect 43587 1056 43603 1120
rect 43667 1056 43673 1120
rect 43357 1055 43673 1056
rect 16481 1050 16547 1053
rect 18137 1050 18203 1053
rect 16481 1048 18203 1050
rect 16481 992 16486 1048
rect 16542 992 18142 1048
rect 18198 992 18203 1048
rect 16481 990 18203 992
rect 16481 987 16547 990
rect 18137 987 18203 990
rect 23749 1050 23815 1053
rect 27153 1050 27219 1053
rect 23749 1048 27219 1050
rect 23749 992 23754 1048
rect 23810 992 27158 1048
rect 27214 992 27219 1048
rect 23749 990 27219 992
rect 23749 987 23815 990
rect 27153 987 27219 990
rect 30230 988 30236 1052
rect 30300 1050 30306 1052
rect 36261 1050 36327 1053
rect 30300 990 32690 1050
rect 30300 988 30306 990
rect 16481 914 16547 917
rect 31937 914 32003 917
rect 16481 912 32003 914
rect 16481 856 16486 912
rect 16542 856 31942 912
rect 31998 856 32003 912
rect 16481 854 32003 856
rect 32630 914 32690 990
rect 33182 1048 36327 1050
rect 33182 992 36266 1048
rect 36322 992 36327 1048
rect 33182 990 36327 992
rect 33182 914 33242 990
rect 36261 987 36327 990
rect 32630 854 33242 914
rect 16481 851 16547 854
rect 31937 851 32003 854
rect 15285 778 15351 781
rect 32581 778 32647 781
rect 15285 776 32647 778
rect 15285 720 15290 776
rect 15346 720 32586 776
rect 32642 720 32647 776
rect 15285 718 32647 720
rect 15285 715 15351 718
rect 32581 715 32647 718
rect 10685 642 10751 645
rect 28993 642 29059 645
rect 10685 640 29059 642
rect 10685 584 10690 640
rect 10746 584 28998 640
rect 29054 584 29059 640
rect 10685 582 29059 584
rect 10685 579 10751 582
rect 28993 579 29059 582
rect 11237 506 11303 509
rect 27981 506 28047 509
rect 38837 506 38903 509
rect 11237 504 25330 506
rect 11237 448 11242 504
rect 11298 448 25330 504
rect 11237 446 25330 448
rect 11237 443 11303 446
rect 12249 370 12315 373
rect 25270 370 25330 446
rect 27981 504 38903 506
rect 27981 448 27986 504
rect 28042 448 38842 504
rect 38898 448 38903 504
rect 27981 446 38903 448
rect 27981 443 28047 446
rect 38837 443 38903 446
rect 28441 370 28507 373
rect 12249 368 25146 370
rect 12249 312 12254 368
rect 12310 312 25146 368
rect 12249 310 25146 312
rect 25270 368 28507 370
rect 25270 312 28446 368
rect 28502 312 28507 368
rect 25270 310 28507 312
rect 12249 307 12315 310
rect 10777 234 10843 237
rect 24894 234 24900 236
rect 10777 232 24900 234
rect 10777 176 10782 232
rect 10838 176 24900 232
rect 10777 174 24900 176
rect 10777 171 10843 174
rect 24894 172 24900 174
rect 24964 172 24970 236
rect 25086 234 25146 310
rect 28441 307 28507 310
rect 28257 234 28323 237
rect 25086 232 28323 234
rect 25086 176 28262 232
rect 28318 176 28323 232
rect 25086 174 28323 176
rect 28257 171 28323 174
<< via3 >>
rect 11554 8732 11618 8736
rect 11554 8676 11558 8732
rect 11558 8676 11614 8732
rect 11614 8676 11618 8732
rect 11554 8672 11618 8676
rect 11634 8732 11698 8736
rect 11634 8676 11638 8732
rect 11638 8676 11694 8732
rect 11694 8676 11698 8732
rect 11634 8672 11698 8676
rect 11714 8732 11778 8736
rect 11714 8676 11718 8732
rect 11718 8676 11774 8732
rect 11774 8676 11778 8732
rect 11714 8672 11778 8676
rect 11794 8732 11858 8736
rect 11794 8676 11798 8732
rect 11798 8676 11854 8732
rect 11854 8676 11858 8732
rect 11794 8672 11858 8676
rect 22157 8732 22221 8736
rect 22157 8676 22161 8732
rect 22161 8676 22217 8732
rect 22217 8676 22221 8732
rect 22157 8672 22221 8676
rect 22237 8732 22301 8736
rect 22237 8676 22241 8732
rect 22241 8676 22297 8732
rect 22297 8676 22301 8732
rect 22237 8672 22301 8676
rect 22317 8732 22381 8736
rect 22317 8676 22321 8732
rect 22321 8676 22377 8732
rect 22377 8676 22381 8732
rect 22317 8672 22381 8676
rect 22397 8732 22461 8736
rect 22397 8676 22401 8732
rect 22401 8676 22457 8732
rect 22457 8676 22461 8732
rect 22397 8672 22461 8676
rect 32760 8732 32824 8736
rect 32760 8676 32764 8732
rect 32764 8676 32820 8732
rect 32820 8676 32824 8732
rect 32760 8672 32824 8676
rect 32840 8732 32904 8736
rect 32840 8676 32844 8732
rect 32844 8676 32900 8732
rect 32900 8676 32904 8732
rect 32840 8672 32904 8676
rect 32920 8732 32984 8736
rect 32920 8676 32924 8732
rect 32924 8676 32980 8732
rect 32980 8676 32984 8732
rect 32920 8672 32984 8676
rect 33000 8732 33064 8736
rect 33000 8676 33004 8732
rect 33004 8676 33060 8732
rect 33060 8676 33064 8732
rect 33000 8672 33064 8676
rect 43363 8732 43427 8736
rect 43363 8676 43367 8732
rect 43367 8676 43423 8732
rect 43423 8676 43427 8732
rect 43363 8672 43427 8676
rect 43443 8732 43507 8736
rect 43443 8676 43447 8732
rect 43447 8676 43503 8732
rect 43503 8676 43507 8732
rect 43443 8672 43507 8676
rect 43523 8732 43587 8736
rect 43523 8676 43527 8732
rect 43527 8676 43583 8732
rect 43583 8676 43587 8732
rect 43523 8672 43587 8676
rect 43603 8732 43667 8736
rect 43603 8676 43607 8732
rect 43607 8676 43663 8732
rect 43663 8676 43667 8732
rect 43603 8672 43667 8676
rect 27844 8468 27908 8532
rect 29500 8332 29564 8396
rect 6253 8188 6317 8192
rect 6253 8132 6257 8188
rect 6257 8132 6313 8188
rect 6313 8132 6317 8188
rect 6253 8128 6317 8132
rect 6333 8188 6397 8192
rect 6333 8132 6337 8188
rect 6337 8132 6393 8188
rect 6393 8132 6397 8188
rect 6333 8128 6397 8132
rect 6413 8188 6477 8192
rect 6413 8132 6417 8188
rect 6417 8132 6473 8188
rect 6473 8132 6477 8188
rect 6413 8128 6477 8132
rect 6493 8188 6557 8192
rect 6493 8132 6497 8188
rect 6497 8132 6553 8188
rect 6553 8132 6557 8188
rect 6493 8128 6557 8132
rect 16856 8188 16920 8192
rect 16856 8132 16860 8188
rect 16860 8132 16916 8188
rect 16916 8132 16920 8188
rect 16856 8128 16920 8132
rect 16936 8188 17000 8192
rect 16936 8132 16940 8188
rect 16940 8132 16996 8188
rect 16996 8132 17000 8188
rect 16936 8128 17000 8132
rect 17016 8188 17080 8192
rect 17016 8132 17020 8188
rect 17020 8132 17076 8188
rect 17076 8132 17080 8188
rect 17016 8128 17080 8132
rect 17096 8188 17160 8192
rect 17096 8132 17100 8188
rect 17100 8132 17156 8188
rect 17156 8132 17160 8188
rect 17096 8128 17160 8132
rect 27459 8188 27523 8192
rect 27459 8132 27463 8188
rect 27463 8132 27519 8188
rect 27519 8132 27523 8188
rect 27459 8128 27523 8132
rect 27539 8188 27603 8192
rect 27539 8132 27543 8188
rect 27543 8132 27599 8188
rect 27599 8132 27603 8188
rect 27539 8128 27603 8132
rect 27619 8188 27683 8192
rect 27619 8132 27623 8188
rect 27623 8132 27679 8188
rect 27679 8132 27683 8188
rect 27619 8128 27683 8132
rect 27699 8188 27763 8192
rect 27699 8132 27703 8188
rect 27703 8132 27759 8188
rect 27759 8132 27763 8188
rect 27699 8128 27763 8132
rect 38062 8188 38126 8192
rect 38062 8132 38066 8188
rect 38066 8132 38122 8188
rect 38122 8132 38126 8188
rect 38062 8128 38126 8132
rect 38142 8188 38206 8192
rect 38142 8132 38146 8188
rect 38146 8132 38202 8188
rect 38202 8132 38206 8188
rect 38142 8128 38206 8132
rect 38222 8188 38286 8192
rect 38222 8132 38226 8188
rect 38226 8132 38282 8188
rect 38282 8132 38286 8188
rect 38222 8128 38286 8132
rect 38302 8188 38366 8192
rect 38302 8132 38306 8188
rect 38306 8132 38362 8188
rect 38362 8132 38366 8188
rect 38302 8128 38366 8132
rect 11554 7644 11618 7648
rect 11554 7588 11558 7644
rect 11558 7588 11614 7644
rect 11614 7588 11618 7644
rect 11554 7584 11618 7588
rect 11634 7644 11698 7648
rect 11634 7588 11638 7644
rect 11638 7588 11694 7644
rect 11694 7588 11698 7644
rect 11634 7584 11698 7588
rect 11714 7644 11778 7648
rect 11714 7588 11718 7644
rect 11718 7588 11774 7644
rect 11774 7588 11778 7644
rect 11714 7584 11778 7588
rect 11794 7644 11858 7648
rect 11794 7588 11798 7644
rect 11798 7588 11854 7644
rect 11854 7588 11858 7644
rect 11794 7584 11858 7588
rect 22157 7644 22221 7648
rect 22157 7588 22161 7644
rect 22161 7588 22217 7644
rect 22217 7588 22221 7644
rect 22157 7584 22221 7588
rect 22237 7644 22301 7648
rect 22237 7588 22241 7644
rect 22241 7588 22297 7644
rect 22297 7588 22301 7644
rect 22237 7584 22301 7588
rect 22317 7644 22381 7648
rect 22317 7588 22321 7644
rect 22321 7588 22377 7644
rect 22377 7588 22381 7644
rect 22317 7584 22381 7588
rect 22397 7644 22461 7648
rect 22397 7588 22401 7644
rect 22401 7588 22457 7644
rect 22457 7588 22461 7644
rect 22397 7584 22461 7588
rect 32760 7644 32824 7648
rect 32760 7588 32764 7644
rect 32764 7588 32820 7644
rect 32820 7588 32824 7644
rect 32760 7584 32824 7588
rect 32840 7644 32904 7648
rect 32840 7588 32844 7644
rect 32844 7588 32900 7644
rect 32900 7588 32904 7644
rect 32840 7584 32904 7588
rect 32920 7644 32984 7648
rect 32920 7588 32924 7644
rect 32924 7588 32980 7644
rect 32980 7588 32984 7644
rect 32920 7584 32984 7588
rect 33000 7644 33064 7648
rect 33000 7588 33004 7644
rect 33004 7588 33060 7644
rect 33060 7588 33064 7644
rect 33000 7584 33064 7588
rect 43363 7644 43427 7648
rect 43363 7588 43367 7644
rect 43367 7588 43423 7644
rect 43423 7588 43427 7644
rect 43363 7584 43427 7588
rect 43443 7644 43507 7648
rect 43443 7588 43447 7644
rect 43447 7588 43503 7644
rect 43503 7588 43507 7644
rect 43443 7584 43507 7588
rect 43523 7644 43587 7648
rect 43523 7588 43527 7644
rect 43527 7588 43583 7644
rect 43583 7588 43587 7644
rect 43523 7584 43587 7588
rect 43603 7644 43667 7648
rect 43603 7588 43607 7644
rect 43607 7588 43663 7644
rect 43663 7588 43667 7644
rect 43603 7584 43667 7588
rect 6253 7100 6317 7104
rect 6253 7044 6257 7100
rect 6257 7044 6313 7100
rect 6313 7044 6317 7100
rect 6253 7040 6317 7044
rect 6333 7100 6397 7104
rect 6333 7044 6337 7100
rect 6337 7044 6393 7100
rect 6393 7044 6397 7100
rect 6333 7040 6397 7044
rect 6413 7100 6477 7104
rect 6413 7044 6417 7100
rect 6417 7044 6473 7100
rect 6473 7044 6477 7100
rect 6413 7040 6477 7044
rect 6493 7100 6557 7104
rect 6493 7044 6497 7100
rect 6497 7044 6553 7100
rect 6553 7044 6557 7100
rect 6493 7040 6557 7044
rect 16856 7100 16920 7104
rect 16856 7044 16860 7100
rect 16860 7044 16916 7100
rect 16916 7044 16920 7100
rect 16856 7040 16920 7044
rect 16936 7100 17000 7104
rect 16936 7044 16940 7100
rect 16940 7044 16996 7100
rect 16996 7044 17000 7100
rect 16936 7040 17000 7044
rect 17016 7100 17080 7104
rect 17016 7044 17020 7100
rect 17020 7044 17076 7100
rect 17076 7044 17080 7100
rect 17016 7040 17080 7044
rect 17096 7100 17160 7104
rect 17096 7044 17100 7100
rect 17100 7044 17156 7100
rect 17156 7044 17160 7100
rect 17096 7040 17160 7044
rect 27459 7100 27523 7104
rect 27459 7044 27463 7100
rect 27463 7044 27519 7100
rect 27519 7044 27523 7100
rect 27459 7040 27523 7044
rect 27539 7100 27603 7104
rect 27539 7044 27543 7100
rect 27543 7044 27599 7100
rect 27599 7044 27603 7100
rect 27539 7040 27603 7044
rect 27619 7100 27683 7104
rect 27619 7044 27623 7100
rect 27623 7044 27679 7100
rect 27679 7044 27683 7100
rect 27619 7040 27683 7044
rect 27699 7100 27763 7104
rect 27699 7044 27703 7100
rect 27703 7044 27759 7100
rect 27759 7044 27763 7100
rect 27699 7040 27763 7044
rect 38062 7100 38126 7104
rect 38062 7044 38066 7100
rect 38066 7044 38122 7100
rect 38122 7044 38126 7100
rect 38062 7040 38126 7044
rect 38142 7100 38206 7104
rect 38142 7044 38146 7100
rect 38146 7044 38202 7100
rect 38202 7044 38206 7100
rect 38142 7040 38206 7044
rect 38222 7100 38286 7104
rect 38222 7044 38226 7100
rect 38226 7044 38282 7100
rect 38282 7044 38286 7100
rect 38222 7040 38286 7044
rect 38302 7100 38366 7104
rect 38302 7044 38306 7100
rect 38306 7044 38362 7100
rect 38362 7044 38366 7100
rect 38302 7040 38366 7044
rect 11554 6556 11618 6560
rect 11554 6500 11558 6556
rect 11558 6500 11614 6556
rect 11614 6500 11618 6556
rect 11554 6496 11618 6500
rect 11634 6556 11698 6560
rect 11634 6500 11638 6556
rect 11638 6500 11694 6556
rect 11694 6500 11698 6556
rect 11634 6496 11698 6500
rect 11714 6556 11778 6560
rect 11714 6500 11718 6556
rect 11718 6500 11774 6556
rect 11774 6500 11778 6556
rect 11714 6496 11778 6500
rect 11794 6556 11858 6560
rect 11794 6500 11798 6556
rect 11798 6500 11854 6556
rect 11854 6500 11858 6556
rect 11794 6496 11858 6500
rect 22157 6556 22221 6560
rect 22157 6500 22161 6556
rect 22161 6500 22217 6556
rect 22217 6500 22221 6556
rect 22157 6496 22221 6500
rect 22237 6556 22301 6560
rect 22237 6500 22241 6556
rect 22241 6500 22297 6556
rect 22297 6500 22301 6556
rect 22237 6496 22301 6500
rect 22317 6556 22381 6560
rect 22317 6500 22321 6556
rect 22321 6500 22377 6556
rect 22377 6500 22381 6556
rect 22317 6496 22381 6500
rect 22397 6556 22461 6560
rect 22397 6500 22401 6556
rect 22401 6500 22457 6556
rect 22457 6500 22461 6556
rect 22397 6496 22461 6500
rect 32760 6556 32824 6560
rect 32760 6500 32764 6556
rect 32764 6500 32820 6556
rect 32820 6500 32824 6556
rect 32760 6496 32824 6500
rect 32840 6556 32904 6560
rect 32840 6500 32844 6556
rect 32844 6500 32900 6556
rect 32900 6500 32904 6556
rect 32840 6496 32904 6500
rect 32920 6556 32984 6560
rect 32920 6500 32924 6556
rect 32924 6500 32980 6556
rect 32980 6500 32984 6556
rect 32920 6496 32984 6500
rect 33000 6556 33064 6560
rect 33000 6500 33004 6556
rect 33004 6500 33060 6556
rect 33060 6500 33064 6556
rect 33000 6496 33064 6500
rect 43363 6556 43427 6560
rect 43363 6500 43367 6556
rect 43367 6500 43423 6556
rect 43423 6500 43427 6556
rect 43363 6496 43427 6500
rect 43443 6556 43507 6560
rect 43443 6500 43447 6556
rect 43447 6500 43503 6556
rect 43503 6500 43507 6556
rect 43443 6496 43507 6500
rect 43523 6556 43587 6560
rect 43523 6500 43527 6556
rect 43527 6500 43583 6556
rect 43583 6500 43587 6556
rect 43523 6496 43587 6500
rect 43603 6556 43667 6560
rect 43603 6500 43607 6556
rect 43607 6500 43663 6556
rect 43663 6500 43667 6556
rect 43603 6496 43667 6500
rect 6253 6012 6317 6016
rect 6253 5956 6257 6012
rect 6257 5956 6313 6012
rect 6313 5956 6317 6012
rect 6253 5952 6317 5956
rect 6333 6012 6397 6016
rect 6333 5956 6337 6012
rect 6337 5956 6393 6012
rect 6393 5956 6397 6012
rect 6333 5952 6397 5956
rect 6413 6012 6477 6016
rect 6413 5956 6417 6012
rect 6417 5956 6473 6012
rect 6473 5956 6477 6012
rect 6413 5952 6477 5956
rect 6493 6012 6557 6016
rect 6493 5956 6497 6012
rect 6497 5956 6553 6012
rect 6553 5956 6557 6012
rect 6493 5952 6557 5956
rect 16856 6012 16920 6016
rect 16856 5956 16860 6012
rect 16860 5956 16916 6012
rect 16916 5956 16920 6012
rect 16856 5952 16920 5956
rect 16936 6012 17000 6016
rect 16936 5956 16940 6012
rect 16940 5956 16996 6012
rect 16996 5956 17000 6012
rect 16936 5952 17000 5956
rect 17016 6012 17080 6016
rect 17016 5956 17020 6012
rect 17020 5956 17076 6012
rect 17076 5956 17080 6012
rect 17016 5952 17080 5956
rect 17096 6012 17160 6016
rect 17096 5956 17100 6012
rect 17100 5956 17156 6012
rect 17156 5956 17160 6012
rect 17096 5952 17160 5956
rect 27459 6012 27523 6016
rect 27459 5956 27463 6012
rect 27463 5956 27519 6012
rect 27519 5956 27523 6012
rect 27459 5952 27523 5956
rect 27539 6012 27603 6016
rect 27539 5956 27543 6012
rect 27543 5956 27599 6012
rect 27599 5956 27603 6012
rect 27539 5952 27603 5956
rect 27619 6012 27683 6016
rect 27619 5956 27623 6012
rect 27623 5956 27679 6012
rect 27679 5956 27683 6012
rect 27619 5952 27683 5956
rect 27699 6012 27763 6016
rect 27699 5956 27703 6012
rect 27703 5956 27759 6012
rect 27759 5956 27763 6012
rect 27699 5952 27763 5956
rect 38062 6012 38126 6016
rect 38062 5956 38066 6012
rect 38066 5956 38122 6012
rect 38122 5956 38126 6012
rect 38062 5952 38126 5956
rect 38142 6012 38206 6016
rect 38142 5956 38146 6012
rect 38146 5956 38202 6012
rect 38202 5956 38206 6012
rect 38142 5952 38206 5956
rect 38222 6012 38286 6016
rect 38222 5956 38226 6012
rect 38226 5956 38282 6012
rect 38282 5956 38286 6012
rect 38222 5952 38286 5956
rect 38302 6012 38366 6016
rect 38302 5956 38306 6012
rect 38306 5956 38362 6012
rect 38362 5956 38366 6012
rect 38302 5952 38366 5956
rect 11554 5468 11618 5472
rect 11554 5412 11558 5468
rect 11558 5412 11614 5468
rect 11614 5412 11618 5468
rect 11554 5408 11618 5412
rect 11634 5468 11698 5472
rect 11634 5412 11638 5468
rect 11638 5412 11694 5468
rect 11694 5412 11698 5468
rect 11634 5408 11698 5412
rect 11714 5468 11778 5472
rect 11714 5412 11718 5468
rect 11718 5412 11774 5468
rect 11774 5412 11778 5468
rect 11714 5408 11778 5412
rect 11794 5468 11858 5472
rect 11794 5412 11798 5468
rect 11798 5412 11854 5468
rect 11854 5412 11858 5468
rect 11794 5408 11858 5412
rect 22157 5468 22221 5472
rect 22157 5412 22161 5468
rect 22161 5412 22217 5468
rect 22217 5412 22221 5468
rect 22157 5408 22221 5412
rect 22237 5468 22301 5472
rect 22237 5412 22241 5468
rect 22241 5412 22297 5468
rect 22297 5412 22301 5468
rect 22237 5408 22301 5412
rect 22317 5468 22381 5472
rect 22317 5412 22321 5468
rect 22321 5412 22377 5468
rect 22377 5412 22381 5468
rect 22317 5408 22381 5412
rect 22397 5468 22461 5472
rect 22397 5412 22401 5468
rect 22401 5412 22457 5468
rect 22457 5412 22461 5468
rect 22397 5408 22461 5412
rect 32760 5468 32824 5472
rect 32760 5412 32764 5468
rect 32764 5412 32820 5468
rect 32820 5412 32824 5468
rect 32760 5408 32824 5412
rect 32840 5468 32904 5472
rect 32840 5412 32844 5468
rect 32844 5412 32900 5468
rect 32900 5412 32904 5468
rect 32840 5408 32904 5412
rect 32920 5468 32984 5472
rect 32920 5412 32924 5468
rect 32924 5412 32980 5468
rect 32980 5412 32984 5468
rect 32920 5408 32984 5412
rect 33000 5468 33064 5472
rect 33000 5412 33004 5468
rect 33004 5412 33060 5468
rect 33060 5412 33064 5468
rect 33000 5408 33064 5412
rect 43363 5468 43427 5472
rect 43363 5412 43367 5468
rect 43367 5412 43423 5468
rect 43423 5412 43427 5468
rect 43363 5408 43427 5412
rect 43443 5468 43507 5472
rect 43443 5412 43447 5468
rect 43447 5412 43503 5468
rect 43503 5412 43507 5468
rect 43443 5408 43507 5412
rect 43523 5468 43587 5472
rect 43523 5412 43527 5468
rect 43527 5412 43583 5468
rect 43583 5412 43587 5468
rect 43523 5408 43587 5412
rect 43603 5468 43667 5472
rect 43603 5412 43607 5468
rect 43607 5412 43663 5468
rect 43663 5412 43667 5468
rect 43603 5408 43667 5412
rect 6253 4924 6317 4928
rect 6253 4868 6257 4924
rect 6257 4868 6313 4924
rect 6313 4868 6317 4924
rect 6253 4864 6317 4868
rect 6333 4924 6397 4928
rect 6333 4868 6337 4924
rect 6337 4868 6393 4924
rect 6393 4868 6397 4924
rect 6333 4864 6397 4868
rect 6413 4924 6477 4928
rect 6413 4868 6417 4924
rect 6417 4868 6473 4924
rect 6473 4868 6477 4924
rect 6413 4864 6477 4868
rect 6493 4924 6557 4928
rect 6493 4868 6497 4924
rect 6497 4868 6553 4924
rect 6553 4868 6557 4924
rect 6493 4864 6557 4868
rect 16856 4924 16920 4928
rect 16856 4868 16860 4924
rect 16860 4868 16916 4924
rect 16916 4868 16920 4924
rect 16856 4864 16920 4868
rect 16936 4924 17000 4928
rect 16936 4868 16940 4924
rect 16940 4868 16996 4924
rect 16996 4868 17000 4924
rect 16936 4864 17000 4868
rect 17016 4924 17080 4928
rect 17016 4868 17020 4924
rect 17020 4868 17076 4924
rect 17076 4868 17080 4924
rect 17016 4864 17080 4868
rect 17096 4924 17160 4928
rect 17096 4868 17100 4924
rect 17100 4868 17156 4924
rect 17156 4868 17160 4924
rect 17096 4864 17160 4868
rect 27459 4924 27523 4928
rect 27459 4868 27463 4924
rect 27463 4868 27519 4924
rect 27519 4868 27523 4924
rect 27459 4864 27523 4868
rect 27539 4924 27603 4928
rect 27539 4868 27543 4924
rect 27543 4868 27599 4924
rect 27599 4868 27603 4924
rect 27539 4864 27603 4868
rect 27619 4924 27683 4928
rect 27619 4868 27623 4924
rect 27623 4868 27679 4924
rect 27679 4868 27683 4924
rect 27619 4864 27683 4868
rect 27699 4924 27763 4928
rect 27699 4868 27703 4924
rect 27703 4868 27759 4924
rect 27759 4868 27763 4924
rect 27699 4864 27763 4868
rect 38062 4924 38126 4928
rect 38062 4868 38066 4924
rect 38066 4868 38122 4924
rect 38122 4868 38126 4924
rect 38062 4864 38126 4868
rect 38142 4924 38206 4928
rect 38142 4868 38146 4924
rect 38146 4868 38202 4924
rect 38202 4868 38206 4924
rect 38142 4864 38206 4868
rect 38222 4924 38286 4928
rect 38222 4868 38226 4924
rect 38226 4868 38282 4924
rect 38282 4868 38286 4924
rect 38222 4864 38286 4868
rect 38302 4924 38366 4928
rect 38302 4868 38306 4924
rect 38306 4868 38362 4924
rect 38362 4868 38366 4924
rect 38302 4864 38366 4868
rect 16068 4524 16132 4588
rect 11554 4380 11618 4384
rect 11554 4324 11558 4380
rect 11558 4324 11614 4380
rect 11614 4324 11618 4380
rect 11554 4320 11618 4324
rect 11634 4380 11698 4384
rect 11634 4324 11638 4380
rect 11638 4324 11694 4380
rect 11694 4324 11698 4380
rect 11634 4320 11698 4324
rect 11714 4380 11778 4384
rect 11714 4324 11718 4380
rect 11718 4324 11774 4380
rect 11774 4324 11778 4380
rect 11714 4320 11778 4324
rect 11794 4380 11858 4384
rect 11794 4324 11798 4380
rect 11798 4324 11854 4380
rect 11854 4324 11858 4380
rect 11794 4320 11858 4324
rect 22157 4380 22221 4384
rect 22157 4324 22161 4380
rect 22161 4324 22217 4380
rect 22217 4324 22221 4380
rect 22157 4320 22221 4324
rect 22237 4380 22301 4384
rect 22237 4324 22241 4380
rect 22241 4324 22297 4380
rect 22297 4324 22301 4380
rect 22237 4320 22301 4324
rect 22317 4380 22381 4384
rect 22317 4324 22321 4380
rect 22321 4324 22377 4380
rect 22377 4324 22381 4380
rect 22317 4320 22381 4324
rect 22397 4380 22461 4384
rect 22397 4324 22401 4380
rect 22401 4324 22457 4380
rect 22457 4324 22461 4380
rect 22397 4320 22461 4324
rect 32760 4380 32824 4384
rect 32760 4324 32764 4380
rect 32764 4324 32820 4380
rect 32820 4324 32824 4380
rect 32760 4320 32824 4324
rect 32840 4380 32904 4384
rect 32840 4324 32844 4380
rect 32844 4324 32900 4380
rect 32900 4324 32904 4380
rect 32840 4320 32904 4324
rect 32920 4380 32984 4384
rect 32920 4324 32924 4380
rect 32924 4324 32980 4380
rect 32980 4324 32984 4380
rect 32920 4320 32984 4324
rect 33000 4380 33064 4384
rect 33000 4324 33004 4380
rect 33004 4324 33060 4380
rect 33060 4324 33064 4380
rect 33000 4320 33064 4324
rect 43363 4380 43427 4384
rect 43363 4324 43367 4380
rect 43367 4324 43423 4380
rect 43423 4324 43427 4380
rect 43363 4320 43427 4324
rect 43443 4380 43507 4384
rect 43443 4324 43447 4380
rect 43447 4324 43503 4380
rect 43503 4324 43507 4380
rect 43443 4320 43507 4324
rect 43523 4380 43587 4384
rect 43523 4324 43527 4380
rect 43527 4324 43583 4380
rect 43583 4324 43587 4380
rect 43523 4320 43587 4324
rect 43603 4380 43667 4384
rect 43603 4324 43607 4380
rect 43607 4324 43663 4380
rect 43663 4324 43667 4380
rect 43603 4320 43667 4324
rect 31708 3844 31772 3908
rect 6253 3836 6317 3840
rect 6253 3780 6257 3836
rect 6257 3780 6313 3836
rect 6313 3780 6317 3836
rect 6253 3776 6317 3780
rect 6333 3836 6397 3840
rect 6333 3780 6337 3836
rect 6337 3780 6393 3836
rect 6393 3780 6397 3836
rect 6333 3776 6397 3780
rect 6413 3836 6477 3840
rect 6413 3780 6417 3836
rect 6417 3780 6473 3836
rect 6473 3780 6477 3836
rect 6413 3776 6477 3780
rect 6493 3836 6557 3840
rect 6493 3780 6497 3836
rect 6497 3780 6553 3836
rect 6553 3780 6557 3836
rect 6493 3776 6557 3780
rect 16856 3836 16920 3840
rect 16856 3780 16860 3836
rect 16860 3780 16916 3836
rect 16916 3780 16920 3836
rect 16856 3776 16920 3780
rect 16936 3836 17000 3840
rect 16936 3780 16940 3836
rect 16940 3780 16996 3836
rect 16996 3780 17000 3836
rect 16936 3776 17000 3780
rect 17016 3836 17080 3840
rect 17016 3780 17020 3836
rect 17020 3780 17076 3836
rect 17076 3780 17080 3836
rect 17016 3776 17080 3780
rect 17096 3836 17160 3840
rect 17096 3780 17100 3836
rect 17100 3780 17156 3836
rect 17156 3780 17160 3836
rect 17096 3776 17160 3780
rect 27459 3836 27523 3840
rect 27459 3780 27463 3836
rect 27463 3780 27519 3836
rect 27519 3780 27523 3836
rect 27459 3776 27523 3780
rect 27539 3836 27603 3840
rect 27539 3780 27543 3836
rect 27543 3780 27599 3836
rect 27599 3780 27603 3836
rect 27539 3776 27603 3780
rect 27619 3836 27683 3840
rect 27619 3780 27623 3836
rect 27623 3780 27679 3836
rect 27679 3780 27683 3836
rect 27619 3776 27683 3780
rect 27699 3836 27763 3840
rect 27699 3780 27703 3836
rect 27703 3780 27759 3836
rect 27759 3780 27763 3836
rect 27699 3776 27763 3780
rect 38062 3836 38126 3840
rect 38062 3780 38066 3836
rect 38066 3780 38122 3836
rect 38122 3780 38126 3836
rect 38062 3776 38126 3780
rect 38142 3836 38206 3840
rect 38142 3780 38146 3836
rect 38146 3780 38202 3836
rect 38202 3780 38206 3836
rect 38142 3776 38206 3780
rect 38222 3836 38286 3840
rect 38222 3780 38226 3836
rect 38226 3780 38282 3836
rect 38282 3780 38286 3836
rect 38222 3776 38286 3780
rect 38302 3836 38366 3840
rect 38302 3780 38306 3836
rect 38306 3780 38362 3836
rect 38362 3780 38366 3836
rect 38302 3776 38366 3780
rect 34652 3436 34716 3500
rect 11554 3292 11618 3296
rect 11554 3236 11558 3292
rect 11558 3236 11614 3292
rect 11614 3236 11618 3292
rect 11554 3232 11618 3236
rect 11634 3292 11698 3296
rect 11634 3236 11638 3292
rect 11638 3236 11694 3292
rect 11694 3236 11698 3292
rect 11634 3232 11698 3236
rect 11714 3292 11778 3296
rect 11714 3236 11718 3292
rect 11718 3236 11774 3292
rect 11774 3236 11778 3292
rect 11714 3232 11778 3236
rect 11794 3292 11858 3296
rect 11794 3236 11798 3292
rect 11798 3236 11854 3292
rect 11854 3236 11858 3292
rect 11794 3232 11858 3236
rect 22157 3292 22221 3296
rect 22157 3236 22161 3292
rect 22161 3236 22217 3292
rect 22217 3236 22221 3292
rect 22157 3232 22221 3236
rect 22237 3292 22301 3296
rect 22237 3236 22241 3292
rect 22241 3236 22297 3292
rect 22297 3236 22301 3292
rect 22237 3232 22301 3236
rect 22317 3292 22381 3296
rect 22317 3236 22321 3292
rect 22321 3236 22377 3292
rect 22377 3236 22381 3292
rect 22317 3232 22381 3236
rect 22397 3292 22461 3296
rect 22397 3236 22401 3292
rect 22401 3236 22457 3292
rect 22457 3236 22461 3292
rect 22397 3232 22461 3236
rect 32760 3292 32824 3296
rect 32760 3236 32764 3292
rect 32764 3236 32820 3292
rect 32820 3236 32824 3292
rect 32760 3232 32824 3236
rect 32840 3292 32904 3296
rect 32840 3236 32844 3292
rect 32844 3236 32900 3292
rect 32900 3236 32904 3292
rect 32840 3232 32904 3236
rect 32920 3292 32984 3296
rect 32920 3236 32924 3292
rect 32924 3236 32980 3292
rect 32980 3236 32984 3292
rect 32920 3232 32984 3236
rect 33000 3292 33064 3296
rect 33000 3236 33004 3292
rect 33004 3236 33060 3292
rect 33060 3236 33064 3292
rect 33000 3232 33064 3236
rect 43363 3292 43427 3296
rect 43363 3236 43367 3292
rect 43367 3236 43423 3292
rect 43423 3236 43427 3292
rect 43363 3232 43427 3236
rect 43443 3292 43507 3296
rect 43443 3236 43447 3292
rect 43447 3236 43503 3292
rect 43503 3236 43507 3292
rect 43443 3232 43507 3236
rect 43523 3292 43587 3296
rect 43523 3236 43527 3292
rect 43527 3236 43583 3292
rect 43583 3236 43587 3292
rect 43523 3232 43587 3236
rect 43603 3292 43667 3296
rect 43603 3236 43607 3292
rect 43607 3236 43663 3292
rect 43663 3236 43667 3292
rect 43603 3232 43667 3236
rect 27292 2756 27356 2820
rect 30236 2816 30300 2820
rect 30236 2760 30250 2816
rect 30250 2760 30300 2816
rect 30236 2756 30300 2760
rect 6253 2748 6317 2752
rect 6253 2692 6257 2748
rect 6257 2692 6313 2748
rect 6313 2692 6317 2748
rect 6253 2688 6317 2692
rect 6333 2748 6397 2752
rect 6333 2692 6337 2748
rect 6337 2692 6393 2748
rect 6393 2692 6397 2748
rect 6333 2688 6397 2692
rect 6413 2748 6477 2752
rect 6413 2692 6417 2748
rect 6417 2692 6473 2748
rect 6473 2692 6477 2748
rect 6413 2688 6477 2692
rect 6493 2748 6557 2752
rect 6493 2692 6497 2748
rect 6497 2692 6553 2748
rect 6553 2692 6557 2748
rect 6493 2688 6557 2692
rect 16856 2748 16920 2752
rect 16856 2692 16860 2748
rect 16860 2692 16916 2748
rect 16916 2692 16920 2748
rect 16856 2688 16920 2692
rect 16936 2748 17000 2752
rect 16936 2692 16940 2748
rect 16940 2692 16996 2748
rect 16996 2692 17000 2748
rect 16936 2688 17000 2692
rect 17016 2748 17080 2752
rect 17016 2692 17020 2748
rect 17020 2692 17076 2748
rect 17076 2692 17080 2748
rect 17016 2688 17080 2692
rect 17096 2748 17160 2752
rect 17096 2692 17100 2748
rect 17100 2692 17156 2748
rect 17156 2692 17160 2748
rect 17096 2688 17160 2692
rect 27459 2748 27523 2752
rect 27459 2692 27463 2748
rect 27463 2692 27519 2748
rect 27519 2692 27523 2748
rect 27459 2688 27523 2692
rect 27539 2748 27603 2752
rect 27539 2692 27543 2748
rect 27543 2692 27599 2748
rect 27599 2692 27603 2748
rect 27539 2688 27603 2692
rect 27619 2748 27683 2752
rect 27619 2692 27623 2748
rect 27623 2692 27679 2748
rect 27679 2692 27683 2748
rect 27619 2688 27683 2692
rect 27699 2748 27763 2752
rect 27699 2692 27703 2748
rect 27703 2692 27759 2748
rect 27759 2692 27763 2748
rect 27699 2688 27763 2692
rect 38062 2748 38126 2752
rect 38062 2692 38066 2748
rect 38066 2692 38122 2748
rect 38122 2692 38126 2748
rect 38062 2688 38126 2692
rect 38142 2748 38206 2752
rect 38142 2692 38146 2748
rect 38146 2692 38202 2748
rect 38202 2692 38206 2748
rect 38142 2688 38206 2692
rect 38222 2748 38286 2752
rect 38222 2692 38226 2748
rect 38226 2692 38282 2748
rect 38282 2692 38286 2748
rect 38222 2688 38286 2692
rect 38302 2748 38366 2752
rect 38302 2692 38306 2748
rect 38306 2692 38362 2748
rect 38362 2692 38366 2748
rect 38302 2688 38366 2692
rect 27844 2680 27908 2684
rect 27844 2624 27894 2680
rect 27894 2624 27908 2680
rect 27844 2620 27908 2624
rect 29500 2620 29564 2684
rect 31708 2620 31772 2684
rect 24900 2484 24964 2548
rect 16068 2212 16132 2276
rect 11554 2204 11618 2208
rect 11554 2148 11558 2204
rect 11558 2148 11614 2204
rect 11614 2148 11618 2204
rect 11554 2144 11618 2148
rect 11634 2204 11698 2208
rect 11634 2148 11638 2204
rect 11638 2148 11694 2204
rect 11694 2148 11698 2204
rect 11634 2144 11698 2148
rect 11714 2204 11778 2208
rect 11714 2148 11718 2204
rect 11718 2148 11774 2204
rect 11774 2148 11778 2204
rect 11714 2144 11778 2148
rect 11794 2204 11858 2208
rect 11794 2148 11798 2204
rect 11798 2148 11854 2204
rect 11854 2148 11858 2204
rect 11794 2144 11858 2148
rect 22157 2204 22221 2208
rect 22157 2148 22161 2204
rect 22161 2148 22217 2204
rect 22217 2148 22221 2204
rect 22157 2144 22221 2148
rect 22237 2204 22301 2208
rect 22237 2148 22241 2204
rect 22241 2148 22297 2204
rect 22297 2148 22301 2204
rect 22237 2144 22301 2148
rect 22317 2204 22381 2208
rect 22317 2148 22321 2204
rect 22321 2148 22377 2204
rect 22377 2148 22381 2204
rect 22317 2144 22381 2148
rect 22397 2204 22461 2208
rect 22397 2148 22401 2204
rect 22401 2148 22457 2204
rect 22457 2148 22461 2204
rect 22397 2144 22461 2148
rect 32760 2204 32824 2208
rect 32760 2148 32764 2204
rect 32764 2148 32820 2204
rect 32820 2148 32824 2204
rect 32760 2144 32824 2148
rect 32840 2204 32904 2208
rect 32840 2148 32844 2204
rect 32844 2148 32900 2204
rect 32900 2148 32904 2204
rect 32840 2144 32904 2148
rect 32920 2204 32984 2208
rect 32920 2148 32924 2204
rect 32924 2148 32980 2204
rect 32980 2148 32984 2204
rect 32920 2144 32984 2148
rect 33000 2204 33064 2208
rect 33000 2148 33004 2204
rect 33004 2148 33060 2204
rect 33060 2148 33064 2204
rect 33000 2144 33064 2148
rect 43363 2204 43427 2208
rect 43363 2148 43367 2204
rect 43367 2148 43423 2204
rect 43423 2148 43427 2204
rect 43363 2144 43427 2148
rect 43443 2204 43507 2208
rect 43443 2148 43447 2204
rect 43447 2148 43503 2204
rect 43503 2148 43507 2204
rect 43443 2144 43507 2148
rect 43523 2204 43587 2208
rect 43523 2148 43527 2204
rect 43527 2148 43583 2204
rect 43583 2148 43587 2204
rect 43523 2144 43587 2148
rect 43603 2204 43667 2208
rect 43603 2148 43607 2204
rect 43607 2148 43663 2204
rect 43663 2148 43667 2204
rect 43603 2144 43667 2148
rect 27292 1940 27356 2004
rect 6253 1660 6317 1664
rect 6253 1604 6257 1660
rect 6257 1604 6313 1660
rect 6313 1604 6317 1660
rect 6253 1600 6317 1604
rect 6333 1660 6397 1664
rect 6333 1604 6337 1660
rect 6337 1604 6393 1660
rect 6393 1604 6397 1660
rect 6333 1600 6397 1604
rect 6413 1660 6477 1664
rect 6413 1604 6417 1660
rect 6417 1604 6473 1660
rect 6473 1604 6477 1660
rect 6413 1600 6477 1604
rect 6493 1660 6557 1664
rect 6493 1604 6497 1660
rect 6497 1604 6553 1660
rect 6553 1604 6557 1660
rect 6493 1600 6557 1604
rect 16856 1660 16920 1664
rect 16856 1604 16860 1660
rect 16860 1604 16916 1660
rect 16916 1604 16920 1660
rect 16856 1600 16920 1604
rect 16936 1660 17000 1664
rect 16936 1604 16940 1660
rect 16940 1604 16996 1660
rect 16996 1604 17000 1660
rect 16936 1600 17000 1604
rect 17016 1660 17080 1664
rect 17016 1604 17020 1660
rect 17020 1604 17076 1660
rect 17076 1604 17080 1660
rect 17016 1600 17080 1604
rect 17096 1660 17160 1664
rect 17096 1604 17100 1660
rect 17100 1604 17156 1660
rect 17156 1604 17160 1660
rect 17096 1600 17160 1604
rect 27459 1660 27523 1664
rect 27459 1604 27463 1660
rect 27463 1604 27519 1660
rect 27519 1604 27523 1660
rect 27459 1600 27523 1604
rect 27539 1660 27603 1664
rect 27539 1604 27543 1660
rect 27543 1604 27599 1660
rect 27599 1604 27603 1660
rect 27539 1600 27603 1604
rect 27619 1660 27683 1664
rect 27619 1604 27623 1660
rect 27623 1604 27679 1660
rect 27679 1604 27683 1660
rect 27619 1600 27683 1604
rect 27699 1660 27763 1664
rect 27699 1604 27703 1660
rect 27703 1604 27759 1660
rect 27759 1604 27763 1660
rect 27699 1600 27763 1604
rect 38062 1660 38126 1664
rect 38062 1604 38066 1660
rect 38066 1604 38122 1660
rect 38122 1604 38126 1660
rect 38062 1600 38126 1604
rect 38142 1660 38206 1664
rect 38142 1604 38146 1660
rect 38146 1604 38202 1660
rect 38202 1604 38206 1660
rect 38142 1600 38206 1604
rect 38222 1660 38286 1664
rect 38222 1604 38226 1660
rect 38226 1604 38282 1660
rect 38282 1604 38286 1660
rect 38222 1600 38286 1604
rect 38302 1660 38366 1664
rect 38302 1604 38306 1660
rect 38306 1604 38362 1660
rect 38362 1604 38366 1660
rect 38302 1600 38366 1604
rect 34652 1260 34716 1324
rect 11554 1116 11618 1120
rect 11554 1060 11558 1116
rect 11558 1060 11614 1116
rect 11614 1060 11618 1116
rect 11554 1056 11618 1060
rect 11634 1116 11698 1120
rect 11634 1060 11638 1116
rect 11638 1060 11694 1116
rect 11694 1060 11698 1116
rect 11634 1056 11698 1060
rect 11714 1116 11778 1120
rect 11714 1060 11718 1116
rect 11718 1060 11774 1116
rect 11774 1060 11778 1116
rect 11714 1056 11778 1060
rect 11794 1116 11858 1120
rect 11794 1060 11798 1116
rect 11798 1060 11854 1116
rect 11854 1060 11858 1116
rect 11794 1056 11858 1060
rect 22157 1116 22221 1120
rect 22157 1060 22161 1116
rect 22161 1060 22217 1116
rect 22217 1060 22221 1116
rect 22157 1056 22221 1060
rect 22237 1116 22301 1120
rect 22237 1060 22241 1116
rect 22241 1060 22297 1116
rect 22297 1060 22301 1116
rect 22237 1056 22301 1060
rect 22317 1116 22381 1120
rect 22317 1060 22321 1116
rect 22321 1060 22377 1116
rect 22377 1060 22381 1116
rect 22317 1056 22381 1060
rect 22397 1116 22461 1120
rect 22397 1060 22401 1116
rect 22401 1060 22457 1116
rect 22457 1060 22461 1116
rect 22397 1056 22461 1060
rect 32760 1116 32824 1120
rect 32760 1060 32764 1116
rect 32764 1060 32820 1116
rect 32820 1060 32824 1116
rect 32760 1056 32824 1060
rect 32840 1116 32904 1120
rect 32840 1060 32844 1116
rect 32844 1060 32900 1116
rect 32900 1060 32904 1116
rect 32840 1056 32904 1060
rect 32920 1116 32984 1120
rect 32920 1060 32924 1116
rect 32924 1060 32980 1116
rect 32980 1060 32984 1116
rect 32920 1056 32984 1060
rect 33000 1116 33064 1120
rect 33000 1060 33004 1116
rect 33004 1060 33060 1116
rect 33060 1060 33064 1116
rect 33000 1056 33064 1060
rect 43363 1116 43427 1120
rect 43363 1060 43367 1116
rect 43367 1060 43423 1116
rect 43423 1060 43427 1116
rect 43363 1056 43427 1060
rect 43443 1116 43507 1120
rect 43443 1060 43447 1116
rect 43447 1060 43503 1116
rect 43503 1060 43507 1116
rect 43443 1056 43507 1060
rect 43523 1116 43587 1120
rect 43523 1060 43527 1116
rect 43527 1060 43583 1116
rect 43583 1060 43587 1116
rect 43523 1056 43587 1060
rect 43603 1116 43667 1120
rect 43603 1060 43607 1116
rect 43607 1060 43663 1116
rect 43663 1060 43667 1116
rect 43603 1056 43667 1060
rect 30236 988 30300 1052
rect 24900 172 24964 236
<< metal4 >>
rect 6245 8192 6565 8752
rect 6245 8128 6253 8192
rect 6317 8128 6333 8192
rect 6397 8128 6413 8192
rect 6477 8128 6493 8192
rect 6557 8128 6565 8192
rect 6245 7104 6565 8128
rect 6245 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6565 7104
rect 6245 6016 6565 7040
rect 6245 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6565 6016
rect 6245 4928 6565 5952
rect 6245 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6565 4928
rect 6245 3840 6565 4864
rect 6245 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6565 3840
rect 6245 2752 6565 3776
rect 6245 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6565 2752
rect 6245 1664 6565 2688
rect 6245 1600 6253 1664
rect 6317 1600 6333 1664
rect 6397 1600 6413 1664
rect 6477 1600 6493 1664
rect 6557 1600 6565 1664
rect 6245 1040 6565 1600
rect 11546 8736 11866 8752
rect 11546 8672 11554 8736
rect 11618 8672 11634 8736
rect 11698 8672 11714 8736
rect 11778 8672 11794 8736
rect 11858 8672 11866 8736
rect 11546 7648 11866 8672
rect 11546 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11866 7648
rect 11546 6560 11866 7584
rect 11546 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11866 6560
rect 11546 5472 11866 6496
rect 11546 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11866 5472
rect 11546 4384 11866 5408
rect 16848 8192 17168 8752
rect 16848 8128 16856 8192
rect 16920 8128 16936 8192
rect 17000 8128 17016 8192
rect 17080 8128 17096 8192
rect 17160 8128 17168 8192
rect 16848 7104 17168 8128
rect 16848 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17168 7104
rect 16848 6016 17168 7040
rect 16848 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17168 6016
rect 16848 4928 17168 5952
rect 16848 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17168 4928
rect 16067 4588 16133 4589
rect 16067 4524 16068 4588
rect 16132 4524 16133 4588
rect 16067 4523 16133 4524
rect 11546 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11866 4384
rect 11546 3296 11866 4320
rect 11546 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11866 3296
rect 11546 2208 11866 3232
rect 16070 2277 16130 4523
rect 16848 3840 17168 4864
rect 16848 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17168 3840
rect 16848 2752 17168 3776
rect 16848 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17168 2752
rect 16067 2276 16133 2277
rect 16067 2212 16068 2276
rect 16132 2212 16133 2276
rect 16067 2211 16133 2212
rect 11546 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11866 2208
rect 11546 1120 11866 2144
rect 11546 1056 11554 1120
rect 11618 1056 11634 1120
rect 11698 1056 11714 1120
rect 11778 1056 11794 1120
rect 11858 1056 11866 1120
rect 11546 1040 11866 1056
rect 16848 1664 17168 2688
rect 16848 1600 16856 1664
rect 16920 1600 16936 1664
rect 17000 1600 17016 1664
rect 17080 1600 17096 1664
rect 17160 1600 17168 1664
rect 16848 1040 17168 1600
rect 22149 8736 22469 8752
rect 22149 8672 22157 8736
rect 22221 8672 22237 8736
rect 22301 8672 22317 8736
rect 22381 8672 22397 8736
rect 22461 8672 22469 8736
rect 22149 7648 22469 8672
rect 22149 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22469 7648
rect 22149 6560 22469 7584
rect 22149 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22469 6560
rect 22149 5472 22469 6496
rect 22149 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22469 5472
rect 22149 4384 22469 5408
rect 22149 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22469 4384
rect 22149 3296 22469 4320
rect 22149 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22469 3296
rect 22149 2208 22469 3232
rect 27451 8192 27771 8752
rect 32752 8736 33072 8752
rect 32752 8672 32760 8736
rect 32824 8672 32840 8736
rect 32904 8672 32920 8736
rect 32984 8672 33000 8736
rect 33064 8672 33072 8736
rect 27843 8532 27909 8533
rect 27843 8468 27844 8532
rect 27908 8468 27909 8532
rect 27843 8467 27909 8468
rect 27451 8128 27459 8192
rect 27523 8128 27539 8192
rect 27603 8128 27619 8192
rect 27683 8128 27699 8192
rect 27763 8128 27771 8192
rect 27451 7104 27771 8128
rect 27451 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27771 7104
rect 27451 6016 27771 7040
rect 27451 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27771 6016
rect 27451 4928 27771 5952
rect 27451 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27771 4928
rect 27451 3840 27771 4864
rect 27451 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27771 3840
rect 27291 2820 27357 2821
rect 27291 2756 27292 2820
rect 27356 2756 27357 2820
rect 27291 2755 27357 2756
rect 24899 2548 24965 2549
rect 24899 2484 24900 2548
rect 24964 2484 24965 2548
rect 24899 2483 24965 2484
rect 22149 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22469 2208
rect 22149 1120 22469 2144
rect 22149 1056 22157 1120
rect 22221 1056 22237 1120
rect 22301 1056 22317 1120
rect 22381 1056 22397 1120
rect 22461 1056 22469 1120
rect 22149 1040 22469 1056
rect 24902 237 24962 2483
rect 27294 2005 27354 2755
rect 27451 2752 27771 3776
rect 27451 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27771 2752
rect 27291 2004 27357 2005
rect 27291 1940 27292 2004
rect 27356 1940 27357 2004
rect 27291 1939 27357 1940
rect 27451 1664 27771 2688
rect 27846 2685 27906 8467
rect 29499 8396 29565 8397
rect 29499 8332 29500 8396
rect 29564 8332 29565 8396
rect 29499 8331 29565 8332
rect 29502 2685 29562 8331
rect 32752 7648 33072 8672
rect 32752 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33072 7648
rect 32752 6560 33072 7584
rect 32752 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33072 6560
rect 32752 5472 33072 6496
rect 32752 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33072 5472
rect 32752 4384 33072 5408
rect 32752 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33072 4384
rect 31707 3908 31773 3909
rect 31707 3844 31708 3908
rect 31772 3844 31773 3908
rect 31707 3843 31773 3844
rect 30235 2820 30301 2821
rect 30235 2756 30236 2820
rect 30300 2756 30301 2820
rect 30235 2755 30301 2756
rect 27843 2684 27909 2685
rect 27843 2620 27844 2684
rect 27908 2620 27909 2684
rect 27843 2619 27909 2620
rect 29499 2684 29565 2685
rect 29499 2620 29500 2684
rect 29564 2620 29565 2684
rect 29499 2619 29565 2620
rect 27451 1600 27459 1664
rect 27523 1600 27539 1664
rect 27603 1600 27619 1664
rect 27683 1600 27699 1664
rect 27763 1600 27771 1664
rect 27451 1040 27771 1600
rect 30238 1053 30298 2755
rect 31710 2685 31770 3843
rect 32752 3296 33072 4320
rect 38054 8192 38374 8752
rect 38054 8128 38062 8192
rect 38126 8128 38142 8192
rect 38206 8128 38222 8192
rect 38286 8128 38302 8192
rect 38366 8128 38374 8192
rect 38054 7104 38374 8128
rect 38054 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38374 7104
rect 38054 6016 38374 7040
rect 38054 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38374 6016
rect 38054 4928 38374 5952
rect 38054 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38374 4928
rect 38054 3840 38374 4864
rect 38054 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38374 3840
rect 34651 3500 34717 3501
rect 34651 3436 34652 3500
rect 34716 3436 34717 3500
rect 34651 3435 34717 3436
rect 32752 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33072 3296
rect 31707 2684 31773 2685
rect 31707 2620 31708 2684
rect 31772 2620 31773 2684
rect 31707 2619 31773 2620
rect 32752 2208 33072 3232
rect 32752 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33072 2208
rect 32752 1120 33072 2144
rect 34654 1325 34714 3435
rect 38054 2752 38374 3776
rect 38054 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38374 2752
rect 38054 1664 38374 2688
rect 38054 1600 38062 1664
rect 38126 1600 38142 1664
rect 38206 1600 38222 1664
rect 38286 1600 38302 1664
rect 38366 1600 38374 1664
rect 34651 1324 34717 1325
rect 34651 1260 34652 1324
rect 34716 1260 34717 1324
rect 34651 1259 34717 1260
rect 32752 1056 32760 1120
rect 32824 1056 32840 1120
rect 32904 1056 32920 1120
rect 32984 1056 33000 1120
rect 33064 1056 33072 1120
rect 30235 1052 30301 1053
rect 30235 988 30236 1052
rect 30300 988 30301 1052
rect 32752 1040 33072 1056
rect 38054 1040 38374 1600
rect 43355 8736 43675 8752
rect 43355 8672 43363 8736
rect 43427 8672 43443 8736
rect 43507 8672 43523 8736
rect 43587 8672 43603 8736
rect 43667 8672 43675 8736
rect 43355 7648 43675 8672
rect 43355 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43675 7648
rect 43355 6560 43675 7584
rect 43355 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43675 6560
rect 43355 5472 43675 6496
rect 43355 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43675 5472
rect 43355 4384 43675 5408
rect 43355 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43675 4384
rect 43355 3296 43675 4320
rect 43355 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43675 3296
rect 43355 2208 43675 3232
rect 43355 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43675 2208
rect 43355 1120 43675 2144
rect 43355 1056 43363 1120
rect 43427 1056 43443 1120
rect 43507 1056 43523 1120
rect 43587 1056 43603 1120
rect 43667 1056 43675 1120
rect 43355 1040 43675 1056
rect 30235 987 30301 988
rect 24899 236 24965 237
rect 24899 172 24900 236
rect 24964 172 24965 236
rect 24899 171 24965 172
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 27140 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 33396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 34500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 35420 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_174
timestamp 1688980957
transform 1 0 17112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_233
timestamp 1688980957
transform 1 0 22540 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_353
timestamp 1688980957
transform 1 0 33580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_371
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1688980957
transform 1 0 36984 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_238
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_266
timestamp 1688980957
transform 1 0 25576 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_285
timestamp 1688980957
transform 1 0 27324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_332
timestamp 1688980957
transform 1 0 31648 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_365
timestamp 1688980957
transform 1 0 34684 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_376
timestamp 1688980957
transform 1 0 35696 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1688980957
transform 1 0 36984 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_398
timestamp 1688980957
transform 1 0 37720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_403
timestamp 1688980957
transform 1 0 38180 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_410
timestamp 1688980957
transform 1 0 38824 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_418
timestamp 1688980957
transform 1 0 39560 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_426
timestamp 1688980957
transform 1 0 40296 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_438
timestamp 1688980957
transform 1 0 41400 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_163
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_172
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_180
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_244
timestamp 1688980957
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_257
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_291
timestamp 1688980957
transform 1 0 27876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_312
timestamp 1688980957
transform 1 0 29808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_322
timestamp 1688980957
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_352
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_371
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_380
timestamp 1688980957
transform 1 0 36064 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_392
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_411
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_427
timestamp 1688980957
transform 1 0 40388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_431
timestamp 1688980957
transform 1 0 40756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_443
timestamp 1688980957
transform 1 0 41860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_452
timestamp 1688980957
transform 1 0 42688 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1688980957
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_228
timestamp 1688980957
transform 1 0 22080 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_240
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_252
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_267
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_297
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_308
timestamp 1688980957
transform 1 0 29440 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_312
timestamp 1688980957
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_324
timestamp 1688980957
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_457
timestamp 1688980957
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_457
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_13
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_74
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_89
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_120
timestamp 1688980957
transform 1 0 12144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_132
timestamp 1688980957
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_147
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_189
timestamp 1688980957
transform 1 0 18492 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_212
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_235
timestamp 1688980957
transform 1 0 22724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_247
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_258
timestamp 1688980957
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_270
timestamp 1688980957
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_285
timestamp 1688980957
transform 1 0 27324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_297
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_304
timestamp 1688980957
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_321
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_327
timestamp 1688980957
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_350
timestamp 1688980957
transform 1 0 33304 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_362
timestamp 1688980957
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_365
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_399
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_419
timestamp 1688980957
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_421
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_433
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_437
timestamp 1688980957
transform 1 0 41308 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_444
timestamp 1688980957
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_453
timestamp 1688980957
transform 1 0 42780 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39192 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 39468 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 40112 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 40388 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 40664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 41768 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 36708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 37536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 37812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 38088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 36708 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 38640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 9108 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 9476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 14628 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 14904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 12052 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 14904 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__00_
timestamp 1688980957
transform 1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__01_
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__02_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__03_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__04_
timestamp 1688980957
transform 1 0 23184 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__05_
timestamp 1688980957
transform 1 0 23460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__06_
timestamp 1688980957
transform 1 0 24748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__07_
timestamp 1688980957
transform 1 0 25024 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__08_
timestamp 1688980957
transform 1 0 18768 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__09_
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__10_
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__11_
timestamp 1688980957
transform 1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__12_
timestamp 1688980957
transform 1 0 19320 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__13_
timestamp 1688980957
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__14_
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__15_
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__16_
timestamp 1688980957
transform 1 0 25300 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__17_
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__18_
timestamp 1688980957
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__19_
timestamp 1688980957
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__20_
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__21_
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__22_
timestamp 1688980957
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__23_
timestamp 1688980957
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__24_
timestamp 1688980957
transform 1 0 25944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__25_
timestamp 1688980957
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__26_
timestamp 1688980957
transform 1 0 27508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__27_
timestamp 1688980957
transform 1 0 26496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__28_
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__29_
timestamp 1688980957
transform 1 0 27048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__30_
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__31_
timestamp 1688980957
transform 1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__32_
timestamp 1688980957
transform 1 0 19596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__33_
timestamp 1688980957
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__34_
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__35_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__36_
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__37_
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__38_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__39_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__40_
timestamp 1688980957
transform 1 0 18216 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__41_
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__42_
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__43_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__44_
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__45_
timestamp 1688980957
transform 1 0 17112 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__46_
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_DSP_switch_matrix__47_
timestamp 1688980957
transform 1 0 16836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__48_
timestamp 1688980957
transform 1 0 17664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__49_
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__50_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_DSP_switch_matrix__51_
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 39284 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 41400 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 17940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1688980957
transform 1 0 19320 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 19688 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 20424 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 22724 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 24748 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 25300 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 25852 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 20056 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 21160 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 20976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 21988 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 22632 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 26404 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 28336 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 29992 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 28888 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 30544 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 29440 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 25668 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 26220 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 27508 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 28060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 27784 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 28612 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 30636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 32660 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 35604 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 36156 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 34868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 31096 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1688980957
transform 1 0 31372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 31188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 33764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43516 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 43516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 43516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 43516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 23736 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 27324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 29532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 31740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 37444 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 36432 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 37904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 38548 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 39744 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 40020 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 27968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 22724 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 27324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 40480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 34150 -300 34206 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 36910 -300 36966 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 37186 -300 37242 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 37462 -300 37518 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 37738 -300 37794 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 38014 -300 38070 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 38290 -300 38346 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 38566 -300 38622 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 38842 -300 38898 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 39118 -300 39174 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 39394 -300 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 34426 -300 34482 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 34702 -300 34758 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 34978 -300 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 35254 -300 35310 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 35530 -300 35586 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 35806 -300 35862 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 36082 -300 36138 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 36358 -300 36414 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 36634 -300 36690 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 3238 9840 3294 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 24398 9840 24454 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 26514 9840 26570 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 28630 9840 28686 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 30746 9840 30802 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 32862 9840 32918 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 34978 9840 35034 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 37094 9840 37150 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 39210 9840 39266 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 41326 9840 41382 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 43442 9840 43498 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 5354 9840 5410 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 7470 9840 7526 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 9586 9840 9642 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 11702 9840 11758 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 13818 9840 13874 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 15934 9840 15990 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 18050 9840 18106 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 20166 9840 20222 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 22282 9840 22338 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 5170 -300 5226 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 5446 -300 5502 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 5722 -300 5778 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 5998 -300 6054 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 8482 -300 8538 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 8758 -300 8814 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 9034 -300 9090 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 9310 -300 9366 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 9586 -300 9642 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 9862 -300 9918 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 10138 -300 10194 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 10414 -300 10470 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 6274 -300 6330 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 6550 -300 6606 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 6826 -300 6882 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 7102 -300 7158 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 7378 -300 7434 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 7654 -300 7710 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 7930 -300 7986 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 8206 -300 8262 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 10690 -300 10746 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 13450 -300 13506 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 13726 -300 13782 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 14002 -300 14058 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 14278 -300 14334 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 14554 -300 14610 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 14830 -300 14886 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 10966 -300 11022 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 11242 -300 11298 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 11518 -300 11574 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 11794 -300 11850 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 12070 -300 12126 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 12346 -300 12402 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 12622 -300 12678 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 12898 -300 12954 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 13174 -300 13230 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 15106 -300 15162 160 0 FreeSans 224 90 0 0 NN4END[0]
port 76 nsew signal input
flabel metal2 s 17866 -300 17922 160 0 FreeSans 224 90 0 0 NN4END[10]
port 77 nsew signal input
flabel metal2 s 18142 -300 18198 160 0 FreeSans 224 90 0 0 NN4END[11]
port 78 nsew signal input
flabel metal2 s 18418 -300 18474 160 0 FreeSans 224 90 0 0 NN4END[12]
port 79 nsew signal input
flabel metal2 s 18694 -300 18750 160 0 FreeSans 224 90 0 0 NN4END[13]
port 80 nsew signal input
flabel metal2 s 18970 -300 19026 160 0 FreeSans 224 90 0 0 NN4END[14]
port 81 nsew signal input
flabel metal2 s 19246 -300 19302 160 0 FreeSans 224 90 0 0 NN4END[15]
port 82 nsew signal input
flabel metal2 s 15382 -300 15438 160 0 FreeSans 224 90 0 0 NN4END[1]
port 83 nsew signal input
flabel metal2 s 15658 -300 15714 160 0 FreeSans 224 90 0 0 NN4END[2]
port 84 nsew signal input
flabel metal2 s 15934 -300 15990 160 0 FreeSans 224 90 0 0 NN4END[3]
port 85 nsew signal input
flabel metal2 s 16210 -300 16266 160 0 FreeSans 224 90 0 0 NN4END[4]
port 86 nsew signal input
flabel metal2 s 16486 -300 16542 160 0 FreeSans 224 90 0 0 NN4END[5]
port 87 nsew signal input
flabel metal2 s 16762 -300 16818 160 0 FreeSans 224 90 0 0 NN4END[6]
port 88 nsew signal input
flabel metal2 s 17038 -300 17094 160 0 FreeSans 224 90 0 0 NN4END[7]
port 89 nsew signal input
flabel metal2 s 17314 -300 17370 160 0 FreeSans 224 90 0 0 NN4END[8]
port 90 nsew signal input
flabel metal2 s 17590 -300 17646 160 0 FreeSans 224 90 0 0 NN4END[9]
port 91 nsew signal input
flabel metal2 s 19522 -300 19578 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 92 nsew signal tristate
flabel metal2 s 19798 -300 19854 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 93 nsew signal tristate
flabel metal2 s 20074 -300 20130 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 94 nsew signal tristate
flabel metal2 s 20350 -300 20406 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 95 nsew signal tristate
flabel metal2 s 22834 -300 22890 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 96 nsew signal tristate
flabel metal2 s 23110 -300 23166 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 97 nsew signal tristate
flabel metal2 s 23386 -300 23442 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 98 nsew signal tristate
flabel metal2 s 23662 -300 23718 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 99 nsew signal tristate
flabel metal2 s 23938 -300 23994 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 100 nsew signal tristate
flabel metal2 s 24214 -300 24270 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 101 nsew signal tristate
flabel metal2 s 24490 -300 24546 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 102 nsew signal tristate
flabel metal2 s 24766 -300 24822 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 103 nsew signal tristate
flabel metal2 s 20626 -300 20682 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 104 nsew signal tristate
flabel metal2 s 20902 -300 20958 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 105 nsew signal tristate
flabel metal2 s 21178 -300 21234 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 106 nsew signal tristate
flabel metal2 s 21454 -300 21510 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 107 nsew signal tristate
flabel metal2 s 21730 -300 21786 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 108 nsew signal tristate
flabel metal2 s 22006 -300 22062 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 109 nsew signal tristate
flabel metal2 s 22282 -300 22338 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 110 nsew signal tristate
flabel metal2 s 22558 -300 22614 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 111 nsew signal tristate
flabel metal2 s 25042 -300 25098 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 112 nsew signal tristate
flabel metal2 s 27802 -300 27858 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 113 nsew signal tristate
flabel metal2 s 28078 -300 28134 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 114 nsew signal tristate
flabel metal2 s 28354 -300 28410 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 115 nsew signal tristate
flabel metal2 s 28630 -300 28686 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 116 nsew signal tristate
flabel metal2 s 28906 -300 28962 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 117 nsew signal tristate
flabel metal2 s 29182 -300 29238 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 118 nsew signal tristate
flabel metal2 s 25318 -300 25374 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 119 nsew signal tristate
flabel metal2 s 25594 -300 25650 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 120 nsew signal tristate
flabel metal2 s 25870 -300 25926 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 121 nsew signal tristate
flabel metal2 s 26146 -300 26202 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 122 nsew signal tristate
flabel metal2 s 26422 -300 26478 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 123 nsew signal tristate
flabel metal2 s 26698 -300 26754 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 124 nsew signal tristate
flabel metal2 s 26974 -300 27030 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 125 nsew signal tristate
flabel metal2 s 27250 -300 27306 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 126 nsew signal tristate
flabel metal2 s 27526 -300 27582 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 127 nsew signal tristate
flabel metal2 s 29458 -300 29514 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 128 nsew signal tristate
flabel metal2 s 32218 -300 32274 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 129 nsew signal tristate
flabel metal2 s 32494 -300 32550 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 130 nsew signal tristate
flabel metal2 s 32770 -300 32826 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 131 nsew signal tristate
flabel metal2 s 33046 -300 33102 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 132 nsew signal tristate
flabel metal2 s 33322 -300 33378 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 133 nsew signal tristate
flabel metal2 s 33598 -300 33654 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 134 nsew signal tristate
flabel metal2 s 29734 -300 29790 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 135 nsew signal tristate
flabel metal2 s 30010 -300 30066 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 136 nsew signal tristate
flabel metal2 s 30286 -300 30342 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 137 nsew signal tristate
flabel metal2 s 30562 -300 30618 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 138 nsew signal tristate
flabel metal2 s 30838 -300 30894 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 139 nsew signal tristate
flabel metal2 s 31114 -300 31170 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 140 nsew signal tristate
flabel metal2 s 31390 -300 31446 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 141 nsew signal tristate
flabel metal2 s 31666 -300 31722 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 142 nsew signal tristate
flabel metal2 s 31942 -300 31998 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 143 nsew signal tristate
flabel metal2 s 33874 -300 33930 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 1122 9840 1178 10300 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6245 1040 6565 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 16848 1040 17168 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 27451 1040 27771 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 38054 1040 38374 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 11546 1040 11866 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 22149 1040 22469 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 32752 1040 33072 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 43355 1040 43675 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 22310 8160 22310 8160 0 vccd1
rlabel via1 22389 8704 22389 8704 0 vssd1
rlabel metal2 34178 551 34178 551 0 FrameStrobe[0]
rlabel metal2 37168 2890 37168 2890 0 FrameStrobe[10]
rlabel metal2 37260 2788 37260 2788 0 FrameStrobe[11]
rlabel metal1 38824 3162 38824 3162 0 FrameStrobe[12]
rlabel metal1 39100 3434 39100 3434 0 FrameStrobe[13]
rlabel metal2 37996 2822 37996 2822 0 FrameStrobe[14]
rlabel metal1 39698 3502 39698 3502 0 FrameStrobe[15]
rlabel metal1 39882 3026 39882 3026 0 FrameStrobe[16]
rlabel metal2 41446 850 41446 850 0 FrameStrobe[17]
rlabel metal2 41722 918 41722 918 0 FrameStrobe[18]
rlabel metal1 41814 1360 41814 1360 0 FrameStrobe[19]
rlabel metal2 34454 670 34454 670 0 FrameStrobe[1]
rlabel metal2 34829 68 34829 68 0 FrameStrobe[2]
rlabel metal2 35105 68 35105 68 0 FrameStrobe[3]
rlabel metal2 35381 68 35381 68 0 FrameStrobe[4]
rlabel metal2 35657 68 35657 68 0 FrameStrobe[5]
rlabel metal2 35834 976 35834 976 0 FrameStrobe[6]
rlabel metal2 36110 534 36110 534 0 FrameStrobe[7]
rlabel metal1 37536 2822 37536 2822 0 FrameStrobe[8]
rlabel metal2 36800 3570 36800 3570 0 FrameStrobe[9]
rlabel metal1 3404 8602 3404 8602 0 FrameStrobe_O[0]
rlabel metal1 24564 8602 24564 8602 0 FrameStrobe_O[10]
rlabel metal1 26864 8602 26864 8602 0 FrameStrobe_O[11]
rlabel metal1 28796 8602 28796 8602 0 FrameStrobe_O[12]
rlabel metal1 30912 8602 30912 8602 0 FrameStrobe_O[13]
rlabel metal2 32890 9445 32890 9445 0 FrameStrobe_O[14]
rlabel metal1 35144 8602 35144 8602 0 FrameStrobe_O[15]
rlabel metal2 37122 9224 37122 9224 0 FrameStrobe_O[16]
rlabel metal1 39376 8602 39376 8602 0 FrameStrobe_O[17]
rlabel metal2 41354 9224 41354 9224 0 FrameStrobe_O[18]
rlabel metal1 43194 8602 43194 8602 0 FrameStrobe_O[19]
rlabel metal2 5382 9445 5382 9445 0 FrameStrobe_O[1]
rlabel metal1 7636 8602 7636 8602 0 FrameStrobe_O[2]
rlabel metal2 9614 9224 9614 9224 0 FrameStrobe_O[3]
rlabel metal1 11960 8602 11960 8602 0 FrameStrobe_O[4]
rlabel metal2 13846 9224 13846 9224 0 FrameStrobe_O[5]
rlabel metal1 16100 8602 16100 8602 0 FrameStrobe_O[6]
rlabel metal2 18078 9224 18078 9224 0 FrameStrobe_O[7]
rlabel metal1 20332 8602 20332 8602 0 FrameStrobe_O[8]
rlabel metal2 22586 9231 22586 9231 0 FrameStrobe_O[9]
rlabel metal1 28842 2346 28842 2346 0 FrameStrobe_O_i\[0\]
rlabel metal1 25070 2380 25070 2380 0 FrameStrobe_O_i\[10\]
rlabel metal2 27462 2414 27462 2414 0 FrameStrobe_O_i\[11\]
rlabel metal1 29486 3026 29486 3026 0 FrameStrobe_O_i\[12\]
rlabel metal2 31326 2244 31326 2244 0 FrameStrobe_O_i\[13\]
rlabel metal1 37490 2040 37490 2040 0 FrameStrobe_O_i\[14\]
rlabel metal1 36248 2074 36248 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 37858 2074 37858 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 39008 2074 39008 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 40250 2074 40250 2074 0 FrameStrobe_O_i\[18\]
rlabel metal1 42642 1938 42642 1938 0 FrameStrobe_O_i\[19\]
rlabel metal2 24058 2210 24058 2210 0 FrameStrobe_O_i\[1\]
rlabel metal1 25162 2448 25162 2448 0 FrameStrobe_O_i\[2\]
rlabel metal1 27738 2822 27738 2822 0 FrameStrobe_O_i\[3\]
rlabel metal1 22218 2380 22218 2380 0 FrameStrobe_O_i\[4\]
rlabel metal1 15548 2414 15548 2414 0 FrameStrobe_O_i\[5\]
rlabel metal1 16376 2414 16376 2414 0 FrameStrobe_O_i\[6\]
rlabel metal1 18722 2414 18722 2414 0 FrameStrobe_O_i\[7\]
rlabel metal1 20700 2414 20700 2414 0 FrameStrobe_O_i\[8\]
rlabel metal2 23782 2278 23782 2278 0 FrameStrobe_O_i\[9\]
rlabel metal2 5198 670 5198 670 0 N1END[0]
rlabel metal2 5474 670 5474 670 0 N1END[1]
rlabel metal2 5750 670 5750 670 0 N1END[2]
rlabel metal2 6026 143 6026 143 0 N1END[3]
rlabel metal2 8510 415 8510 415 0 N2END[0]
rlabel metal2 8687 68 8687 68 0 N2END[1]
rlabel metal2 9115 68 9115 68 0 N2END[2]
rlabel metal2 9338 398 9338 398 0 N2END[3]
rlabel metal2 9614 670 9614 670 0 N2END[4]
rlabel metal2 9791 68 9791 68 0 N2END[5]
rlabel metal2 10067 68 10067 68 0 N2END[6]
rlabel metal2 10442 670 10442 670 0 N2END[7]
rlabel metal2 6302 670 6302 670 0 N2MID[0]
rlabel metal2 6479 68 6479 68 0 N2MID[1]
rlabel metal2 6755 68 6755 68 0 N2MID[2]
rlabel metal2 6762 544 6762 544 0 N2MID[3]
rlabel metal2 7353 68 7353 68 0 N2MID[4]
rlabel metal2 7583 68 7583 68 0 N2MID[5]
rlabel metal2 7859 68 7859 68 0 N2MID[6]
rlabel metal2 8135 68 8135 68 0 N2MID[7]
rlabel metal2 10619 68 10619 68 0 N4END[0]
rlabel metal2 13478 415 13478 415 0 N4END[10]
rlabel metal2 13754 398 13754 398 0 N4END[11]
rlabel metal2 13931 68 13931 68 0 N4END[12]
rlabel metal2 14306 551 14306 551 0 N4END[13]
rlabel metal2 14582 551 14582 551 0 N4END[14]
rlabel metal2 14858 551 14858 551 0 N4END[15]
rlabel metal2 10994 398 10994 398 0 N4END[1]
rlabel metal2 11171 68 11171 68 0 N4END[2]
rlabel metal2 11546 415 11546 415 0 N4END[3]
rlabel metal2 11822 398 11822 398 0 N4END[4]
rlabel metal2 12098 415 12098 415 0 N4END[5]
rlabel metal2 12374 636 12374 636 0 N4END[6]
rlabel metal1 12282 1360 12282 1360 0 N4END[7]
rlabel metal2 12926 483 12926 483 0 N4END[8]
rlabel metal2 13202 347 13202 347 0 N4END[9]
rlabel metal2 15134 1044 15134 1044 0 NN4END[0]
rlabel metal2 17894 347 17894 347 0 NN4END[10]
rlabel metal2 18170 551 18170 551 0 NN4END[11]
rlabel metal2 18446 466 18446 466 0 NN4END[12]
rlabel metal2 18722 347 18722 347 0 NN4END[13]
rlabel metal2 18998 364 18998 364 0 NN4END[14]
rlabel metal2 19274 211 19274 211 0 NN4END[15]
rlabel metal2 15410 211 15410 211 0 NN4END[1]
rlabel metal2 15686 347 15686 347 0 NN4END[2]
rlabel metal2 15962 347 15962 347 0 NN4END[3]
rlabel metal2 16238 755 16238 755 0 NN4END[4]
rlabel metal2 16514 279 16514 279 0 NN4END[5]
rlabel metal2 16691 68 16691 68 0 NN4END[6]
rlabel metal2 17066 398 17066 398 0 NN4END[7]
rlabel metal2 17342 1248 17342 1248 0 NN4END[8]
rlabel metal2 17618 415 17618 415 0 NN4END[9]
rlabel metal2 19550 364 19550 364 0 S1BEG[0]
rlabel metal2 19826 636 19826 636 0 S1BEG[1]
rlabel metal2 20102 636 20102 636 0 S1BEG[2]
rlabel metal2 20378 959 20378 959 0 S1BEG[3]
rlabel metal2 22915 68 22915 68 0 S2BEG[0]
rlabel metal2 23138 636 23138 636 0 S2BEG[1]
rlabel metal2 23414 806 23414 806 0 S2BEG[2]
rlabel metal2 23690 636 23690 636 0 S2BEG[3]
rlabel metal2 23966 908 23966 908 0 S2BEG[4]
rlabel metal2 24242 806 24242 806 0 S2BEG[5]
rlabel metal2 24617 68 24617 68 0 S2BEG[6]
rlabel metal2 24794 636 24794 636 0 S2BEG[7]
rlabel metal2 20654 347 20654 347 0 S2BEGb[0]
rlabel metal2 20930 772 20930 772 0 S2BEGb[1]
rlabel metal2 21305 68 21305 68 0 S2BEGb[2]
rlabel metal2 21482 1180 21482 1180 0 S2BEGb[3]
rlabel metal2 21758 636 21758 636 0 S2BEGb[4]
rlabel metal2 22034 908 22034 908 0 S2BEGb[5]
rlabel metal2 22409 68 22409 68 0 S2BEGb[6]
rlabel metal2 22685 68 22685 68 0 S2BEGb[7]
rlabel metal2 25070 364 25070 364 0 S4BEG[0]
rlabel metal2 27830 942 27830 942 0 S4BEG[10]
rlabel metal2 28106 1010 28106 1010 0 S4BEG[11]
rlabel metal2 28481 68 28481 68 0 S4BEG[12]
rlabel metal1 29762 2822 29762 2822 0 S4BEG[13]
rlabel metal2 28934 755 28934 755 0 S4BEG[14]
rlabel metal2 29309 68 29309 68 0 S4BEG[15]
rlabel metal2 25445 68 25445 68 0 S4BEG[1]
rlabel metal2 25622 908 25622 908 0 S4BEG[2]
rlabel metal2 25898 908 25898 908 0 S4BEG[3]
rlabel metal2 26174 279 26174 279 0 S4BEG[4]
rlabel metal2 26450 636 26450 636 0 S4BEG[5]
rlabel metal2 26726 483 26726 483 0 S4BEG[6]
rlabel metal2 27002 347 27002 347 0 S4BEG[7]
rlabel metal2 27278 279 27278 279 0 S4BEG[8]
rlabel metal2 27554 228 27554 228 0 S4BEG[9]
rlabel metal2 29585 68 29585 68 0 SS4BEG[0]
rlabel metal2 32345 68 32345 68 0 SS4BEG[10]
rlabel metal2 32621 68 32621 68 0 SS4BEG[11]
rlabel metal2 32798 534 32798 534 0 SS4BEG[12]
rlabel metal2 33074 500 33074 500 0 SS4BEG[13]
rlabel metal2 33449 68 33449 68 0 SS4BEG[14]
rlabel metal2 33626 942 33626 942 0 SS4BEG[15]
rlabel metal2 29762 160 29762 160 0 SS4BEG[1]
rlabel metal2 30137 68 30137 68 0 SS4BEG[2]
rlabel metal2 30413 68 30413 68 0 SS4BEG[3]
rlabel metal2 30590 1180 30590 1180 0 SS4BEG[4]
rlabel metal2 30866 806 30866 806 0 SS4BEG[5]
rlabel metal2 31241 68 31241 68 0 SS4BEG[6]
rlabel metal1 33442 1768 33442 1768 0 SS4BEG[7]
rlabel metal2 31694 262 31694 262 0 SS4BEG[8]
rlabel metal2 31970 415 31970 415 0 SS4BEG[9]
rlabel metal2 33902 704 33902 704 0 UserCLK
rlabel metal2 1150 9445 1150 9445 0 UserCLKo
rlabel metal2 35466 2210 35466 2210 0 net1
rlabel metal2 40158 1734 40158 1734 0 net10
rlabel metal1 22678 2822 22678 2822 0 net100
rlabel metal2 21850 1462 21850 1462 0 net101
rlabel metal1 24426 2006 24426 2006 0 net102
rlabel metal2 24886 1530 24886 1530 0 net103
rlabel metal1 25116 1326 25116 1326 0 net104
rlabel metal1 25530 1258 25530 1258 0 net105
rlabel metal1 20194 1360 20194 1360 0 net106
rlabel metal2 19274 1530 19274 1530 0 net107
rlabel metal1 21022 2006 21022 2006 0 net108
rlabel metal1 21022 2346 21022 2346 0 net109
rlabel metal2 41814 1734 41814 1734 0 net11
rlabel metal1 20884 1326 20884 1326 0 net110
rlabel metal1 21988 2006 21988 2006 0 net111
rlabel metal2 21574 1802 21574 1802 0 net112
rlabel metal1 20194 1836 20194 1836 0 net113
rlabel metal1 26358 1326 26358 1326 0 net114
rlabel metal1 28428 2006 28428 2006 0 net115
rlabel metal1 29946 2006 29946 2006 0 net116
rlabel metal1 28980 2006 28980 2006 0 net117
rlabel metal1 30682 2040 30682 2040 0 net118
rlabel metal1 29348 1530 29348 1530 0 net119
rlabel metal2 36938 782 36938 782 0 net12
rlabel metal2 31050 1938 31050 1938 0 net120
rlabel metal1 26634 1258 26634 1258 0 net121
rlabel metal1 25852 2006 25852 2006 0 net122
rlabel metal1 25852 2822 25852 2822 0 net123
rlabel metal1 27508 1326 27508 1326 0 net124
rlabel metal1 27738 1258 27738 1258 0 net125
rlabel metal1 27370 2006 27370 2006 0 net126
rlabel metal1 28336 1326 28336 1326 0 net127
rlabel metal1 29256 1258 29256 1258 0 net128
rlabel metal1 29164 3094 29164 3094 0 net129
rlabel metal2 26818 2550 26818 2550 0 net13
rlabel metal2 20286 1360 20286 1360 0 net130
rlabel metal3 22057 2924 22057 2924 0 net131
rlabel metal2 18354 935 18354 935 0 net132
rlabel metal2 16744 3468 16744 3468 0 net133
rlabel metal2 30222 3111 30222 3111 0 net134
rlabel metal2 15686 2159 15686 2159 0 net135
rlabel metal1 33580 2074 33580 2074 0 net136
rlabel metal1 32246 646 32246 646 0 net137
rlabel metal2 29302 1989 29302 1989 0 net138
rlabel metal2 18814 1088 18814 1088 0 net139
rlabel metal3 31786 2924 31786 2924 0 net14
rlabel metal1 18262 952 18262 952 0 net140
rlabel metal2 30958 952 30958 952 0 net141
rlabel metal2 30222 2125 30222 2125 0 net142
rlabel via2 17158 2091 17158 2091 0 net143
rlabel metal1 34822 1224 34822 1224 0 net144
rlabel metal2 17710 2788 17710 2788 0 net145
rlabel via2 2254 8347 2254 8347 0 net146
rlabel metal1 37858 238 37858 238 0 net15
rlabel metal2 16606 3196 16606 3196 0 net16
rlabel metal2 17296 3876 17296 3876 0 net17
rlabel metal1 21298 3162 21298 3162 0 net18
rlabel metal2 20930 1989 20930 1989 0 net19
rlabel metal1 39376 1190 39376 1190 0 net2
rlabel metal1 34730 748 34730 748 0 net20
rlabel metal1 4830 952 4830 952 0 net21
rlabel metal1 4922 374 4922 374 0 net22
rlabel metal2 5842 1156 5842 1156 0 net23
rlabel metal1 6118 408 6118 408 0 net24
rlabel metal1 8280 1190 8280 1190 0 net25
rlabel metal1 8694 680 8694 680 0 net26
rlabel metal1 10166 2074 10166 2074 0 net27
rlabel metal2 19458 1156 19458 1156 0 net28
rlabel metal1 9246 1190 9246 1190 0 net29
rlabel via2 27554 3043 27554 3043 0 net3
rlabel metal2 20010 1853 20010 1853 0 net30
rlabel metal1 9706 1496 9706 1496 0 net31
rlabel metal2 10258 238 10258 238 0 net32
rlabel metal2 7222 2856 7222 2856 0 net33
rlabel metal1 6348 1190 6348 1190 0 net34
rlabel metal2 6578 1088 6578 1088 0 net35
rlabel metal2 8602 2992 8602 2992 0 net36
rlabel metal1 7222 204 7222 204 0 net37
rlabel metal1 22034 2992 22034 2992 0 net38
rlabel metal2 7682 986 7682 986 0 net39
rlabel metal1 37766 2958 37766 2958 0 net4
rlabel metal1 8050 1190 8050 1190 0 net40
rlabel metal2 31970 1105 31970 1105 0 net41
rlabel metal1 13018 340 13018 340 0 net42
rlabel metal2 17710 3009 17710 3009 0 net43
rlabel metal2 25622 3264 25622 3264 0 net44
rlabel metal2 17986 3060 17986 3060 0 net45
rlabel metal1 18538 2414 18538 2414 0 net46
rlabel metal1 18078 1972 18078 1972 0 net47
rlabel metal2 10718 901 10718 901 0 net48
rlabel metal2 10810 697 10810 697 0 net49
rlabel metal1 31878 884 31878 884 0 net5
rlabel metal2 11086 2040 11086 2040 0 net50
rlabel metal2 11362 2890 11362 2890 0 net51
rlabel metal2 11270 833 11270 833 0 net52
rlabel metal2 12006 2550 12006 2550 0 net53
rlabel metal2 12282 765 12282 765 0 net54
rlabel metal2 26910 527 26910 527 0 net55
rlabel metal2 12834 1819 12834 1819 0 net56
rlabel metal1 15226 1904 15226 1904 0 net57
rlabel metal1 16606 1462 16606 1462 0 net58
rlabel metal1 18078 1360 18078 1360 0 net59
rlabel metal1 40434 1224 40434 1224 0 net6
rlabel metal1 18630 1360 18630 1360 0 net60
rlabel metal1 18262 1904 18262 1904 0 net61
rlabel metal2 17802 986 17802 986 0 net62
rlabel metal1 18538 1190 18538 1190 0 net63
rlabel metal1 13984 1190 13984 1190 0 net64
rlabel metal1 14306 1530 14306 1530 0 net65
rlabel metal2 14398 1088 14398 1088 0 net66
rlabel metal1 14766 1462 14766 1462 0 net67
rlabel metal1 14996 1190 14996 1190 0 net68
rlabel metal1 16882 1292 16882 1292 0 net69
rlabel metal2 40710 952 40710 952 0 net7
rlabel metal1 15962 1530 15962 1530 0 net70
rlabel metal1 17112 1938 17112 1938 0 net71
rlabel metal2 15778 1020 15778 1020 0 net72
rlabel metal1 33764 1462 33764 1462 0 net73
rlabel metal1 3358 8500 3358 8500 0 net74
rlabel metal1 24702 8466 24702 8466 0 net75
rlabel metal2 27094 6900 27094 6900 0 net76
rlabel metal1 28980 3162 28980 3162 0 net77
rlabel metal1 31004 2618 31004 2618 0 net78
rlabel metal1 33074 8466 33074 8466 0 net79
rlabel metal2 40986 1734 40986 1734 0 net8
rlabel metal1 35466 2618 35466 2618 0 net80
rlabel metal1 37490 2618 37490 2618 0 net81
rlabel metal1 39284 2618 39284 2618 0 net82
rlabel metal1 41032 8466 41032 8466 0 net83
rlabel metal1 42688 2618 42688 2618 0 net84
rlabel metal1 6141 8466 6141 8466 0 net85
rlabel metal2 7590 8636 7590 8636 0 net86
rlabel via2 9614 8483 9614 8483 0 net87
rlabel via1 14306 8347 14306 8347 0 net88
rlabel metal1 14766 8466 14766 8466 0 net89
rlabel metal2 41262 1666 41262 1666 0 net9
rlabel metal1 15962 2618 15962 2618 0 net90
rlabel metal1 18262 2618 18262 2618 0 net91
rlabel metal1 20378 2550 20378 2550 0 net92
rlabel metal1 22586 8466 22586 8466 0 net93
rlabel metal3 18400 1836 18400 1836 0 net94
rlabel metal1 19366 1394 19366 1394 0 net95
rlabel metal1 18906 1224 18906 1224 0 net96
rlabel metal1 20240 2006 20240 2006 0 net97
rlabel metal2 21942 1768 21942 1768 0 net98
rlabel metal1 23046 1326 23046 1326 0 net99
<< properties >>
string FIXED_BBOX 0 0 44700 10000
<< end >>
