magic
tech sky130A
magscale 1 2
timestamp 1734825390
<< viali >>
rect 33609 86377 33643 86411
rect 41981 86377 42015 86411
rect 47317 86377 47351 86411
rect 49525 86377 49559 86411
rect 50353 86377 50387 86411
rect 50721 86377 50755 86411
rect 52469 86377 52503 86411
rect 61209 86377 61243 86411
rect 24501 86309 24535 86343
rect 29929 86309 29963 86343
rect 37381 86309 37415 86343
rect 44833 86309 44867 86343
rect 47869 86309 47903 86343
rect 25053 86241 25087 86275
rect 39221 86241 39255 86275
rect 39589 86241 39623 86275
rect 40049 86241 40083 86275
rect 40417 86241 40451 86275
rect 40601 86241 40635 86275
rect 27629 86173 27663 86207
rect 35081 86173 35115 86207
rect 43453 86173 43487 86207
rect 46581 86173 46615 86207
rect 49224 86173 49258 86207
rect 55321 86173 55355 86207
rect 108037 86173 108071 86207
rect 19423 86105 19457 86139
rect 19717 86105 19751 86139
rect 19901 86105 19935 86139
rect 19993 86105 20027 86139
rect 24777 86105 24811 86139
rect 27353 86105 27387 86139
rect 30205 86105 30239 86139
rect 30481 86105 30515 86139
rect 33885 86105 33919 86139
rect 34069 86105 34103 86139
rect 34161 86105 34195 86139
rect 35348 86105 35382 86139
rect 37657 86105 37691 86139
rect 37933 86105 37967 86139
rect 38853 86105 38887 86139
rect 40868 86105 40902 86139
rect 43720 86105 43754 86139
rect 45017 86105 45051 86139
rect 48982 86105 49016 86139
rect 53389 86105 53423 86139
rect 55588 86105 55622 86139
rect 24961 86037 24995 86071
rect 27059 86037 27093 86071
rect 27537 86037 27571 86071
rect 30389 86037 30423 86071
rect 36461 86037 36495 86071
rect 37841 86037 37875 86071
rect 42901 86037 42935 86071
rect 43269 86037 43303 86071
rect 49893 86037 49927 86071
rect 51181 86037 51215 86071
rect 51641 86037 51675 86071
rect 52009 86037 52043 86071
rect 53021 86037 53055 86071
rect 54677 86037 54711 86071
rect 56701 86037 56735 86071
rect 1501 84609 1535 84643
rect 1685 84473 1719 84507
rect 1501 83521 1535 83555
rect 1685 83385 1719 83419
rect 1501 82841 1535 82875
rect 1685 82841 1719 82875
rect 1501 81753 1535 81787
rect 1685 81753 1719 81787
rect 1501 80665 1535 80699
rect 1685 80665 1719 80699
rect 1501 79577 1535 79611
rect 1685 79577 1719 79611
rect 1409 79169 1443 79203
rect 1593 78965 1627 78999
rect 1409 78081 1443 78115
rect 1593 77877 1627 77911
rect 9321 77129 9355 77163
rect 1501 76993 1535 77027
rect 9229 76993 9263 77027
rect 9413 76925 9447 76959
rect 1685 76857 1719 76891
rect 8861 76789 8895 76823
rect 8677 76449 8711 76483
rect 8401 76381 8435 76415
rect 8493 76381 8527 76415
rect 8033 76245 8067 76279
rect 1501 75905 1535 75939
rect 1685 75769 1719 75803
rect 9229 75293 9263 75327
rect 9321 75293 9355 75327
rect 9413 75293 9447 75327
rect 9597 75293 9631 75327
rect 1501 75225 1535 75259
rect 1685 75225 1719 75259
rect 8953 75157 8987 75191
rect 8401 74817 8435 74851
rect 8493 74817 8527 74851
rect 8585 74817 8619 74851
rect 8769 74817 8803 74851
rect 9229 74817 9263 74851
rect 9321 74749 9355 74783
rect 9413 74749 9447 74783
rect 8125 74613 8159 74647
rect 8861 74613 8895 74647
rect 8677 74341 8711 74375
rect 1409 74205 1443 74239
rect 8493 74205 8527 74239
rect 9229 74205 9263 74239
rect 9321 74205 9355 74239
rect 9413 74205 9447 74239
rect 9597 74205 9631 74239
rect 1593 74069 1627 74103
rect 8953 74069 8987 74103
rect 6653 73729 6687 73763
rect 7849 73729 7883 73763
rect 7941 73729 7975 73763
rect 8125 73729 8159 73763
rect 8217 73729 8251 73763
rect 8769 73729 8803 73763
rect 6929 73661 6963 73695
rect 9045 73661 9079 73695
rect 7573 73593 7607 73627
rect 6837 73525 6871 73559
rect 7205 73525 7239 73559
rect 7665 73525 7699 73559
rect 7113 73321 7147 73355
rect 8953 73321 8987 73355
rect 5779 73253 5813 73287
rect 5549 73185 5583 73219
rect 7297 73185 7331 73219
rect 7941 73185 7975 73219
rect 7021 73117 7055 73151
rect 8125 73117 8159 73151
rect 8217 73117 8251 73151
rect 8401 73117 8435 73151
rect 8493 73117 8527 73151
rect 9137 73117 9171 73151
rect 9229 73117 9263 73151
rect 9413 73117 9447 73151
rect 9505 73117 9539 73151
rect 1501 73049 1535 73083
rect 1593 72981 1627 73015
rect 7573 72981 7607 73015
rect 6469 72641 6503 72675
rect 7389 72641 7423 72675
rect 7481 72641 7515 72675
rect 7573 72641 7607 72675
rect 7757 72641 7791 72675
rect 8125 72641 8159 72675
rect 8217 72641 8251 72675
rect 8401 72641 8435 72675
rect 8493 72641 8527 72675
rect 8769 72641 8803 72675
rect 8861 72641 8895 72675
rect 9045 72641 9079 72675
rect 9137 72641 9171 72675
rect 9229 72641 9263 72675
rect 6745 72573 6779 72607
rect 6837 72437 6871 72471
rect 7021 72437 7055 72471
rect 7113 72437 7147 72471
rect 7941 72437 7975 72471
rect 8585 72437 8619 72471
rect 9413 72437 9447 72471
rect 7389 72233 7423 72267
rect 7849 72233 7883 72267
rect 5365 72029 5399 72063
rect 5641 72029 5675 72063
rect 6377 72029 6411 72063
rect 6653 72029 6687 72063
rect 7297 72029 7331 72063
rect 7573 72029 7607 72063
rect 8125 72029 8159 72063
rect 1501 71961 1535 71995
rect 1593 71893 1627 71927
rect 8309 71893 8343 71927
rect 7849 71621 7883 71655
rect 9229 71621 9263 71655
rect 9321 71621 9355 71655
rect 1501 71553 1535 71587
rect 6377 71553 6411 71587
rect 6644 71553 6678 71587
rect 8125 71553 8159 71587
rect 8217 71553 8251 71587
rect 8309 71553 8343 71587
rect 8493 71553 8527 71587
rect 9505 71485 9539 71519
rect 1593 71349 1627 71383
rect 7757 71349 7791 71383
rect 8861 71349 8895 71383
rect 9137 71145 9171 71179
rect 8033 71077 8067 71111
rect 8493 71009 8527 71043
rect 8677 71009 8711 71043
rect 6561 70941 6595 70975
rect 6837 70941 6871 70975
rect 9045 70941 9079 70975
rect 7757 70805 7791 70839
rect 8401 70805 8435 70839
rect 1593 70601 1627 70635
rect 8769 70601 8803 70635
rect 8861 70601 8895 70635
rect 9229 70601 9263 70635
rect 1409 70465 1443 70499
rect 7113 70465 7147 70499
rect 7205 70465 7239 70499
rect 7297 70465 7331 70499
rect 7481 70465 7515 70499
rect 7941 70465 7975 70499
rect 8033 70468 8067 70502
rect 8125 70465 8159 70499
rect 8309 70465 8343 70499
rect 8585 70465 8619 70499
rect 6837 70397 6871 70431
rect 9321 70397 9355 70431
rect 9413 70397 9447 70431
rect 7665 70261 7699 70295
rect 5733 70057 5767 70091
rect 6377 70057 6411 70091
rect 7021 70057 7055 70091
rect 9229 70057 9263 70091
rect 5917 69989 5951 70023
rect 6561 69989 6595 70023
rect 5641 69921 5675 69955
rect 6285 69921 6319 69955
rect 5365 69853 5399 69887
rect 5998 69855 6032 69889
rect 6653 69853 6687 69887
rect 7021 69853 7055 69887
rect 7297 69853 7331 69887
rect 7481 69853 7515 69887
rect 7573 69853 7607 69887
rect 7757 69853 7791 69887
rect 7849 69853 7883 69887
rect 8125 69853 8159 69887
rect 8290 69853 8324 69887
rect 8401 69853 8435 69887
rect 8503 69853 8537 69887
rect 7941 69785 7975 69819
rect 7205 69717 7239 69751
rect 6745 69513 6779 69547
rect 6837 69513 6871 69547
rect 8401 69513 8435 69547
rect 7573 69445 7607 69479
rect 8493 69445 8527 69479
rect 1501 69377 1535 69411
rect 9045 69377 9079 69411
rect 9137 69377 9171 69411
rect 9321 69377 9355 69411
rect 9413 69377 9447 69411
rect 6929 69309 6963 69343
rect 8585 69309 8619 69343
rect 1685 69241 1719 69275
rect 6377 69173 6411 69207
rect 8033 69173 8067 69207
rect 8861 69173 8895 69207
rect 4261 68969 4295 69003
rect 7205 68969 7239 69003
rect 5733 68901 5767 68935
rect 8309 68901 8343 68935
rect 6653 68833 6687 68867
rect 7849 68833 7883 68867
rect 4077 68765 4111 68799
rect 4353 68765 4387 68799
rect 4620 68765 4654 68799
rect 6101 68765 6135 68799
rect 6377 68765 6411 68799
rect 6560 68765 6594 68799
rect 6791 68765 6825 68799
rect 6929 68765 6963 68799
rect 7113 68765 7147 68799
rect 8953 68765 8987 68799
rect 7573 68697 7607 68731
rect 7665 68629 7699 68663
rect 9137 68629 9171 68663
rect 4997 68425 5031 68459
rect 1501 68289 1535 68323
rect 4169 68289 4203 68323
rect 4813 68289 4847 68323
rect 6653 68289 6687 68323
rect 6836 68295 6870 68329
rect 6929 68289 6963 68323
rect 7205 68289 7239 68323
rect 7757 68289 7791 68323
rect 7940 68292 7974 68326
rect 8033 68289 8067 68323
rect 8309 68289 8343 68323
rect 4629 68221 4663 68255
rect 7021 68221 7055 68255
rect 8125 68221 8159 68255
rect 8493 68153 8527 68187
rect 1593 68085 1627 68119
rect 4445 68085 4479 68119
rect 7297 68085 7331 68119
rect 4813 67813 4847 67847
rect 6837 67813 6871 67847
rect 7849 67745 7883 67779
rect 7573 67677 7607 67711
rect 7721 67677 7755 67711
rect 7941 67677 7975 67711
rect 8125 67677 8159 67711
rect 1501 67609 1535 67643
rect 1685 67609 1719 67643
rect 4537 67609 4571 67643
rect 6653 67609 6687 67643
rect 8309 67609 8343 67643
rect 4997 67541 5031 67575
rect 4721 67337 4755 67371
rect 7205 67337 7239 67371
rect 8677 67337 8711 67371
rect 9045 67337 9079 67371
rect 8217 67269 8251 67303
rect 4813 67201 4847 67235
rect 5069 67201 5103 67235
rect 6653 67201 6687 67235
rect 6929 67201 6963 67235
rect 8309 67201 8343 67235
rect 4261 67133 4295 67167
rect 8401 67133 8435 67167
rect 9137 67133 9171 67167
rect 9229 67133 9263 67167
rect 4629 67065 4663 67099
rect 7573 67065 7607 67099
rect 7849 67065 7883 67099
rect 6193 66997 6227 67031
rect 7021 66997 7055 67031
rect 8033 66793 8067 66827
rect 1685 66657 1719 66691
rect 6377 66657 6411 66691
rect 7481 66657 7515 66691
rect 7573 66657 7607 66691
rect 8677 66657 8711 66691
rect 6101 66589 6135 66623
rect 7205 66589 7239 66623
rect 7388 66589 7422 66623
rect 7757 66589 7791 66623
rect 8401 66589 8435 66623
rect 9209 66589 9243 66623
rect 9321 66589 9355 66623
rect 9413 66589 9447 66623
rect 9597 66589 9631 66623
rect 1501 66521 1535 66555
rect 4813 66521 4847 66555
rect 7941 66521 7975 66555
rect 4905 66453 4939 66487
rect 8493 66453 8527 66487
rect 8953 66453 8987 66487
rect 7021 66249 7055 66283
rect 8125 66249 8159 66283
rect 8493 66249 8527 66283
rect 5917 66181 5951 66215
rect 8585 66181 8619 66215
rect 5181 66113 5215 66147
rect 5365 66113 5399 66147
rect 5825 66113 5859 66147
rect 7294 66113 7328 66147
rect 7445 66116 7479 66150
rect 7849 66113 7883 66147
rect 6101 66045 6135 66079
rect 7573 66045 7607 66079
rect 7665 66045 7699 66079
rect 8769 66045 8803 66079
rect 5457 65977 5491 66011
rect 8033 65977 8067 66011
rect 5181 65909 5215 65943
rect 5549 65705 5583 65739
rect 5917 65569 5951 65603
rect 1501 65433 1535 65467
rect 1685 65433 1719 65467
rect 5089 65433 5123 65467
rect 5457 65433 5491 65467
rect 6184 65433 6218 65467
rect 5181 65365 5215 65399
rect 7297 65365 7331 65399
rect 8861 65161 8895 65195
rect 9229 65161 9263 65195
rect 4629 65093 4663 65127
rect 8585 65093 8619 65127
rect 4445 65025 4479 65059
rect 5549 65025 5583 65059
rect 7481 65025 7515 65059
rect 7665 65025 7699 65059
rect 7757 65025 7791 65059
rect 8033 65025 8067 65059
rect 4261 64957 4295 64991
rect 5273 64957 5307 64991
rect 7849 64957 7883 64991
rect 9321 64957 9355 64991
rect 9505 64957 9539 64991
rect 8217 64889 8251 64923
rect 5733 64481 5767 64515
rect 8585 64481 8619 64515
rect 5989 64413 6023 64447
rect 8401 64413 8435 64447
rect 1501 64345 1535 64379
rect 8493 64345 8527 64379
rect 1593 64277 1627 64311
rect 7113 64277 7147 64311
rect 8033 64277 8067 64311
rect 8217 64073 8251 64107
rect 8861 64073 8895 64107
rect 1501 63937 1535 63971
rect 6469 63937 6503 63971
rect 6736 63937 6770 63971
rect 8953 63869 8987 63903
rect 9045 63869 9079 63903
rect 7849 63801 7883 63835
rect 1593 63733 1627 63767
rect 8493 63733 8527 63767
rect 6929 63393 6963 63427
rect 7113 63393 7147 63427
rect 8309 63393 8343 63427
rect 8401 63393 8435 63427
rect 6837 63325 6871 63359
rect 8033 63325 8067 63359
rect 8217 63325 8251 63359
rect 8585 63325 8619 63359
rect 6469 63189 6503 63223
rect 7757 63189 7791 63223
rect 8769 63189 8803 63223
rect 4997 62985 5031 63019
rect 8033 62985 8067 63019
rect 8493 62985 8527 63019
rect 1501 62849 1535 62883
rect 4905 62849 4939 62883
rect 6561 62849 6595 62883
rect 6828 62849 6862 62883
rect 8401 62849 8435 62883
rect 8861 62849 8895 62883
rect 8585 62781 8619 62815
rect 1777 62645 1811 62679
rect 7941 62645 7975 62679
rect 9045 62645 9079 62679
rect 7481 62441 7515 62475
rect 7205 62305 7239 62339
rect 7941 62305 7975 62339
rect 8033 62305 8067 62339
rect 2329 62237 2363 62271
rect 7021 62237 7055 62271
rect 7113 62237 7147 62271
rect 7849 62237 7883 62271
rect 8309 62237 8343 62271
rect 2145 62101 2179 62135
rect 6653 62101 6687 62135
rect 8493 62101 8527 62135
rect 1685 61829 1719 61863
rect 8493 61829 8527 61863
rect 1501 61761 1535 61795
rect 6653 61761 6687 61795
rect 6920 61761 6954 61795
rect 8585 61693 8619 61727
rect 8677 61693 8711 61727
rect 8033 61557 8067 61591
rect 8125 61557 8159 61591
rect 7665 61217 7699 61251
rect 7849 61217 7883 61251
rect 8493 61217 8527 61251
rect 8677 61217 8711 61251
rect 7573 61149 7607 61183
rect 8401 61149 8435 61183
rect 8953 61149 8987 61183
rect 7205 61013 7239 61047
rect 8033 61013 8067 61047
rect 9137 61013 9171 61047
rect 5181 60741 5215 60775
rect 7012 60741 7046 60775
rect 1409 60673 1443 60707
rect 4077 60673 4111 60707
rect 4445 60673 4479 60707
rect 4905 60673 4939 60707
rect 6745 60673 6779 60707
rect 8125 60537 8159 60571
rect 1593 60469 1627 60503
rect 7297 60129 7331 60163
rect 7564 60061 7598 60095
rect 1501 59993 1535 60027
rect 1593 59925 1627 59959
rect 8677 59925 8711 59959
rect 4169 59721 4203 59755
rect 9137 59721 9171 59755
rect 3985 59585 4019 59619
rect 4353 59585 4387 59619
rect 5089 59585 5123 59619
rect 7849 59585 7883 59619
rect 4905 59517 4939 59551
rect 3801 59381 3835 59415
rect 5273 59381 5307 59415
rect 6837 59177 6871 59211
rect 1501 58973 1535 59007
rect 4997 58973 5031 59007
rect 5181 58973 5215 59007
rect 5457 58973 5491 59007
rect 7113 58973 7147 59007
rect 7380 58973 7414 59007
rect 5702 58905 5736 58939
rect 1593 58837 1627 58871
rect 5365 58837 5399 58871
rect 8493 58837 8527 58871
rect 8217 58633 8251 58667
rect 6009 58497 6043 58531
rect 6745 58497 6779 58531
rect 7205 58497 7239 58531
rect 8125 58497 8159 58531
rect 8585 58497 8619 58531
rect 6561 58429 6595 58463
rect 7021 58429 7055 58463
rect 8309 58429 8343 58463
rect 6929 58361 6963 58395
rect 6193 58293 6227 58327
rect 7389 58293 7423 58327
rect 7757 58293 7791 58327
rect 8769 58293 8803 58327
rect 7113 58089 7147 58123
rect 7665 58089 7699 58123
rect 7205 57953 7239 57987
rect 8217 57953 8251 57987
rect 1501 57885 1535 57919
rect 6929 57885 6963 57919
rect 7389 57885 7423 57919
rect 8033 57885 8067 57919
rect 8125 57885 8159 57919
rect 8585 57885 8619 57919
rect 8953 57885 8987 57919
rect 1593 57749 1627 57783
rect 7573 57749 7607 57783
rect 8677 57749 8711 57783
rect 9137 57749 9171 57783
rect 4353 57545 4387 57579
rect 3893 57409 3927 57443
rect 4721 57409 4755 57443
rect 6377 57409 6411 57443
rect 6633 57409 6667 57443
rect 8033 57409 8067 57443
rect 7849 57341 7883 57375
rect 8217 57273 8251 57307
rect 4077 57205 4111 57239
rect 4537 57205 4571 57239
rect 7757 57205 7791 57239
rect 1501 56797 1535 56831
rect 4169 56797 4203 56831
rect 7573 56797 7607 56831
rect 1593 56661 1627 56695
rect 4353 56661 4387 56695
rect 7757 56661 7791 56695
rect 7573 56457 7607 56491
rect 1501 56389 1535 56423
rect 4261 56321 4295 56355
rect 4721 56321 4755 56355
rect 7481 56321 7515 56355
rect 4537 56185 4571 56219
rect 1593 56117 1627 56151
rect 4445 56117 4479 56151
rect 4169 55913 4203 55947
rect 7113 55709 7147 55743
rect 7205 55709 7239 55743
rect 7573 55709 7607 55743
rect 7665 55709 7699 55743
rect 4077 55641 4111 55675
rect 7389 55573 7423 55607
rect 7849 55573 7883 55607
rect 1501 55301 1535 55335
rect 1593 55029 1627 55063
rect 4445 54621 4479 54655
rect 6745 54621 6779 54655
rect 6929 54553 6963 54587
rect 4261 54485 4295 54519
rect 1501 54213 1535 54247
rect 7389 54213 7423 54247
rect 4445 54145 4479 54179
rect 4537 54145 4571 54179
rect 7205 54145 7239 54179
rect 7665 54145 7699 54179
rect 7847 54145 7881 54179
rect 4721 54009 4755 54043
rect 1593 53941 1627 53975
rect 4261 53941 4295 53975
rect 7573 53941 7607 53975
rect 8033 53941 8067 53975
rect 4997 53737 5031 53771
rect 4905 53533 4939 53567
rect 7205 53533 7239 53567
rect 7757 53533 7791 53567
rect 7021 53465 7055 53499
rect 7389 53397 7423 53431
rect 7941 53397 7975 53431
rect 1501 53125 1535 53159
rect 4537 53125 4571 53159
rect 4353 53057 4387 53091
rect 4813 53057 4847 53091
rect 4997 53057 5031 53091
rect 7021 53057 7055 53091
rect 7205 53057 7239 53091
rect 7665 53057 7699 53091
rect 7941 53057 7975 53091
rect 8217 53057 8251 53091
rect 4721 52989 4755 53023
rect 7389 52989 7423 53023
rect 8033 52921 8067 52955
rect 1593 52853 1627 52887
rect 5181 52853 5215 52887
rect 7481 52853 7515 52887
rect 7757 52853 7791 52887
rect 6009 52581 6043 52615
rect 8125 52581 8159 52615
rect 6193 52445 6227 52479
rect 6745 52445 6779 52479
rect 7001 52445 7035 52479
rect 1501 52377 1535 52411
rect 1593 52309 1627 52343
rect 7012 52037 7046 52071
rect 4353 51969 4387 52003
rect 6745 51901 6779 51935
rect 4537 51765 4571 51799
rect 8125 51765 8159 51799
rect 8125 51493 8159 51527
rect 1501 51357 1535 51391
rect 6285 51357 6319 51391
rect 6745 51357 6779 51391
rect 8401 51357 8435 51391
rect 8493 51357 8527 51391
rect 6469 51289 6503 51323
rect 7012 51289 7046 51323
rect 1593 51221 1627 51255
rect 6653 51221 6687 51255
rect 8217 51221 8251 51255
rect 8677 51221 8711 51255
rect 6920 50949 6954 50983
rect 6561 50881 6595 50915
rect 6653 50881 6687 50915
rect 6377 50677 6411 50711
rect 8033 50677 8067 50711
rect 1501 50269 1535 50303
rect 1593 50133 1627 50167
rect 8125 49929 8159 49963
rect 4261 49861 4295 49895
rect 4997 49861 5031 49895
rect 6920 49861 6954 49895
rect 4813 49793 4847 49827
rect 6653 49793 6687 49827
rect 8309 49793 8343 49827
rect 4721 49725 4755 49759
rect 4537 49657 4571 49691
rect 5181 49589 5215 49623
rect 8033 49589 8067 49623
rect 6469 49385 6503 49419
rect 8309 49385 8343 49419
rect 1501 49181 1535 49215
rect 6193 49181 6227 49215
rect 6745 49181 6779 49215
rect 8217 49181 8251 49215
rect 7012 49113 7046 49147
rect 1593 49045 1627 49079
rect 6653 49045 6687 49079
rect 8125 49045 8159 49079
rect 8677 49045 8711 49079
rect 1501 48773 1535 48807
rect 6920 48773 6954 48807
rect 4721 48705 4755 48739
rect 5365 48705 5399 48739
rect 5641 48705 5675 48739
rect 6653 48705 6687 48739
rect 1593 48501 1627 48535
rect 4537 48501 4571 48535
rect 8033 48501 8067 48535
rect 6653 48093 6687 48127
rect 6920 48093 6954 48127
rect 8033 47957 8067 47991
rect 1501 47685 1535 47719
rect 6929 47617 6963 47651
rect 7389 47481 7423 47515
rect 1593 47413 1627 47447
rect 7205 47413 7239 47447
rect 3801 47005 3835 47039
rect 6745 47005 6779 47039
rect 4068 46937 4102 46971
rect 7012 46937 7046 46971
rect 5181 46869 5215 46903
rect 8125 46869 8159 46903
rect 9137 46665 9171 46699
rect 1501 46597 1535 46631
rect 7849 46597 7883 46631
rect 5733 46529 5767 46563
rect 6644 46529 6678 46563
rect 6377 46461 6411 46495
rect 1593 46325 1627 46359
rect 5825 46325 5859 46359
rect 6193 46325 6227 46359
rect 7757 46325 7791 46359
rect 8309 46121 8343 46155
rect 9045 46121 9079 46155
rect 6653 45985 6687 46019
rect 8217 45917 8251 45951
rect 8953 45917 8987 45951
rect 6909 45849 6943 45883
rect 8033 45781 8067 45815
rect 8677 45781 8711 45815
rect 9413 45781 9447 45815
rect 1501 45509 1535 45543
rect 4629 45441 4663 45475
rect 4905 45441 4939 45475
rect 7205 45441 7239 45475
rect 8217 45441 8251 45475
rect 4813 45373 4847 45407
rect 4721 45305 4755 45339
rect 8401 45305 8435 45339
rect 1593 45237 1627 45271
rect 4445 45237 4479 45271
rect 7481 45237 7515 45271
rect 7665 45237 7699 45271
rect 4353 45033 4387 45067
rect 4721 44965 4755 44999
rect 4813 44965 4847 44999
rect 5365 44965 5399 44999
rect 6745 44965 6779 44999
rect 4445 44897 4479 44931
rect 7389 44897 7423 44931
rect 1409 44829 1443 44863
rect 4195 44829 4229 44863
rect 4629 44829 4663 44863
rect 4917 44829 4951 44863
rect 5273 44829 5307 44863
rect 5457 44829 5491 44863
rect 5549 44829 5583 44863
rect 7205 44829 7239 44863
rect 7113 44761 7147 44795
rect 1593 44693 1627 44727
rect 5089 44693 5123 44727
rect 4169 44489 4203 44523
rect 4343 44353 4377 44387
rect 4629 44353 4663 44387
rect 4997 44353 5031 44387
rect 5089 44353 5123 44387
rect 5181 44353 5215 44387
rect 5273 44353 5307 44387
rect 6745 44353 6779 44387
rect 7012 44353 7046 44387
rect 4445 44285 4479 44319
rect 4537 44285 4571 44319
rect 4813 44149 4847 44183
rect 8125 44149 8159 44183
rect 4353 43945 4387 43979
rect 6745 43809 6779 43843
rect 1409 43741 1443 43775
rect 4261 43741 4295 43775
rect 7012 43741 7046 43775
rect 1593 43605 1627 43639
rect 4721 43605 4755 43639
rect 8125 43605 8159 43639
rect 7012 43333 7046 43367
rect 6745 43265 6779 43299
rect 8125 43061 8159 43095
rect 4813 42789 4847 42823
rect 4905 42721 4939 42755
rect 5549 42721 5583 42755
rect 7113 42721 7147 42755
rect 4077 42653 4111 42687
rect 4261 42653 4295 42687
rect 4721 42653 4755 42687
rect 4997 42653 5031 42687
rect 5365 42653 5399 42687
rect 5457 42653 5491 42687
rect 5641 42653 5675 42687
rect 1501 42585 1535 42619
rect 1869 42585 1903 42619
rect 4445 42585 4479 42619
rect 6837 42585 6871 42619
rect 4537 42517 4571 42551
rect 5181 42517 5215 42551
rect 6469 42517 6503 42551
rect 6929 42517 6963 42551
rect 7012 42245 7046 42279
rect 6745 42177 6779 42211
rect 8125 41973 8159 42007
rect 4445 41701 4479 41735
rect 4537 41701 4571 41735
rect 4353 41565 4387 41599
rect 4629 41565 4663 41599
rect 1501 41497 1535 41531
rect 1869 41497 1903 41531
rect 4169 41429 4203 41463
rect 1501 41089 1535 41123
rect 1777 40885 1811 40919
rect 7665 40545 7699 40579
rect 7389 40477 7423 40511
rect 4537 40409 4571 40443
rect 4721 40409 4755 40443
rect 7481 40409 7515 40443
rect 7021 40341 7055 40375
rect 6929 40137 6963 40171
rect 7389 40137 7423 40171
rect 8125 40137 8159 40171
rect 8585 40137 8619 40171
rect 8953 40137 8987 40171
rect 1501 40069 1535 40103
rect 7297 40069 7331 40103
rect 9045 40001 9079 40035
rect 7573 39933 7607 39967
rect 8217 39933 8251 39967
rect 8309 39933 8343 39967
rect 9229 39933 9263 39967
rect 1777 39797 1811 39831
rect 7757 39797 7791 39831
rect 4445 39593 4479 39627
rect 7389 39525 7423 39559
rect 7205 39457 7239 39491
rect 7849 39457 7883 39491
rect 7941 39457 7975 39491
rect 4353 39389 4387 39423
rect 6929 39389 6963 39423
rect 7021 39321 7055 39355
rect 4813 39253 4847 39287
rect 6561 39253 6595 39287
rect 7757 39253 7791 39287
rect 6653 39049 6687 39083
rect 7481 39049 7515 39083
rect 7849 38981 7883 39015
rect 1501 38913 1535 38947
rect 7389 38913 7423 38947
rect 7665 38845 7699 38879
rect 1777 38709 1811 38743
rect 7021 38709 7055 38743
rect 9321 38709 9355 38743
rect 7573 38437 7607 38471
rect 8125 38301 8159 38335
rect 7849 38233 7883 38267
rect 8033 38165 8067 38199
rect 7021 37961 7055 37995
rect 8033 37961 8067 37995
rect 7113 37893 7147 37927
rect 1501 37825 1535 37859
rect 7297 37757 7331 37791
rect 7941 37757 7975 37791
rect 8125 37757 8159 37791
rect 1777 37621 1811 37655
rect 6653 37621 6687 37655
rect 7573 37621 7607 37655
rect 6929 37281 6963 37315
rect 7665 37281 7699 37315
rect 7757 37281 7791 37315
rect 1409 37213 1443 37247
rect 1685 37145 1719 37179
rect 7205 37077 7239 37111
rect 7573 37077 7607 37111
rect 8585 36873 8619 36907
rect 8585 36669 8619 36703
rect 8677 36669 8711 36703
rect 8125 36533 8159 36567
rect 8769 36193 8803 36227
rect 1409 36125 1443 36159
rect 8033 36125 8067 36159
rect 8125 36125 8159 36159
rect 8309 36125 8343 36159
rect 1685 36057 1719 36091
rect 7389 36057 7423 36091
rect 7481 35989 7515 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 8115 34697 8149 34731
rect 8585 34629 8619 34663
rect 8585 34493 8619 34527
rect 8677 34493 8711 34527
rect 8125 34085 8159 34119
rect 8585 34017 8619 34051
rect 1409 33949 1443 33983
rect 8585 33881 8619 33915
rect 8677 33881 8711 33915
rect 1593 33813 1627 33847
rect 8585 33609 8619 33643
rect 1501 33473 1535 33507
rect 8401 33473 8435 33507
rect 8677 33473 8711 33507
rect 8125 33337 8159 33371
rect 1777 33269 1811 33303
rect 8033 32997 8067 33031
rect 8585 32929 8619 32963
rect 8309 32793 8343 32827
rect 8493 32725 8527 32759
rect 7205 32521 7239 32555
rect 6469 32453 6503 32487
rect 1501 32385 1535 32419
rect 7297 32385 7331 32419
rect 7389 32317 7423 32351
rect 1777 32181 1811 32215
rect 6561 32181 6595 32215
rect 6837 32181 6871 32215
rect 8033 31977 8067 32011
rect 7021 31909 7055 31943
rect 7573 31841 7607 31875
rect 7481 31773 7515 31807
rect 8309 31773 8343 31807
rect 8585 31773 8619 31807
rect 7389 31705 7423 31739
rect 8493 31705 8527 31739
rect 1593 31297 1627 31331
rect 1409 31093 1443 31127
rect 7665 30277 7699 30311
rect 1593 30209 1627 30243
rect 7481 30209 7515 30243
rect 1409 30005 1443 30039
rect 1593 29597 1627 29631
rect 1409 29461 1443 29495
rect 8769 29257 8803 29291
rect 7481 29189 7515 29223
rect 8861 29189 8895 29223
rect 7297 29121 7331 29155
rect 8769 29053 8803 29087
rect 8309 28985 8343 29019
rect 7113 28713 7147 28747
rect 8125 28645 8159 28679
rect 7665 28577 7699 28611
rect 8585 28577 8619 28611
rect 1593 28509 1627 28543
rect 7481 28509 7515 28543
rect 8677 28509 8711 28543
rect 8585 28441 8619 28475
rect 1409 28373 1443 28407
rect 7573 28373 7607 28407
rect 7389 27625 7423 27659
rect 1409 27421 1443 27455
rect 1685 27353 1719 27387
rect 7297 27353 7331 27387
rect 7665 27081 7699 27115
rect 7757 27081 7791 27115
rect 7021 27013 7055 27047
rect 7849 26877 7883 26911
rect 7297 26741 7331 26775
rect 6561 26537 6595 26571
rect 9505 26537 9539 26571
rect 7297 26469 7331 26503
rect 7849 26401 7883 26435
rect 1409 26333 1443 26367
rect 3985 26333 4019 26367
rect 6837 26333 6871 26367
rect 6929 26333 6963 26367
rect 7021 26333 7055 26367
rect 7205 26333 7239 26367
rect 9229 26333 9263 26367
rect 1685 26265 1719 26299
rect 7665 26265 7699 26299
rect 7757 26265 7791 26299
rect 4169 26197 4203 26231
rect 1593 25993 1627 26027
rect 7573 25993 7607 26027
rect 8401 25993 8435 26027
rect 9137 25993 9171 26027
rect 9045 25925 9079 25959
rect 1501 25857 1535 25891
rect 4169 25857 4203 25891
rect 5825 25857 5859 25891
rect 6003 25857 6037 25891
rect 6929 25789 6963 25823
rect 7665 25789 7699 25823
rect 7757 25789 7791 25823
rect 8493 25789 8527 25823
rect 8585 25789 8619 25823
rect 5825 25721 5859 25755
rect 4353 25653 4387 25687
rect 7205 25653 7239 25687
rect 8033 25653 8067 25687
rect 7573 25449 7607 25483
rect 7481 25245 7515 25279
rect 1409 24769 1443 24803
rect 1593 24565 1627 24599
rect 9321 24361 9355 24395
rect 7297 24293 7331 24327
rect 8125 24293 8159 24327
rect 7849 24225 7883 24259
rect 4169 24157 4203 24191
rect 7113 24157 7147 24191
rect 7757 24157 7791 24191
rect 8309 24157 8343 24191
rect 8401 24157 8435 24191
rect 9229 24157 9263 24191
rect 6929 24089 6963 24123
rect 8125 24089 8159 24123
rect 4353 24021 4387 24055
rect 7665 24021 7699 24055
rect 1593 23817 1627 23851
rect 1409 23681 1443 23715
rect 4353 23681 4387 23715
rect 4537 23477 4571 23511
rect 8677 23273 8711 23307
rect 9505 23205 9539 23239
rect 4169 23069 4203 23103
rect 8493 23069 8527 23103
rect 9229 23069 9263 23103
rect 4353 22933 4387 22967
rect 1685 22661 1719 22695
rect 7757 22661 7791 22695
rect 1501 22593 1535 22627
rect 4077 22593 4111 22627
rect 4353 22593 4387 22627
rect 4261 22389 4295 22423
rect 4537 22389 4571 22423
rect 7849 22389 7883 22423
rect 1409 21981 1443 22015
rect 4077 21981 4111 22015
rect 9321 21981 9355 22015
rect 1685 21913 1719 21947
rect 4261 21845 4295 21879
rect 9505 21845 9539 21879
rect 7205 21505 7239 21539
rect 7389 21505 7423 21539
rect 7573 21301 7607 21335
rect 1409 20893 1443 20927
rect 1685 20825 1719 20859
rect 9321 20417 9355 20451
rect 9505 20213 9539 20247
rect 1409 19805 1443 19839
rect 9321 19805 9355 19839
rect 1685 19737 1719 19771
rect 9505 19669 9539 19703
rect 2237 18785 2271 18819
rect 7389 18717 7423 18751
rect 7481 18717 7515 18751
rect 7665 18717 7699 18751
rect 7757 18717 7791 18751
rect 1409 18649 1443 18683
rect 7205 18581 7239 18615
rect 1501 18309 1535 18343
rect 1593 18037 1627 18071
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 7849 17493 7883 17527
rect 1501 17221 1535 17255
rect 7481 17153 7515 17187
rect 1593 16949 1627 16983
rect 7665 16949 7699 16983
rect 7297 16745 7331 16779
rect 8125 16677 8159 16711
rect 8217 16677 8251 16711
rect 7573 16541 7607 16575
rect 7757 16541 7791 16575
rect 8033 16541 8067 16575
rect 8309 16541 8343 16575
rect 9321 16541 9355 16575
rect 7481 16405 7515 16439
rect 7849 16405 7883 16439
rect 9505 16405 9539 16439
rect 1501 16133 1535 16167
rect 9229 16133 9263 16167
rect 9413 16133 9447 16167
rect 9505 15997 9539 16031
rect 1593 15861 1627 15895
rect 8953 15861 8987 15895
rect 9321 15453 9355 15487
rect 9505 15317 9539 15351
rect 1501 15045 1535 15079
rect 1593 14773 1627 14807
rect 8125 14501 8159 14535
rect 8585 14433 8619 14467
rect 1501 14365 1535 14399
rect 8677 14365 8711 14399
rect 9321 14365 9355 14399
rect 8585 14297 8619 14331
rect 1593 14229 1627 14263
rect 9505 14229 9539 14263
rect 7757 13345 7791 13379
rect 1501 13277 1535 13311
rect 8033 13277 8067 13311
rect 1593 13141 1627 13175
rect 8769 13141 8803 13175
rect 1501 12189 1535 12223
rect 1593 12053 1627 12087
rect 8861 11713 8895 11747
rect 8585 11645 8619 11679
rect 9597 11509 9631 11543
rect 1593 11305 1627 11339
rect 8769 11237 8803 11271
rect 7757 11169 7791 11203
rect 1501 11101 1535 11135
rect 8033 11101 8067 11135
rect 1501 10693 1535 10727
rect 1593 10421 1627 10455
rect 1501 9605 1535 9639
rect 8861 9537 8895 9571
rect 8585 9469 8619 9503
rect 1593 9333 1627 9367
rect 9597 9333 9631 9367
rect 1501 8517 1535 8551
rect 1685 8313 1719 8347
rect 1501 7429 1535 7463
rect 1593 7157 1627 7191
rect 1501 6749 1535 6783
rect 1593 6613 1627 6647
rect 1501 5661 1535 5695
rect 1593 5525 1627 5559
rect 1501 4573 1535 4607
rect 1593 4437 1627 4471
rect 1501 3485 1535 3519
rect 1593 3349 1627 3383
rect 27537 1377 27571 1411
rect 34713 1377 34747 1411
rect 35817 1377 35851 1411
rect 22845 1309 22879 1343
rect 26157 1309 26191 1343
rect 27813 1309 27847 1343
rect 28457 1309 28491 1343
rect 29653 1309 29687 1343
rect 32137 1309 32171 1343
rect 32413 1309 32447 1343
rect 33609 1309 33643 1343
rect 33885 1309 33919 1343
rect 34989 1309 35023 1343
rect 37473 1309 37507 1343
rect 37749 1309 37783 1343
rect 23213 1241 23247 1275
rect 23397 1241 23431 1275
rect 24501 1241 24535 1275
rect 24685 1241 24719 1275
rect 27077 1241 27111 1275
rect 27261 1241 27295 1275
rect 30573 1241 30607 1275
rect 22937 1173 22971 1207
rect 26341 1173 26375 1207
rect 28641 1173 28675 1207
rect 29745 1173 29779 1207
rect 30113 1173 30147 1207
rect 30665 1173 30699 1207
rect 38577 1173 38611 1207
<< metal1 >>
rect 36538 87592 36544 87644
rect 36596 87632 36602 87644
rect 47302 87632 47308 87644
rect 36596 87604 47308 87632
rect 36596 87592 36602 87604
rect 47302 87592 47308 87604
rect 47360 87592 47366 87644
rect 27522 87524 27528 87576
rect 27580 87564 27586 87576
rect 41690 87564 41696 87576
rect 27580 87536 41696 87564
rect 27580 87524 27586 87536
rect 41690 87524 41696 87536
rect 41748 87524 41754 87576
rect 33870 87456 33876 87508
rect 33928 87496 33934 87508
rect 47854 87496 47860 87508
rect 33928 87468 47860 87496
rect 33928 87456 33934 87468
rect 47854 87456 47860 87468
rect 47912 87456 47918 87508
rect 37642 87388 37648 87440
rect 37700 87428 37706 87440
rect 53558 87428 53564 87440
rect 37700 87400 53564 87428
rect 37700 87388 37706 87400
rect 53558 87388 53564 87400
rect 53616 87388 53622 87440
rect 3418 87320 3424 87372
rect 3476 87360 3482 87372
rect 91278 87360 91284 87372
rect 3476 87332 91284 87360
rect 3476 87320 3482 87332
rect 91278 87320 91284 87332
rect 91336 87320 91342 87372
rect 11330 87252 11336 87304
rect 11388 87292 11394 87304
rect 30190 87292 30196 87304
rect 11388 87264 30196 87292
rect 11388 87252 11394 87264
rect 30190 87252 30196 87264
rect 30248 87252 30254 87304
rect 30374 87252 30380 87304
rect 30432 87292 30438 87304
rect 44818 87292 44824 87304
rect 30432 87264 44824 87292
rect 30432 87252 30438 87264
rect 44818 87252 44824 87264
rect 44876 87252 44882 87304
rect 1302 87184 1308 87236
rect 1360 87224 1366 87236
rect 17310 87224 17316 87236
rect 1360 87196 17316 87224
rect 1360 87184 1366 87196
rect 17310 87184 17316 87196
rect 17368 87184 17374 87236
rect 30208 87224 30236 87252
rect 44910 87224 44916 87236
rect 30208 87196 44916 87224
rect 44910 87184 44916 87196
rect 44968 87184 44974 87236
rect 45094 87184 45100 87236
rect 45152 87224 45158 87236
rect 63494 87224 63500 87236
rect 45152 87196 63500 87224
rect 45152 87184 45158 87196
rect 63494 87184 63500 87196
rect 63552 87184 63558 87236
rect 9030 87116 9036 87168
rect 9088 87156 9094 87168
rect 24762 87156 24768 87168
rect 9088 87128 24768 87156
rect 9088 87116 9094 87128
rect 24762 87116 24768 87128
rect 24820 87156 24826 87168
rect 35342 87156 35348 87168
rect 24820 87128 35348 87156
rect 24820 87116 24826 87128
rect 35342 87116 35348 87128
rect 35400 87156 35406 87168
rect 72142 87156 72148 87168
rect 35400 87128 44588 87156
rect 35400 87116 35406 87128
rect 10778 87048 10784 87100
rect 10836 87088 10842 87100
rect 41782 87088 41788 87100
rect 10836 87060 41788 87088
rect 10836 87048 10842 87060
rect 41782 87048 41788 87060
rect 41840 87048 41846 87100
rect 44560 87088 44588 87128
rect 44744 87128 72148 87156
rect 44744 87088 44772 87128
rect 72142 87116 72148 87128
rect 72200 87116 72206 87168
rect 77662 87088 77668 87100
rect 44560 87060 44772 87088
rect 51046 87060 77668 87088
rect 10410 86980 10416 87032
rect 10468 87020 10474 87032
rect 36538 87020 36544 87032
rect 10468 86992 36544 87020
rect 10468 86980 10474 86992
rect 36538 86980 36544 86992
rect 36596 86980 36602 87032
rect 44910 86980 44916 87032
rect 44968 87020 44974 87032
rect 51046 87020 51074 87060
rect 77662 87048 77668 87060
rect 77720 87048 77726 87100
rect 44968 86992 51074 87020
rect 44968 86980 44974 86992
rect 11422 86912 11428 86964
rect 11480 86952 11486 86964
rect 50798 86952 50804 86964
rect 11480 86924 50804 86952
rect 11480 86912 11486 86924
rect 50798 86912 50804 86924
rect 50856 86912 50862 86964
rect 10502 86844 10508 86896
rect 10560 86884 10566 86896
rect 62482 86884 62488 86896
rect 10560 86856 62488 86884
rect 10560 86844 10566 86856
rect 62482 86844 62488 86856
rect 62540 86844 62546 86896
rect 4890 86776 4896 86828
rect 4948 86816 4954 86828
rect 58342 86816 58348 86828
rect 4948 86788 58348 86816
rect 4948 86776 4954 86788
rect 58342 86776 58348 86788
rect 58400 86776 58406 86828
rect 5534 86708 5540 86760
rect 5592 86748 5598 86760
rect 61010 86748 61016 86760
rect 5592 86720 61016 86748
rect 5592 86708 5598 86720
rect 61010 86708 61016 86720
rect 61068 86708 61074 86760
rect 11514 86640 11520 86692
rect 11572 86680 11578 86692
rect 68094 86680 68100 86692
rect 11572 86652 68100 86680
rect 11572 86640 11578 86652
rect 68094 86640 68100 86652
rect 68152 86640 68158 86692
rect 10594 86572 10600 86624
rect 10652 86612 10658 86624
rect 68002 86612 68008 86624
rect 10652 86584 68008 86612
rect 10652 86572 10658 86584
rect 68002 86572 68008 86584
rect 68060 86572 68066 86624
rect 1104 86522 108836 86544
rect 1104 86470 3610 86522
rect 3662 86470 3674 86522
rect 3726 86470 3738 86522
rect 3790 86470 3802 86522
rect 3854 86470 3866 86522
rect 3918 86470 5210 86522
rect 5262 86470 5274 86522
rect 5326 86470 5338 86522
rect 5390 86470 5402 86522
rect 5454 86470 5466 86522
rect 5518 86470 6810 86522
rect 6862 86470 6874 86522
rect 6926 86470 6938 86522
rect 6990 86470 7002 86522
rect 7054 86470 7066 86522
rect 7118 86470 8410 86522
rect 8462 86470 8474 86522
rect 8526 86470 8538 86522
rect 8590 86470 8602 86522
rect 8654 86470 8666 86522
rect 8718 86470 10010 86522
rect 10062 86470 10074 86522
rect 10126 86470 10138 86522
rect 10190 86470 10202 86522
rect 10254 86470 10266 86522
rect 10318 86470 11610 86522
rect 11662 86470 11674 86522
rect 11726 86470 11738 86522
rect 11790 86470 11802 86522
rect 11854 86470 11866 86522
rect 11918 86470 13210 86522
rect 13262 86470 13274 86522
rect 13326 86470 13338 86522
rect 13390 86470 13402 86522
rect 13454 86470 13466 86522
rect 13518 86470 14810 86522
rect 14862 86470 14874 86522
rect 14926 86470 14938 86522
rect 14990 86470 15002 86522
rect 15054 86470 15066 86522
rect 15118 86470 16410 86522
rect 16462 86470 16474 86522
rect 16526 86470 16538 86522
rect 16590 86470 16602 86522
rect 16654 86470 16666 86522
rect 16718 86470 18010 86522
rect 18062 86470 18074 86522
rect 18126 86470 18138 86522
rect 18190 86470 18202 86522
rect 18254 86470 18266 86522
rect 18318 86470 19610 86522
rect 19662 86470 19674 86522
rect 19726 86470 19738 86522
rect 19790 86470 19802 86522
rect 19854 86470 19866 86522
rect 19918 86470 21210 86522
rect 21262 86470 21274 86522
rect 21326 86470 21338 86522
rect 21390 86470 21402 86522
rect 21454 86470 21466 86522
rect 21518 86470 22810 86522
rect 22862 86470 22874 86522
rect 22926 86470 22938 86522
rect 22990 86470 23002 86522
rect 23054 86470 23066 86522
rect 23118 86470 24410 86522
rect 24462 86470 24474 86522
rect 24526 86470 24538 86522
rect 24590 86470 24602 86522
rect 24654 86470 24666 86522
rect 24718 86470 26010 86522
rect 26062 86470 26074 86522
rect 26126 86470 26138 86522
rect 26190 86470 26202 86522
rect 26254 86470 26266 86522
rect 26318 86470 27610 86522
rect 27662 86470 27674 86522
rect 27726 86470 27738 86522
rect 27790 86470 27802 86522
rect 27854 86470 27866 86522
rect 27918 86470 29210 86522
rect 29262 86470 29274 86522
rect 29326 86470 29338 86522
rect 29390 86470 29402 86522
rect 29454 86470 29466 86522
rect 29518 86470 30810 86522
rect 30862 86470 30874 86522
rect 30926 86470 30938 86522
rect 30990 86470 31002 86522
rect 31054 86470 31066 86522
rect 31118 86470 32410 86522
rect 32462 86470 32474 86522
rect 32526 86470 32538 86522
rect 32590 86470 32602 86522
rect 32654 86470 32666 86522
rect 32718 86470 34010 86522
rect 34062 86470 34074 86522
rect 34126 86470 34138 86522
rect 34190 86470 34202 86522
rect 34254 86470 34266 86522
rect 34318 86470 35610 86522
rect 35662 86470 35674 86522
rect 35726 86470 35738 86522
rect 35790 86470 35802 86522
rect 35854 86470 35866 86522
rect 35918 86470 37210 86522
rect 37262 86470 37274 86522
rect 37326 86470 37338 86522
rect 37390 86470 37402 86522
rect 37454 86470 37466 86522
rect 37518 86470 38810 86522
rect 38862 86470 38874 86522
rect 38926 86470 38938 86522
rect 38990 86470 39002 86522
rect 39054 86470 39066 86522
rect 39118 86470 40410 86522
rect 40462 86470 40474 86522
rect 40526 86470 40538 86522
rect 40590 86470 40602 86522
rect 40654 86470 40666 86522
rect 40718 86470 42010 86522
rect 42062 86470 42074 86522
rect 42126 86470 42138 86522
rect 42190 86470 42202 86522
rect 42254 86470 42266 86522
rect 42318 86470 43610 86522
rect 43662 86470 43674 86522
rect 43726 86470 43738 86522
rect 43790 86470 43802 86522
rect 43854 86470 43866 86522
rect 43918 86470 45210 86522
rect 45262 86470 45274 86522
rect 45326 86470 45338 86522
rect 45390 86470 45402 86522
rect 45454 86470 45466 86522
rect 45518 86470 46810 86522
rect 46862 86470 46874 86522
rect 46926 86470 46938 86522
rect 46990 86470 47002 86522
rect 47054 86470 47066 86522
rect 47118 86470 48410 86522
rect 48462 86470 48474 86522
rect 48526 86470 48538 86522
rect 48590 86470 48602 86522
rect 48654 86470 48666 86522
rect 48718 86470 50010 86522
rect 50062 86470 50074 86522
rect 50126 86470 50138 86522
rect 50190 86470 50202 86522
rect 50254 86470 50266 86522
rect 50318 86470 51610 86522
rect 51662 86470 51674 86522
rect 51726 86470 51738 86522
rect 51790 86470 51802 86522
rect 51854 86470 51866 86522
rect 51918 86470 53210 86522
rect 53262 86470 53274 86522
rect 53326 86470 53338 86522
rect 53390 86470 53402 86522
rect 53454 86470 53466 86522
rect 53518 86470 54810 86522
rect 54862 86470 54874 86522
rect 54926 86470 54938 86522
rect 54990 86470 55002 86522
rect 55054 86470 55066 86522
rect 55118 86470 56410 86522
rect 56462 86470 56474 86522
rect 56526 86470 56538 86522
rect 56590 86470 56602 86522
rect 56654 86470 56666 86522
rect 56718 86470 58010 86522
rect 58062 86470 58074 86522
rect 58126 86470 58138 86522
rect 58190 86470 58202 86522
rect 58254 86470 58266 86522
rect 58318 86470 59610 86522
rect 59662 86470 59674 86522
rect 59726 86470 59738 86522
rect 59790 86470 59802 86522
rect 59854 86470 59866 86522
rect 59918 86470 61210 86522
rect 61262 86470 61274 86522
rect 61326 86470 61338 86522
rect 61390 86470 61402 86522
rect 61454 86470 61466 86522
rect 61518 86470 62810 86522
rect 62862 86470 62874 86522
rect 62926 86470 62938 86522
rect 62990 86470 63002 86522
rect 63054 86470 63066 86522
rect 63118 86470 64410 86522
rect 64462 86470 64474 86522
rect 64526 86470 64538 86522
rect 64590 86470 64602 86522
rect 64654 86470 64666 86522
rect 64718 86470 66010 86522
rect 66062 86470 66074 86522
rect 66126 86470 66138 86522
rect 66190 86470 66202 86522
rect 66254 86470 66266 86522
rect 66318 86470 67610 86522
rect 67662 86470 67674 86522
rect 67726 86470 67738 86522
rect 67790 86470 67802 86522
rect 67854 86470 67866 86522
rect 67918 86470 69210 86522
rect 69262 86470 69274 86522
rect 69326 86470 69338 86522
rect 69390 86470 69402 86522
rect 69454 86470 69466 86522
rect 69518 86470 70810 86522
rect 70862 86470 70874 86522
rect 70926 86470 70938 86522
rect 70990 86470 71002 86522
rect 71054 86470 71066 86522
rect 71118 86470 72410 86522
rect 72462 86470 72474 86522
rect 72526 86470 72538 86522
rect 72590 86470 72602 86522
rect 72654 86470 72666 86522
rect 72718 86470 74010 86522
rect 74062 86470 74074 86522
rect 74126 86470 74138 86522
rect 74190 86470 74202 86522
rect 74254 86470 74266 86522
rect 74318 86470 75610 86522
rect 75662 86470 75674 86522
rect 75726 86470 75738 86522
rect 75790 86470 75802 86522
rect 75854 86470 75866 86522
rect 75918 86470 77210 86522
rect 77262 86470 77274 86522
rect 77326 86470 77338 86522
rect 77390 86470 77402 86522
rect 77454 86470 77466 86522
rect 77518 86470 78810 86522
rect 78862 86470 78874 86522
rect 78926 86470 78938 86522
rect 78990 86470 79002 86522
rect 79054 86470 79066 86522
rect 79118 86470 80410 86522
rect 80462 86470 80474 86522
rect 80526 86470 80538 86522
rect 80590 86470 80602 86522
rect 80654 86470 80666 86522
rect 80718 86470 82010 86522
rect 82062 86470 82074 86522
rect 82126 86470 82138 86522
rect 82190 86470 82202 86522
rect 82254 86470 82266 86522
rect 82318 86470 83610 86522
rect 83662 86470 83674 86522
rect 83726 86470 83738 86522
rect 83790 86470 83802 86522
rect 83854 86470 83866 86522
rect 83918 86470 85210 86522
rect 85262 86470 85274 86522
rect 85326 86470 85338 86522
rect 85390 86470 85402 86522
rect 85454 86470 85466 86522
rect 85518 86470 86810 86522
rect 86862 86470 86874 86522
rect 86926 86470 86938 86522
rect 86990 86470 87002 86522
rect 87054 86470 87066 86522
rect 87118 86470 88410 86522
rect 88462 86470 88474 86522
rect 88526 86470 88538 86522
rect 88590 86470 88602 86522
rect 88654 86470 88666 86522
rect 88718 86470 90010 86522
rect 90062 86470 90074 86522
rect 90126 86470 90138 86522
rect 90190 86470 90202 86522
rect 90254 86470 90266 86522
rect 90318 86470 91610 86522
rect 91662 86470 91674 86522
rect 91726 86470 91738 86522
rect 91790 86470 91802 86522
rect 91854 86470 91866 86522
rect 91918 86470 93210 86522
rect 93262 86470 93274 86522
rect 93326 86470 93338 86522
rect 93390 86470 93402 86522
rect 93454 86470 93466 86522
rect 93518 86470 94810 86522
rect 94862 86470 94874 86522
rect 94926 86470 94938 86522
rect 94990 86470 95002 86522
rect 95054 86470 95066 86522
rect 95118 86470 96410 86522
rect 96462 86470 96474 86522
rect 96526 86470 96538 86522
rect 96590 86470 96602 86522
rect 96654 86470 96666 86522
rect 96718 86470 98010 86522
rect 98062 86470 98074 86522
rect 98126 86470 98138 86522
rect 98190 86470 98202 86522
rect 98254 86470 98266 86522
rect 98318 86470 99610 86522
rect 99662 86470 99674 86522
rect 99726 86470 99738 86522
rect 99790 86470 99802 86522
rect 99854 86470 99866 86522
rect 99918 86470 101210 86522
rect 101262 86470 101274 86522
rect 101326 86470 101338 86522
rect 101390 86470 101402 86522
rect 101454 86470 101466 86522
rect 101518 86470 102810 86522
rect 102862 86470 102874 86522
rect 102926 86470 102938 86522
rect 102990 86470 103002 86522
rect 103054 86470 103066 86522
rect 103118 86470 104410 86522
rect 104462 86470 104474 86522
rect 104526 86470 104538 86522
rect 104590 86470 104602 86522
rect 104654 86470 104666 86522
rect 104718 86470 106010 86522
rect 106062 86470 106074 86522
rect 106126 86470 106138 86522
rect 106190 86470 106202 86522
rect 106254 86470 106266 86522
rect 106318 86470 107610 86522
rect 107662 86470 107674 86522
rect 107726 86470 107738 86522
rect 107790 86470 107802 86522
rect 107854 86470 107866 86522
rect 107918 86470 108836 86522
rect 1104 86448 108836 86470
rect 5994 86368 6000 86420
rect 6052 86408 6058 86420
rect 13722 86408 13728 86420
rect 6052 86380 13728 86408
rect 6052 86368 6058 86380
rect 13722 86368 13728 86380
rect 13780 86368 13786 86420
rect 33597 86411 33655 86417
rect 33597 86408 33609 86411
rect 13832 86380 33609 86408
rect 5902 86300 5908 86352
rect 5960 86340 5966 86352
rect 13832 86340 13860 86380
rect 33597 86377 33609 86380
rect 33643 86377 33655 86411
rect 33597 86371 33655 86377
rect 34808 86380 40632 86408
rect 34808 86352 34836 86380
rect 24489 86343 24547 86349
rect 24489 86340 24501 86343
rect 5960 86312 13860 86340
rect 17144 86312 24501 86340
rect 5960 86300 5966 86312
rect 4338 86232 4344 86284
rect 4396 86272 4402 86284
rect 16942 86272 16948 86284
rect 4396 86244 16948 86272
rect 4396 86232 4402 86244
rect 16942 86232 16948 86244
rect 17000 86232 17006 86284
rect 4982 86164 4988 86216
rect 5040 86204 5046 86216
rect 17144 86204 17172 86312
rect 24489 86309 24501 86312
rect 24535 86309 24547 86343
rect 29917 86343 29975 86349
rect 29917 86340 29929 86343
rect 24489 86303 24547 86309
rect 24964 86312 29929 86340
rect 17218 86232 17224 86284
rect 17276 86272 17282 86284
rect 24964 86272 24992 86312
rect 29917 86309 29929 86312
rect 29963 86309 29975 86343
rect 29917 86303 29975 86309
rect 34790 86300 34796 86352
rect 34848 86300 34854 86352
rect 37366 86300 37372 86352
rect 37424 86300 37430 86352
rect 17276 86244 24992 86272
rect 17276 86232 17282 86244
rect 25038 86232 25044 86284
rect 25096 86232 25102 86284
rect 27154 86232 27160 86284
rect 27212 86272 27218 86284
rect 27212 86244 35204 86272
rect 27212 86232 27218 86244
rect 26786 86204 26792 86216
rect 5040 86176 17172 86204
rect 17236 86176 26792 86204
rect 5040 86164 5046 86176
rect 11974 86096 11980 86148
rect 12032 86136 12038 86148
rect 17236 86136 17264 86176
rect 26786 86164 26792 86176
rect 26844 86164 26850 86216
rect 26896 86176 27476 86204
rect 12032 86108 17264 86136
rect 12032 86096 12038 86108
rect 17310 86096 17316 86148
rect 17368 86136 17374 86148
rect 19411 86139 19469 86145
rect 19411 86136 19423 86139
rect 17368 86108 19423 86136
rect 17368 86096 17374 86108
rect 19411 86105 19423 86108
rect 19457 86105 19469 86139
rect 19411 86099 19469 86105
rect 19702 86096 19708 86148
rect 19760 86096 19766 86148
rect 19794 86096 19800 86148
rect 19852 86136 19858 86148
rect 19889 86139 19947 86145
rect 19889 86136 19901 86139
rect 19852 86108 19901 86136
rect 19852 86096 19858 86108
rect 19889 86105 19901 86108
rect 19935 86105 19947 86139
rect 19889 86099 19947 86105
rect 19978 86096 19984 86148
rect 20036 86096 20042 86148
rect 24762 86096 24768 86148
rect 24820 86096 24826 86148
rect 26896 86136 26924 86176
rect 27341 86139 27399 86145
rect 27341 86136 27353 86139
rect 24872 86108 26924 86136
rect 26988 86108 27353 86136
rect 8754 86028 8760 86080
rect 8812 86068 8818 86080
rect 24872 86068 24900 86108
rect 8812 86040 24900 86068
rect 8812 86028 8818 86040
rect 24946 86028 24952 86080
rect 25004 86028 25010 86080
rect 26786 86028 26792 86080
rect 26844 86068 26850 86080
rect 26988 86068 27016 86108
rect 27341 86105 27353 86108
rect 27387 86105 27399 86139
rect 27448 86136 27476 86176
rect 27614 86164 27620 86216
rect 27672 86164 27678 86216
rect 30006 86204 30012 86216
rect 27724 86176 30012 86204
rect 27724 86136 27752 86176
rect 30006 86164 30012 86176
rect 30064 86164 30070 86216
rect 30668 86176 34192 86204
rect 27448 86108 27752 86136
rect 27341 86099 27399 86105
rect 30190 86096 30196 86148
rect 30248 86096 30254 86148
rect 30469 86139 30527 86145
rect 30469 86136 30481 86139
rect 30300 86108 30481 86136
rect 26844 86040 27016 86068
rect 27047 86071 27105 86077
rect 26844 86028 26850 86040
rect 27047 86037 27059 86071
rect 27093 86068 27105 86071
rect 27246 86068 27252 86080
rect 27093 86040 27252 86068
rect 27093 86037 27105 86040
rect 27047 86031 27105 86037
rect 27246 86028 27252 86040
rect 27304 86028 27310 86080
rect 27522 86028 27528 86080
rect 27580 86028 27586 86080
rect 27614 86028 27620 86080
rect 27672 86068 27678 86080
rect 30300 86068 30328 86108
rect 30469 86105 30481 86108
rect 30515 86136 30527 86139
rect 30668 86136 30696 86176
rect 30515 86108 30696 86136
rect 30515 86105 30527 86108
rect 30469 86099 30527 86105
rect 33870 86096 33876 86148
rect 33928 86096 33934 86148
rect 33962 86096 33968 86148
rect 34020 86136 34026 86148
rect 34164 86145 34192 86176
rect 34790 86164 34796 86216
rect 34848 86204 34854 86216
rect 35069 86207 35127 86213
rect 35069 86204 35081 86207
rect 34848 86176 35081 86204
rect 34848 86164 34854 86176
rect 35069 86173 35081 86176
rect 35115 86173 35127 86207
rect 35176 86204 35204 86244
rect 36078 86232 36084 86284
rect 36136 86272 36142 86284
rect 39209 86275 39267 86281
rect 39209 86272 39221 86275
rect 36136 86244 39221 86272
rect 36136 86232 36142 86244
rect 39209 86241 39221 86244
rect 39255 86272 39267 86275
rect 39577 86275 39635 86281
rect 39577 86272 39589 86275
rect 39255 86244 39589 86272
rect 39255 86241 39267 86244
rect 39209 86235 39267 86241
rect 39577 86241 39589 86244
rect 39623 86272 39635 86275
rect 40037 86275 40095 86281
rect 40037 86272 40049 86275
rect 39623 86244 40049 86272
rect 39623 86241 39635 86244
rect 39577 86235 39635 86241
rect 40037 86241 40049 86244
rect 40083 86272 40095 86275
rect 40402 86272 40408 86284
rect 40083 86244 40408 86272
rect 40083 86241 40095 86244
rect 40037 86235 40095 86241
rect 40402 86232 40408 86244
rect 40460 86232 40466 86284
rect 40604 86281 40632 86380
rect 40770 86368 40776 86420
rect 40828 86408 40834 86420
rect 40828 86380 41644 86408
rect 40828 86368 40834 86380
rect 41616 86340 41644 86380
rect 41690 86368 41696 86420
rect 41748 86408 41754 86420
rect 41969 86411 42027 86417
rect 41969 86408 41981 86411
rect 41748 86380 41981 86408
rect 41748 86368 41754 86380
rect 41969 86377 41981 86380
rect 42015 86377 42027 86411
rect 47305 86411 47363 86417
rect 47305 86408 47317 86411
rect 41969 86371 42027 86377
rect 42812 86380 47317 86408
rect 41616 86312 42748 86340
rect 42720 86284 42748 86312
rect 42812 86284 42840 86380
rect 47305 86377 47317 86380
rect 47351 86408 47363 86411
rect 48958 86408 48964 86420
rect 47351 86380 48964 86408
rect 47351 86377 47363 86380
rect 47305 86371 47363 86377
rect 48958 86368 48964 86380
rect 49016 86408 49022 86420
rect 49513 86411 49571 86417
rect 49513 86408 49525 86411
rect 49016 86380 49525 86408
rect 49016 86368 49022 86380
rect 49513 86377 49525 86380
rect 49559 86408 49571 86411
rect 50341 86411 50399 86417
rect 50341 86408 50353 86411
rect 49559 86380 50353 86408
rect 49559 86377 49571 86380
rect 49513 86371 49571 86377
rect 50341 86377 50353 86380
rect 50387 86408 50399 86411
rect 50706 86408 50712 86420
rect 50387 86380 50712 86408
rect 50387 86377 50399 86380
rect 50341 86371 50399 86377
rect 50706 86368 50712 86380
rect 50764 86368 50770 86420
rect 50798 86368 50804 86420
rect 50856 86408 50862 86420
rect 52457 86411 52515 86417
rect 52457 86408 52469 86411
rect 50856 86380 52469 86408
rect 50856 86368 50862 86380
rect 52457 86377 52469 86380
rect 52503 86377 52515 86411
rect 52457 86371 52515 86377
rect 58342 86368 58348 86420
rect 58400 86408 58406 86420
rect 61197 86411 61255 86417
rect 61197 86408 61209 86411
rect 58400 86380 61209 86408
rect 58400 86368 58406 86380
rect 61197 86377 61209 86380
rect 61243 86377 61255 86411
rect 61197 86371 61255 86377
rect 44818 86300 44824 86352
rect 44876 86300 44882 86352
rect 47854 86300 47860 86352
rect 47912 86300 47918 86352
rect 40589 86275 40647 86281
rect 40589 86241 40601 86275
rect 40635 86241 40647 86275
rect 40589 86235 40647 86241
rect 40604 86204 40632 86235
rect 42702 86232 42708 86284
rect 42760 86232 42766 86284
rect 42794 86232 42800 86284
rect 42852 86232 42858 86284
rect 43441 86207 43499 86213
rect 43441 86204 43453 86207
rect 35176 86176 40540 86204
rect 40604 86176 43453 86204
rect 35069 86167 35127 86173
rect 35342 86145 35348 86148
rect 34057 86139 34115 86145
rect 34057 86136 34069 86139
rect 34020 86108 34069 86136
rect 34020 86096 34026 86108
rect 34057 86105 34069 86108
rect 34103 86105 34115 86139
rect 34057 86099 34115 86105
rect 34149 86139 34207 86145
rect 34149 86105 34161 86139
rect 34195 86105 34207 86139
rect 35336 86136 35348 86145
rect 35303 86108 35348 86136
rect 34149 86099 34207 86105
rect 35336 86099 35348 86108
rect 27672 86040 30328 86068
rect 27672 86028 27678 86040
rect 30374 86028 30380 86080
rect 30432 86028 30438 86080
rect 34164 86068 34192 86099
rect 35342 86096 35348 86099
rect 35400 86096 35406 86148
rect 35452 86108 36584 86136
rect 35452 86068 35480 86108
rect 34164 86040 35480 86068
rect 36446 86028 36452 86080
rect 36504 86028 36510 86080
rect 36556 86068 36584 86108
rect 37642 86096 37648 86148
rect 37700 86096 37706 86148
rect 37921 86139 37979 86145
rect 37921 86136 37933 86139
rect 37752 86108 37933 86136
rect 37752 86068 37780 86108
rect 37921 86105 37933 86108
rect 37967 86105 37979 86139
rect 37921 86099 37979 86105
rect 38838 86096 38844 86148
rect 38896 86096 38902 86148
rect 36556 86040 37780 86068
rect 37826 86028 37832 86080
rect 37884 86028 37890 86080
rect 40512 86068 40540 86176
rect 43441 86173 43453 86176
rect 43487 86204 43499 86207
rect 46569 86207 46627 86213
rect 46569 86204 46581 86207
rect 43487 86176 46581 86204
rect 43487 86173 43499 86176
rect 43441 86167 43499 86173
rect 46569 86173 46581 86176
rect 46615 86204 46627 86207
rect 49212 86207 49270 86213
rect 49212 86204 49224 86207
rect 46615 86176 49224 86204
rect 46615 86173 46627 86176
rect 46569 86167 46627 86173
rect 48884 86148 48912 86176
rect 49212 86173 49224 86176
rect 49258 86173 49270 86207
rect 49212 86167 49270 86173
rect 49528 86176 53512 86204
rect 40862 86145 40868 86148
rect 40856 86136 40868 86145
rect 40823 86108 40868 86136
rect 40856 86099 40868 86108
rect 40862 86096 40868 86099
rect 40920 86096 40926 86148
rect 43708 86139 43766 86145
rect 41386 86108 43392 86136
rect 41386 86068 41414 86108
rect 40512 86040 41414 86068
rect 42794 86028 42800 86080
rect 42852 86068 42858 86080
rect 42889 86071 42947 86077
rect 42889 86068 42901 86071
rect 42852 86040 42901 86068
rect 42852 86028 42858 86040
rect 42889 86037 42901 86040
rect 42935 86068 42947 86071
rect 43257 86071 43315 86077
rect 43257 86068 43269 86071
rect 42935 86040 43269 86068
rect 42935 86037 42947 86040
rect 42889 86031 42947 86037
rect 43257 86037 43269 86040
rect 43303 86037 43315 86071
rect 43364 86068 43392 86108
rect 43708 86105 43720 86139
rect 43754 86136 43766 86139
rect 44910 86136 44916 86148
rect 43754 86108 44916 86136
rect 43754 86105 43766 86108
rect 43708 86099 43766 86105
rect 44910 86096 44916 86108
rect 44968 86096 44974 86148
rect 45005 86139 45063 86145
rect 45005 86105 45017 86139
rect 45051 86105 45063 86139
rect 45005 86099 45063 86105
rect 45020 86068 45048 86099
rect 48866 86096 48872 86148
rect 48924 86096 48930 86148
rect 48958 86096 48964 86148
rect 49016 86145 49022 86148
rect 49016 86136 49028 86145
rect 49528 86136 49556 86176
rect 49016 86108 49061 86136
rect 49160 86108 49556 86136
rect 49804 86108 50016 86136
rect 49016 86099 49028 86108
rect 49016 86096 49022 86099
rect 49160 86068 49188 86108
rect 43364 86040 49188 86068
rect 43257 86031 43315 86037
rect 49234 86028 49240 86080
rect 49292 86068 49298 86080
rect 49804 86068 49832 86108
rect 49292 86040 49832 86068
rect 49292 86028 49298 86040
rect 49878 86028 49884 86080
rect 49936 86028 49942 86080
rect 49988 86068 50016 86108
rect 50706 86096 50712 86148
rect 50764 86136 50770 86148
rect 53377 86139 53435 86145
rect 53377 86136 53389 86139
rect 50764 86108 51672 86136
rect 50764 86096 50770 86108
rect 51644 86077 51672 86108
rect 53024 86108 53389 86136
rect 53024 86080 53052 86108
rect 53377 86105 53389 86108
rect 53423 86105 53435 86139
rect 53377 86099 53435 86105
rect 51169 86071 51227 86077
rect 51169 86068 51181 86071
rect 49988 86040 51181 86068
rect 51169 86037 51181 86040
rect 51215 86037 51227 86071
rect 51169 86031 51227 86037
rect 51629 86071 51687 86077
rect 51629 86037 51641 86071
rect 51675 86068 51687 86071
rect 51994 86068 52000 86080
rect 51675 86040 52000 86068
rect 51675 86037 51687 86040
rect 51629 86031 51687 86037
rect 51994 86028 52000 86040
rect 52052 86028 52058 86080
rect 53006 86028 53012 86080
rect 53064 86028 53070 86080
rect 53484 86068 53512 86176
rect 55306 86164 55312 86216
rect 55364 86204 55370 86216
rect 100938 86204 100944 86216
rect 55364 86176 100944 86204
rect 55364 86164 55370 86176
rect 100938 86164 100944 86176
rect 100996 86164 101002 86216
rect 108022 86164 108028 86216
rect 108080 86164 108086 86216
rect 53558 86096 53564 86148
rect 53616 86136 53622 86148
rect 55576 86139 55634 86145
rect 55576 86136 55588 86139
rect 53616 86108 55588 86136
rect 53616 86096 53622 86108
rect 55576 86105 55588 86108
rect 55622 86136 55634 86139
rect 74626 86136 74632 86148
rect 55622 86108 74632 86136
rect 55622 86105 55634 86108
rect 55576 86099 55634 86105
rect 74626 86096 74632 86108
rect 74684 86096 74690 86148
rect 54665 86071 54723 86077
rect 54665 86068 54677 86071
rect 53484 86040 54677 86068
rect 54665 86037 54677 86040
rect 54711 86037 54723 86071
rect 54665 86031 54723 86037
rect 56686 86028 56692 86080
rect 56744 86028 56750 86080
rect 1104 85978 108864 86000
rect 1104 85926 2950 85978
rect 3002 85926 3014 85978
rect 3066 85926 3078 85978
rect 3130 85926 3142 85978
rect 3194 85926 3206 85978
rect 3258 85926 4550 85978
rect 4602 85926 4614 85978
rect 4666 85926 4678 85978
rect 4730 85926 4742 85978
rect 4794 85926 4806 85978
rect 4858 85926 6150 85978
rect 6202 85926 6214 85978
rect 6266 85926 6278 85978
rect 6330 85926 6342 85978
rect 6394 85926 6406 85978
rect 6458 85926 7750 85978
rect 7802 85926 7814 85978
rect 7866 85926 7878 85978
rect 7930 85926 7942 85978
rect 7994 85926 8006 85978
rect 8058 85926 9350 85978
rect 9402 85926 9414 85978
rect 9466 85926 9478 85978
rect 9530 85926 9542 85978
rect 9594 85926 9606 85978
rect 9658 85926 10950 85978
rect 11002 85926 11014 85978
rect 11066 85926 11078 85978
rect 11130 85926 11142 85978
rect 11194 85926 11206 85978
rect 11258 85926 12550 85978
rect 12602 85926 12614 85978
rect 12666 85926 12678 85978
rect 12730 85926 12742 85978
rect 12794 85926 12806 85978
rect 12858 85926 14150 85978
rect 14202 85926 14214 85978
rect 14266 85926 14278 85978
rect 14330 85926 14342 85978
rect 14394 85926 14406 85978
rect 14458 85926 15750 85978
rect 15802 85926 15814 85978
rect 15866 85926 15878 85978
rect 15930 85926 15942 85978
rect 15994 85926 16006 85978
rect 16058 85926 17350 85978
rect 17402 85926 17414 85978
rect 17466 85926 17478 85978
rect 17530 85926 17542 85978
rect 17594 85926 17606 85978
rect 17658 85926 18950 85978
rect 19002 85926 19014 85978
rect 19066 85926 19078 85978
rect 19130 85926 19142 85978
rect 19194 85926 19206 85978
rect 19258 85926 20550 85978
rect 20602 85926 20614 85978
rect 20666 85926 20678 85978
rect 20730 85926 20742 85978
rect 20794 85926 20806 85978
rect 20858 85926 22150 85978
rect 22202 85926 22214 85978
rect 22266 85926 22278 85978
rect 22330 85926 22342 85978
rect 22394 85926 22406 85978
rect 22458 85926 23750 85978
rect 23802 85926 23814 85978
rect 23866 85926 23878 85978
rect 23930 85926 23942 85978
rect 23994 85926 24006 85978
rect 24058 85926 25350 85978
rect 25402 85926 25414 85978
rect 25466 85926 25478 85978
rect 25530 85926 25542 85978
rect 25594 85926 25606 85978
rect 25658 85926 26950 85978
rect 27002 85926 27014 85978
rect 27066 85926 27078 85978
rect 27130 85926 27142 85978
rect 27194 85926 27206 85978
rect 27258 85926 28550 85978
rect 28602 85926 28614 85978
rect 28666 85926 28678 85978
rect 28730 85926 28742 85978
rect 28794 85926 28806 85978
rect 28858 85926 30150 85978
rect 30202 85926 30214 85978
rect 30266 85926 30278 85978
rect 30330 85926 30342 85978
rect 30394 85926 30406 85978
rect 30458 85926 31750 85978
rect 31802 85926 31814 85978
rect 31866 85926 31878 85978
rect 31930 85926 31942 85978
rect 31994 85926 32006 85978
rect 32058 85926 33350 85978
rect 33402 85926 33414 85978
rect 33466 85926 33478 85978
rect 33530 85926 33542 85978
rect 33594 85926 33606 85978
rect 33658 85926 34950 85978
rect 35002 85926 35014 85978
rect 35066 85926 35078 85978
rect 35130 85926 35142 85978
rect 35194 85926 35206 85978
rect 35258 85926 36550 85978
rect 36602 85926 36614 85978
rect 36666 85926 36678 85978
rect 36730 85926 36742 85978
rect 36794 85926 36806 85978
rect 36858 85926 38150 85978
rect 38202 85926 38214 85978
rect 38266 85926 38278 85978
rect 38330 85926 38342 85978
rect 38394 85926 38406 85978
rect 38458 85926 39750 85978
rect 39802 85926 39814 85978
rect 39866 85926 39878 85978
rect 39930 85926 39942 85978
rect 39994 85926 40006 85978
rect 40058 85926 41350 85978
rect 41402 85926 41414 85978
rect 41466 85926 41478 85978
rect 41530 85926 41542 85978
rect 41594 85926 41606 85978
rect 41658 85926 42950 85978
rect 43002 85926 43014 85978
rect 43066 85926 43078 85978
rect 43130 85926 43142 85978
rect 43194 85926 43206 85978
rect 43258 85926 44550 85978
rect 44602 85926 44614 85978
rect 44666 85926 44678 85978
rect 44730 85926 44742 85978
rect 44794 85926 44806 85978
rect 44858 85926 46150 85978
rect 46202 85926 46214 85978
rect 46266 85926 46278 85978
rect 46330 85926 46342 85978
rect 46394 85926 46406 85978
rect 46458 85926 47750 85978
rect 47802 85926 47814 85978
rect 47866 85926 47878 85978
rect 47930 85926 47942 85978
rect 47994 85926 48006 85978
rect 48058 85926 49350 85978
rect 49402 85926 49414 85978
rect 49466 85926 49478 85978
rect 49530 85926 49542 85978
rect 49594 85926 49606 85978
rect 49658 85926 50950 85978
rect 51002 85926 51014 85978
rect 51066 85926 51078 85978
rect 51130 85926 51142 85978
rect 51194 85926 51206 85978
rect 51258 85926 52550 85978
rect 52602 85926 52614 85978
rect 52666 85926 52678 85978
rect 52730 85926 52742 85978
rect 52794 85926 52806 85978
rect 52858 85926 54150 85978
rect 54202 85926 54214 85978
rect 54266 85926 54278 85978
rect 54330 85926 54342 85978
rect 54394 85926 54406 85978
rect 54458 85926 55750 85978
rect 55802 85926 55814 85978
rect 55866 85926 55878 85978
rect 55930 85926 55942 85978
rect 55994 85926 56006 85978
rect 56058 85926 57350 85978
rect 57402 85926 57414 85978
rect 57466 85926 57478 85978
rect 57530 85926 57542 85978
rect 57594 85926 57606 85978
rect 57658 85926 58950 85978
rect 59002 85926 59014 85978
rect 59066 85926 59078 85978
rect 59130 85926 59142 85978
rect 59194 85926 59206 85978
rect 59258 85926 60550 85978
rect 60602 85926 60614 85978
rect 60666 85926 60678 85978
rect 60730 85926 60742 85978
rect 60794 85926 60806 85978
rect 60858 85926 62150 85978
rect 62202 85926 62214 85978
rect 62266 85926 62278 85978
rect 62330 85926 62342 85978
rect 62394 85926 62406 85978
rect 62458 85926 63750 85978
rect 63802 85926 63814 85978
rect 63866 85926 63878 85978
rect 63930 85926 63942 85978
rect 63994 85926 64006 85978
rect 64058 85926 65350 85978
rect 65402 85926 65414 85978
rect 65466 85926 65478 85978
rect 65530 85926 65542 85978
rect 65594 85926 65606 85978
rect 65658 85926 66950 85978
rect 67002 85926 67014 85978
rect 67066 85926 67078 85978
rect 67130 85926 67142 85978
rect 67194 85926 67206 85978
rect 67258 85926 68550 85978
rect 68602 85926 68614 85978
rect 68666 85926 68678 85978
rect 68730 85926 68742 85978
rect 68794 85926 68806 85978
rect 68858 85926 70150 85978
rect 70202 85926 70214 85978
rect 70266 85926 70278 85978
rect 70330 85926 70342 85978
rect 70394 85926 70406 85978
rect 70458 85926 71750 85978
rect 71802 85926 71814 85978
rect 71866 85926 71878 85978
rect 71930 85926 71942 85978
rect 71994 85926 72006 85978
rect 72058 85926 73350 85978
rect 73402 85926 73414 85978
rect 73466 85926 73478 85978
rect 73530 85926 73542 85978
rect 73594 85926 73606 85978
rect 73658 85926 74950 85978
rect 75002 85926 75014 85978
rect 75066 85926 75078 85978
rect 75130 85926 75142 85978
rect 75194 85926 75206 85978
rect 75258 85926 76550 85978
rect 76602 85926 76614 85978
rect 76666 85926 76678 85978
rect 76730 85926 76742 85978
rect 76794 85926 76806 85978
rect 76858 85926 78150 85978
rect 78202 85926 78214 85978
rect 78266 85926 78278 85978
rect 78330 85926 78342 85978
rect 78394 85926 78406 85978
rect 78458 85926 79750 85978
rect 79802 85926 79814 85978
rect 79866 85926 79878 85978
rect 79930 85926 79942 85978
rect 79994 85926 80006 85978
rect 80058 85926 81350 85978
rect 81402 85926 81414 85978
rect 81466 85926 81478 85978
rect 81530 85926 81542 85978
rect 81594 85926 81606 85978
rect 81658 85926 82950 85978
rect 83002 85926 83014 85978
rect 83066 85926 83078 85978
rect 83130 85926 83142 85978
rect 83194 85926 83206 85978
rect 83258 85926 84550 85978
rect 84602 85926 84614 85978
rect 84666 85926 84678 85978
rect 84730 85926 84742 85978
rect 84794 85926 84806 85978
rect 84858 85926 86150 85978
rect 86202 85926 86214 85978
rect 86266 85926 86278 85978
rect 86330 85926 86342 85978
rect 86394 85926 86406 85978
rect 86458 85926 87750 85978
rect 87802 85926 87814 85978
rect 87866 85926 87878 85978
rect 87930 85926 87942 85978
rect 87994 85926 88006 85978
rect 88058 85926 89350 85978
rect 89402 85926 89414 85978
rect 89466 85926 89478 85978
rect 89530 85926 89542 85978
rect 89594 85926 89606 85978
rect 89658 85926 90950 85978
rect 91002 85926 91014 85978
rect 91066 85926 91078 85978
rect 91130 85926 91142 85978
rect 91194 85926 91206 85978
rect 91258 85926 92550 85978
rect 92602 85926 92614 85978
rect 92666 85926 92678 85978
rect 92730 85926 92742 85978
rect 92794 85926 92806 85978
rect 92858 85926 94150 85978
rect 94202 85926 94214 85978
rect 94266 85926 94278 85978
rect 94330 85926 94342 85978
rect 94394 85926 94406 85978
rect 94458 85926 95750 85978
rect 95802 85926 95814 85978
rect 95866 85926 95878 85978
rect 95930 85926 95942 85978
rect 95994 85926 96006 85978
rect 96058 85926 97350 85978
rect 97402 85926 97414 85978
rect 97466 85926 97478 85978
rect 97530 85926 97542 85978
rect 97594 85926 97606 85978
rect 97658 85926 98950 85978
rect 99002 85926 99014 85978
rect 99066 85926 99078 85978
rect 99130 85926 99142 85978
rect 99194 85926 99206 85978
rect 99258 85926 100550 85978
rect 100602 85926 100614 85978
rect 100666 85926 100678 85978
rect 100730 85926 100742 85978
rect 100794 85926 100806 85978
rect 100858 85926 102150 85978
rect 102202 85926 102214 85978
rect 102266 85926 102278 85978
rect 102330 85926 102342 85978
rect 102394 85926 102406 85978
rect 102458 85926 103750 85978
rect 103802 85926 103814 85978
rect 103866 85926 103878 85978
rect 103930 85926 103942 85978
rect 103994 85926 104006 85978
rect 104058 85926 105350 85978
rect 105402 85926 105414 85978
rect 105466 85926 105478 85978
rect 105530 85926 105542 85978
rect 105594 85926 105606 85978
rect 105658 85926 106950 85978
rect 107002 85926 107014 85978
rect 107066 85926 107078 85978
rect 107130 85926 107142 85978
rect 107194 85926 107206 85978
rect 107258 85926 108550 85978
rect 108602 85926 108614 85978
rect 108666 85926 108678 85978
rect 108730 85926 108742 85978
rect 108794 85926 108806 85978
rect 108858 85926 108864 85978
rect 1104 85904 108864 85926
rect 4430 85824 4436 85876
rect 4488 85864 4494 85876
rect 25038 85864 25044 85876
rect 4488 85836 25044 85864
rect 4488 85824 4494 85836
rect 25038 85824 25044 85836
rect 25096 85864 25102 85876
rect 27614 85864 27620 85876
rect 25096 85836 27620 85864
rect 25096 85824 25102 85836
rect 27614 85824 27620 85836
rect 27672 85824 27678 85876
rect 30006 85824 30012 85876
rect 30064 85864 30070 85876
rect 33870 85864 33876 85876
rect 30064 85836 33876 85864
rect 30064 85824 30070 85836
rect 33870 85824 33876 85836
rect 33928 85864 33934 85876
rect 36078 85864 36084 85876
rect 33928 85836 36084 85864
rect 33928 85824 33934 85836
rect 36078 85824 36084 85836
rect 36136 85824 36142 85876
rect 40402 85824 40408 85876
rect 40460 85864 40466 85876
rect 42794 85864 42800 85876
rect 40460 85836 42800 85864
rect 40460 85824 40466 85836
rect 42794 85824 42800 85836
rect 42852 85824 42858 85876
rect 75914 85864 75920 85876
rect 43088 85836 75920 85864
rect 9214 85756 9220 85808
rect 9272 85796 9278 85808
rect 19794 85796 19800 85808
rect 9272 85768 19800 85796
rect 9272 85756 9278 85768
rect 19794 85756 19800 85768
rect 19852 85796 19858 85808
rect 37642 85796 37648 85808
rect 19852 85768 37648 85796
rect 19852 85756 19858 85768
rect 37642 85756 37648 85768
rect 37700 85756 37706 85808
rect 40862 85796 40868 85808
rect 37752 85768 40868 85796
rect 8938 85688 8944 85740
rect 8996 85728 9002 85740
rect 19978 85728 19984 85740
rect 8996 85700 19984 85728
rect 8996 85688 9002 85700
rect 19978 85688 19984 85700
rect 20036 85688 20042 85740
rect 24946 85688 24952 85740
rect 25004 85728 25010 85740
rect 36446 85728 36452 85740
rect 25004 85700 36452 85728
rect 25004 85688 25010 85700
rect 36446 85688 36452 85700
rect 36504 85688 36510 85740
rect 13722 85620 13728 85672
rect 13780 85660 13786 85672
rect 19702 85660 19708 85672
rect 13780 85632 19708 85660
rect 13780 85620 13786 85632
rect 19702 85620 19708 85632
rect 19760 85660 19766 85672
rect 19760 85632 26924 85660
rect 19760 85620 19766 85632
rect 9122 85552 9128 85604
rect 9180 85592 9186 85604
rect 26786 85592 26792 85604
rect 9180 85564 26792 85592
rect 9180 85552 9186 85564
rect 26786 85552 26792 85564
rect 26844 85552 26850 85604
rect 26896 85592 26924 85632
rect 26970 85620 26976 85672
rect 27028 85660 27034 85672
rect 37752 85660 37780 85768
rect 40862 85756 40868 85768
rect 40920 85796 40926 85808
rect 43088 85796 43116 85836
rect 75914 85824 75920 85836
rect 75972 85824 75978 85876
rect 40920 85768 43116 85796
rect 40920 85756 40926 85768
rect 46566 85756 46572 85808
rect 46624 85796 46630 85808
rect 49878 85796 49884 85808
rect 46624 85768 49884 85796
rect 46624 85756 46630 85768
rect 49878 85756 49884 85768
rect 49936 85756 49942 85808
rect 56686 85796 56692 85808
rect 51046 85768 56692 85796
rect 37826 85688 37832 85740
rect 37884 85728 37890 85740
rect 51046 85728 51074 85768
rect 56686 85756 56692 85768
rect 56744 85756 56750 85808
rect 37884 85700 51074 85728
rect 37884 85688 37890 85700
rect 51994 85688 52000 85740
rect 52052 85728 52058 85740
rect 73154 85728 73160 85740
rect 52052 85700 73160 85728
rect 52052 85688 52058 85700
rect 73154 85688 73160 85700
rect 73212 85688 73218 85740
rect 40770 85660 40776 85672
rect 27028 85632 37780 85660
rect 37844 85632 40776 85660
rect 27028 85620 27034 85632
rect 37844 85592 37872 85632
rect 40770 85620 40776 85632
rect 40828 85620 40834 85672
rect 42702 85620 42708 85672
rect 42760 85660 42766 85672
rect 55214 85660 55220 85672
rect 42760 85632 55220 85660
rect 42760 85620 42766 85632
rect 55214 85620 55220 85632
rect 55272 85620 55278 85672
rect 26896 85564 37872 85592
rect 38838 85552 38844 85604
rect 38896 85592 38902 85604
rect 42794 85592 42800 85604
rect 38896 85564 42800 85592
rect 38896 85552 38902 85564
rect 42794 85552 42800 85564
rect 42852 85552 42858 85604
rect 46934 85552 46940 85604
rect 46992 85592 46998 85604
rect 55674 85592 55680 85604
rect 46992 85564 55680 85592
rect 46992 85552 46998 85564
rect 55674 85552 55680 85564
rect 55732 85552 55738 85604
rect 1026 85484 1032 85536
rect 1084 85524 1090 85536
rect 40034 85524 40040 85536
rect 1084 85496 40040 85524
rect 1084 85484 1090 85496
rect 40034 85484 40040 85496
rect 40092 85484 40098 85536
rect 1104 85434 9936 85456
rect 1104 85382 3610 85434
rect 3662 85382 3674 85434
rect 3726 85382 3738 85434
rect 3790 85382 3802 85434
rect 3854 85382 3866 85434
rect 3918 85382 5210 85434
rect 5262 85382 5274 85434
rect 5326 85382 5338 85434
rect 5390 85382 5402 85434
rect 5454 85382 5466 85434
rect 5518 85382 6810 85434
rect 6862 85382 6874 85434
rect 6926 85382 6938 85434
rect 6990 85382 7002 85434
rect 7054 85382 7066 85434
rect 7118 85382 8410 85434
rect 8462 85382 8474 85434
rect 8526 85382 8538 85434
rect 8590 85382 8602 85434
rect 8654 85382 8666 85434
rect 8718 85382 9936 85434
rect 10318 85416 10324 85468
rect 10376 85456 10382 85468
rect 46566 85456 46572 85468
rect 10376 85428 46572 85456
rect 10376 85416 10382 85428
rect 46566 85416 46572 85428
rect 46624 85416 46630 85468
rect 1104 85360 9936 85382
rect 11698 85348 11704 85400
rect 11756 85388 11762 85400
rect 49234 85388 49240 85400
rect 11756 85360 49240 85388
rect 11756 85348 11762 85360
rect 49234 85348 49240 85360
rect 49292 85348 49298 85400
rect 10134 85280 10140 85332
rect 10192 85320 10198 85332
rect 52454 85320 52460 85332
rect 10192 85292 52460 85320
rect 10192 85280 10198 85292
rect 52454 85280 52460 85292
rect 52512 85280 52518 85332
rect 8202 85212 8208 85264
rect 8260 85252 8266 85264
rect 53834 85252 53840 85264
rect 8260 85224 53840 85252
rect 8260 85212 8266 85224
rect 53834 85212 53840 85224
rect 53892 85212 53898 85264
rect 8110 85144 8116 85196
rect 8168 85184 8174 85196
rect 51166 85184 51172 85196
rect 8168 85156 51172 85184
rect 8168 85144 8174 85156
rect 51166 85144 51172 85156
rect 51224 85144 51230 85196
rect 7466 85076 7472 85128
rect 7524 85116 7530 85128
rect 66254 85116 66260 85128
rect 7524 85088 66260 85116
rect 7524 85076 7530 85088
rect 66254 85076 66260 85088
rect 66312 85076 66318 85128
rect 7190 85008 7196 85060
rect 7248 85048 7254 85060
rect 71222 85048 71228 85060
rect 7248 85020 71228 85048
rect 7248 85008 7254 85020
rect 71222 85008 71228 85020
rect 71280 85008 71286 85060
rect 6546 84940 6552 84992
rect 6604 84980 6610 84992
rect 34790 84980 34796 84992
rect 6604 84952 34796 84980
rect 6604 84940 6610 84952
rect 34790 84940 34796 84952
rect 34848 84940 34854 84992
rect 1104 84890 9936 84912
rect 1104 84838 2950 84890
rect 3002 84838 3014 84890
rect 3066 84838 3078 84890
rect 3130 84838 3142 84890
rect 3194 84838 3206 84890
rect 3258 84838 4550 84890
rect 4602 84838 4614 84890
rect 4666 84838 4678 84890
rect 4730 84838 4742 84890
rect 4794 84838 4806 84890
rect 4858 84838 6150 84890
rect 6202 84838 6214 84890
rect 6266 84838 6278 84890
rect 6330 84838 6342 84890
rect 6394 84838 6406 84890
rect 6458 84838 7750 84890
rect 7802 84838 7814 84890
rect 7866 84838 7878 84890
rect 7930 84838 7942 84890
rect 7994 84838 8006 84890
rect 8058 84838 9350 84890
rect 9402 84838 9414 84890
rect 9466 84838 9478 84890
rect 9530 84838 9542 84890
rect 9594 84838 9606 84890
rect 9658 84838 9936 84890
rect 10870 84872 10876 84924
rect 10928 84912 10934 84924
rect 57606 84912 57612 84924
rect 10928 84884 57612 84912
rect 10928 84872 10934 84884
rect 57606 84872 57612 84884
rect 57664 84872 57670 84924
rect 1104 84816 9936 84838
rect 10686 84804 10692 84856
rect 10744 84844 10750 84856
rect 78674 84844 78680 84856
rect 10744 84816 78680 84844
rect 10744 84804 10750 84816
rect 78674 84804 78680 84816
rect 78732 84804 78738 84856
rect 11790 84736 11796 84788
rect 11848 84776 11854 84788
rect 44726 84776 44732 84788
rect 11848 84748 44732 84776
rect 11848 84736 11854 84748
rect 44726 84736 44732 84748
rect 44784 84736 44790 84788
rect 11882 84668 11888 84720
rect 11940 84708 11946 84720
rect 42518 84708 42524 84720
rect 11940 84680 42524 84708
rect 11940 84668 11946 84680
rect 42518 84668 42524 84680
rect 42576 84668 42582 84720
rect 934 84600 940 84652
rect 992 84640 998 84652
rect 1489 84643 1547 84649
rect 1489 84640 1501 84643
rect 992 84612 1501 84640
rect 992 84600 998 84612
rect 1489 84609 1501 84612
rect 1535 84609 1547 84643
rect 1489 84603 1547 84609
rect 4154 84600 4160 84652
rect 4212 84640 4218 84652
rect 27338 84640 27344 84652
rect 4212 84612 27344 84640
rect 4212 84600 4218 84612
rect 27338 84600 27344 84612
rect 27396 84600 27402 84652
rect 1670 84464 1676 84516
rect 1728 84464 1734 84516
rect 1104 84346 9936 84368
rect 1104 84294 3610 84346
rect 3662 84294 3674 84346
rect 3726 84294 3738 84346
rect 3790 84294 3802 84346
rect 3854 84294 3866 84346
rect 3918 84294 5210 84346
rect 5262 84294 5274 84346
rect 5326 84294 5338 84346
rect 5390 84294 5402 84346
rect 5454 84294 5466 84346
rect 5518 84294 6810 84346
rect 6862 84294 6874 84346
rect 6926 84294 6938 84346
rect 6990 84294 7002 84346
rect 7054 84294 7066 84346
rect 7118 84294 8410 84346
rect 8462 84294 8474 84346
rect 8526 84294 8538 84346
rect 8590 84294 8602 84346
rect 8654 84294 8666 84346
rect 8718 84294 9936 84346
rect 1104 84272 9936 84294
rect 6638 83852 6644 83904
rect 6696 83892 6702 83904
rect 37366 83892 37372 83904
rect 6696 83864 37372 83892
rect 6696 83852 6702 83864
rect 37366 83852 37372 83864
rect 37424 83852 37430 83904
rect 1104 83802 9936 83824
rect 1104 83750 2950 83802
rect 3002 83750 3014 83802
rect 3066 83750 3078 83802
rect 3130 83750 3142 83802
rect 3194 83750 3206 83802
rect 3258 83750 4550 83802
rect 4602 83750 4614 83802
rect 4666 83750 4678 83802
rect 4730 83750 4742 83802
rect 4794 83750 4806 83802
rect 4858 83750 6150 83802
rect 6202 83750 6214 83802
rect 6266 83750 6278 83802
rect 6330 83750 6342 83802
rect 6394 83750 6406 83802
rect 6458 83750 7750 83802
rect 7802 83750 7814 83802
rect 7866 83750 7878 83802
rect 7930 83750 7942 83802
rect 7994 83750 8006 83802
rect 8058 83750 9350 83802
rect 9402 83750 9414 83802
rect 9466 83750 9478 83802
rect 9530 83750 9542 83802
rect 9594 83750 9606 83802
rect 9658 83750 9936 83802
rect 1104 83728 9936 83750
rect 7374 83648 7380 83700
rect 7432 83688 7438 83700
rect 45094 83688 45100 83700
rect 7432 83660 45100 83688
rect 7432 83648 7438 83660
rect 45094 83648 45100 83660
rect 45152 83648 45158 83700
rect 8294 83580 8300 83632
rect 8352 83620 8358 83632
rect 46934 83620 46940 83632
rect 8352 83592 46940 83620
rect 8352 83580 8358 83592
rect 46934 83580 46940 83592
rect 46992 83580 46998 83632
rect 934 83512 940 83564
rect 992 83552 998 83564
rect 1489 83555 1547 83561
rect 1489 83552 1501 83555
rect 992 83524 1501 83552
rect 992 83512 998 83524
rect 1489 83521 1501 83524
rect 1535 83521 1547 83555
rect 1489 83515 1547 83521
rect 10962 83512 10968 83564
rect 11020 83552 11026 83564
rect 59906 83552 59912 83564
rect 11020 83524 59912 83552
rect 11020 83512 11026 83524
rect 59906 83512 59912 83524
rect 59964 83512 59970 83564
rect 10226 83444 10232 83496
rect 10284 83484 10290 83496
rect 70210 83484 70216 83496
rect 10284 83456 70216 83484
rect 10284 83444 10290 83456
rect 70210 83444 70216 83456
rect 70268 83444 70274 83496
rect 1673 83419 1731 83425
rect 1673 83385 1685 83419
rect 1719 83416 1731 83419
rect 3970 83416 3976 83428
rect 1719 83388 3976 83416
rect 1719 83385 1731 83388
rect 1673 83379 1731 83385
rect 3970 83376 3976 83388
rect 4028 83376 4034 83428
rect 1104 83258 9936 83280
rect 1104 83206 3610 83258
rect 3662 83206 3674 83258
rect 3726 83206 3738 83258
rect 3790 83206 3802 83258
rect 3854 83206 3866 83258
rect 3918 83206 5210 83258
rect 5262 83206 5274 83258
rect 5326 83206 5338 83258
rect 5390 83206 5402 83258
rect 5454 83206 5466 83258
rect 5518 83206 6810 83258
rect 6862 83206 6874 83258
rect 6926 83206 6938 83258
rect 6990 83206 7002 83258
rect 7054 83206 7066 83258
rect 7118 83206 8410 83258
rect 8462 83206 8474 83258
rect 8526 83206 8538 83258
rect 8590 83206 8602 83258
rect 8654 83206 8666 83258
rect 8718 83206 9936 83258
rect 1104 83184 9936 83206
rect 1486 82832 1492 82884
rect 1544 82832 1550 82884
rect 1673 82875 1731 82881
rect 1673 82841 1685 82875
rect 1719 82872 1731 82875
rect 2222 82872 2228 82884
rect 1719 82844 2228 82872
rect 1719 82841 1731 82844
rect 1673 82835 1731 82841
rect 2222 82832 2228 82844
rect 2280 82832 2286 82884
rect 1104 82714 9936 82736
rect 1104 82662 2950 82714
rect 3002 82662 3014 82714
rect 3066 82662 3078 82714
rect 3130 82662 3142 82714
rect 3194 82662 3206 82714
rect 3258 82662 4550 82714
rect 4602 82662 4614 82714
rect 4666 82662 4678 82714
rect 4730 82662 4742 82714
rect 4794 82662 4806 82714
rect 4858 82662 6150 82714
rect 6202 82662 6214 82714
rect 6266 82662 6278 82714
rect 6330 82662 6342 82714
rect 6394 82662 6406 82714
rect 6458 82662 7750 82714
rect 7802 82662 7814 82714
rect 7866 82662 7878 82714
rect 7930 82662 7942 82714
rect 7994 82662 8006 82714
rect 8058 82662 9350 82714
rect 9402 82662 9414 82714
rect 9466 82662 9478 82714
rect 9530 82662 9542 82714
rect 9594 82662 9606 82714
rect 9658 82662 9936 82714
rect 1104 82640 9936 82662
rect 1104 82170 9936 82192
rect 1104 82118 3610 82170
rect 3662 82118 3674 82170
rect 3726 82118 3738 82170
rect 3790 82118 3802 82170
rect 3854 82118 3866 82170
rect 3918 82118 5210 82170
rect 5262 82118 5274 82170
rect 5326 82118 5338 82170
rect 5390 82118 5402 82170
rect 5454 82118 5466 82170
rect 5518 82118 6810 82170
rect 6862 82118 6874 82170
rect 6926 82118 6938 82170
rect 6990 82118 7002 82170
rect 7054 82118 7066 82170
rect 7118 82118 8410 82170
rect 8462 82118 8474 82170
rect 8526 82118 8538 82170
rect 8590 82118 8602 82170
rect 8654 82118 8666 82170
rect 8718 82118 9936 82170
rect 1104 82096 9936 82118
rect 934 81744 940 81796
rect 992 81784 998 81796
rect 1489 81787 1547 81793
rect 1489 81784 1501 81787
rect 992 81756 1501 81784
rect 992 81744 998 81756
rect 1489 81753 1501 81756
rect 1535 81753 1547 81787
rect 1489 81747 1547 81753
rect 1673 81787 1731 81793
rect 1673 81753 1685 81787
rect 1719 81784 1731 81787
rect 1762 81784 1768 81796
rect 1719 81756 1768 81784
rect 1719 81753 1731 81756
rect 1673 81747 1731 81753
rect 1762 81744 1768 81756
rect 1820 81744 1826 81796
rect 1104 81626 9936 81648
rect 1104 81574 2950 81626
rect 3002 81574 3014 81626
rect 3066 81574 3078 81626
rect 3130 81574 3142 81626
rect 3194 81574 3206 81626
rect 3258 81574 4550 81626
rect 4602 81574 4614 81626
rect 4666 81574 4678 81626
rect 4730 81574 4742 81626
rect 4794 81574 4806 81626
rect 4858 81574 6150 81626
rect 6202 81574 6214 81626
rect 6266 81574 6278 81626
rect 6330 81574 6342 81626
rect 6394 81574 6406 81626
rect 6458 81574 7750 81626
rect 7802 81574 7814 81626
rect 7866 81574 7878 81626
rect 7930 81574 7942 81626
rect 7994 81574 8006 81626
rect 8058 81574 9350 81626
rect 9402 81574 9414 81626
rect 9466 81574 9478 81626
rect 9530 81574 9542 81626
rect 9594 81574 9606 81626
rect 9658 81574 9936 81626
rect 1104 81552 9936 81574
rect 1104 81082 9936 81104
rect 1104 81030 3610 81082
rect 3662 81030 3674 81082
rect 3726 81030 3738 81082
rect 3790 81030 3802 81082
rect 3854 81030 3866 81082
rect 3918 81030 5210 81082
rect 5262 81030 5274 81082
rect 5326 81030 5338 81082
rect 5390 81030 5402 81082
rect 5454 81030 5466 81082
rect 5518 81030 6810 81082
rect 6862 81030 6874 81082
rect 6926 81030 6938 81082
rect 6990 81030 7002 81082
rect 7054 81030 7066 81082
rect 7118 81030 8410 81082
rect 8462 81030 8474 81082
rect 8526 81030 8538 81082
rect 8590 81030 8602 81082
rect 8654 81030 8666 81082
rect 8718 81030 9936 81082
rect 1104 81008 9936 81030
rect 934 80656 940 80708
rect 992 80696 998 80708
rect 1489 80699 1547 80705
rect 1489 80696 1501 80699
rect 992 80668 1501 80696
rect 992 80656 998 80668
rect 1489 80665 1501 80668
rect 1535 80665 1547 80699
rect 1489 80659 1547 80665
rect 1673 80699 1731 80705
rect 1673 80665 1685 80699
rect 1719 80696 1731 80699
rect 1854 80696 1860 80708
rect 1719 80668 1860 80696
rect 1719 80665 1731 80668
rect 1673 80659 1731 80665
rect 1854 80656 1860 80668
rect 1912 80656 1918 80708
rect 1104 80538 9936 80560
rect 1104 80486 2950 80538
rect 3002 80486 3014 80538
rect 3066 80486 3078 80538
rect 3130 80486 3142 80538
rect 3194 80486 3206 80538
rect 3258 80486 4550 80538
rect 4602 80486 4614 80538
rect 4666 80486 4678 80538
rect 4730 80486 4742 80538
rect 4794 80486 4806 80538
rect 4858 80486 6150 80538
rect 6202 80486 6214 80538
rect 6266 80486 6278 80538
rect 6330 80486 6342 80538
rect 6394 80486 6406 80538
rect 6458 80486 7750 80538
rect 7802 80486 7814 80538
rect 7866 80486 7878 80538
rect 7930 80486 7942 80538
rect 7994 80486 8006 80538
rect 8058 80486 9350 80538
rect 9402 80486 9414 80538
rect 9466 80486 9478 80538
rect 9530 80486 9542 80538
rect 9594 80486 9606 80538
rect 9658 80486 9936 80538
rect 1104 80464 9936 80486
rect 1104 79994 9936 80016
rect 1104 79942 3610 79994
rect 3662 79942 3674 79994
rect 3726 79942 3738 79994
rect 3790 79942 3802 79994
rect 3854 79942 3866 79994
rect 3918 79942 5210 79994
rect 5262 79942 5274 79994
rect 5326 79942 5338 79994
rect 5390 79942 5402 79994
rect 5454 79942 5466 79994
rect 5518 79942 6810 79994
rect 6862 79942 6874 79994
rect 6926 79942 6938 79994
rect 6990 79942 7002 79994
rect 7054 79942 7066 79994
rect 7118 79942 8410 79994
rect 8462 79942 8474 79994
rect 8526 79942 8538 79994
rect 8590 79942 8602 79994
rect 8654 79942 8666 79994
rect 8718 79942 9936 79994
rect 1104 79920 9936 79942
rect 934 79568 940 79620
rect 992 79608 998 79620
rect 1489 79611 1547 79617
rect 1489 79608 1501 79611
rect 992 79580 1501 79608
rect 992 79568 998 79580
rect 1489 79577 1501 79580
rect 1535 79577 1547 79611
rect 1489 79571 1547 79577
rect 1673 79611 1731 79617
rect 1673 79577 1685 79611
rect 1719 79608 1731 79611
rect 2038 79608 2044 79620
rect 1719 79580 2044 79608
rect 1719 79577 1731 79580
rect 1673 79571 1731 79577
rect 2038 79568 2044 79580
rect 2096 79568 2102 79620
rect 4154 79500 4160 79552
rect 4212 79540 4218 79552
rect 4982 79540 4988 79552
rect 4212 79512 4988 79540
rect 4212 79500 4218 79512
rect 4982 79500 4988 79512
rect 5040 79500 5046 79552
rect 1104 79450 9936 79472
rect 1104 79398 2950 79450
rect 3002 79398 3014 79450
rect 3066 79398 3078 79450
rect 3130 79398 3142 79450
rect 3194 79398 3206 79450
rect 3258 79398 4550 79450
rect 4602 79398 4614 79450
rect 4666 79398 4678 79450
rect 4730 79398 4742 79450
rect 4794 79398 4806 79450
rect 4858 79398 6150 79450
rect 6202 79398 6214 79450
rect 6266 79398 6278 79450
rect 6330 79398 6342 79450
rect 6394 79398 6406 79450
rect 6458 79398 7750 79450
rect 7802 79398 7814 79450
rect 7866 79398 7878 79450
rect 7930 79398 7942 79450
rect 7994 79398 8006 79450
rect 8058 79398 9350 79450
rect 9402 79398 9414 79450
rect 9466 79398 9478 79450
rect 9530 79398 9542 79450
rect 9594 79398 9606 79450
rect 9658 79398 9936 79450
rect 1104 79376 9936 79398
rect 934 79160 940 79212
rect 992 79200 998 79212
rect 1397 79203 1455 79209
rect 1397 79200 1409 79203
rect 992 79172 1409 79200
rect 992 79160 998 79172
rect 1397 79169 1409 79172
rect 1443 79169 1455 79203
rect 1397 79163 1455 79169
rect 1210 78956 1216 79008
rect 1268 78996 1274 79008
rect 1581 78999 1639 79005
rect 1581 78996 1593 78999
rect 1268 78968 1593 78996
rect 1268 78956 1274 78968
rect 1581 78965 1593 78968
rect 1627 78965 1639 78999
rect 1581 78959 1639 78965
rect 1104 78906 9936 78928
rect 1104 78854 3610 78906
rect 3662 78854 3674 78906
rect 3726 78854 3738 78906
rect 3790 78854 3802 78906
rect 3854 78854 3866 78906
rect 3918 78854 5210 78906
rect 5262 78854 5274 78906
rect 5326 78854 5338 78906
rect 5390 78854 5402 78906
rect 5454 78854 5466 78906
rect 5518 78854 6810 78906
rect 6862 78854 6874 78906
rect 6926 78854 6938 78906
rect 6990 78854 7002 78906
rect 7054 78854 7066 78906
rect 7118 78854 8410 78906
rect 8462 78854 8474 78906
rect 8526 78854 8538 78906
rect 8590 78854 8602 78906
rect 8654 78854 8666 78906
rect 8718 78854 9936 78906
rect 1104 78832 9936 78854
rect 1104 78362 9936 78384
rect 1104 78310 2950 78362
rect 3002 78310 3014 78362
rect 3066 78310 3078 78362
rect 3130 78310 3142 78362
rect 3194 78310 3206 78362
rect 3258 78310 4550 78362
rect 4602 78310 4614 78362
rect 4666 78310 4678 78362
rect 4730 78310 4742 78362
rect 4794 78310 4806 78362
rect 4858 78310 6150 78362
rect 6202 78310 6214 78362
rect 6266 78310 6278 78362
rect 6330 78310 6342 78362
rect 6394 78310 6406 78362
rect 6458 78310 7750 78362
rect 7802 78310 7814 78362
rect 7866 78310 7878 78362
rect 7930 78310 7942 78362
rect 7994 78310 8006 78362
rect 8058 78310 9350 78362
rect 9402 78310 9414 78362
rect 9466 78310 9478 78362
rect 9530 78310 9542 78362
rect 9594 78310 9606 78362
rect 9658 78310 9936 78362
rect 1104 78288 9936 78310
rect 934 78072 940 78124
rect 992 78112 998 78124
rect 1397 78115 1455 78121
rect 1397 78112 1409 78115
rect 992 78084 1409 78112
rect 992 78072 998 78084
rect 1397 78081 1409 78084
rect 1443 78081 1455 78115
rect 1397 78075 1455 78081
rect 1581 77911 1639 77917
rect 1581 77877 1593 77911
rect 1627 77908 1639 77911
rect 3326 77908 3332 77920
rect 1627 77880 3332 77908
rect 1627 77877 1639 77880
rect 1581 77871 1639 77877
rect 3326 77868 3332 77880
rect 3384 77868 3390 77920
rect 1104 77818 9936 77840
rect 1104 77766 3610 77818
rect 3662 77766 3674 77818
rect 3726 77766 3738 77818
rect 3790 77766 3802 77818
rect 3854 77766 3866 77818
rect 3918 77766 5210 77818
rect 5262 77766 5274 77818
rect 5326 77766 5338 77818
rect 5390 77766 5402 77818
rect 5454 77766 5466 77818
rect 5518 77766 6810 77818
rect 6862 77766 6874 77818
rect 6926 77766 6938 77818
rect 6990 77766 7002 77818
rect 7054 77766 7066 77818
rect 7118 77766 8410 77818
rect 8462 77766 8474 77818
rect 8526 77766 8538 77818
rect 8590 77766 8602 77818
rect 8654 77766 8666 77818
rect 8718 77766 9936 77818
rect 1104 77744 9936 77766
rect 1104 77274 9936 77296
rect 1104 77222 2950 77274
rect 3002 77222 3014 77274
rect 3066 77222 3078 77274
rect 3130 77222 3142 77274
rect 3194 77222 3206 77274
rect 3258 77222 4550 77274
rect 4602 77222 4614 77274
rect 4666 77222 4678 77274
rect 4730 77222 4742 77274
rect 4794 77222 4806 77274
rect 4858 77222 6150 77274
rect 6202 77222 6214 77274
rect 6266 77222 6278 77274
rect 6330 77222 6342 77274
rect 6394 77222 6406 77274
rect 6458 77222 7750 77274
rect 7802 77222 7814 77274
rect 7866 77222 7878 77274
rect 7930 77222 7942 77274
rect 7994 77222 8006 77274
rect 8058 77222 9350 77274
rect 9402 77222 9414 77274
rect 9466 77222 9478 77274
rect 9530 77222 9542 77274
rect 9594 77222 9606 77274
rect 9658 77222 9936 77274
rect 1104 77200 9936 77222
rect 9030 77120 9036 77172
rect 9088 77160 9094 77172
rect 9309 77163 9367 77169
rect 9309 77160 9321 77163
rect 9088 77132 9321 77160
rect 9088 77120 9094 77132
rect 9309 77129 9321 77132
rect 9355 77129 9367 77163
rect 9309 77123 9367 77129
rect 934 76984 940 77036
rect 992 77024 998 77036
rect 1489 77027 1547 77033
rect 1489 77024 1501 77027
rect 992 76996 1501 77024
rect 992 76984 998 76996
rect 1489 76993 1501 76996
rect 1535 76993 1547 77027
rect 1489 76987 1547 76993
rect 7650 76984 7656 77036
rect 7708 77024 7714 77036
rect 9217 77027 9275 77033
rect 9217 77024 9229 77027
rect 7708 76996 9229 77024
rect 7708 76984 7714 76996
rect 9217 76993 9229 76996
rect 9263 77024 9275 77027
rect 10134 77024 10140 77036
rect 9263 76996 10140 77024
rect 9263 76993 9275 76996
rect 9217 76987 9275 76993
rect 10134 76984 10140 76996
rect 10192 76984 10198 77036
rect 8938 76916 8944 76968
rect 8996 76956 9002 76968
rect 9401 76959 9459 76965
rect 9401 76956 9413 76959
rect 8996 76928 9413 76956
rect 8996 76916 9002 76928
rect 9401 76925 9413 76928
rect 9447 76925 9459 76959
rect 9401 76919 9459 76925
rect 1673 76891 1731 76897
rect 1673 76857 1685 76891
rect 1719 76888 1731 76891
rect 2590 76888 2596 76900
rect 1719 76860 2596 76888
rect 1719 76857 1731 76860
rect 1673 76851 1731 76857
rect 2590 76848 2596 76860
rect 2648 76848 2654 76900
rect 2498 76780 2504 76832
rect 2556 76820 2562 76832
rect 8849 76823 8907 76829
rect 8849 76820 8861 76823
rect 2556 76792 8861 76820
rect 2556 76780 2562 76792
rect 8849 76789 8861 76792
rect 8895 76789 8907 76823
rect 8849 76783 8907 76789
rect 1104 76730 9936 76752
rect 1104 76678 3610 76730
rect 3662 76678 3674 76730
rect 3726 76678 3738 76730
rect 3790 76678 3802 76730
rect 3854 76678 3866 76730
rect 3918 76678 5210 76730
rect 5262 76678 5274 76730
rect 5326 76678 5338 76730
rect 5390 76678 5402 76730
rect 5454 76678 5466 76730
rect 5518 76678 6810 76730
rect 6862 76678 6874 76730
rect 6926 76678 6938 76730
rect 6990 76678 7002 76730
rect 7054 76678 7066 76730
rect 7118 76678 8410 76730
rect 8462 76678 8474 76730
rect 8526 76678 8538 76730
rect 8590 76678 8602 76730
rect 8654 76678 8666 76730
rect 8718 76678 9936 76730
rect 1104 76656 9936 76678
rect 8680 76520 8984 76548
rect 8680 76489 8708 76520
rect 8956 76492 8984 76520
rect 8665 76483 8723 76489
rect 8665 76449 8677 76483
rect 8711 76449 8723 76483
rect 8665 76443 8723 76449
rect 8754 76440 8760 76492
rect 8812 76440 8818 76492
rect 8938 76440 8944 76492
rect 8996 76440 9002 76492
rect 8202 76372 8208 76424
rect 8260 76412 8266 76424
rect 8389 76415 8447 76421
rect 8389 76412 8401 76415
rect 8260 76384 8401 76412
rect 8260 76372 8266 76384
rect 8389 76381 8401 76384
rect 8435 76381 8447 76415
rect 8389 76375 8447 76381
rect 8481 76415 8539 76421
rect 8481 76381 8493 76415
rect 8527 76412 8539 76415
rect 8772 76412 8800 76440
rect 8527 76384 8800 76412
rect 8527 76381 8539 76384
rect 8481 76375 8539 76381
rect 8404 76344 8432 76375
rect 8846 76344 8852 76356
rect 8404 76316 8852 76344
rect 8846 76304 8852 76316
rect 8904 76304 8910 76356
rect 1118 76236 1124 76288
rect 1176 76276 1182 76288
rect 8021 76279 8079 76285
rect 8021 76276 8033 76279
rect 1176 76248 8033 76276
rect 1176 76236 1182 76248
rect 8021 76245 8033 76248
rect 8067 76245 8079 76279
rect 8021 76239 8079 76245
rect 1104 76186 9936 76208
rect 1104 76134 2950 76186
rect 3002 76134 3014 76186
rect 3066 76134 3078 76186
rect 3130 76134 3142 76186
rect 3194 76134 3206 76186
rect 3258 76134 4550 76186
rect 4602 76134 4614 76186
rect 4666 76134 4678 76186
rect 4730 76134 4742 76186
rect 4794 76134 4806 76186
rect 4858 76134 6150 76186
rect 6202 76134 6214 76186
rect 6266 76134 6278 76186
rect 6330 76134 6342 76186
rect 6394 76134 6406 76186
rect 6458 76134 7750 76186
rect 7802 76134 7814 76186
rect 7866 76134 7878 76186
rect 7930 76134 7942 76186
rect 7994 76134 8006 76186
rect 8058 76134 9350 76186
rect 9402 76134 9414 76186
rect 9466 76134 9478 76186
rect 9530 76134 9542 76186
rect 9594 76134 9606 76186
rect 9658 76134 9936 76186
rect 1104 76112 9936 76134
rect 1486 75896 1492 75948
rect 1544 75896 1550 75948
rect 1673 75803 1731 75809
rect 1673 75769 1685 75803
rect 1719 75800 1731 75803
rect 4062 75800 4068 75812
rect 1719 75772 4068 75800
rect 1719 75769 1731 75772
rect 1673 75763 1731 75769
rect 4062 75760 4068 75772
rect 4120 75760 4126 75812
rect 1104 75642 9936 75664
rect 1104 75590 3610 75642
rect 3662 75590 3674 75642
rect 3726 75590 3738 75642
rect 3790 75590 3802 75642
rect 3854 75590 3866 75642
rect 3918 75590 5210 75642
rect 5262 75590 5274 75642
rect 5326 75590 5338 75642
rect 5390 75590 5402 75642
rect 5454 75590 5466 75642
rect 5518 75590 6810 75642
rect 6862 75590 6874 75642
rect 6926 75590 6938 75642
rect 6990 75590 7002 75642
rect 7054 75590 7066 75642
rect 7118 75590 8410 75642
rect 8462 75590 8474 75642
rect 8526 75590 8538 75642
rect 8590 75590 8602 75642
rect 8654 75590 8666 75642
rect 8718 75590 9936 75642
rect 1104 75568 9936 75590
rect 4430 75352 4436 75404
rect 4488 75392 4494 75404
rect 5718 75392 5724 75404
rect 4488 75364 5724 75392
rect 4488 75352 4494 75364
rect 5718 75352 5724 75364
rect 5776 75352 5782 75404
rect 8478 75352 8484 75404
rect 8536 75392 8542 75404
rect 8536 75364 9352 75392
rect 8536 75352 8542 75364
rect 9214 75284 9220 75336
rect 9272 75284 9278 75336
rect 9324 75333 9352 75364
rect 9309 75327 9367 75333
rect 9309 75293 9321 75327
rect 9355 75293 9367 75327
rect 9309 75287 9367 75293
rect 9401 75327 9459 75333
rect 9401 75293 9413 75327
rect 9447 75293 9459 75327
rect 9401 75287 9459 75293
rect 934 75216 940 75268
rect 992 75256 998 75268
rect 1489 75259 1547 75265
rect 1489 75256 1501 75259
rect 992 75228 1501 75256
rect 992 75216 998 75228
rect 1489 75225 1501 75228
rect 1535 75225 1547 75259
rect 1489 75219 1547 75225
rect 1673 75259 1731 75265
rect 1673 75225 1685 75259
rect 1719 75256 1731 75259
rect 2682 75256 2688 75268
rect 1719 75228 2688 75256
rect 1719 75225 1731 75228
rect 1673 75219 1731 75225
rect 2682 75216 2688 75228
rect 2740 75216 2746 75268
rect 7190 75216 7196 75268
rect 7248 75256 7254 75268
rect 9416 75256 9444 75287
rect 9490 75284 9496 75336
rect 9548 75324 9554 75336
rect 9585 75327 9643 75333
rect 9585 75324 9597 75327
rect 9548 75296 9597 75324
rect 9548 75284 9554 75296
rect 9585 75293 9597 75296
rect 9631 75293 9643 75327
rect 9585 75287 9643 75293
rect 7248 75228 9444 75256
rect 7248 75216 7254 75228
rect 4430 75148 4436 75200
rect 4488 75188 4494 75200
rect 4890 75188 4896 75200
rect 4488 75160 4896 75188
rect 4488 75148 4494 75160
rect 4890 75148 4896 75160
rect 4948 75148 4954 75200
rect 5626 75148 5632 75200
rect 5684 75188 5690 75200
rect 8941 75191 8999 75197
rect 8941 75188 8953 75191
rect 5684 75160 8953 75188
rect 5684 75148 5690 75160
rect 8941 75157 8953 75160
rect 8987 75157 8999 75191
rect 8941 75151 8999 75157
rect 1104 75098 9936 75120
rect 1104 75046 2950 75098
rect 3002 75046 3014 75098
rect 3066 75046 3078 75098
rect 3130 75046 3142 75098
rect 3194 75046 3206 75098
rect 3258 75046 4550 75098
rect 4602 75046 4614 75098
rect 4666 75046 4678 75098
rect 4730 75046 4742 75098
rect 4794 75046 4806 75098
rect 4858 75046 6150 75098
rect 6202 75046 6214 75098
rect 6266 75046 6278 75098
rect 6330 75046 6342 75098
rect 6394 75046 6406 75098
rect 6458 75046 7750 75098
rect 7802 75046 7814 75098
rect 7866 75046 7878 75098
rect 7930 75046 7942 75098
rect 7994 75046 8006 75098
rect 8058 75046 9350 75098
rect 9402 75046 9414 75098
rect 9466 75046 9478 75098
rect 9530 75046 9542 75098
rect 9594 75046 9606 75098
rect 9658 75046 9936 75098
rect 1104 75024 9936 75046
rect 4246 74944 4252 74996
rect 4304 74984 4310 74996
rect 4890 74984 4896 74996
rect 4304 74956 4896 74984
rect 4304 74944 4310 74956
rect 4890 74944 4896 74956
rect 4948 74944 4954 74996
rect 8754 74944 8760 74996
rect 8812 74944 8818 74996
rect 8772 74916 8800 74944
rect 9582 74916 9588 74928
rect 8404 74888 8800 74916
rect 8864 74888 9588 74916
rect 8404 74857 8432 74888
rect 8389 74851 8447 74857
rect 8389 74817 8401 74851
rect 8435 74817 8447 74851
rect 8389 74811 8447 74817
rect 8478 74808 8484 74860
rect 8536 74808 8542 74860
rect 8573 74851 8631 74857
rect 8573 74817 8585 74851
rect 8619 74817 8631 74851
rect 8573 74811 8631 74817
rect 8757 74851 8815 74857
rect 8757 74817 8769 74851
rect 8803 74848 8815 74851
rect 8864 74848 8892 74888
rect 9582 74876 9588 74888
rect 9640 74876 9646 74928
rect 9217 74851 9275 74857
rect 9217 74848 9229 74851
rect 8803 74820 8892 74848
rect 8956 74820 9229 74848
rect 8803 74817 8815 74820
rect 8757 74811 8815 74817
rect 7558 74740 7564 74792
rect 7616 74780 7622 74792
rect 8588 74780 8616 74811
rect 7616 74752 8616 74780
rect 7616 74740 7622 74752
rect 8294 74672 8300 74724
rect 8352 74712 8358 74724
rect 8754 74712 8760 74724
rect 8352 74684 8760 74712
rect 8352 74672 8358 74684
rect 8754 74672 8760 74684
rect 8812 74712 8818 74724
rect 8956 74712 8984 74820
rect 9217 74817 9229 74820
rect 9263 74817 9275 74851
rect 9217 74811 9275 74817
rect 9306 74740 9312 74792
rect 9364 74740 9370 74792
rect 9398 74740 9404 74792
rect 9456 74740 9462 74792
rect 8812 74684 8984 74712
rect 8812 74672 8818 74684
rect 5902 74604 5908 74656
rect 5960 74644 5966 74656
rect 8113 74647 8171 74653
rect 8113 74644 8125 74647
rect 5960 74616 8125 74644
rect 5960 74604 5966 74616
rect 8113 74613 8125 74616
rect 8159 74613 8171 74647
rect 8113 74607 8171 74613
rect 8202 74604 8208 74656
rect 8260 74644 8266 74656
rect 8478 74644 8484 74656
rect 8260 74616 8484 74644
rect 8260 74604 8266 74616
rect 8478 74604 8484 74616
rect 8536 74604 8542 74656
rect 8849 74647 8907 74653
rect 8849 74613 8861 74647
rect 8895 74644 8907 74647
rect 9674 74644 9680 74656
rect 8895 74616 9680 74644
rect 8895 74613 8907 74616
rect 8849 74607 8907 74613
rect 9674 74604 9680 74616
rect 9732 74604 9738 74656
rect 1104 74554 9936 74576
rect 1104 74502 3610 74554
rect 3662 74502 3674 74554
rect 3726 74502 3738 74554
rect 3790 74502 3802 74554
rect 3854 74502 3866 74554
rect 3918 74502 5210 74554
rect 5262 74502 5274 74554
rect 5326 74502 5338 74554
rect 5390 74502 5402 74554
rect 5454 74502 5466 74554
rect 5518 74502 6810 74554
rect 6862 74502 6874 74554
rect 6926 74502 6938 74554
rect 6990 74502 7002 74554
rect 7054 74502 7066 74554
rect 7118 74502 8410 74554
rect 8462 74502 8474 74554
rect 8526 74502 8538 74554
rect 8590 74502 8602 74554
rect 8654 74502 8666 74554
rect 8718 74502 9936 74554
rect 1104 74480 9936 74502
rect 7282 74400 7288 74452
rect 7340 74440 7346 74452
rect 9306 74440 9312 74452
rect 7340 74412 9312 74440
rect 7340 74400 7346 74412
rect 9306 74400 9312 74412
rect 9364 74400 9370 74452
rect 8665 74375 8723 74381
rect 8665 74341 8677 74375
rect 8711 74372 8723 74375
rect 8938 74372 8944 74384
rect 8711 74344 8944 74372
rect 8711 74341 8723 74344
rect 8665 74335 8723 74341
rect 8938 74332 8944 74344
rect 8996 74372 9002 74384
rect 9214 74372 9220 74384
rect 8996 74344 9220 74372
rect 8996 74332 9002 74344
rect 9214 74332 9220 74344
rect 9272 74332 9278 74384
rect 8220 74276 9352 74304
rect 8220 74248 8248 74276
rect 934 74196 940 74248
rect 992 74236 998 74248
rect 1397 74239 1455 74245
rect 1397 74236 1409 74239
rect 992 74208 1409 74236
rect 992 74196 998 74208
rect 1397 74205 1409 74208
rect 1443 74205 1455 74239
rect 1397 74199 1455 74205
rect 6914 74196 6920 74248
rect 6972 74236 6978 74248
rect 7190 74236 7196 74248
rect 6972 74208 7196 74236
rect 6972 74196 6978 74208
rect 7190 74196 7196 74208
rect 7248 74196 7254 74248
rect 8202 74196 8208 74248
rect 8260 74196 8266 74248
rect 8481 74239 8539 74245
rect 8481 74205 8493 74239
rect 8527 74205 8539 74239
rect 8481 74199 8539 74205
rect 8496 74168 8524 74199
rect 9030 74196 9036 74248
rect 9088 74236 9094 74248
rect 9324 74245 9352 74276
rect 9217 74239 9275 74245
rect 9217 74236 9229 74239
rect 9088 74208 9229 74236
rect 9088 74196 9094 74208
rect 9217 74205 9229 74208
rect 9263 74205 9275 74239
rect 9217 74199 9275 74205
rect 9309 74239 9367 74245
rect 9309 74205 9321 74239
rect 9355 74205 9367 74239
rect 9309 74199 9367 74205
rect 9401 74239 9459 74245
rect 9401 74205 9413 74239
rect 9447 74205 9459 74239
rect 9582 74236 9588 74248
rect 9543 74208 9588 74236
rect 9401 74199 9459 74205
rect 8496 74140 9076 74168
rect 9048 74112 9076 74140
rect 9122 74128 9128 74180
rect 9180 74168 9186 74180
rect 9416 74168 9444 74199
rect 9582 74196 9588 74208
rect 9640 74196 9646 74248
rect 9180 74140 9444 74168
rect 9180 74128 9186 74140
rect 1581 74103 1639 74109
rect 1581 74069 1593 74103
rect 1627 74100 1639 74103
rect 1946 74100 1952 74112
rect 1627 74072 1952 74100
rect 1627 74069 1639 74072
rect 1581 74063 1639 74069
rect 1946 74060 1952 74072
rect 2004 74060 2010 74112
rect 8938 74060 8944 74112
rect 8996 74060 9002 74112
rect 9030 74060 9036 74112
rect 9088 74100 9094 74112
rect 9398 74100 9404 74112
rect 9088 74072 9404 74100
rect 9088 74060 9094 74072
rect 9398 74060 9404 74072
rect 9456 74060 9462 74112
rect 9600 74100 9628 74196
rect 9766 74100 9772 74112
rect 9600 74072 9772 74100
rect 9766 74060 9772 74072
rect 9824 74060 9830 74112
rect 1104 74010 9936 74032
rect 1104 73958 2950 74010
rect 3002 73958 3014 74010
rect 3066 73958 3078 74010
rect 3130 73958 3142 74010
rect 3194 73958 3206 74010
rect 3258 73958 4550 74010
rect 4602 73958 4614 74010
rect 4666 73958 4678 74010
rect 4730 73958 4742 74010
rect 4794 73958 4806 74010
rect 4858 73958 6150 74010
rect 6202 73958 6214 74010
rect 6266 73958 6278 74010
rect 6330 73958 6342 74010
rect 6394 73958 6406 74010
rect 6458 73958 7750 74010
rect 7802 73958 7814 74010
rect 7866 73958 7878 74010
rect 7930 73958 7942 74010
rect 7994 73958 8006 74010
rect 8058 73958 9350 74010
rect 9402 73958 9414 74010
rect 9466 73958 9478 74010
rect 9530 73958 9542 74010
rect 9594 73958 9606 74010
rect 9658 73958 9936 74010
rect 1104 73936 9936 73958
rect 3510 73856 3516 73908
rect 3568 73896 3574 73908
rect 3568 73868 9076 73896
rect 3568 73856 3574 73868
rect 6822 73788 6828 73840
rect 6880 73828 6886 73840
rect 6880 73800 8800 73828
rect 6880 73788 6886 73800
rect 6641 73763 6699 73769
rect 6641 73729 6653 73763
rect 6687 73760 6699 73763
rect 6730 73760 6736 73772
rect 6687 73732 6736 73760
rect 6687 73729 6699 73732
rect 6641 73723 6699 73729
rect 6730 73720 6736 73732
rect 6788 73720 6794 73772
rect 7834 73720 7840 73772
rect 7892 73720 7898 73772
rect 7929 73763 7987 73769
rect 7929 73729 7941 73763
rect 7975 73760 7987 73763
rect 8018 73760 8024 73772
rect 7975 73732 8024 73760
rect 7975 73729 7987 73732
rect 7929 73723 7987 73729
rect 8018 73720 8024 73732
rect 8076 73720 8082 73772
rect 8110 73720 8116 73772
rect 8168 73720 8174 73772
rect 8205 73763 8263 73769
rect 8205 73729 8217 73763
rect 8251 73760 8263 73763
rect 8386 73760 8392 73772
rect 8251 73732 8392 73760
rect 8251 73729 8263 73732
rect 8205 73723 8263 73729
rect 8386 73720 8392 73732
rect 8444 73720 8450 73772
rect 8772 73769 8800 73800
rect 8757 73763 8815 73769
rect 8757 73729 8769 73763
rect 8803 73729 8815 73763
rect 8757 73723 8815 73729
rect 6454 73652 6460 73704
rect 6512 73692 6518 73704
rect 6917 73695 6975 73701
rect 6917 73692 6929 73695
rect 6512 73664 6929 73692
rect 6512 73652 6518 73664
rect 6917 73661 6929 73664
rect 6963 73661 6975 73695
rect 6917 73655 6975 73661
rect 7190 73652 7196 73704
rect 7248 73692 7254 73704
rect 7466 73692 7472 73704
rect 7248 73664 7472 73692
rect 7248 73652 7254 73664
rect 7466 73652 7472 73664
rect 7524 73652 7530 73704
rect 9048 73701 9076 73868
rect 9033 73695 9091 73701
rect 9033 73661 9045 73695
rect 9079 73661 9091 73695
rect 9033 73655 9091 73661
rect 7561 73627 7619 73633
rect 7561 73624 7573 73627
rect 6840 73596 7573 73624
rect 6840 73565 6868 73596
rect 7561 73593 7573 73596
rect 7607 73624 7619 73627
rect 9950 73624 9956 73636
rect 7607 73596 9956 73624
rect 7607 73593 7619 73596
rect 7561 73587 7619 73593
rect 9950 73584 9956 73596
rect 10008 73584 10014 73636
rect 6825 73559 6883 73565
rect 6825 73525 6837 73559
rect 6871 73525 6883 73559
rect 6825 73519 6883 73525
rect 6914 73516 6920 73568
rect 6972 73556 6978 73568
rect 7193 73559 7251 73565
rect 7193 73556 7205 73559
rect 6972 73528 7205 73556
rect 6972 73516 6978 73528
rect 7193 73525 7205 73528
rect 7239 73525 7251 73559
rect 7193 73519 7251 73525
rect 7653 73559 7711 73565
rect 7653 73525 7665 73559
rect 7699 73556 7711 73559
rect 8294 73556 8300 73568
rect 7699 73528 8300 73556
rect 7699 73525 7711 73528
rect 7653 73519 7711 73525
rect 8294 73516 8300 73528
rect 8352 73516 8358 73568
rect 8386 73516 8392 73568
rect 8444 73556 8450 73568
rect 9306 73556 9312 73568
rect 8444 73528 9312 73556
rect 8444 73516 8450 73528
rect 9306 73516 9312 73528
rect 9364 73516 9370 73568
rect 1104 73466 9936 73488
rect 1104 73414 3610 73466
rect 3662 73414 3674 73466
rect 3726 73414 3738 73466
rect 3790 73414 3802 73466
rect 3854 73414 3866 73466
rect 3918 73414 5210 73466
rect 5262 73414 5274 73466
rect 5326 73414 5338 73466
rect 5390 73414 5402 73466
rect 5454 73414 5466 73466
rect 5518 73414 6810 73466
rect 6862 73414 6874 73466
rect 6926 73414 6938 73466
rect 6990 73414 7002 73466
rect 7054 73414 7066 73466
rect 7118 73414 8410 73466
rect 8462 73414 8474 73466
rect 8526 73414 8538 73466
rect 8590 73414 8602 73466
rect 8654 73414 8666 73466
rect 8718 73414 9936 73466
rect 1104 73392 9936 73414
rect 4982 73312 4988 73364
rect 5040 73352 5046 73364
rect 7101 73355 7159 73361
rect 7101 73352 7113 73355
rect 5040 73324 7113 73352
rect 5040 73312 5046 73324
rect 7101 73321 7113 73324
rect 7147 73352 7159 73355
rect 7374 73352 7380 73364
rect 7147 73324 7380 73352
rect 7147 73321 7159 73324
rect 7101 73315 7159 73321
rect 7374 73312 7380 73324
rect 7432 73312 7438 73364
rect 8110 73312 8116 73364
rect 8168 73352 8174 73364
rect 8168 73324 8432 73352
rect 8168 73312 8174 73324
rect 8404 73296 8432 73324
rect 8478 73312 8484 73364
rect 8536 73352 8542 73364
rect 8941 73355 8999 73361
rect 8941 73352 8953 73355
rect 8536 73324 8953 73352
rect 8536 73312 8542 73324
rect 8941 73321 8953 73324
rect 8987 73321 8999 73355
rect 8941 73315 8999 73321
rect 5767 73287 5825 73293
rect 5767 73253 5779 73287
rect 5813 73284 5825 73287
rect 7834 73284 7840 73296
rect 5813 73256 7840 73284
rect 5813 73253 5825 73256
rect 5767 73247 5825 73253
rect 7834 73244 7840 73256
rect 7892 73284 7898 73296
rect 8202 73284 8208 73296
rect 7892 73256 8208 73284
rect 7892 73244 7898 73256
rect 5537 73219 5595 73225
rect 5537 73185 5549 73219
rect 5583 73216 5595 73219
rect 6638 73216 6644 73228
rect 5583 73188 6644 73216
rect 5583 73185 5595 73188
rect 5537 73179 5595 73185
rect 6638 73176 6644 73188
rect 6696 73176 6702 73228
rect 6914 73216 6920 73228
rect 6748 73188 6920 73216
rect 6454 73108 6460 73160
rect 6512 73148 6518 73160
rect 6748 73148 6776 73188
rect 6914 73176 6920 73188
rect 6972 73216 6978 73228
rect 7285 73219 7343 73225
rect 7285 73216 7297 73219
rect 6972 73188 7297 73216
rect 6972 73176 6978 73188
rect 7285 73185 7297 73188
rect 7331 73185 7343 73219
rect 7742 73216 7748 73228
rect 7285 73179 7343 73185
rect 7484 73188 7748 73216
rect 6512 73120 6776 73148
rect 6512 73108 6518 73120
rect 6822 73108 6828 73160
rect 6880 73148 6886 73160
rect 7009 73151 7067 73157
rect 7009 73148 7021 73151
rect 6880 73120 7021 73148
rect 6880 73108 6886 73120
rect 7009 73117 7021 73120
rect 7055 73117 7067 73151
rect 7009 73111 7067 73117
rect 7484 73092 7512 73188
rect 7742 73176 7748 73188
rect 7800 73176 7806 73228
rect 7926 73176 7932 73228
rect 7984 73176 7990 73228
rect 8128 73216 8156 73256
rect 8202 73244 8208 73256
rect 8260 73244 8266 73296
rect 8386 73244 8392 73296
rect 8444 73284 8450 73296
rect 8444 73256 9444 73284
rect 8444 73244 8450 73256
rect 8128 73188 9168 73216
rect 7558 73108 7564 73160
rect 7616 73108 7622 73160
rect 8128 73157 8156 73188
rect 8113 73151 8171 73157
rect 8113 73117 8125 73151
rect 8159 73117 8171 73151
rect 8113 73111 8171 73117
rect 8205 73151 8263 73157
rect 8205 73117 8217 73151
rect 8251 73117 8263 73151
rect 8205 73111 8263 73117
rect 934 73040 940 73092
rect 992 73080 998 73092
rect 1489 73083 1547 73089
rect 1489 73080 1501 73083
rect 992 73052 1501 73080
rect 992 73040 998 73052
rect 1489 73049 1501 73052
rect 1535 73049 1547 73083
rect 1489 73043 1547 73049
rect 4338 73040 4344 73092
rect 4396 73080 4402 73092
rect 7098 73080 7104 73092
rect 4396 73052 7104 73080
rect 4396 73040 4402 73052
rect 7098 73040 7104 73052
rect 7156 73040 7162 73092
rect 7466 73040 7472 73092
rect 7524 73040 7530 73092
rect 1578 72972 1584 73024
rect 1636 72972 1642 73024
rect 7576 73021 7604 73108
rect 7650 73040 7656 73092
rect 7708 73080 7714 73092
rect 8220 73080 8248 73111
rect 8386 73108 8392 73160
rect 8444 73108 8450 73160
rect 8481 73151 8539 73157
rect 8481 73117 8493 73151
rect 8527 73117 8539 73151
rect 8481 73111 8539 73117
rect 7708 73052 8248 73080
rect 7708 73040 7714 73052
rect 8496 73024 8524 73111
rect 8846 73108 8852 73160
rect 8904 73108 8910 73160
rect 9140 73157 9168 73188
rect 9416 73157 9444 73256
rect 9125 73151 9183 73157
rect 9125 73117 9137 73151
rect 9171 73117 9183 73151
rect 9125 73111 9183 73117
rect 9217 73151 9275 73157
rect 9217 73117 9229 73151
rect 9263 73117 9275 73151
rect 9217 73111 9275 73117
rect 9401 73151 9459 73157
rect 9401 73117 9413 73151
rect 9447 73117 9459 73151
rect 9401 73111 9459 73117
rect 9493 73151 9551 73157
rect 9493 73117 9505 73151
rect 9539 73117 9551 73151
rect 9493 73111 9551 73117
rect 8864 73080 8892 73108
rect 9232 73080 9260 73111
rect 9508 73080 9536 73111
rect 10134 73108 10140 73160
rect 10192 73148 10198 73160
rect 10502 73148 10508 73160
rect 10192 73120 10508 73148
rect 10192 73108 10198 73120
rect 10502 73108 10508 73120
rect 10560 73108 10566 73160
rect 8864 73052 9260 73080
rect 9416 73052 9536 73080
rect 7561 73015 7619 73021
rect 7561 72981 7573 73015
rect 7607 72981 7619 73015
rect 7561 72975 7619 72981
rect 8478 72972 8484 73024
rect 8536 73012 8542 73024
rect 9306 73012 9312 73024
rect 8536 72984 9312 73012
rect 8536 72972 8542 72984
rect 9306 72972 9312 72984
rect 9364 73012 9370 73024
rect 9416 73012 9444 73052
rect 9364 72984 9444 73012
rect 9364 72972 9370 72984
rect 1104 72922 9936 72944
rect 1104 72870 2950 72922
rect 3002 72870 3014 72922
rect 3066 72870 3078 72922
rect 3130 72870 3142 72922
rect 3194 72870 3206 72922
rect 3258 72870 4550 72922
rect 4602 72870 4614 72922
rect 4666 72870 4678 72922
rect 4730 72870 4742 72922
rect 4794 72870 4806 72922
rect 4858 72870 6150 72922
rect 6202 72870 6214 72922
rect 6266 72870 6278 72922
rect 6330 72870 6342 72922
rect 6394 72870 6406 72922
rect 6458 72870 7750 72922
rect 7802 72870 7814 72922
rect 7866 72870 7878 72922
rect 7930 72870 7942 72922
rect 7994 72870 8006 72922
rect 8058 72870 9350 72922
rect 9402 72870 9414 72922
rect 9466 72870 9478 72922
rect 9530 72870 9542 72922
rect 9594 72870 9606 72922
rect 9658 72870 9936 72922
rect 1104 72848 9936 72870
rect 8478 72808 8484 72820
rect 2056 72780 8484 72808
rect 2056 72684 2084 72780
rect 8478 72768 8484 72780
rect 8536 72808 8542 72820
rect 8536 72780 9168 72808
rect 8536 72768 8542 72780
rect 5994 72700 6000 72752
rect 6052 72740 6058 72752
rect 6052 72712 8248 72740
rect 6052 72700 6058 72712
rect 2038 72632 2044 72684
rect 2096 72632 2102 72684
rect 4246 72632 4252 72684
rect 4304 72672 4310 72684
rect 6454 72672 6460 72684
rect 4304 72644 6460 72672
rect 4304 72632 4310 72644
rect 6454 72632 6460 72644
rect 6512 72672 6518 72684
rect 6822 72672 6828 72684
rect 6512 72644 6828 72672
rect 6512 72632 6518 72644
rect 6822 72632 6828 72644
rect 6880 72632 6886 72684
rect 7190 72632 7196 72684
rect 7248 72672 7254 72684
rect 7374 72672 7380 72684
rect 7248 72644 7380 72672
rect 7248 72632 7254 72644
rect 7374 72632 7380 72644
rect 7432 72632 7438 72684
rect 7466 72632 7472 72684
rect 7524 72632 7530 72684
rect 7561 72675 7619 72681
rect 7561 72641 7573 72675
rect 7607 72672 7619 72675
rect 7650 72672 7656 72684
rect 7607 72644 7656 72672
rect 7607 72641 7619 72644
rect 7561 72635 7619 72641
rect 7650 72632 7656 72644
rect 7708 72632 7714 72684
rect 7745 72675 7803 72681
rect 7745 72641 7757 72675
rect 7791 72672 7803 72675
rect 7926 72672 7932 72684
rect 7791 72644 7932 72672
rect 7791 72641 7803 72644
rect 7745 72635 7803 72641
rect 7926 72632 7932 72644
rect 7984 72632 7990 72684
rect 8220 72681 8248 72712
rect 8404 72712 9076 72740
rect 8404 72684 8432 72712
rect 8113 72675 8171 72681
rect 8113 72641 8125 72675
rect 8159 72641 8171 72675
rect 8113 72635 8171 72641
rect 8205 72675 8263 72681
rect 8205 72641 8217 72675
rect 8251 72641 8263 72675
rect 8205 72635 8263 72641
rect 5994 72564 6000 72616
rect 6052 72604 6058 72616
rect 6733 72607 6791 72613
rect 6733 72604 6745 72607
rect 6052 72576 6745 72604
rect 6052 72564 6058 72576
rect 6733 72573 6745 72576
rect 6779 72604 6791 72607
rect 6914 72604 6920 72616
rect 6779 72576 6920 72604
rect 6779 72573 6791 72576
rect 6733 72567 6791 72573
rect 6914 72564 6920 72576
rect 6972 72564 6978 72616
rect 7098 72564 7104 72616
rect 7156 72604 7162 72616
rect 8018 72604 8024 72616
rect 7156 72576 8024 72604
rect 7156 72564 7162 72576
rect 8018 72564 8024 72576
rect 8076 72564 8082 72616
rect 8128 72604 8156 72635
rect 8386 72632 8392 72684
rect 8444 72632 8450 72684
rect 8478 72632 8484 72684
rect 8536 72632 8542 72684
rect 8757 72675 8815 72681
rect 8757 72641 8769 72675
rect 8803 72641 8815 72675
rect 8757 72635 8815 72641
rect 8772 72604 8800 72635
rect 8846 72632 8852 72684
rect 8904 72632 8910 72684
rect 9048 72681 9076 72712
rect 9140 72681 9168 72780
rect 9033 72675 9091 72681
rect 9033 72641 9045 72675
rect 9079 72641 9091 72675
rect 9033 72635 9091 72641
rect 9125 72675 9183 72681
rect 9125 72641 9137 72675
rect 9171 72641 9183 72675
rect 9125 72635 9183 72641
rect 9217 72675 9275 72681
rect 9217 72641 9229 72675
rect 9263 72641 9275 72675
rect 9217 72635 9275 72641
rect 8128 72576 8800 72604
rect 8220 72548 8248 72576
rect 4890 72496 4896 72548
rect 4948 72536 4954 72548
rect 4948 72508 8061 72536
rect 4948 72496 4954 72508
rect 6822 72428 6828 72480
rect 6880 72428 6886 72480
rect 7006 72428 7012 72480
rect 7064 72428 7070 72480
rect 7101 72471 7159 72477
rect 7101 72437 7113 72471
rect 7147 72468 7159 72471
rect 7466 72468 7472 72480
rect 7147 72440 7472 72468
rect 7147 72437 7159 72440
rect 7101 72431 7159 72437
rect 7466 72428 7472 72440
rect 7524 72428 7530 72480
rect 7742 72428 7748 72480
rect 7800 72468 7806 72480
rect 7929 72471 7987 72477
rect 7929 72468 7941 72471
rect 7800 72440 7941 72468
rect 7800 72428 7806 72440
rect 7929 72437 7941 72440
rect 7975 72437 7987 72471
rect 8033 72468 8061 72508
rect 8202 72496 8208 72548
rect 8260 72496 8266 72548
rect 9232 72536 9260 72635
rect 9398 72564 9404 72616
rect 9456 72604 9462 72616
rect 10134 72604 10140 72616
rect 9456 72576 10140 72604
rect 9456 72564 9462 72576
rect 10134 72564 10140 72576
rect 10192 72564 10198 72616
rect 8312 72508 9260 72536
rect 8312 72468 8340 72508
rect 8033 72440 8340 72468
rect 7929 72431 7987 72437
rect 8570 72428 8576 72480
rect 8628 72428 8634 72480
rect 9398 72428 9404 72480
rect 9456 72428 9462 72480
rect 1104 72378 9936 72400
rect 1104 72326 3610 72378
rect 3662 72326 3674 72378
rect 3726 72326 3738 72378
rect 3790 72326 3802 72378
rect 3854 72326 3866 72378
rect 3918 72326 5210 72378
rect 5262 72326 5274 72378
rect 5326 72326 5338 72378
rect 5390 72326 5402 72378
rect 5454 72326 5466 72378
rect 5518 72326 6810 72378
rect 6862 72326 6874 72378
rect 6926 72326 6938 72378
rect 6990 72326 7002 72378
rect 7054 72326 7066 72378
rect 7118 72326 8410 72378
rect 8462 72326 8474 72378
rect 8526 72326 8538 72378
rect 8590 72326 8602 72378
rect 8654 72326 8666 72378
rect 8718 72326 9936 72378
rect 1104 72304 9936 72326
rect 5534 72224 5540 72276
rect 5592 72264 5598 72276
rect 7377 72267 7435 72273
rect 7377 72264 7389 72267
rect 5592 72236 7389 72264
rect 5592 72224 5598 72236
rect 7377 72233 7389 72236
rect 7423 72264 7435 72267
rect 7423 72236 7604 72264
rect 7423 72233 7435 72236
rect 7377 72227 7435 72233
rect 6454 72088 6460 72140
rect 6512 72088 6518 72140
rect 7190 72128 7196 72140
rect 6656 72100 7196 72128
rect 5353 72063 5411 72069
rect 5353 72029 5365 72063
rect 5399 72060 5411 72063
rect 5534 72060 5540 72072
rect 5399 72032 5540 72060
rect 5399 72029 5411 72032
rect 5353 72023 5411 72029
rect 5534 72020 5540 72032
rect 5592 72020 5598 72072
rect 5629 72063 5687 72069
rect 5629 72029 5641 72063
rect 5675 72029 5687 72063
rect 5629 72023 5687 72029
rect 934 71952 940 72004
rect 992 71992 998 72004
rect 1489 71995 1547 72001
rect 1489 71992 1501 71995
rect 992 71964 1501 71992
rect 992 71952 998 71964
rect 1489 71961 1501 71964
rect 1535 71961 1547 71995
rect 5644 71992 5672 72023
rect 5718 72020 5724 72072
rect 5776 72060 5782 72072
rect 6365 72063 6423 72069
rect 6365 72060 6377 72063
rect 5776 72032 6377 72060
rect 5776 72020 5782 72032
rect 6365 72029 6377 72032
rect 6411 72029 6423 72063
rect 6365 72023 6423 72029
rect 6270 71992 6276 72004
rect 5644 71964 6276 71992
rect 1489 71955 1547 71961
rect 6270 71952 6276 71964
rect 6328 71952 6334 72004
rect 6472 71992 6500 72088
rect 6656 72069 6684 72100
rect 7190 72088 7196 72100
rect 7248 72088 7254 72140
rect 7576 72128 7604 72236
rect 7650 72224 7656 72276
rect 7708 72264 7714 72276
rect 7837 72267 7895 72273
rect 7837 72264 7849 72267
rect 7708 72236 7849 72264
rect 7708 72224 7714 72236
rect 7837 72233 7849 72236
rect 7883 72233 7895 72267
rect 7837 72227 7895 72233
rect 7926 72156 7932 72208
rect 7984 72196 7990 72208
rect 9766 72196 9772 72208
rect 7984 72168 9772 72196
rect 7984 72156 7990 72168
rect 9766 72156 9772 72168
rect 9824 72156 9830 72208
rect 8570 72128 8576 72140
rect 7576 72100 8576 72128
rect 8570 72088 8576 72100
rect 8628 72088 8634 72140
rect 6641 72063 6699 72069
rect 6641 72029 6653 72063
rect 6687 72029 6699 72063
rect 6641 72023 6699 72029
rect 7285 72063 7343 72069
rect 7285 72029 7297 72063
rect 7331 72029 7343 72063
rect 7285 72023 7343 72029
rect 7561 72063 7619 72069
rect 7561 72029 7573 72063
rect 7607 72029 7619 72063
rect 7561 72023 7619 72029
rect 7300 71992 7328 72023
rect 6472 71964 7328 71992
rect 1578 71884 1584 71936
rect 1636 71884 1642 71936
rect 5994 71884 6000 71936
rect 6052 71924 6058 71936
rect 7576 71924 7604 72023
rect 8018 72020 8024 72072
rect 8076 72060 8082 72072
rect 8113 72063 8171 72069
rect 8113 72060 8125 72063
rect 8076 72032 8125 72060
rect 8076 72020 8082 72032
rect 8113 72029 8125 72032
rect 8159 72029 8171 72063
rect 8113 72023 8171 72029
rect 6052 71896 7604 71924
rect 8297 71927 8355 71933
rect 6052 71884 6058 71896
rect 8297 71893 8309 71927
rect 8343 71924 8355 71927
rect 8386 71924 8392 71936
rect 8343 71896 8392 71924
rect 8343 71893 8355 71896
rect 8297 71887 8355 71893
rect 8386 71884 8392 71896
rect 8444 71884 8450 71936
rect 1104 71834 9936 71856
rect 1104 71782 2950 71834
rect 3002 71782 3014 71834
rect 3066 71782 3078 71834
rect 3130 71782 3142 71834
rect 3194 71782 3206 71834
rect 3258 71782 4550 71834
rect 4602 71782 4614 71834
rect 4666 71782 4678 71834
rect 4730 71782 4742 71834
rect 4794 71782 4806 71834
rect 4858 71782 6150 71834
rect 6202 71782 6214 71834
rect 6266 71782 6278 71834
rect 6330 71782 6342 71834
rect 6394 71782 6406 71834
rect 6458 71782 7750 71834
rect 7802 71782 7814 71834
rect 7866 71782 7878 71834
rect 7930 71782 7942 71834
rect 7994 71782 8006 71834
rect 8058 71782 9350 71834
rect 9402 71782 9414 71834
rect 9466 71782 9478 71834
rect 9530 71782 9542 71834
rect 9594 71782 9606 71834
rect 9658 71782 9936 71834
rect 1104 71760 9936 71782
rect 4338 71680 4344 71732
rect 4396 71720 4402 71732
rect 6822 71720 6828 71732
rect 4396 71692 6828 71720
rect 4396 71680 4402 71692
rect 6822 71680 6828 71692
rect 6880 71680 6886 71732
rect 7282 71680 7288 71732
rect 7340 71720 7346 71732
rect 10870 71720 10876 71732
rect 7340 71692 8156 71720
rect 7340 71680 7346 71692
rect 658 71612 664 71664
rect 716 71652 722 71664
rect 1118 71652 1124 71664
rect 716 71624 1124 71652
rect 716 71612 722 71624
rect 1118 71612 1124 71624
rect 1176 71612 1182 71664
rect 4890 71612 4896 71664
rect 4948 71652 4954 71664
rect 7837 71655 7895 71661
rect 7837 71652 7849 71655
rect 4948 71624 7849 71652
rect 4948 71612 4954 71624
rect 7837 71621 7849 71624
rect 7883 71621 7895 71655
rect 7837 71615 7895 71621
rect 934 71544 940 71596
rect 992 71584 998 71596
rect 1489 71587 1547 71593
rect 1489 71584 1501 71587
rect 992 71556 1501 71584
rect 992 71544 998 71556
rect 1489 71553 1501 71556
rect 1535 71553 1547 71587
rect 1489 71547 1547 71553
rect 6362 71544 6368 71596
rect 6420 71544 6426 71596
rect 6454 71544 6460 71596
rect 6512 71584 6518 71596
rect 6632 71587 6690 71593
rect 6632 71584 6644 71587
rect 6512 71556 6644 71584
rect 6512 71544 6518 71556
rect 6632 71553 6644 71556
rect 6678 71584 6690 71587
rect 7098 71584 7104 71596
rect 6678 71556 7104 71584
rect 6678 71553 6690 71556
rect 6632 71547 6690 71553
rect 7098 71544 7104 71556
rect 7156 71544 7162 71596
rect 7190 71544 7196 71596
rect 7248 71584 7254 71596
rect 7742 71584 7748 71596
rect 7248 71556 7748 71584
rect 7248 71544 7254 71556
rect 7742 71544 7748 71556
rect 7800 71544 7806 71596
rect 8128 71593 8156 71692
rect 9232 71692 10876 71720
rect 9122 71612 9128 71664
rect 9180 71652 9186 71664
rect 9232 71661 9260 71692
rect 10870 71680 10876 71692
rect 10928 71680 10934 71732
rect 11330 71680 11336 71732
rect 11388 71680 11394 71732
rect 9217 71655 9275 71661
rect 9217 71652 9229 71655
rect 9180 71624 9229 71652
rect 9180 71612 9186 71624
rect 9217 71621 9229 71624
rect 9263 71621 9275 71655
rect 9217 71615 9275 71621
rect 9309 71655 9367 71661
rect 9309 71621 9321 71655
rect 9355 71652 9367 71655
rect 11348 71652 11376 71680
rect 9355 71624 11376 71652
rect 9355 71621 9367 71624
rect 9309 71615 9367 71621
rect 8113 71587 8171 71593
rect 8113 71553 8125 71587
rect 8159 71553 8171 71587
rect 8113 71547 8171 71553
rect 8202 71544 8208 71596
rect 8260 71544 8266 71596
rect 8297 71587 8355 71593
rect 8297 71553 8309 71587
rect 8343 71553 8355 71587
rect 8297 71547 8355 71553
rect 8481 71587 8539 71593
rect 8481 71553 8493 71587
rect 8527 71553 8539 71587
rect 8481 71547 8539 71553
rect 1118 71476 1124 71528
rect 1176 71516 1182 71528
rect 1302 71516 1308 71528
rect 1176 71488 1308 71516
rect 1176 71476 1182 71488
rect 1302 71476 1308 71488
rect 1360 71476 1366 71528
rect 7374 71476 7380 71528
rect 7432 71516 7438 71528
rect 8312 71516 8340 71547
rect 7432 71488 8340 71516
rect 7432 71476 7438 71488
rect 8496 71448 8524 71547
rect 9030 71544 9036 71596
rect 9088 71584 9094 71596
rect 9088 71556 9444 71584
rect 9088 71544 9094 71556
rect 8570 71476 8576 71528
rect 8628 71516 8634 71528
rect 9416 71516 9444 71556
rect 9493 71519 9551 71525
rect 9493 71516 9505 71519
rect 8628 71488 9076 71516
rect 9416 71488 9505 71516
rect 8628 71476 8634 71488
rect 9048 71460 9076 71488
rect 9493 71485 9505 71488
rect 9539 71516 9551 71519
rect 11146 71516 11152 71528
rect 9539 71488 11152 71516
rect 9539 71485 9551 71488
rect 9493 71479 9551 71485
rect 11146 71476 11152 71488
rect 11204 71476 11210 71528
rect 7944 71420 8524 71448
rect 7944 71392 7972 71420
rect 9030 71408 9036 71460
rect 9088 71408 9094 71460
rect 566 71340 572 71392
rect 624 71380 630 71392
rect 1581 71383 1639 71389
rect 1581 71380 1593 71383
rect 624 71352 1593 71380
rect 624 71340 630 71352
rect 1581 71349 1593 71352
rect 1627 71349 1639 71383
rect 1581 71343 1639 71349
rect 5534 71340 5540 71392
rect 5592 71380 5598 71392
rect 6730 71380 6736 71392
rect 5592 71352 6736 71380
rect 5592 71340 5598 71352
rect 6730 71340 6736 71352
rect 6788 71340 6794 71392
rect 7098 71340 7104 71392
rect 7156 71380 7162 71392
rect 7745 71383 7803 71389
rect 7745 71380 7757 71383
rect 7156 71352 7757 71380
rect 7156 71340 7162 71352
rect 7745 71349 7757 71352
rect 7791 71349 7803 71383
rect 7745 71343 7803 71349
rect 7926 71340 7932 71392
rect 7984 71340 7990 71392
rect 8849 71383 8907 71389
rect 8849 71349 8861 71383
rect 8895 71380 8907 71383
rect 11238 71380 11244 71392
rect 8895 71352 11244 71380
rect 8895 71349 8907 71352
rect 8849 71343 8907 71349
rect 11238 71340 11244 71352
rect 11296 71340 11302 71392
rect 1104 71290 9936 71312
rect 1104 71238 3610 71290
rect 3662 71238 3674 71290
rect 3726 71238 3738 71290
rect 3790 71238 3802 71290
rect 3854 71238 3866 71290
rect 3918 71238 5210 71290
rect 5262 71238 5274 71290
rect 5326 71238 5338 71290
rect 5390 71238 5402 71290
rect 5454 71238 5466 71290
rect 5518 71238 6810 71290
rect 6862 71238 6874 71290
rect 6926 71238 6938 71290
rect 6990 71238 7002 71290
rect 7054 71238 7066 71290
rect 7118 71238 8410 71290
rect 8462 71238 8474 71290
rect 8526 71238 8538 71290
rect 8590 71238 8602 71290
rect 8654 71238 8666 71290
rect 8718 71238 9936 71290
rect 1104 71216 9936 71238
rect 6454 71136 6460 71188
rect 6512 71176 6518 71188
rect 6914 71176 6920 71188
rect 6512 71148 6920 71176
rect 6512 71136 6518 71148
rect 6914 71136 6920 71148
rect 6972 71136 6978 71188
rect 7006 71136 7012 71188
rect 7064 71176 7070 71188
rect 7282 71176 7288 71188
rect 7064 71148 7288 71176
rect 7064 71136 7070 71148
rect 7282 71136 7288 71148
rect 7340 71136 7346 71188
rect 7834 71136 7840 71188
rect 7892 71176 7898 71188
rect 9125 71179 9183 71185
rect 9125 71176 9137 71179
rect 7892 71148 9137 71176
rect 7892 71136 7898 71148
rect 9125 71145 9137 71148
rect 9171 71145 9183 71179
rect 9125 71139 9183 71145
rect 6822 71068 6828 71120
rect 6880 71108 6886 71120
rect 7558 71108 7564 71120
rect 6880 71080 7564 71108
rect 6880 71068 6886 71080
rect 7558 71068 7564 71080
rect 7616 71068 7622 71120
rect 8021 71111 8079 71117
rect 8021 71077 8033 71111
rect 8067 71108 8079 71111
rect 9766 71108 9772 71120
rect 8067 71080 9772 71108
rect 8067 71077 8079 71080
rect 8021 71071 8079 71077
rect 9766 71068 9772 71080
rect 9824 71068 9830 71120
rect 5718 71000 5724 71052
rect 5776 71040 5782 71052
rect 7926 71040 7932 71052
rect 5776 71012 7932 71040
rect 5776 71000 5782 71012
rect 7926 71000 7932 71012
rect 7984 71040 7990 71052
rect 8386 71040 8392 71052
rect 7984 71012 8392 71040
rect 7984 71000 7990 71012
rect 8386 71000 8392 71012
rect 8444 71000 8450 71052
rect 8478 71000 8484 71052
rect 8536 71000 8542 71052
rect 8665 71043 8723 71049
rect 8665 71009 8677 71043
rect 8711 71040 8723 71043
rect 9214 71040 9220 71052
rect 8711 71012 9220 71040
rect 8711 71009 8723 71012
rect 8665 71003 8723 71009
rect 9214 71000 9220 71012
rect 9272 71000 9278 71052
rect 5534 70932 5540 70984
rect 5592 70972 5598 70984
rect 6546 70972 6552 70984
rect 5592 70944 6552 70972
rect 5592 70932 5598 70944
rect 6546 70932 6552 70944
rect 6604 70932 6610 70984
rect 6825 70975 6883 70981
rect 6825 70941 6837 70975
rect 6871 70972 6883 70975
rect 7006 70972 7012 70984
rect 6871 70944 7012 70972
rect 6871 70941 6883 70944
rect 6825 70935 6883 70941
rect 7006 70932 7012 70944
rect 7064 70932 7070 70984
rect 7098 70932 7104 70984
rect 7156 70972 7162 70984
rect 8496 70972 8524 71000
rect 7156 70944 8524 70972
rect 9033 70975 9091 70981
rect 7156 70932 7162 70944
rect 9033 70941 9045 70975
rect 9079 70972 9091 70975
rect 10226 70972 10232 70984
rect 9079 70944 10232 70972
rect 9079 70941 9091 70944
rect 9033 70935 9091 70941
rect 10226 70932 10232 70944
rect 10284 70932 10290 70984
rect 2774 70864 2780 70916
rect 2832 70904 2838 70916
rect 8570 70904 8576 70916
rect 2832 70876 8576 70904
rect 2832 70864 2838 70876
rect 8570 70864 8576 70876
rect 8628 70864 8634 70916
rect 2406 70796 2412 70848
rect 2464 70836 2470 70848
rect 3510 70836 3516 70848
rect 2464 70808 3516 70836
rect 2464 70796 2470 70808
rect 3510 70796 3516 70808
rect 3568 70796 3574 70848
rect 7190 70796 7196 70848
rect 7248 70836 7254 70848
rect 7374 70836 7380 70848
rect 7248 70808 7380 70836
rect 7248 70796 7254 70808
rect 7374 70796 7380 70808
rect 7432 70796 7438 70848
rect 7745 70839 7803 70845
rect 7745 70805 7757 70839
rect 7791 70836 7803 70839
rect 8389 70839 8447 70845
rect 8389 70836 8401 70839
rect 7791 70808 8401 70836
rect 7791 70805 7803 70808
rect 7745 70799 7803 70805
rect 8389 70805 8401 70808
rect 8435 70836 8447 70839
rect 8478 70836 8484 70848
rect 8435 70808 8484 70836
rect 8435 70805 8447 70808
rect 8389 70799 8447 70805
rect 8478 70796 8484 70808
rect 8536 70796 8542 70848
rect 8846 70796 8852 70848
rect 8904 70836 8910 70848
rect 9122 70836 9128 70848
rect 8904 70808 9128 70836
rect 8904 70796 8910 70808
rect 9122 70796 9128 70808
rect 9180 70796 9186 70848
rect 1104 70746 9936 70768
rect 1104 70694 2950 70746
rect 3002 70694 3014 70746
rect 3066 70694 3078 70746
rect 3130 70694 3142 70746
rect 3194 70694 3206 70746
rect 3258 70694 4550 70746
rect 4602 70694 4614 70746
rect 4666 70694 4678 70746
rect 4730 70694 4742 70746
rect 4794 70694 4806 70746
rect 4858 70694 6150 70746
rect 6202 70694 6214 70746
rect 6266 70694 6278 70746
rect 6330 70694 6342 70746
rect 6394 70694 6406 70746
rect 6458 70694 7750 70746
rect 7802 70694 7814 70746
rect 7866 70694 7878 70746
rect 7930 70694 7942 70746
rect 7994 70694 8006 70746
rect 8058 70694 9350 70746
rect 9402 70694 9414 70746
rect 9466 70694 9478 70746
rect 9530 70694 9542 70746
rect 9594 70694 9606 70746
rect 9658 70694 9936 70746
rect 1104 70672 9936 70694
rect 658 70592 664 70644
rect 716 70632 722 70644
rect 1581 70635 1639 70641
rect 1581 70632 1593 70635
rect 716 70604 1593 70632
rect 716 70592 722 70604
rect 1581 70601 1593 70604
rect 1627 70601 1639 70635
rect 1581 70595 1639 70601
rect 6362 70592 6368 70644
rect 6420 70632 6426 70644
rect 6822 70632 6828 70644
rect 6420 70604 6828 70632
rect 6420 70592 6426 70604
rect 6822 70592 6828 70604
rect 6880 70592 6886 70644
rect 6932 70604 7420 70632
rect 6546 70524 6552 70576
rect 6604 70564 6610 70576
rect 6932 70564 6960 70604
rect 6604 70536 6960 70564
rect 6604 70524 6610 70536
rect 7006 70524 7012 70576
rect 7064 70564 7070 70576
rect 7064 70536 7236 70564
rect 7064 70524 7070 70536
rect 1394 70456 1400 70508
rect 1452 70456 1458 70508
rect 2038 70456 2044 70508
rect 2096 70456 2102 70508
rect 3510 70456 3516 70508
rect 3568 70496 3574 70508
rect 4338 70496 4344 70508
rect 3568 70468 4344 70496
rect 3568 70456 3574 70468
rect 4338 70456 4344 70468
rect 4396 70456 4402 70508
rect 6454 70456 6460 70508
rect 6512 70496 6518 70508
rect 6914 70496 6920 70508
rect 6512 70468 6920 70496
rect 6512 70456 6518 70468
rect 6914 70456 6920 70468
rect 6972 70456 6978 70508
rect 7098 70456 7104 70508
rect 7156 70456 7162 70508
rect 7208 70505 7236 70536
rect 7392 70508 7420 70604
rect 7742 70592 7748 70644
rect 7800 70632 7806 70644
rect 7800 70604 8321 70632
rect 7800 70592 7806 70604
rect 8293 70564 8321 70604
rect 8570 70592 8576 70644
rect 8628 70632 8634 70644
rect 8757 70635 8815 70641
rect 8757 70632 8769 70635
rect 8628 70604 8769 70632
rect 8628 70592 8634 70604
rect 8757 70601 8769 70604
rect 8803 70601 8815 70635
rect 8757 70595 8815 70601
rect 8849 70635 8907 70641
rect 8849 70601 8861 70635
rect 8895 70601 8907 70635
rect 8849 70595 8907 70601
rect 8864 70564 8892 70595
rect 9122 70592 9128 70644
rect 9180 70632 9186 70644
rect 9217 70635 9275 70641
rect 9217 70632 9229 70635
rect 9180 70604 9229 70632
rect 9180 70592 9186 70604
rect 9217 70601 9229 70604
rect 9263 70601 9275 70635
rect 10042 70632 10048 70644
rect 9217 70595 9275 70601
rect 9324 70604 10048 70632
rect 9324 70564 9352 70604
rect 10042 70592 10048 70604
rect 10100 70592 10106 70644
rect 8036 70536 8248 70564
rect 8293 70536 8708 70564
rect 8864 70536 9352 70564
rect 8036 70508 8064 70536
rect 8220 70508 8248 70536
rect 7193 70499 7251 70505
rect 7193 70465 7205 70499
rect 7239 70465 7251 70499
rect 7193 70459 7251 70465
rect 7285 70499 7343 70505
rect 7285 70465 7297 70499
rect 7331 70465 7343 70499
rect 7285 70459 7343 70465
rect 2056 70428 2084 70456
rect 1320 70400 2084 70428
rect 1320 70304 1348 70400
rect 5994 70388 6000 70440
rect 6052 70428 6058 70440
rect 6825 70431 6883 70437
rect 6825 70428 6837 70431
rect 6052 70400 6837 70428
rect 6052 70388 6058 70400
rect 6825 70397 6837 70400
rect 6871 70397 6883 70431
rect 6825 70391 6883 70397
rect 5718 70360 5724 70372
rect 4448 70332 5724 70360
rect 4448 70304 4476 70332
rect 5718 70320 5724 70332
rect 5776 70320 5782 70372
rect 5810 70320 5816 70372
rect 5868 70360 5874 70372
rect 7116 70360 7144 70456
rect 5868 70332 7144 70360
rect 5868 70320 5874 70332
rect 1302 70252 1308 70304
rect 1360 70252 1366 70304
rect 4430 70252 4436 70304
rect 4488 70252 4494 70304
rect 4706 70252 4712 70304
rect 4764 70292 4770 70304
rect 6086 70292 6092 70304
rect 4764 70264 6092 70292
rect 4764 70252 4770 70264
rect 6086 70252 6092 70264
rect 6144 70252 6150 70304
rect 6178 70252 6184 70304
rect 6236 70292 6242 70304
rect 7300 70292 7328 70459
rect 7374 70456 7380 70508
rect 7432 70456 7438 70508
rect 7469 70499 7527 70505
rect 7469 70465 7481 70499
rect 7515 70496 7527 70499
rect 7650 70496 7656 70508
rect 7515 70468 7656 70496
rect 7515 70465 7527 70468
rect 7469 70459 7527 70465
rect 7650 70456 7656 70468
rect 7708 70456 7714 70508
rect 7929 70499 7987 70505
rect 7929 70465 7941 70499
rect 7975 70465 7987 70499
rect 7929 70459 7987 70465
rect 8021 70502 8079 70508
rect 8021 70468 8033 70502
rect 8067 70468 8079 70502
rect 8021 70462 8079 70468
rect 8113 70499 8171 70505
rect 8113 70465 8125 70499
rect 8159 70465 8171 70499
rect 8113 70459 8171 70465
rect 6236 70264 7328 70292
rect 6236 70252 6242 70264
rect 7650 70252 7656 70304
rect 7708 70252 7714 70304
rect 7943 70292 7971 70459
rect 8018 70320 8024 70372
rect 8076 70360 8082 70372
rect 8128 70360 8156 70459
rect 8202 70456 8208 70508
rect 8260 70456 8266 70508
rect 8297 70499 8355 70505
rect 8297 70465 8309 70499
rect 8343 70496 8355 70499
rect 8386 70496 8392 70508
rect 8343 70468 8392 70496
rect 8343 70465 8355 70468
rect 8297 70459 8355 70465
rect 8386 70456 8392 70468
rect 8444 70456 8450 70508
rect 8570 70456 8576 70508
rect 8628 70456 8634 70508
rect 8680 70496 8708 70536
rect 9398 70524 9404 70576
rect 9456 70564 9462 70576
rect 11422 70564 11428 70576
rect 9456 70536 11428 70564
rect 9456 70524 9462 70536
rect 11422 70524 11428 70536
rect 11480 70524 11486 70576
rect 8680 70468 9076 70496
rect 9048 70428 9076 70468
rect 9214 70456 9220 70508
rect 9272 70496 9278 70508
rect 11330 70496 11336 70508
rect 9272 70468 9444 70496
rect 9272 70456 9278 70468
rect 9416 70437 9444 70468
rect 9508 70468 11336 70496
rect 9309 70431 9367 70437
rect 9309 70428 9321 70431
rect 8076 70332 8156 70360
rect 8772 70400 8984 70428
rect 9048 70400 9321 70428
rect 8076 70320 8082 70332
rect 8772 70292 8800 70400
rect 8956 70360 8984 70400
rect 9309 70397 9321 70400
rect 9355 70397 9367 70431
rect 9309 70391 9367 70397
rect 9401 70431 9459 70437
rect 9401 70397 9413 70431
rect 9447 70397 9459 70431
rect 9401 70391 9459 70397
rect 9508 70360 9536 70468
rect 11330 70456 11336 70468
rect 11388 70456 11394 70508
rect 8956 70332 9536 70360
rect 9582 70320 9588 70372
rect 9640 70360 9646 70372
rect 11514 70360 11520 70372
rect 9640 70332 11520 70360
rect 9640 70320 9646 70332
rect 11514 70320 11520 70332
rect 11572 70320 11578 70372
rect 7943 70264 8800 70292
rect 1104 70202 9936 70224
rect 1104 70150 3610 70202
rect 3662 70150 3674 70202
rect 3726 70150 3738 70202
rect 3790 70150 3802 70202
rect 3854 70150 3866 70202
rect 3918 70150 5210 70202
rect 5262 70150 5274 70202
rect 5326 70150 5338 70202
rect 5390 70150 5402 70202
rect 5454 70150 5466 70202
rect 5518 70150 6810 70202
rect 6862 70150 6874 70202
rect 6926 70150 6938 70202
rect 6990 70150 7002 70202
rect 7054 70150 7066 70202
rect 7118 70150 8410 70202
rect 8462 70150 8474 70202
rect 8526 70150 8538 70202
rect 8590 70150 8602 70202
rect 8654 70150 8666 70202
rect 8718 70150 9936 70202
rect 1104 70128 9936 70150
rect 4982 70048 4988 70100
rect 5040 70088 5046 70100
rect 5166 70088 5172 70100
rect 5040 70060 5172 70088
rect 5040 70048 5046 70060
rect 5166 70048 5172 70060
rect 5224 70048 5230 70100
rect 5718 70048 5724 70100
rect 5776 70048 5782 70100
rect 6178 70048 6184 70100
rect 6236 70048 6242 70100
rect 6362 70048 6368 70100
rect 6420 70088 6426 70100
rect 6914 70088 6920 70100
rect 6420 70060 6920 70088
rect 6420 70048 6426 70060
rect 6914 70048 6920 70060
rect 6972 70048 6978 70100
rect 7009 70091 7067 70097
rect 7009 70057 7021 70091
rect 7055 70088 7067 70091
rect 9030 70088 9036 70100
rect 7055 70060 9036 70088
rect 7055 70057 7067 70060
rect 7009 70051 7067 70057
rect 9030 70048 9036 70060
rect 9088 70088 9094 70100
rect 9217 70091 9275 70097
rect 9088 70060 9168 70088
rect 9088 70048 9094 70060
rect 5905 70023 5963 70029
rect 4632 69992 5672 70020
rect 4632 69964 4660 69992
rect 4614 69912 4620 69964
rect 4672 69912 4678 69964
rect 5644 69961 5672 69992
rect 5905 69989 5917 70023
rect 5951 70020 5963 70023
rect 6196 70020 6224 70048
rect 5951 69992 6224 70020
rect 6549 70023 6607 70029
rect 5951 69989 5963 69992
rect 5905 69983 5963 69989
rect 6549 69989 6561 70023
rect 6595 70020 6607 70023
rect 7190 70020 7196 70032
rect 6595 69992 7196 70020
rect 6595 69989 6607 69992
rect 6549 69983 6607 69989
rect 7190 69980 7196 69992
rect 7248 69980 7254 70032
rect 7282 69980 7288 70032
rect 7340 69980 7346 70032
rect 7484 69992 8156 70020
rect 5629 69955 5687 69961
rect 5629 69921 5641 69955
rect 5675 69921 5687 69955
rect 5629 69915 5687 69921
rect 6178 69912 6184 69964
rect 6236 69952 6242 69964
rect 6273 69955 6331 69961
rect 6273 69952 6285 69955
rect 6236 69924 6285 69952
rect 6236 69912 6242 69924
rect 6273 69921 6285 69924
rect 6319 69921 6331 69955
rect 6273 69915 6331 69921
rect 6822 69912 6828 69964
rect 6880 69952 6886 69964
rect 7300 69952 7328 69980
rect 6880 69924 7328 69952
rect 6880 69912 6886 69924
rect 5353 69887 5411 69893
rect 5353 69884 5365 69887
rect 4264 69856 5365 69884
rect 4264 69828 4292 69856
rect 5353 69853 5365 69856
rect 5399 69853 5411 69887
rect 5353 69847 5411 69853
rect 5442 69844 5448 69896
rect 5500 69884 5506 69896
rect 5986 69889 6044 69895
rect 5986 69886 5998 69889
rect 5828 69884 5998 69886
rect 5500 69858 5998 69884
rect 5500 69856 5856 69858
rect 5500 69844 5506 69856
rect 5986 69855 5998 69858
rect 6032 69855 6044 69889
rect 5986 69849 6044 69855
rect 6641 69887 6699 69893
rect 6641 69853 6653 69887
rect 6687 69853 6699 69887
rect 6641 69847 6699 69853
rect 7009 69887 7067 69893
rect 7009 69853 7021 69887
rect 7055 69884 7067 69887
rect 7190 69884 7196 69896
rect 7055 69856 7196 69884
rect 7055 69853 7067 69856
rect 7009 69847 7067 69853
rect 4246 69776 4252 69828
rect 4304 69776 4310 69828
rect 4706 69776 4712 69828
rect 4764 69816 4770 69828
rect 4982 69816 4988 69828
rect 4764 69788 4988 69816
rect 4764 69776 4770 69788
rect 4982 69776 4988 69788
rect 5040 69776 5046 69828
rect 6656 69816 6684 69847
rect 7190 69844 7196 69856
rect 7248 69844 7254 69896
rect 7282 69844 7288 69896
rect 7340 69844 7346 69896
rect 7374 69844 7380 69896
rect 7432 69884 7438 69896
rect 7484 69893 7512 69992
rect 7926 69952 7932 69964
rect 7576 69924 7932 69952
rect 7576 69893 7604 69924
rect 7926 69912 7932 69924
rect 7984 69912 7990 69964
rect 8128 69893 8156 69992
rect 8202 69980 8208 70032
rect 8260 70020 8266 70032
rect 8260 69992 8340 70020
rect 8260 69980 8266 69992
rect 8312 69893 8340 69992
rect 8386 69980 8392 70032
rect 8444 69980 8450 70032
rect 9140 70020 9168 70060
rect 9217 70057 9229 70091
rect 9263 70088 9275 70091
rect 9306 70088 9312 70100
rect 9263 70060 9312 70088
rect 9263 70057 9275 70060
rect 9217 70051 9275 70057
rect 9306 70048 9312 70060
rect 9364 70048 9370 70100
rect 9582 70048 9588 70100
rect 9640 70048 9646 70100
rect 9600 70020 9628 70048
rect 9140 69992 9628 70020
rect 8404 69893 8432 69980
rect 8662 69912 8668 69964
rect 8720 69952 8726 69964
rect 9214 69952 9220 69964
rect 8720 69924 9220 69952
rect 8720 69912 8726 69924
rect 9214 69912 9220 69924
rect 9272 69912 9278 69964
rect 9674 69912 9680 69964
rect 9732 69952 9738 69964
rect 10870 69952 10876 69964
rect 9732 69924 10876 69952
rect 9732 69912 9738 69924
rect 10870 69912 10876 69924
rect 10928 69912 10934 69964
rect 7469 69887 7527 69893
rect 7469 69884 7481 69887
rect 7432 69856 7481 69884
rect 7432 69844 7438 69856
rect 7469 69853 7481 69856
rect 7515 69853 7527 69887
rect 7469 69847 7527 69853
rect 7561 69887 7619 69893
rect 7561 69853 7573 69887
rect 7607 69853 7619 69887
rect 7561 69847 7619 69853
rect 7745 69887 7803 69893
rect 7745 69853 7757 69887
rect 7791 69853 7803 69887
rect 7745 69847 7803 69853
rect 7837 69887 7895 69893
rect 7837 69853 7849 69887
rect 7883 69853 7895 69887
rect 7837 69847 7895 69853
rect 8113 69887 8171 69893
rect 8113 69853 8125 69887
rect 8159 69853 8171 69887
rect 8113 69847 8171 69853
rect 8278 69887 8340 69893
rect 8278 69853 8290 69887
rect 8324 69856 8340 69887
rect 8389 69887 8447 69893
rect 8324 69853 8336 69856
rect 8278 69847 8336 69853
rect 8389 69853 8401 69887
rect 8435 69853 8447 69887
rect 8389 69847 8447 69853
rect 6288 69788 6684 69816
rect 6288 69760 6316 69788
rect 6730 69776 6736 69828
rect 6788 69816 6794 69828
rect 7760 69816 7788 69847
rect 6788 69788 7788 69816
rect 6788 69776 6794 69788
rect 7116 69760 7144 69788
rect 5442 69708 5448 69760
rect 5500 69748 5506 69760
rect 6086 69748 6092 69760
rect 5500 69720 6092 69748
rect 5500 69708 5506 69720
rect 6086 69708 6092 69720
rect 6144 69708 6150 69760
rect 6270 69708 6276 69760
rect 6328 69708 6334 69760
rect 7098 69708 7104 69760
rect 7156 69708 7162 69760
rect 7193 69751 7251 69757
rect 7193 69717 7205 69751
rect 7239 69748 7251 69751
rect 7742 69748 7748 69760
rect 7239 69720 7748 69748
rect 7239 69717 7251 69720
rect 7193 69711 7251 69717
rect 7742 69708 7748 69720
rect 7800 69708 7806 69760
rect 7852 69748 7880 69847
rect 8478 69844 8484 69896
rect 8536 69893 8542 69896
rect 8536 69887 8549 69893
rect 8537 69884 8549 69887
rect 8537 69856 8581 69884
rect 8537 69853 8549 69856
rect 8536 69847 8549 69853
rect 8536 69844 8542 69847
rect 7929 69819 7987 69825
rect 7929 69785 7941 69819
rect 7975 69816 7987 69819
rect 9674 69816 9680 69828
rect 7975 69788 9680 69816
rect 7975 69785 7987 69788
rect 7929 69779 7987 69785
rect 9674 69776 9680 69788
rect 9732 69776 9738 69828
rect 8478 69748 8484 69760
rect 7852 69720 8484 69748
rect 8478 69708 8484 69720
rect 8536 69748 8542 69760
rect 9214 69748 9220 69760
rect 8536 69720 9220 69748
rect 8536 69708 8542 69720
rect 9214 69708 9220 69720
rect 9272 69708 9278 69760
rect 9582 69708 9588 69760
rect 9640 69748 9646 69760
rect 10962 69748 10968 69760
rect 9640 69720 10968 69748
rect 9640 69708 9646 69720
rect 10962 69708 10968 69720
rect 11020 69708 11026 69760
rect 1104 69658 9936 69680
rect 1104 69606 2950 69658
rect 3002 69606 3014 69658
rect 3066 69606 3078 69658
rect 3130 69606 3142 69658
rect 3194 69606 3206 69658
rect 3258 69606 4550 69658
rect 4602 69606 4614 69658
rect 4666 69606 4678 69658
rect 4730 69606 4742 69658
rect 4794 69606 4806 69658
rect 4858 69606 6150 69658
rect 6202 69606 6214 69658
rect 6266 69606 6278 69658
rect 6330 69606 6342 69658
rect 6394 69606 6406 69658
rect 6458 69606 7750 69658
rect 7802 69606 7814 69658
rect 7866 69606 7878 69658
rect 7930 69606 7942 69658
rect 7994 69606 8006 69658
rect 8058 69606 9350 69658
rect 9402 69606 9414 69658
rect 9466 69606 9478 69658
rect 9530 69606 9542 69658
rect 9594 69606 9606 69658
rect 9658 69606 9936 69658
rect 1104 69584 9936 69606
rect 4338 69504 4344 69556
rect 4396 69504 4402 69556
rect 4798 69504 4804 69556
rect 4856 69544 4862 69556
rect 5166 69544 5172 69556
rect 4856 69516 5172 69544
rect 4856 69504 4862 69516
rect 5166 69504 5172 69516
rect 5224 69504 5230 69556
rect 6546 69504 6552 69556
rect 6604 69544 6610 69556
rect 6733 69547 6791 69553
rect 6733 69544 6745 69547
rect 6604 69516 6745 69544
rect 6604 69504 6610 69516
rect 6733 69513 6745 69516
rect 6779 69513 6791 69547
rect 6733 69507 6791 69513
rect 6822 69504 6828 69556
rect 6880 69504 6886 69556
rect 6914 69504 6920 69556
rect 6972 69544 6978 69556
rect 7742 69544 7748 69556
rect 6972 69516 7748 69544
rect 6972 69504 6978 69516
rect 7742 69504 7748 69516
rect 7800 69504 7806 69556
rect 8389 69547 8447 69553
rect 8389 69513 8401 69547
rect 8435 69544 8447 69547
rect 8754 69544 8760 69556
rect 8435 69516 8760 69544
rect 8435 69513 8447 69516
rect 8389 69507 8447 69513
rect 8754 69504 8760 69516
rect 8812 69544 8818 69556
rect 10778 69544 10784 69556
rect 8812 69516 10784 69544
rect 8812 69504 8818 69516
rect 10778 69504 10784 69516
rect 10836 69504 10842 69556
rect 4356 69476 4384 69504
rect 7561 69479 7619 69485
rect 7561 69476 7573 69479
rect 4356 69448 7573 69476
rect 7561 69445 7573 69448
rect 7607 69476 7619 69479
rect 8018 69476 8024 69488
rect 7607 69448 8024 69476
rect 7607 69445 7619 69448
rect 7561 69439 7619 69445
rect 8018 69436 8024 69448
rect 8076 69476 8082 69488
rect 8202 69476 8208 69488
rect 8076 69448 8208 69476
rect 8076 69436 8082 69448
rect 8202 69436 8208 69448
rect 8260 69436 8266 69488
rect 8481 69479 8539 69485
rect 8481 69445 8493 69479
rect 8527 69476 8539 69479
rect 8570 69476 8576 69488
rect 8527 69448 8576 69476
rect 8527 69445 8539 69448
rect 8481 69439 8539 69445
rect 8570 69436 8576 69448
rect 8628 69476 8634 69488
rect 8628 69448 9674 69476
rect 8628 69436 8634 69448
rect 934 69368 940 69420
rect 992 69408 998 69420
rect 1489 69411 1547 69417
rect 1489 69408 1501 69411
rect 992 69380 1501 69408
rect 992 69368 998 69380
rect 1489 69377 1501 69380
rect 1535 69377 1547 69411
rect 1489 69371 1547 69377
rect 1578 69368 1584 69420
rect 1636 69408 1642 69420
rect 6362 69408 6368 69420
rect 1636 69380 6368 69408
rect 1636 69368 1642 69380
rect 6362 69368 6368 69380
rect 6420 69368 6426 69420
rect 7098 69408 7104 69420
rect 6472 69380 7104 69408
rect 1673 69275 1731 69281
rect 1673 69241 1685 69275
rect 1719 69272 1731 69275
rect 2130 69272 2136 69284
rect 1719 69244 2136 69272
rect 1719 69241 1731 69244
rect 1673 69235 1731 69241
rect 2130 69232 2136 69244
rect 2188 69232 2194 69284
rect 6472 69272 6500 69380
rect 7098 69368 7104 69380
rect 7156 69408 7162 69420
rect 7156 69380 7333 69408
rect 7156 69368 7162 69380
rect 6914 69300 6920 69352
rect 6972 69300 6978 69352
rect 7305 69340 7333 69380
rect 7374 69368 7380 69420
rect 7432 69408 7438 69420
rect 9033 69411 9091 69417
rect 9033 69408 9045 69411
rect 7432 69380 9045 69408
rect 7432 69368 7438 69380
rect 9033 69377 9045 69380
rect 9079 69377 9091 69411
rect 9033 69371 9091 69377
rect 9122 69368 9128 69420
rect 9180 69368 9186 69420
rect 9306 69368 9312 69420
rect 9364 69368 9370 69420
rect 9398 69368 9404 69420
rect 9456 69368 9462 69420
rect 9646 69408 9674 69448
rect 9950 69408 9956 69420
rect 9646 69380 9956 69408
rect 9950 69368 9956 69380
rect 10008 69368 10014 69420
rect 7926 69340 7932 69352
rect 7305 69312 7932 69340
rect 7926 69300 7932 69312
rect 7984 69340 7990 69352
rect 8386 69340 8392 69352
rect 7984 69312 8392 69340
rect 7984 69300 7990 69312
rect 8386 69300 8392 69312
rect 8444 69300 8450 69352
rect 8573 69343 8631 69349
rect 8573 69309 8585 69343
rect 8619 69309 8631 69343
rect 8573 69303 8631 69309
rect 4632 69244 6500 69272
rect 4632 69216 4660 69244
rect 6546 69232 6552 69284
rect 6604 69272 6610 69284
rect 8588 69272 8616 69303
rect 6604 69244 8064 69272
rect 8588 69244 9076 69272
rect 6604 69232 6610 69244
rect 4614 69164 4620 69216
rect 4672 69164 4678 69216
rect 4706 69164 4712 69216
rect 4764 69204 4770 69216
rect 5442 69204 5448 69216
rect 4764 69176 5448 69204
rect 4764 69164 4770 69176
rect 5442 69164 5448 69176
rect 5500 69164 5506 69216
rect 6086 69164 6092 69216
rect 6144 69204 6150 69216
rect 6365 69207 6423 69213
rect 6365 69204 6377 69207
rect 6144 69176 6377 69204
rect 6144 69164 6150 69176
rect 6365 69173 6377 69176
rect 6411 69173 6423 69207
rect 6365 69167 6423 69173
rect 6454 69164 6460 69216
rect 6512 69204 6518 69216
rect 6914 69204 6920 69216
rect 6512 69176 6920 69204
rect 6512 69164 6518 69176
rect 6914 69164 6920 69176
rect 6972 69164 6978 69216
rect 8036 69213 8064 69244
rect 9048 69216 9076 69244
rect 8021 69207 8079 69213
rect 8021 69173 8033 69207
rect 8067 69173 8079 69207
rect 8021 69167 8079 69173
rect 8202 69164 8208 69216
rect 8260 69204 8266 69216
rect 8849 69207 8907 69213
rect 8849 69204 8861 69207
rect 8260 69176 8861 69204
rect 8260 69164 8266 69176
rect 8849 69173 8861 69176
rect 8895 69173 8907 69207
rect 8849 69167 8907 69173
rect 9030 69164 9036 69216
rect 9088 69164 9094 69216
rect 1104 69114 9936 69136
rect 1104 69062 3610 69114
rect 3662 69062 3674 69114
rect 3726 69062 3738 69114
rect 3790 69062 3802 69114
rect 3854 69062 3866 69114
rect 3918 69062 5210 69114
rect 5262 69062 5274 69114
rect 5326 69062 5338 69114
rect 5390 69062 5402 69114
rect 5454 69062 5466 69114
rect 5518 69062 6810 69114
rect 6862 69062 6874 69114
rect 6926 69062 6938 69114
rect 6990 69062 7002 69114
rect 7054 69062 7066 69114
rect 7118 69062 8410 69114
rect 8462 69062 8474 69114
rect 8526 69062 8538 69114
rect 8590 69062 8602 69114
rect 8654 69062 8666 69114
rect 8718 69062 9936 69114
rect 1104 69040 9936 69062
rect 4246 68960 4252 69012
rect 4304 68960 4310 69012
rect 4338 68960 4344 69012
rect 4396 69000 4402 69012
rect 7193 69003 7251 69009
rect 7193 69000 7205 69003
rect 4396 68972 7205 69000
rect 4396 68960 4402 68972
rect 7193 68969 7205 68972
rect 7239 68969 7251 69003
rect 7558 69000 7564 69012
rect 7193 68963 7251 68969
rect 7297 68972 7564 69000
rect 5350 68892 5356 68944
rect 5408 68932 5414 68944
rect 5721 68935 5779 68941
rect 5721 68932 5733 68935
rect 5408 68904 5733 68932
rect 5408 68892 5414 68904
rect 5721 68901 5733 68904
rect 5767 68901 5779 68935
rect 5721 68895 5779 68901
rect 5902 68892 5908 68944
rect 5960 68892 5966 68944
rect 7006 68892 7012 68944
rect 7064 68892 7070 68944
rect 7098 68892 7104 68944
rect 7156 68932 7162 68944
rect 7297 68932 7325 68972
rect 7558 68960 7564 68972
rect 7616 68960 7622 69012
rect 8478 68960 8484 69012
rect 8536 69000 8542 69012
rect 9398 69000 9404 69012
rect 8536 68972 9404 69000
rect 8536 68960 8542 68972
rect 9398 68960 9404 68972
rect 9456 68960 9462 69012
rect 8297 68935 8355 68941
rect 8297 68932 8309 68935
rect 7156 68904 7325 68932
rect 7576 68904 8309 68932
rect 7156 68892 7162 68904
rect 3878 68824 3884 68876
rect 3936 68864 3942 68876
rect 5920 68864 5948 68892
rect 6641 68867 6699 68873
rect 3936 68836 4476 68864
rect 5920 68836 6592 68864
rect 3936 68824 3942 68836
rect 4065 68799 4123 68805
rect 4065 68765 4077 68799
rect 4111 68796 4123 68799
rect 4111 68768 4292 68796
rect 4111 68765 4123 68768
rect 4065 68759 4123 68765
rect 4264 68672 4292 68768
rect 4338 68756 4344 68808
rect 4396 68756 4402 68808
rect 4448 68728 4476 68836
rect 4608 68799 4666 68805
rect 4608 68765 4620 68799
rect 4654 68796 4666 68799
rect 5810 68796 5816 68808
rect 4654 68768 5816 68796
rect 4654 68765 4666 68768
rect 4608 68759 4666 68765
rect 5810 68756 5816 68768
rect 5868 68756 5874 68808
rect 6454 68806 6460 68808
rect 6380 68805 6460 68806
rect 6089 68799 6147 68805
rect 6089 68765 6101 68799
rect 6135 68796 6147 68799
rect 6365 68799 6460 68805
rect 6135 68768 6224 68796
rect 6135 68765 6147 68768
rect 6089 68759 6147 68765
rect 4706 68728 4712 68740
rect 4448 68700 4712 68728
rect 4706 68688 4712 68700
rect 4764 68688 4770 68740
rect 4798 68688 4804 68740
rect 4856 68728 4862 68740
rect 5258 68728 5264 68740
rect 4856 68700 5264 68728
rect 4856 68688 4862 68700
rect 5258 68688 5264 68700
rect 5316 68688 5322 68740
rect 4246 68620 4252 68672
rect 4304 68620 4310 68672
rect 4614 68620 4620 68672
rect 4672 68660 4678 68672
rect 5166 68660 5172 68672
rect 4672 68632 5172 68660
rect 4672 68620 4678 68632
rect 5166 68620 5172 68632
rect 5224 68620 5230 68672
rect 5534 68620 5540 68672
rect 5592 68660 5598 68672
rect 6086 68660 6092 68672
rect 5592 68632 6092 68660
rect 5592 68620 5598 68632
rect 6086 68620 6092 68632
rect 6144 68620 6150 68672
rect 6196 68660 6224 68768
rect 6365 68765 6377 68799
rect 6411 68778 6460 68799
rect 6411 68765 6423 68778
rect 6365 68759 6423 68765
rect 6454 68756 6460 68778
rect 6512 68756 6518 68808
rect 6564 68805 6592 68836
rect 6641 68833 6653 68867
rect 6687 68864 6699 68867
rect 7024 68864 7052 68892
rect 6687 68836 7052 68864
rect 6687 68833 6699 68836
rect 6641 68827 6699 68833
rect 6548 68799 6606 68805
rect 6548 68765 6560 68799
rect 6594 68765 6606 68799
rect 6548 68759 6606 68765
rect 6730 68756 6736 68808
rect 6788 68805 6794 68808
rect 6788 68799 6837 68805
rect 6788 68765 6791 68799
rect 6825 68765 6837 68799
rect 6788 68759 6837 68765
rect 6917 68799 6975 68805
rect 6917 68765 6929 68799
rect 6963 68765 6975 68799
rect 6917 68759 6975 68765
rect 6788 68756 6794 68759
rect 6932 68728 6960 68759
rect 7006 68756 7012 68808
rect 7064 68796 7070 68808
rect 7101 68799 7159 68805
rect 7101 68796 7113 68799
rect 7064 68768 7113 68796
rect 7064 68756 7070 68768
rect 7101 68765 7113 68768
rect 7147 68765 7159 68799
rect 7101 68759 7159 68765
rect 7576 68737 7604 68904
rect 8297 68901 8309 68904
rect 8343 68932 8355 68935
rect 8570 68932 8576 68944
rect 8343 68904 8576 68932
rect 8343 68901 8355 68904
rect 8297 68895 8355 68901
rect 8570 68892 8576 68904
rect 8628 68892 8634 68944
rect 7837 68867 7895 68873
rect 7837 68833 7849 68867
rect 7883 68864 7895 68867
rect 9030 68864 9036 68876
rect 7883 68836 9036 68864
rect 7883 68833 7895 68836
rect 7837 68827 7895 68833
rect 9030 68824 9036 68836
rect 9088 68824 9094 68876
rect 8386 68756 8392 68808
rect 8444 68796 8450 68808
rect 8941 68799 8999 68805
rect 8941 68796 8953 68799
rect 8444 68768 8953 68796
rect 8444 68756 8450 68768
rect 8941 68765 8953 68768
rect 8987 68765 8999 68799
rect 8941 68759 8999 68765
rect 7561 68731 7619 68737
rect 7561 68728 7573 68731
rect 6656 68700 7573 68728
rect 6656 68660 6684 68700
rect 7561 68697 7573 68700
rect 7607 68697 7619 68731
rect 7561 68691 7619 68697
rect 7926 68688 7932 68740
rect 7984 68728 7990 68740
rect 9306 68728 9312 68740
rect 7984 68700 9312 68728
rect 7984 68688 7990 68700
rect 9306 68688 9312 68700
rect 9364 68688 9370 68740
rect 6196 68632 6684 68660
rect 6730 68620 6736 68672
rect 6788 68660 6794 68672
rect 7653 68663 7711 68669
rect 7653 68660 7665 68663
rect 6788 68632 7665 68660
rect 6788 68620 6794 68632
rect 7653 68629 7665 68632
rect 7699 68629 7711 68663
rect 7653 68623 7711 68629
rect 8018 68620 8024 68672
rect 8076 68660 8082 68672
rect 8386 68660 8392 68672
rect 8076 68632 8392 68660
rect 8076 68620 8082 68632
rect 8386 68620 8392 68632
rect 8444 68620 8450 68672
rect 9122 68620 9128 68672
rect 9180 68620 9186 68672
rect 1104 68570 9936 68592
rect 1104 68518 2950 68570
rect 3002 68518 3014 68570
rect 3066 68518 3078 68570
rect 3130 68518 3142 68570
rect 3194 68518 3206 68570
rect 3258 68518 4550 68570
rect 4602 68518 4614 68570
rect 4666 68518 4678 68570
rect 4730 68518 4742 68570
rect 4794 68518 4806 68570
rect 4858 68518 6150 68570
rect 6202 68518 6214 68570
rect 6266 68518 6278 68570
rect 6330 68518 6342 68570
rect 6394 68518 6406 68570
rect 6458 68518 7750 68570
rect 7802 68518 7814 68570
rect 7866 68518 7878 68570
rect 7930 68518 7942 68570
rect 7994 68518 8006 68570
rect 8058 68518 9350 68570
rect 9402 68518 9414 68570
rect 9466 68518 9478 68570
rect 9530 68518 9542 68570
rect 9594 68518 9606 68570
rect 9658 68518 9936 68570
rect 1104 68496 9936 68518
rect 4982 68416 4988 68468
rect 5040 68416 5046 68468
rect 5258 68416 5264 68468
rect 5316 68456 5322 68468
rect 6270 68456 6276 68468
rect 5316 68428 6276 68456
rect 5316 68416 5322 68428
rect 6270 68416 6276 68428
rect 6328 68456 6334 68468
rect 6730 68456 6736 68468
rect 6328 68428 6736 68456
rect 6328 68416 6334 68428
rect 6730 68416 6736 68428
rect 6788 68416 6794 68468
rect 7926 68416 7932 68468
rect 7984 68456 7990 68468
rect 8938 68456 8944 68468
rect 7984 68428 8944 68456
rect 7984 68416 7990 68428
rect 8938 68416 8944 68428
rect 8996 68416 9002 68468
rect 5074 68348 5080 68400
rect 5132 68388 5138 68400
rect 5132 68360 5212 68388
rect 5132 68348 5138 68360
rect 934 68280 940 68332
rect 992 68320 998 68332
rect 1489 68323 1547 68329
rect 1489 68320 1501 68323
rect 992 68292 1501 68320
rect 992 68280 998 68292
rect 1489 68289 1501 68292
rect 1535 68289 1547 68323
rect 1489 68283 1547 68289
rect 4157 68323 4215 68329
rect 4157 68289 4169 68323
rect 4203 68320 4215 68323
rect 4522 68320 4528 68332
rect 4203 68292 4528 68320
rect 4203 68289 4215 68292
rect 4157 68283 4215 68289
rect 4522 68280 4528 68292
rect 4580 68280 4586 68332
rect 4798 68280 4804 68332
rect 4856 68280 4862 68332
rect 5184 68320 5212 68360
rect 5626 68348 5632 68400
rect 5684 68388 5690 68400
rect 7006 68388 7012 68400
rect 5684 68360 6776 68388
rect 5684 68348 5690 68360
rect 6454 68320 6460 68332
rect 5184 68292 6460 68320
rect 6454 68280 6460 68292
rect 6512 68280 6518 68332
rect 6641 68323 6699 68329
rect 6641 68320 6653 68323
rect 6564 68292 6653 68320
rect 4430 68212 4436 68264
rect 4488 68252 4494 68264
rect 4617 68255 4675 68261
rect 4617 68252 4629 68255
rect 4488 68224 4629 68252
rect 4488 68212 4494 68224
rect 4617 68221 4629 68224
rect 4663 68252 4675 68255
rect 6178 68252 6184 68264
rect 4663 68224 6184 68252
rect 4663 68221 4675 68224
rect 4617 68215 4675 68221
rect 6178 68212 6184 68224
rect 6236 68212 6242 68264
rect 6564 68196 6592 68292
rect 6641 68289 6653 68292
rect 6687 68289 6699 68323
rect 6748 68320 6776 68360
rect 6932 68360 7012 68388
rect 6824 68329 6882 68335
rect 6932 68329 6960 68360
rect 7006 68348 7012 68360
rect 7064 68348 7070 68400
rect 7116 68360 7328 68388
rect 6824 68320 6836 68329
rect 6748 68295 6836 68320
rect 6870 68295 6882 68329
rect 6748 68292 6882 68295
rect 6824 68289 6882 68292
rect 6917 68323 6975 68329
rect 6917 68289 6929 68323
rect 6963 68289 6975 68323
rect 6641 68283 6699 68289
rect 6917 68283 6975 68289
rect 7009 68255 7067 68261
rect 7009 68252 7021 68255
rect 6886 68224 7021 68252
rect 6886 68196 6914 68224
rect 7009 68221 7021 68224
rect 7055 68252 7067 68255
rect 7116 68252 7144 68360
rect 7193 68323 7251 68329
rect 7193 68289 7205 68323
rect 7239 68289 7251 68323
rect 7193 68283 7251 68289
rect 7055 68224 7144 68252
rect 7055 68221 7067 68224
rect 7009 68215 7067 68221
rect 842 68144 848 68196
rect 900 68184 906 68196
rect 900 68156 4752 68184
rect 900 68144 906 68156
rect 290 68076 296 68128
rect 348 68116 354 68128
rect 1581 68119 1639 68125
rect 1581 68116 1593 68119
rect 348 68088 1593 68116
rect 348 68076 354 68088
rect 1581 68085 1593 68088
rect 1627 68085 1639 68119
rect 1581 68079 1639 68085
rect 2498 68076 2504 68128
rect 2556 68116 2562 68128
rect 2866 68116 2872 68128
rect 2556 68088 2872 68116
rect 2556 68076 2562 68088
rect 2866 68076 2872 68088
rect 2924 68076 2930 68128
rect 3878 68076 3884 68128
rect 3936 68116 3942 68128
rect 4430 68116 4436 68128
rect 3936 68088 4436 68116
rect 3936 68076 3942 68088
rect 4430 68076 4436 68088
rect 4488 68076 4494 68128
rect 4724 68116 4752 68156
rect 5350 68144 5356 68196
rect 5408 68184 5414 68196
rect 5718 68184 5724 68196
rect 5408 68156 5724 68184
rect 5408 68144 5414 68156
rect 5718 68144 5724 68156
rect 5776 68144 5782 68196
rect 6546 68144 6552 68196
rect 6604 68144 6610 68196
rect 6822 68144 6828 68196
rect 6880 68156 6914 68196
rect 7208 68184 7236 68283
rect 7300 68252 7328 68360
rect 7374 68280 7380 68332
rect 7432 68320 7438 68332
rect 7745 68323 7803 68329
rect 7745 68320 7757 68323
rect 7432 68292 7757 68320
rect 7432 68280 7438 68292
rect 7745 68289 7757 68292
rect 7791 68289 7803 68323
rect 7745 68283 7803 68289
rect 7926 68280 7932 68332
rect 7984 68280 7990 68332
rect 8018 68280 8024 68332
rect 8076 68280 8082 68332
rect 8297 68323 8355 68329
rect 8297 68289 8309 68323
rect 8343 68320 8355 68323
rect 8938 68320 8944 68332
rect 8343 68292 8944 68320
rect 8343 68289 8355 68292
rect 8297 68283 8355 68289
rect 8938 68280 8944 68292
rect 8996 68320 9002 68332
rect 11882 68320 11888 68332
rect 8996 68292 11888 68320
rect 8996 68280 9002 68292
rect 11882 68280 11888 68292
rect 11940 68280 11946 68332
rect 8113 68255 8171 68261
rect 8113 68252 8125 68255
rect 7300 68224 8125 68252
rect 8113 68221 8125 68224
rect 8159 68221 8171 68255
rect 9122 68252 9128 68264
rect 8113 68215 8171 68221
rect 8404 68224 9128 68252
rect 8404 68184 8432 68224
rect 9122 68212 9128 68224
rect 9180 68252 9186 68264
rect 11790 68252 11796 68264
rect 9180 68224 11796 68252
rect 9180 68212 9186 68224
rect 11790 68212 11796 68224
rect 11848 68212 11854 68264
rect 7208 68156 7788 68184
rect 6880 68144 6886 68156
rect 7285 68119 7343 68125
rect 7285 68116 7297 68119
rect 4724 68088 7297 68116
rect 7285 68085 7297 68088
rect 7331 68085 7343 68119
rect 7760 68116 7788 68156
rect 7943 68156 8432 68184
rect 8481 68187 8539 68193
rect 7943 68116 7971 68156
rect 8481 68153 8493 68187
rect 8527 68184 8539 68187
rect 11514 68184 11520 68196
rect 8527 68156 11520 68184
rect 8527 68153 8539 68156
rect 8481 68147 8539 68153
rect 11514 68144 11520 68156
rect 11572 68144 11578 68196
rect 7760 68088 7971 68116
rect 7285 68079 7343 68085
rect 8018 68076 8024 68128
rect 8076 68116 8082 68128
rect 8386 68116 8392 68128
rect 8076 68088 8392 68116
rect 8076 68076 8082 68088
rect 8386 68076 8392 68088
rect 8444 68076 8450 68128
rect 1104 68026 9936 68048
rect 1104 67974 3610 68026
rect 3662 67974 3674 68026
rect 3726 67974 3738 68026
rect 3790 67974 3802 68026
rect 3854 67974 3866 68026
rect 3918 67974 5210 68026
rect 5262 67974 5274 68026
rect 5326 67974 5338 68026
rect 5390 67974 5402 68026
rect 5454 67974 5466 68026
rect 5518 67974 6810 68026
rect 6862 67974 6874 68026
rect 6926 67974 6938 68026
rect 6990 67974 7002 68026
rect 7054 67974 7066 68026
rect 7118 67974 8410 68026
rect 8462 67974 8474 68026
rect 8526 67974 8538 68026
rect 8590 67974 8602 68026
rect 8654 67974 8666 68026
rect 8718 67974 9936 68026
rect 1104 67952 9936 67974
rect 4890 67872 4896 67924
rect 4948 67912 4954 67924
rect 5074 67912 5080 67924
rect 4948 67884 5080 67912
rect 4948 67872 4954 67884
rect 5074 67872 5080 67884
rect 5132 67872 5138 67924
rect 5258 67872 5264 67924
rect 5316 67872 5322 67924
rect 5350 67872 5356 67924
rect 5408 67912 5414 67924
rect 7926 67912 7932 67924
rect 5408 67884 7932 67912
rect 5408 67872 5414 67884
rect 7926 67872 7932 67884
rect 7984 67872 7990 67924
rect 9030 67872 9036 67924
rect 9088 67872 9094 67924
rect 4246 67804 4252 67856
rect 4304 67844 4310 67856
rect 4801 67847 4859 67853
rect 4801 67844 4813 67847
rect 4304 67816 4813 67844
rect 4304 67804 4310 67816
rect 4801 67813 4813 67816
rect 4847 67813 4859 67847
rect 5276 67844 5304 67872
rect 5902 67844 5908 67856
rect 5276 67816 5908 67844
rect 4801 67807 4859 67813
rect 5902 67804 5908 67816
rect 5960 67804 5966 67856
rect 6825 67847 6883 67853
rect 6825 67813 6837 67847
rect 6871 67844 6883 67847
rect 9048 67844 9076 67872
rect 6871 67816 9076 67844
rect 6871 67813 6883 67816
rect 6825 67807 6883 67813
rect 750 67736 756 67788
rect 808 67776 814 67788
rect 4614 67776 4620 67788
rect 808 67748 4620 67776
rect 808 67736 814 67748
rect 4614 67736 4620 67748
rect 4672 67736 4678 67788
rect 6546 67736 6552 67788
rect 6604 67776 6610 67788
rect 6604 67748 7052 67776
rect 6604 67736 6610 67748
rect 5534 67668 5540 67720
rect 5592 67708 5598 67720
rect 6086 67708 6092 67720
rect 5592 67680 6092 67708
rect 5592 67668 5598 67680
rect 6086 67668 6092 67680
rect 6144 67708 6150 67720
rect 7024 67708 7052 67748
rect 7466 67736 7472 67788
rect 7524 67776 7530 67788
rect 7837 67779 7895 67785
rect 7524 67748 7752 67776
rect 7524 67736 7530 67748
rect 7374 67708 7380 67720
rect 6144 67680 6684 67708
rect 6144 67668 6150 67680
rect 1486 67600 1492 67652
rect 1544 67600 1550 67652
rect 1673 67643 1731 67649
rect 1673 67609 1685 67643
rect 1719 67640 1731 67643
rect 2314 67640 2320 67652
rect 1719 67612 2320 67640
rect 1719 67609 1731 67612
rect 1673 67603 1731 67609
rect 2314 67600 2320 67612
rect 2372 67600 2378 67652
rect 4525 67643 4583 67649
rect 4525 67609 4537 67643
rect 4571 67640 4583 67643
rect 4798 67640 4804 67652
rect 4571 67612 4804 67640
rect 4571 67609 4583 67612
rect 4525 67603 4583 67609
rect 4798 67600 4804 67612
rect 4856 67640 4862 67652
rect 5074 67640 5080 67652
rect 4856 67612 5080 67640
rect 4856 67600 4862 67612
rect 5074 67600 5080 67612
rect 5132 67600 5138 67652
rect 5442 67600 5448 67652
rect 5500 67600 5506 67652
rect 6656 67649 6684 67680
rect 7024 67680 7380 67708
rect 7024 67652 7052 67680
rect 7374 67668 7380 67680
rect 7432 67708 7438 67720
rect 7724 67717 7752 67748
rect 7837 67745 7849 67779
rect 7883 67776 7895 67779
rect 8294 67776 8300 67788
rect 7883 67748 8300 67776
rect 7883 67745 7895 67748
rect 7837 67739 7895 67745
rect 8294 67736 8300 67748
rect 8352 67736 8358 67788
rect 8386 67736 8392 67788
rect 8444 67776 8450 67788
rect 9214 67776 9220 67788
rect 8444 67748 9220 67776
rect 8444 67736 8450 67748
rect 9214 67736 9220 67748
rect 9272 67736 9278 67788
rect 7561 67711 7619 67717
rect 7561 67708 7573 67711
rect 7432 67680 7573 67708
rect 7432 67668 7438 67680
rect 7561 67677 7573 67680
rect 7607 67677 7619 67711
rect 7561 67671 7619 67677
rect 7709 67711 7767 67717
rect 7709 67677 7721 67711
rect 7755 67677 7767 67711
rect 7709 67671 7767 67677
rect 7929 67711 7987 67717
rect 7929 67677 7941 67711
rect 7975 67677 7987 67711
rect 7929 67671 7987 67677
rect 8113 67711 8171 67717
rect 8113 67677 8125 67711
rect 8159 67708 8171 67711
rect 8754 67708 8760 67720
rect 8159 67680 8760 67708
rect 8159 67677 8171 67680
rect 8113 67671 8171 67677
rect 6641 67643 6699 67649
rect 6641 67609 6653 67643
rect 6687 67640 6699 67643
rect 6914 67640 6920 67652
rect 6687 67612 6920 67640
rect 6687 67609 6699 67612
rect 6641 67603 6699 67609
rect 6914 67600 6920 67612
rect 6972 67600 6978 67652
rect 7006 67600 7012 67652
rect 7064 67600 7070 67652
rect 7098 67600 7104 67652
rect 7156 67640 7162 67652
rect 7944 67640 7972 67671
rect 8754 67668 8760 67680
rect 8812 67668 8818 67720
rect 7156 67612 7972 67640
rect 8297 67643 8355 67649
rect 7156 67600 7162 67612
rect 8297 67609 8309 67643
rect 8343 67640 8355 67643
rect 10778 67640 10784 67652
rect 8343 67612 10784 67640
rect 8343 67609 8355 67612
rect 8297 67603 8355 67609
rect 10778 67600 10784 67612
rect 10836 67600 10842 67652
rect 4985 67575 5043 67581
rect 4985 67541 4997 67575
rect 5031 67572 5043 67575
rect 5460 67572 5488 67600
rect 8570 67572 8576 67584
rect 5031 67544 8576 67572
rect 5031 67541 5043 67544
rect 4985 67535 5043 67541
rect 8570 67532 8576 67544
rect 8628 67532 8634 67584
rect 1104 67482 9936 67504
rect 1104 67430 2950 67482
rect 3002 67430 3014 67482
rect 3066 67430 3078 67482
rect 3130 67430 3142 67482
rect 3194 67430 3206 67482
rect 3258 67430 4550 67482
rect 4602 67430 4614 67482
rect 4666 67430 4678 67482
rect 4730 67430 4742 67482
rect 4794 67430 4806 67482
rect 4858 67430 6150 67482
rect 6202 67430 6214 67482
rect 6266 67430 6278 67482
rect 6330 67430 6342 67482
rect 6394 67430 6406 67482
rect 6458 67430 7750 67482
rect 7802 67430 7814 67482
rect 7866 67430 7878 67482
rect 7930 67430 7942 67482
rect 7994 67430 8006 67482
rect 8058 67430 9350 67482
rect 9402 67430 9414 67482
rect 9466 67430 9478 67482
rect 9530 67430 9542 67482
rect 9594 67430 9606 67482
rect 9658 67430 9936 67482
rect 1104 67408 9936 67430
rect 4709 67371 4767 67377
rect 4709 67337 4721 67371
rect 4755 67368 4767 67371
rect 5258 67368 5264 67380
rect 4755 67340 5264 67368
rect 4755 67337 4767 67340
rect 4709 67331 4767 67337
rect 5258 67328 5264 67340
rect 5316 67328 5322 67380
rect 5902 67328 5908 67380
rect 5960 67368 5966 67380
rect 6454 67368 6460 67380
rect 5960 67340 6460 67368
rect 5960 67328 5966 67340
rect 6454 67328 6460 67340
rect 6512 67328 6518 67380
rect 6546 67328 6552 67380
rect 6604 67368 6610 67380
rect 7006 67368 7012 67380
rect 6604 67340 7012 67368
rect 6604 67328 6610 67340
rect 7006 67328 7012 67340
rect 7064 67328 7070 67380
rect 7193 67371 7251 67377
rect 7193 67337 7205 67371
rect 7239 67368 7251 67371
rect 8665 67371 8723 67377
rect 8665 67368 8677 67371
rect 7239 67340 7333 67368
rect 7239 67337 7251 67340
rect 7193 67331 7251 67337
rect 4338 67260 4344 67312
rect 4396 67300 4402 67312
rect 4396 67272 6960 67300
rect 4396 67260 4402 67272
rect 3878 67192 3884 67244
rect 3936 67232 3942 67244
rect 4614 67232 4620 67244
rect 3936 67204 4620 67232
rect 3936 67192 3942 67204
rect 4614 67192 4620 67204
rect 4672 67232 4678 67244
rect 4801 67235 4859 67241
rect 4801 67232 4813 67235
rect 4672 67204 4813 67232
rect 4672 67192 4678 67204
rect 4801 67201 4813 67204
rect 4847 67201 4859 67235
rect 5057 67235 5115 67241
rect 5057 67232 5069 67235
rect 4801 67195 4859 67201
rect 4908 67204 5069 67232
rect 4246 67124 4252 67176
rect 4304 67124 4310 67176
rect 4706 67124 4712 67176
rect 4764 67164 4770 67176
rect 4908 67164 4936 67204
rect 5057 67201 5069 67204
rect 5103 67232 5115 67235
rect 5350 67232 5356 67244
rect 5103 67204 5356 67232
rect 5103 67201 5115 67204
rect 5057 67195 5115 67201
rect 5350 67192 5356 67204
rect 5408 67192 5414 67244
rect 6932 67241 6960 67272
rect 6641 67235 6699 67241
rect 6641 67232 6653 67235
rect 6104 67204 6653 67232
rect 6104 67176 6132 67204
rect 6641 67201 6653 67204
rect 6687 67201 6699 67235
rect 6641 67195 6699 67201
rect 6917 67235 6975 67241
rect 6917 67201 6929 67235
rect 6963 67232 6975 67235
rect 7190 67232 7196 67244
rect 6963 67204 7196 67232
rect 6963 67201 6975 67204
rect 6917 67195 6975 67201
rect 7190 67192 7196 67204
rect 7248 67192 7254 67244
rect 4764 67136 4936 67164
rect 4764 67124 4770 67136
rect 6086 67124 6092 67176
rect 6144 67124 6150 67176
rect 6730 67124 6736 67176
rect 6788 67124 6794 67176
rect 7305 67164 7333 67340
rect 7392 67340 8677 67368
rect 7392 67312 7420 67340
rect 8665 67337 8677 67340
rect 8711 67337 8723 67371
rect 8665 67331 8723 67337
rect 9033 67371 9091 67377
rect 9033 67337 9045 67371
rect 9079 67368 9091 67371
rect 9122 67368 9128 67380
rect 9079 67340 9128 67368
rect 9079 67337 9091 67340
rect 9033 67331 9091 67337
rect 9122 67328 9128 67340
rect 9180 67328 9186 67380
rect 10318 67328 10324 67380
rect 10376 67328 10382 67380
rect 7374 67260 7380 67312
rect 7432 67260 7438 67312
rect 8205 67303 8263 67309
rect 8205 67300 8217 67303
rect 7668 67272 8217 67300
rect 7668 67244 7696 67272
rect 8205 67269 8217 67272
rect 8251 67300 8263 67303
rect 10336 67300 10364 67328
rect 8251 67272 10364 67300
rect 8251 67269 8263 67272
rect 8205 67263 8263 67269
rect 7650 67192 7656 67244
rect 7708 67192 7714 67244
rect 7742 67192 7748 67244
rect 7800 67232 7806 67244
rect 8297 67235 8355 67241
rect 8297 67232 8309 67235
rect 7800 67204 8309 67232
rect 7800 67192 7806 67204
rect 8297 67201 8309 67204
rect 8343 67201 8355 67235
rect 8297 67195 8355 67201
rect 8754 67192 8760 67244
rect 8812 67232 8818 67244
rect 10134 67232 10140 67244
rect 8812 67204 10140 67232
rect 8812 67192 8818 67204
rect 10134 67192 10140 67204
rect 10192 67192 10198 67244
rect 7926 67164 7932 67176
rect 7305 67136 7932 67164
rect 7926 67124 7932 67136
rect 7984 67124 7990 67176
rect 8389 67167 8447 67173
rect 8389 67133 8401 67167
rect 8435 67164 8447 67167
rect 8478 67164 8484 67176
rect 8435 67136 8484 67164
rect 8435 67133 8447 67136
rect 8389 67127 8447 67133
rect 8478 67124 8484 67136
rect 8536 67124 8542 67176
rect 9030 67124 9036 67176
rect 9088 67124 9094 67176
rect 9122 67124 9128 67176
rect 9180 67124 9186 67176
rect 9217 67167 9275 67173
rect 9217 67133 9229 67167
rect 9263 67133 9275 67167
rect 9217 67127 9275 67133
rect 4617 67099 4675 67105
rect 4617 67065 4629 67099
rect 4663 67096 4675 67099
rect 4663 67068 4844 67096
rect 4663 67065 4675 67068
rect 4617 67059 4675 67065
rect 4816 67028 4844 67068
rect 5994 67056 6000 67108
rect 6052 67096 6058 67108
rect 6748 67096 6776 67124
rect 7561 67099 7619 67105
rect 6052 67068 6776 67096
rect 7024 67068 7325 67096
rect 6052 67056 6058 67068
rect 5074 67028 5080 67040
rect 4816 67000 5080 67028
rect 5074 66988 5080 67000
rect 5132 66988 5138 67040
rect 5442 66988 5448 67040
rect 5500 67028 5506 67040
rect 5902 67028 5908 67040
rect 5500 67000 5908 67028
rect 5500 66988 5506 67000
rect 5902 66988 5908 67000
rect 5960 66988 5966 67040
rect 6181 67031 6239 67037
rect 6181 66997 6193 67031
rect 6227 67028 6239 67031
rect 6730 67028 6736 67040
rect 6227 67000 6736 67028
rect 6227 66997 6239 67000
rect 6181 66991 6239 66997
rect 6730 66988 6736 67000
rect 6788 66988 6794 67040
rect 7024 67037 7052 67068
rect 7009 67031 7067 67037
rect 7009 66997 7021 67031
rect 7055 66997 7067 67031
rect 7297 67028 7325 67068
rect 7561 67065 7573 67099
rect 7607 67096 7619 67099
rect 7650 67096 7656 67108
rect 7607 67068 7656 67096
rect 7607 67065 7619 67068
rect 7561 67059 7619 67065
rect 7650 67056 7656 67068
rect 7708 67056 7714 67108
rect 7834 67056 7840 67108
rect 7892 67056 7898 67108
rect 9048 67096 9076 67124
rect 9232 67096 9260 67127
rect 9398 67124 9404 67176
rect 9456 67164 9462 67176
rect 9858 67164 9864 67176
rect 9456 67136 9864 67164
rect 9456 67124 9462 67136
rect 9858 67124 9864 67136
rect 9916 67124 9922 67176
rect 9048 67068 9260 67096
rect 9858 67028 9864 67040
rect 7297 67000 9864 67028
rect 7009 66991 7067 66997
rect 9858 66988 9864 67000
rect 9916 67028 9922 67040
rect 10594 67028 10600 67040
rect 9916 67000 10600 67028
rect 9916 66988 9922 67000
rect 10594 66988 10600 67000
rect 10652 66988 10658 67040
rect 1104 66938 9936 66960
rect 1104 66886 3610 66938
rect 3662 66886 3674 66938
rect 3726 66886 3738 66938
rect 3790 66886 3802 66938
rect 3854 66886 3866 66938
rect 3918 66886 5210 66938
rect 5262 66886 5274 66938
rect 5326 66886 5338 66938
rect 5390 66886 5402 66938
rect 5454 66886 5466 66938
rect 5518 66886 6810 66938
rect 6862 66886 6874 66938
rect 6926 66886 6938 66938
rect 6990 66886 7002 66938
rect 7054 66886 7066 66938
rect 7118 66886 8410 66938
rect 8462 66886 8474 66938
rect 8526 66886 8538 66938
rect 8590 66886 8602 66938
rect 8654 66886 8666 66938
rect 8718 66886 9936 66938
rect 1104 66864 9936 66886
rect 1026 66784 1032 66836
rect 1084 66824 1090 66836
rect 8021 66827 8079 66833
rect 1084 66796 7788 66824
rect 1084 66784 1090 66796
rect 4890 66716 4896 66768
rect 4948 66756 4954 66768
rect 5166 66756 5172 66768
rect 4948 66728 5172 66756
rect 4948 66716 4954 66728
rect 5166 66716 5172 66728
rect 5224 66716 5230 66768
rect 5350 66716 5356 66768
rect 5408 66756 5414 66768
rect 5902 66756 5908 66768
rect 5408 66728 5908 66756
rect 5408 66716 5414 66728
rect 5902 66716 5908 66728
rect 5960 66716 5966 66768
rect 7190 66756 7196 66768
rect 6380 66728 7196 66756
rect 1673 66691 1731 66697
rect 1673 66657 1685 66691
rect 1719 66688 1731 66691
rect 4522 66688 4528 66700
rect 1719 66660 4528 66688
rect 1719 66657 1731 66660
rect 1673 66651 1731 66657
rect 4522 66648 4528 66660
rect 4580 66648 4586 66700
rect 6380 66697 6408 66728
rect 7190 66716 7196 66728
rect 7248 66756 7254 66768
rect 7248 66728 7604 66756
rect 7248 66716 7254 66728
rect 6365 66691 6423 66697
rect 6365 66657 6377 66691
rect 6411 66657 6423 66691
rect 6365 66651 6423 66657
rect 6454 66648 6460 66700
rect 6512 66688 6518 66700
rect 7576 66697 7604 66728
rect 7469 66691 7527 66697
rect 7469 66688 7481 66691
rect 6512 66660 7481 66688
rect 6512 66648 6518 66660
rect 7469 66657 7481 66660
rect 7515 66657 7527 66691
rect 7469 66651 7527 66657
rect 7561 66691 7619 66697
rect 7561 66657 7573 66691
rect 7607 66657 7619 66691
rect 7561 66651 7619 66657
rect 3970 66580 3976 66632
rect 4028 66620 4034 66632
rect 5902 66620 5908 66632
rect 4028 66592 5908 66620
rect 4028 66580 4034 66592
rect 5902 66580 5908 66592
rect 5960 66580 5966 66632
rect 6089 66623 6147 66629
rect 6089 66589 6101 66623
rect 6135 66620 6147 66623
rect 7006 66620 7012 66632
rect 6135 66592 7012 66620
rect 6135 66589 6147 66592
rect 6089 66583 6147 66589
rect 7006 66580 7012 66592
rect 7064 66580 7070 66632
rect 7193 66623 7251 66629
rect 7193 66589 7205 66623
rect 7239 66589 7251 66623
rect 7374 66620 7380 66632
rect 7335 66592 7380 66620
rect 7193 66583 7251 66589
rect 934 66512 940 66564
rect 992 66552 998 66564
rect 1489 66555 1547 66561
rect 1489 66552 1501 66555
rect 992 66524 1501 66552
rect 992 66512 998 66524
rect 1489 66521 1501 66524
rect 1535 66521 1547 66555
rect 1489 66515 1547 66521
rect 4246 66512 4252 66564
rect 4304 66552 4310 66564
rect 4801 66555 4859 66561
rect 4801 66552 4813 66555
rect 4304 66524 4813 66552
rect 4304 66512 4310 66524
rect 4801 66521 4813 66524
rect 4847 66521 4859 66555
rect 4801 66515 4859 66521
rect 5258 66512 5264 66564
rect 5316 66552 5322 66564
rect 6178 66552 6184 66564
rect 5316 66524 6184 66552
rect 5316 66512 5322 66524
rect 6178 66512 6184 66524
rect 6236 66512 6242 66564
rect 6546 66512 6552 66564
rect 6604 66552 6610 66564
rect 7208 66552 7236 66583
rect 7374 66580 7380 66592
rect 7432 66580 7438 66632
rect 7760 66629 7788 66796
rect 8021 66793 8033 66827
rect 8067 66824 8079 66827
rect 8478 66824 8484 66836
rect 8067 66796 8484 66824
rect 8067 66793 8079 66796
rect 8021 66787 8079 66793
rect 8478 66784 8484 66796
rect 8536 66784 8542 66836
rect 9214 66784 9220 66836
rect 9272 66824 9278 66836
rect 9272 66796 9536 66824
rect 9272 66784 9278 66796
rect 7926 66716 7932 66768
rect 7984 66756 7990 66768
rect 7984 66728 9444 66756
rect 7984 66716 7990 66728
rect 8110 66648 8116 66700
rect 8168 66688 8174 66700
rect 8570 66688 8576 66700
rect 8168 66660 8576 66688
rect 8168 66648 8174 66660
rect 8570 66648 8576 66660
rect 8628 66648 8634 66700
rect 8665 66691 8723 66697
rect 8665 66657 8677 66691
rect 8711 66688 8723 66691
rect 9030 66688 9036 66700
rect 8711 66660 9036 66688
rect 8711 66657 8723 66660
rect 8665 66651 8723 66657
rect 9030 66648 9036 66660
rect 9088 66648 9094 66700
rect 7745 66623 7803 66629
rect 7745 66589 7757 66623
rect 7791 66620 7803 66623
rect 8389 66623 8447 66629
rect 7791 66592 7880 66620
rect 7791 66589 7803 66592
rect 7745 66583 7803 66589
rect 6604 66524 7236 66552
rect 6604 66512 6610 66524
rect 4430 66444 4436 66496
rect 4488 66484 4494 66496
rect 4893 66487 4951 66493
rect 4893 66484 4905 66487
rect 4488 66456 4905 66484
rect 4488 66444 4494 66456
rect 4893 66453 4905 66456
rect 4939 66484 4951 66487
rect 6086 66484 6092 66496
rect 4939 66456 6092 66484
rect 4939 66453 4951 66456
rect 4893 66447 4951 66453
rect 6086 66444 6092 66456
rect 6144 66444 6150 66496
rect 7190 66444 7196 66496
rect 7248 66484 7254 66496
rect 7742 66484 7748 66496
rect 7248 66456 7748 66484
rect 7248 66444 7254 66456
rect 7742 66444 7748 66456
rect 7800 66444 7806 66496
rect 7852 66484 7880 66592
rect 8389 66589 8401 66623
rect 8435 66620 8447 66623
rect 8938 66620 8944 66632
rect 8435 66592 8944 66620
rect 8435 66589 8447 66592
rect 8389 66583 8447 66589
rect 8938 66580 8944 66592
rect 8996 66580 9002 66632
rect 9214 66629 9220 66632
rect 9197 66623 9220 66629
rect 9197 66589 9209 66623
rect 9197 66583 9220 66589
rect 9214 66580 9220 66583
rect 9272 66580 9278 66632
rect 9306 66580 9312 66632
rect 9364 66580 9370 66632
rect 9416 66629 9444 66728
rect 9401 66623 9459 66629
rect 9401 66589 9413 66623
rect 9447 66589 9459 66623
rect 9401 66583 9459 66589
rect 7929 66555 7987 66561
rect 7929 66521 7941 66555
rect 7975 66552 7987 66555
rect 9508 66552 9536 66796
rect 9582 66580 9588 66632
rect 9640 66580 9646 66632
rect 10686 66580 10692 66632
rect 10744 66580 10750 66632
rect 10704 66552 10732 66580
rect 7975 66524 9076 66552
rect 9508 66524 10732 66552
rect 7975 66521 7987 66524
rect 7929 66515 7987 66521
rect 8386 66484 8392 66496
rect 7852 66456 8392 66484
rect 8386 66444 8392 66456
rect 8444 66444 8450 66496
rect 8481 66487 8539 66493
rect 8481 66453 8493 66487
rect 8527 66484 8539 66487
rect 8754 66484 8760 66496
rect 8527 66456 8760 66484
rect 8527 66453 8539 66456
rect 8481 66447 8539 66453
rect 8754 66444 8760 66456
rect 8812 66444 8818 66496
rect 8938 66444 8944 66496
rect 8996 66444 9002 66496
rect 9048 66484 9076 66524
rect 11422 66484 11428 66496
rect 9048 66456 11428 66484
rect 11422 66444 11428 66456
rect 11480 66444 11486 66496
rect 1104 66394 9936 66416
rect 1104 66342 2950 66394
rect 3002 66342 3014 66394
rect 3066 66342 3078 66394
rect 3130 66342 3142 66394
rect 3194 66342 3206 66394
rect 3258 66342 4550 66394
rect 4602 66342 4614 66394
rect 4666 66342 4678 66394
rect 4730 66342 4742 66394
rect 4794 66342 4806 66394
rect 4858 66342 6150 66394
rect 6202 66342 6214 66394
rect 6266 66342 6278 66394
rect 6330 66342 6342 66394
rect 6394 66342 6406 66394
rect 6458 66342 7750 66394
rect 7802 66342 7814 66394
rect 7866 66342 7878 66394
rect 7930 66342 7942 66394
rect 7994 66342 8006 66394
rect 8058 66342 9350 66394
rect 9402 66342 9414 66394
rect 9466 66342 9478 66394
rect 9530 66342 9542 66394
rect 9594 66342 9606 66394
rect 9658 66342 9936 66394
rect 1104 66320 9936 66342
rect 4338 66240 4344 66292
rect 4396 66280 4402 66292
rect 5534 66280 5540 66292
rect 4396 66252 5540 66280
rect 4396 66240 4402 66252
rect 5534 66240 5540 66252
rect 5592 66240 5598 66292
rect 7009 66283 7067 66289
rect 5644 66252 6040 66280
rect 4982 66172 4988 66224
rect 5040 66212 5046 66224
rect 5644 66212 5672 66252
rect 5040 66184 5672 66212
rect 5040 66172 5046 66184
rect 5718 66172 5724 66224
rect 5776 66212 5782 66224
rect 5905 66215 5963 66221
rect 5905 66212 5917 66215
rect 5776 66184 5917 66212
rect 5776 66172 5782 66184
rect 5905 66181 5917 66184
rect 5951 66181 5963 66215
rect 6012 66212 6040 66252
rect 7009 66249 7021 66283
rect 7055 66280 7067 66283
rect 7650 66280 7656 66292
rect 7055 66252 7656 66280
rect 7055 66249 7067 66252
rect 7009 66243 7067 66249
rect 7650 66240 7656 66252
rect 7708 66280 7714 66292
rect 7834 66280 7840 66292
rect 7708 66252 7840 66280
rect 7708 66240 7714 66252
rect 7834 66240 7840 66252
rect 7892 66240 7898 66292
rect 8018 66240 8024 66292
rect 8076 66280 8082 66292
rect 8113 66283 8171 66289
rect 8113 66280 8125 66283
rect 8076 66252 8125 66280
rect 8076 66240 8082 66252
rect 8113 66249 8125 66252
rect 8159 66249 8171 66283
rect 8113 66243 8171 66249
rect 8386 66240 8392 66292
rect 8444 66280 8450 66292
rect 8481 66283 8539 66289
rect 8481 66280 8493 66283
rect 8444 66252 8493 66280
rect 8444 66240 8450 66252
rect 8481 66249 8493 66252
rect 8527 66249 8539 66283
rect 8481 66243 8539 66249
rect 8662 66240 8668 66292
rect 8720 66280 8726 66292
rect 9122 66280 9128 66292
rect 8720 66252 9128 66280
rect 8720 66240 8726 66252
rect 9122 66240 9128 66252
rect 9180 66240 9186 66292
rect 9306 66240 9312 66292
rect 9364 66280 9370 66292
rect 9858 66280 9864 66292
rect 9364 66252 9864 66280
rect 9364 66240 9370 66252
rect 9858 66240 9864 66252
rect 9916 66240 9922 66292
rect 6012 66184 6592 66212
rect 5905 66175 5963 66181
rect 5166 66144 5172 66156
rect 5000 66116 5172 66144
rect 5000 66088 5028 66116
rect 5166 66104 5172 66116
rect 5224 66104 5230 66156
rect 5350 66104 5356 66156
rect 5408 66104 5414 66156
rect 5810 66104 5816 66156
rect 5868 66104 5874 66156
rect 5994 66104 6000 66156
rect 6052 66104 6058 66156
rect 4982 66036 4988 66088
rect 5040 66036 5046 66088
rect 5258 66036 5264 66088
rect 5316 66076 5322 66088
rect 6012 66076 6040 66104
rect 6089 66079 6147 66085
rect 6089 66076 6101 66079
rect 5316 66048 5856 66076
rect 6012 66048 6101 66076
rect 5316 66036 5322 66048
rect 5828 66020 5856 66048
rect 6089 66045 6101 66048
rect 6135 66076 6147 66079
rect 6270 66076 6276 66088
rect 6135 66048 6276 66076
rect 6135 66045 6147 66048
rect 6089 66039 6147 66045
rect 6270 66036 6276 66048
rect 6328 66036 6334 66088
rect 6564 66076 6592 66184
rect 7926 66172 7932 66224
rect 7984 66212 7990 66224
rect 8573 66215 8631 66221
rect 7984 66184 8432 66212
rect 7984 66172 7990 66184
rect 7282 66144 7288 66156
rect 7243 66116 7288 66144
rect 7282 66104 7288 66116
rect 7340 66104 7346 66156
rect 7433 66150 7491 66156
rect 7433 66116 7445 66150
rect 7479 66116 7491 66150
rect 7433 66110 7491 66116
rect 7448 66076 7476 66110
rect 7834 66104 7840 66156
rect 7892 66104 7898 66156
rect 8036 66119 8294 66147
rect 6564 66048 7476 66076
rect 7558 66036 7564 66088
rect 7616 66036 7622 66088
rect 7653 66079 7711 66085
rect 7653 66045 7665 66079
rect 7699 66045 7711 66079
rect 8036 66076 8064 66119
rect 7653 66039 7711 66045
rect 7944 66048 8064 66076
rect 8266 66088 8294 66119
rect 8266 66048 8300 66088
rect 3970 65968 3976 66020
rect 4028 66008 4034 66020
rect 5445 66011 5503 66017
rect 5445 66008 5457 66011
rect 4028 65980 5457 66008
rect 4028 65968 4034 65980
rect 5445 65977 5457 65980
rect 5491 65977 5503 66011
rect 5445 65971 5503 65977
rect 5810 65968 5816 66020
rect 5868 65968 5874 66020
rect 7668 66008 7696 66039
rect 7944 66008 7972 66048
rect 8294 66036 8300 66048
rect 8352 66036 8358 66088
rect 8404 66076 8432 66184
rect 8573 66181 8585 66215
rect 8619 66212 8631 66215
rect 10962 66212 10968 66224
rect 8619 66184 10968 66212
rect 8619 66181 8631 66184
rect 8573 66175 8631 66181
rect 8846 66144 8852 66156
rect 8680 66116 8852 66144
rect 8680 66076 8708 66116
rect 8846 66104 8852 66116
rect 8904 66104 8910 66156
rect 9030 66104 9036 66156
rect 9088 66104 9094 66156
rect 8404 66048 8708 66076
rect 8757 66079 8815 66085
rect 8757 66045 8769 66079
rect 8803 66076 8815 66079
rect 9048 66076 9076 66104
rect 8803 66048 9076 66076
rect 8803 66045 8815 66048
rect 8757 66039 8815 66045
rect 7668 65980 7972 66008
rect 8021 66011 8079 66017
rect 5169 65943 5227 65949
rect 5169 65909 5181 65943
rect 5215 65940 5227 65943
rect 7006 65940 7012 65952
rect 5215 65912 7012 65940
rect 5215 65909 5227 65912
rect 5169 65903 5227 65909
rect 7006 65900 7012 65912
rect 7064 65940 7070 65952
rect 7724 65940 7752 65980
rect 8021 65977 8033 66011
rect 8067 66008 8079 66011
rect 8067 65980 8248 66008
rect 8067 65977 8079 65980
rect 8021 65971 8079 65977
rect 7064 65912 7752 65940
rect 8220 65940 8248 65980
rect 8386 65968 8392 66020
rect 8444 66008 8450 66020
rect 8846 66008 8852 66020
rect 8444 65980 8852 66008
rect 8444 65968 8450 65980
rect 8846 65968 8852 65980
rect 8904 65968 8910 66020
rect 9030 65968 9036 66020
rect 9088 66008 9094 66020
rect 9646 66008 9674 66184
rect 10962 66172 10968 66184
rect 11020 66172 11026 66224
rect 9088 65980 9674 66008
rect 9088 65968 9094 65980
rect 9858 65940 9864 65952
rect 8220 65912 9864 65940
rect 7064 65900 7070 65912
rect 9858 65900 9864 65912
rect 9916 65900 9922 65952
rect 1104 65850 9936 65872
rect 1104 65798 3610 65850
rect 3662 65798 3674 65850
rect 3726 65798 3738 65850
rect 3790 65798 3802 65850
rect 3854 65798 3866 65850
rect 3918 65798 5210 65850
rect 5262 65798 5274 65850
rect 5326 65798 5338 65850
rect 5390 65798 5402 65850
rect 5454 65798 5466 65850
rect 5518 65798 6810 65850
rect 6862 65798 6874 65850
rect 6926 65798 6938 65850
rect 6990 65798 7002 65850
rect 7054 65798 7066 65850
rect 7118 65798 8410 65850
rect 8462 65798 8474 65850
rect 8526 65798 8538 65850
rect 8590 65798 8602 65850
rect 8654 65798 8666 65850
rect 8718 65798 9936 65850
rect 1104 65776 9936 65798
rect 3326 65736 3332 65748
rect 2332 65708 3332 65736
rect 2332 65532 2360 65708
rect 3326 65696 3332 65708
rect 3384 65696 3390 65748
rect 5537 65739 5595 65745
rect 5537 65705 5549 65739
rect 5583 65736 5595 65739
rect 5626 65736 5632 65748
rect 5583 65708 5632 65736
rect 5583 65705 5595 65708
rect 5537 65699 5595 65705
rect 5626 65696 5632 65708
rect 5684 65736 5690 65748
rect 7098 65736 7104 65748
rect 5684 65708 7104 65736
rect 5684 65696 5690 65708
rect 7098 65696 7104 65708
rect 7156 65696 7162 65748
rect 7466 65696 7472 65748
rect 7524 65696 7530 65748
rect 7558 65696 7564 65748
rect 7616 65736 7622 65748
rect 7926 65736 7932 65748
rect 7616 65708 7932 65736
rect 7616 65696 7622 65708
rect 7926 65696 7932 65708
rect 7984 65696 7990 65748
rect 2406 65628 2412 65680
rect 2464 65668 2470 65680
rect 3602 65668 3608 65680
rect 2464 65640 3608 65668
rect 2464 65628 2470 65640
rect 3602 65628 3608 65640
rect 3660 65628 3666 65680
rect 7484 65668 7512 65696
rect 6923 65640 7512 65668
rect 4890 65560 4896 65612
rect 4948 65600 4954 65612
rect 5718 65600 5724 65612
rect 4948 65572 5724 65600
rect 4948 65560 4954 65572
rect 5718 65560 5724 65572
rect 5776 65600 5782 65612
rect 5905 65603 5963 65609
rect 5905 65600 5917 65603
rect 5776 65572 5917 65600
rect 5776 65560 5782 65572
rect 5905 65569 5917 65572
rect 5951 65569 5963 65603
rect 5905 65563 5963 65569
rect 2406 65532 2412 65544
rect 2332 65504 2412 65532
rect 2406 65492 2412 65504
rect 2464 65492 2470 65544
rect 2682 65492 2688 65544
rect 2740 65532 2746 65544
rect 3510 65532 3516 65544
rect 2740 65504 3516 65532
rect 2740 65492 2746 65504
rect 3510 65492 3516 65504
rect 3568 65492 3574 65544
rect 5994 65492 6000 65544
rect 6052 65532 6058 65544
rect 6923 65532 6951 65640
rect 7282 65560 7288 65612
rect 7340 65600 7346 65612
rect 7466 65600 7472 65612
rect 7340 65572 7472 65600
rect 7340 65560 7346 65572
rect 7466 65560 7472 65572
rect 7524 65560 7530 65612
rect 6052 65504 6951 65532
rect 6052 65492 6058 65504
rect 934 65424 940 65476
rect 992 65464 998 65476
rect 1489 65467 1547 65473
rect 1489 65464 1501 65467
rect 992 65436 1501 65464
rect 992 65424 998 65436
rect 1489 65433 1501 65436
rect 1535 65433 1547 65467
rect 1489 65427 1547 65433
rect 1673 65467 1731 65473
rect 1673 65433 1685 65467
rect 1719 65464 1731 65467
rect 2130 65464 2136 65476
rect 1719 65436 2136 65464
rect 1719 65433 1731 65436
rect 1673 65427 1731 65433
rect 2130 65424 2136 65436
rect 2188 65424 2194 65476
rect 2774 65424 2780 65476
rect 2832 65464 2838 65476
rect 3326 65464 3332 65476
rect 2832 65436 3332 65464
rect 2832 65424 2838 65436
rect 3326 65424 3332 65436
rect 3384 65424 3390 65476
rect 5074 65424 5080 65476
rect 5132 65464 5138 65476
rect 5445 65467 5503 65473
rect 5445 65464 5457 65467
rect 5132 65436 5457 65464
rect 5132 65424 5138 65436
rect 5445 65433 5457 65436
rect 5491 65464 5503 65467
rect 5626 65464 5632 65476
rect 5491 65436 5632 65464
rect 5491 65433 5503 65436
rect 5445 65427 5503 65433
rect 5626 65424 5632 65436
rect 5684 65424 5690 65476
rect 6172 65467 6230 65473
rect 6172 65433 6184 65467
rect 6218 65464 6230 65467
rect 7006 65464 7012 65476
rect 6218 65436 7012 65464
rect 6218 65433 6230 65436
rect 6172 65427 6230 65433
rect 7006 65424 7012 65436
rect 7064 65464 7070 65476
rect 9950 65464 9956 65476
rect 7064 65436 9956 65464
rect 7064 65424 7070 65436
rect 9950 65424 9956 65436
rect 10008 65424 10014 65476
rect 290 65356 296 65408
rect 348 65396 354 65408
rect 1210 65396 1216 65408
rect 348 65368 1216 65396
rect 348 65356 354 65368
rect 1210 65356 1216 65368
rect 1268 65356 1274 65408
rect 4614 65356 4620 65408
rect 4672 65396 4678 65408
rect 5166 65396 5172 65408
rect 4672 65368 5172 65396
rect 4672 65356 4678 65368
rect 5166 65356 5172 65368
rect 5224 65356 5230 65408
rect 6270 65356 6276 65408
rect 6328 65396 6334 65408
rect 6822 65396 6828 65408
rect 6328 65368 6828 65396
rect 6328 65356 6334 65368
rect 6822 65356 6828 65368
rect 6880 65356 6886 65408
rect 7282 65356 7288 65408
rect 7340 65356 7346 65408
rect 7558 65356 7564 65408
rect 7616 65396 7622 65408
rect 8018 65396 8024 65408
rect 7616 65368 8024 65396
rect 7616 65356 7622 65368
rect 8018 65356 8024 65368
rect 8076 65356 8082 65408
rect 8478 65356 8484 65408
rect 8536 65396 8542 65408
rect 9306 65396 9312 65408
rect 8536 65368 9312 65396
rect 8536 65356 8542 65368
rect 9306 65356 9312 65368
rect 9364 65356 9370 65408
rect 1104 65306 9936 65328
rect 1104 65254 2950 65306
rect 3002 65254 3014 65306
rect 3066 65254 3078 65306
rect 3130 65254 3142 65306
rect 3194 65254 3206 65306
rect 3258 65254 4550 65306
rect 4602 65254 4614 65306
rect 4666 65254 4678 65306
rect 4730 65254 4742 65306
rect 4794 65254 4806 65306
rect 4858 65254 6150 65306
rect 6202 65254 6214 65306
rect 6266 65254 6278 65306
rect 6330 65254 6342 65306
rect 6394 65254 6406 65306
rect 6458 65254 7750 65306
rect 7802 65254 7814 65306
rect 7866 65254 7878 65306
rect 7930 65254 7942 65306
rect 7994 65254 8006 65306
rect 8058 65254 9350 65306
rect 9402 65254 9414 65306
rect 9466 65254 9478 65306
rect 9530 65254 9542 65306
rect 9594 65254 9606 65306
rect 9658 65254 9936 65306
rect 10042 65288 10048 65340
rect 10100 65328 10106 65340
rect 10318 65328 10324 65340
rect 10100 65300 10324 65328
rect 10100 65288 10106 65300
rect 10318 65288 10324 65300
rect 10376 65288 10382 65340
rect 1104 65232 9936 65254
rect 5074 65152 5080 65204
rect 5132 65192 5138 65204
rect 8849 65195 8907 65201
rect 8849 65192 8861 65195
rect 5132 65164 8861 65192
rect 5132 65152 5138 65164
rect 8849 65161 8861 65164
rect 8895 65161 8907 65195
rect 8849 65155 8907 65161
rect 9122 65152 9128 65204
rect 9180 65192 9186 65204
rect 9217 65195 9275 65201
rect 9217 65192 9229 65195
rect 9180 65164 9229 65192
rect 9180 65152 9186 65164
rect 9217 65161 9229 65164
rect 9263 65161 9275 65195
rect 9217 65155 9275 65161
rect 2498 65084 2504 65136
rect 2556 65124 2562 65136
rect 4617 65127 4675 65133
rect 2556 65096 2912 65124
rect 2556 65084 2562 65096
rect 2590 65016 2596 65068
rect 2648 65016 2654 65068
rect 2130 64948 2136 65000
rect 2188 64988 2194 65000
rect 2608 64988 2636 65016
rect 2188 64960 2636 64988
rect 2188 64948 2194 64960
rect 2884 64864 2912 65096
rect 4617 65093 4629 65127
rect 4663 65124 4675 65127
rect 8573 65127 8631 65133
rect 4663 65096 7604 65124
rect 4663 65093 4675 65096
rect 4617 65087 4675 65093
rect 4433 65059 4491 65065
rect 4433 65025 4445 65059
rect 4479 65056 4491 65059
rect 4706 65056 4712 65068
rect 4479 65028 4712 65056
rect 4479 65025 4491 65028
rect 4433 65019 4491 65025
rect 4706 65016 4712 65028
rect 4764 65016 4770 65068
rect 5537 65059 5595 65065
rect 5537 65025 5549 65059
rect 5583 65056 5595 65059
rect 6546 65056 6552 65068
rect 5583 65028 6552 65056
rect 5583 65025 5595 65028
rect 5537 65019 5595 65025
rect 6546 65016 6552 65028
rect 6604 65016 6610 65068
rect 7466 65016 7472 65068
rect 7524 65016 7530 65068
rect 3234 64948 3240 65000
rect 3292 64988 3298 65000
rect 4249 64991 4307 64997
rect 4249 64988 4261 64991
rect 3292 64960 4261 64988
rect 3292 64948 3298 64960
rect 4249 64957 4261 64960
rect 4295 64988 4307 64991
rect 5166 64988 5172 65000
rect 4295 64960 5172 64988
rect 4295 64957 4307 64960
rect 4249 64951 4307 64957
rect 5166 64948 5172 64960
rect 5224 64948 5230 65000
rect 5261 64991 5319 64997
rect 5261 64957 5273 64991
rect 5307 64988 5319 64991
rect 7484 64988 7512 65016
rect 5307 64960 7512 64988
rect 7576 64988 7604 65096
rect 7760 65096 8248 65124
rect 7650 65016 7656 65068
rect 7708 65016 7714 65068
rect 7760 65065 7788 65096
rect 8220 65068 8248 65096
rect 8573 65093 8585 65127
rect 8619 65124 8631 65127
rect 9140 65124 9168 65152
rect 8619 65096 9168 65124
rect 8619 65093 8631 65096
rect 8573 65087 8631 65093
rect 7745 65059 7803 65065
rect 7745 65025 7757 65059
rect 7791 65025 7803 65059
rect 7745 65019 7803 65025
rect 8018 65016 8024 65068
rect 8076 65016 8082 65068
rect 8202 65016 8208 65068
rect 8260 65016 8266 65068
rect 8478 65016 8484 65068
rect 8536 65056 8542 65068
rect 8536 65028 9076 65056
rect 8536 65016 8542 65028
rect 9048 65000 9076 65028
rect 9858 65016 9864 65068
rect 9916 65056 9922 65068
rect 10226 65056 10232 65068
rect 9916 65028 10232 65056
rect 9916 65016 9922 65028
rect 10226 65016 10232 65028
rect 10284 65016 10290 65068
rect 7837 64991 7895 64997
rect 7576 64960 7788 64988
rect 5307 64957 5319 64960
rect 5261 64951 5319 64957
rect 5276 64920 5304 64951
rect 5092 64892 5304 64920
rect 5092 64864 5120 64892
rect 5350 64880 5356 64932
rect 5408 64920 5414 64932
rect 6086 64920 6092 64932
rect 5408 64892 6092 64920
rect 5408 64880 5414 64892
rect 6086 64880 6092 64892
rect 6144 64880 6150 64932
rect 7098 64880 7104 64932
rect 7156 64880 7162 64932
rect 7484 64920 7512 64960
rect 7650 64920 7656 64932
rect 7484 64892 7656 64920
rect 7650 64880 7656 64892
rect 7708 64880 7714 64932
rect 2866 64812 2872 64864
rect 2924 64812 2930 64864
rect 4154 64812 4160 64864
rect 4212 64852 4218 64864
rect 4890 64852 4896 64864
rect 4212 64824 4896 64852
rect 4212 64812 4218 64824
rect 4890 64812 4896 64824
rect 4948 64812 4954 64864
rect 5074 64812 5080 64864
rect 5132 64812 5138 64864
rect 6546 64812 6552 64864
rect 6604 64852 6610 64864
rect 6822 64852 6828 64864
rect 6604 64824 6828 64852
rect 6604 64812 6610 64824
rect 6822 64812 6828 64824
rect 6880 64812 6886 64864
rect 7116 64852 7144 64880
rect 7466 64852 7472 64864
rect 7116 64824 7472 64852
rect 7466 64812 7472 64824
rect 7524 64812 7530 64864
rect 7760 64852 7788 64960
rect 7837 64957 7849 64991
rect 7883 64988 7895 64991
rect 8294 64988 8300 65000
rect 7883 64960 8300 64988
rect 7883 64957 7895 64960
rect 7837 64951 7895 64957
rect 8294 64948 8300 64960
rect 8352 64988 8358 65000
rect 8754 64988 8760 65000
rect 8352 64960 8760 64988
rect 8352 64948 8358 64960
rect 8754 64948 8760 64960
rect 8812 64948 8818 65000
rect 9030 64948 9036 65000
rect 9088 64948 9094 65000
rect 9306 64948 9312 65000
rect 9364 64948 9370 65000
rect 9490 64948 9496 65000
rect 9548 64988 9554 65000
rect 11146 64988 11152 65000
rect 9548 64960 11152 64988
rect 9548 64948 9554 64960
rect 11146 64948 11152 64960
rect 11204 64948 11210 65000
rect 8205 64923 8263 64929
rect 8205 64889 8217 64923
rect 8251 64920 8263 64923
rect 10134 64920 10140 64932
rect 8251 64892 10140 64920
rect 8251 64889 8263 64892
rect 8205 64883 8263 64889
rect 10134 64880 10140 64892
rect 10192 64880 10198 64932
rect 9490 64852 9496 64864
rect 7760 64824 9496 64852
rect 9490 64812 9496 64824
rect 9548 64812 9554 64864
rect 1104 64762 9936 64784
rect 1104 64710 3610 64762
rect 3662 64710 3674 64762
rect 3726 64710 3738 64762
rect 3790 64710 3802 64762
rect 3854 64710 3866 64762
rect 3918 64710 5210 64762
rect 5262 64710 5274 64762
rect 5326 64710 5338 64762
rect 5390 64710 5402 64762
rect 5454 64710 5466 64762
rect 5518 64710 6810 64762
rect 6862 64710 6874 64762
rect 6926 64710 6938 64762
rect 6990 64710 7002 64762
rect 7054 64710 7066 64762
rect 7118 64710 8410 64762
rect 8462 64710 8474 64762
rect 8526 64710 8538 64762
rect 8590 64710 8602 64762
rect 8654 64710 8666 64762
rect 8718 64710 9936 64762
rect 1104 64688 9936 64710
rect 2406 64608 2412 64660
rect 2464 64648 2470 64660
rect 2774 64648 2780 64660
rect 2464 64620 2780 64648
rect 2464 64608 2470 64620
rect 2774 64608 2780 64620
rect 2832 64608 2838 64660
rect 4798 64608 4804 64660
rect 4856 64648 4862 64660
rect 5166 64648 5172 64660
rect 4856 64620 5172 64648
rect 4856 64608 4862 64620
rect 5166 64608 5172 64620
rect 5224 64608 5230 64660
rect 4154 64472 4160 64524
rect 4212 64512 4218 64524
rect 5074 64512 5080 64524
rect 4212 64484 5080 64512
rect 4212 64472 4218 64484
rect 5074 64472 5080 64484
rect 5132 64472 5138 64524
rect 5718 64472 5724 64524
rect 5776 64472 5782 64524
rect 7466 64472 7472 64524
rect 7524 64512 7530 64524
rect 8570 64512 8576 64524
rect 7524 64484 8576 64512
rect 7524 64472 7530 64484
rect 8570 64472 8576 64484
rect 8628 64472 8634 64524
rect 8662 64472 8668 64524
rect 8720 64512 8726 64524
rect 9030 64512 9036 64524
rect 8720 64484 9036 64512
rect 8720 64472 8726 64484
rect 9030 64472 9036 64484
rect 9088 64472 9094 64524
rect 2682 64404 2688 64456
rect 2740 64444 2746 64456
rect 3234 64444 3240 64456
rect 2740 64416 3240 64444
rect 2740 64404 2746 64416
rect 3234 64404 3240 64416
rect 3292 64404 3298 64456
rect 5810 64404 5816 64456
rect 5868 64444 5874 64456
rect 5977 64447 6035 64453
rect 5977 64444 5989 64447
rect 5868 64416 5989 64444
rect 5868 64404 5874 64416
rect 5977 64413 5989 64416
rect 6023 64444 6035 64447
rect 7098 64444 7104 64456
rect 6023 64416 7104 64444
rect 6023 64413 6035 64416
rect 5977 64407 6035 64413
rect 7098 64404 7104 64416
rect 7156 64404 7162 64456
rect 8018 64404 8024 64456
rect 8076 64444 8082 64456
rect 8389 64447 8447 64453
rect 8389 64444 8401 64447
rect 8076 64416 8401 64444
rect 8076 64404 8082 64416
rect 8389 64413 8401 64416
rect 8435 64444 8447 64447
rect 10410 64444 10416 64456
rect 8435 64416 10416 64444
rect 8435 64413 8447 64416
rect 8389 64407 8447 64413
rect 10410 64404 10416 64416
rect 10468 64404 10474 64456
rect 934 64336 940 64388
rect 992 64376 998 64388
rect 1489 64379 1547 64385
rect 1489 64376 1501 64379
rect 992 64348 1501 64376
rect 992 64336 998 64348
rect 1489 64345 1501 64348
rect 1535 64345 1547 64379
rect 1489 64339 1547 64345
rect 8481 64379 8539 64385
rect 8481 64345 8493 64379
rect 8527 64376 8539 64379
rect 8846 64376 8852 64388
rect 8527 64348 8852 64376
rect 8527 64345 8539 64348
rect 8481 64339 8539 64345
rect 8846 64336 8852 64348
rect 8904 64376 8910 64388
rect 9030 64376 9036 64388
rect 8904 64348 9036 64376
rect 8904 64336 8910 64348
rect 9030 64336 9036 64348
rect 9088 64336 9094 64388
rect 1578 64268 1584 64320
rect 1636 64268 1642 64320
rect 4706 64268 4712 64320
rect 4764 64308 4770 64320
rect 5074 64308 5080 64320
rect 4764 64280 5080 64308
rect 4764 64268 4770 64280
rect 5074 64268 5080 64280
rect 5132 64268 5138 64320
rect 5810 64268 5816 64320
rect 5868 64308 5874 64320
rect 6086 64308 6092 64320
rect 5868 64280 6092 64308
rect 5868 64268 5874 64280
rect 6086 64268 6092 64280
rect 6144 64268 6150 64320
rect 7101 64311 7159 64317
rect 7101 64277 7113 64311
rect 7147 64308 7159 64311
rect 7558 64308 7564 64320
rect 7147 64280 7564 64308
rect 7147 64277 7159 64280
rect 7101 64271 7159 64277
rect 7558 64268 7564 64280
rect 7616 64268 7622 64320
rect 8018 64268 8024 64320
rect 8076 64268 8082 64320
rect 9122 64268 9128 64320
rect 9180 64308 9186 64320
rect 9858 64308 9864 64320
rect 9180 64280 9864 64308
rect 9180 64268 9186 64280
rect 9858 64268 9864 64280
rect 9916 64268 9922 64320
rect 1104 64218 9936 64240
rect 1104 64166 2950 64218
rect 3002 64166 3014 64218
rect 3066 64166 3078 64218
rect 3130 64166 3142 64218
rect 3194 64166 3206 64218
rect 3258 64166 4550 64218
rect 4602 64166 4614 64218
rect 4666 64166 4678 64218
rect 4730 64166 4742 64218
rect 4794 64166 4806 64218
rect 4858 64166 6150 64218
rect 6202 64166 6214 64218
rect 6266 64166 6278 64218
rect 6330 64166 6342 64218
rect 6394 64166 6406 64218
rect 6458 64166 7750 64218
rect 7802 64166 7814 64218
rect 7866 64166 7878 64218
rect 7930 64166 7942 64218
rect 7994 64166 8006 64218
rect 8058 64166 9350 64218
rect 9402 64166 9414 64218
rect 9466 64166 9478 64218
rect 9530 64166 9542 64218
rect 9594 64166 9606 64218
rect 9658 64166 9936 64218
rect 1104 64144 9936 64166
rect 1578 64064 1584 64116
rect 1636 64104 1642 64116
rect 1636 64076 2774 64104
rect 1636 64064 1642 64076
rect 2746 64036 2774 64076
rect 4798 64064 4804 64116
rect 4856 64104 4862 64116
rect 5166 64104 5172 64116
rect 4856 64076 5172 64104
rect 4856 64064 4862 64076
rect 5166 64064 5172 64076
rect 5224 64064 5230 64116
rect 5810 64064 5816 64116
rect 5868 64104 5874 64116
rect 6270 64104 6276 64116
rect 5868 64076 6276 64104
rect 5868 64064 5874 64076
rect 6270 64064 6276 64076
rect 6328 64064 6334 64116
rect 8205 64107 8263 64113
rect 8205 64073 8217 64107
rect 8251 64104 8263 64107
rect 8846 64104 8852 64116
rect 8251 64076 8852 64104
rect 8251 64073 8263 64076
rect 8205 64067 8263 64073
rect 8846 64064 8852 64076
rect 8904 64104 8910 64116
rect 11698 64104 11704 64116
rect 8904 64076 11704 64104
rect 8904 64064 8910 64076
rect 11698 64064 11704 64076
rect 11756 64064 11762 64116
rect 2746 64008 10640 64036
rect 10612 63980 10640 64008
rect 1486 63928 1492 63980
rect 1544 63928 1550 63980
rect 5718 63928 5724 63980
rect 5776 63968 5782 63980
rect 6086 63968 6092 63980
rect 5776 63940 6092 63968
rect 5776 63928 5782 63940
rect 6086 63928 6092 63940
rect 6144 63968 6150 63980
rect 6457 63971 6515 63977
rect 6457 63968 6469 63971
rect 6144 63940 6469 63968
rect 6144 63928 6150 63940
rect 6457 63937 6469 63940
rect 6503 63937 6515 63971
rect 6457 63931 6515 63937
rect 6724 63971 6782 63977
rect 6724 63937 6736 63971
rect 6770 63968 6782 63971
rect 7190 63968 7196 63980
rect 6770 63940 7196 63968
rect 6770 63937 6782 63940
rect 6724 63931 6782 63937
rect 7190 63928 7196 63940
rect 7248 63968 7254 63980
rect 7742 63968 7748 63980
rect 7248 63940 7748 63968
rect 7248 63928 7254 63940
rect 7742 63928 7748 63940
rect 7800 63928 7806 63980
rect 7926 63928 7932 63980
rect 7984 63968 7990 63980
rect 8294 63968 8300 63980
rect 7984 63940 8300 63968
rect 7984 63928 7990 63940
rect 8294 63928 8300 63940
rect 8352 63928 8358 63980
rect 8588 63940 9076 63968
rect 8588 63912 8616 63940
rect 8570 63860 8576 63912
rect 8628 63860 8634 63912
rect 8662 63860 8668 63912
rect 8720 63900 8726 63912
rect 9048 63909 9076 63940
rect 10594 63928 10600 63980
rect 10652 63928 10658 63980
rect 8941 63903 8999 63909
rect 8941 63900 8953 63903
rect 8720 63872 8953 63900
rect 8720 63860 8726 63872
rect 8941 63869 8953 63872
rect 8987 63869 8999 63903
rect 8941 63863 8999 63869
rect 9033 63903 9091 63909
rect 9033 63869 9045 63903
rect 9079 63869 9091 63903
rect 9033 63863 9091 63869
rect 7837 63835 7895 63841
rect 7837 63801 7849 63835
rect 7883 63832 7895 63835
rect 8294 63832 8300 63844
rect 7883 63804 8300 63832
rect 7883 63801 7895 63804
rect 7837 63795 7895 63801
rect 8294 63792 8300 63804
rect 8352 63792 8358 63844
rect 8680 63832 8708 63860
rect 8404 63804 8708 63832
rect 1578 63724 1584 63776
rect 1636 63724 1642 63776
rect 5534 63724 5540 63776
rect 5592 63764 5598 63776
rect 5810 63764 5816 63776
rect 5592 63736 5816 63764
rect 5592 63724 5598 63736
rect 5810 63724 5816 63736
rect 5868 63724 5874 63776
rect 6362 63724 6368 63776
rect 6420 63764 6426 63776
rect 6822 63764 6828 63776
rect 6420 63736 6828 63764
rect 6420 63724 6426 63736
rect 6822 63724 6828 63736
rect 6880 63724 6886 63776
rect 8110 63724 8116 63776
rect 8168 63764 8174 63776
rect 8404 63764 8432 63804
rect 8168 63736 8432 63764
rect 8481 63767 8539 63773
rect 8168 63724 8174 63736
rect 8481 63733 8493 63767
rect 8527 63764 8539 63767
rect 9214 63764 9220 63776
rect 8527 63736 9220 63764
rect 8527 63733 8539 63736
rect 8481 63727 8539 63733
rect 9214 63724 9220 63736
rect 9272 63724 9278 63776
rect 1104 63674 9936 63696
rect 1104 63622 3610 63674
rect 3662 63622 3674 63674
rect 3726 63622 3738 63674
rect 3790 63622 3802 63674
rect 3854 63622 3866 63674
rect 3918 63622 5210 63674
rect 5262 63622 5274 63674
rect 5326 63622 5338 63674
rect 5390 63622 5402 63674
rect 5454 63622 5466 63674
rect 5518 63622 6810 63674
rect 6862 63622 6874 63674
rect 6926 63622 6938 63674
rect 6990 63622 7002 63674
rect 7054 63622 7066 63674
rect 7118 63622 8410 63674
rect 8462 63622 8474 63674
rect 8526 63622 8538 63674
rect 8590 63622 8602 63674
rect 8654 63622 8666 63674
rect 8718 63622 9936 63674
rect 1104 63600 9936 63622
rect 1578 63520 1584 63572
rect 1636 63560 1642 63572
rect 10410 63560 10416 63572
rect 1636 63532 10416 63560
rect 1636 63520 1642 63532
rect 10410 63520 10416 63532
rect 10468 63520 10474 63572
rect 2130 63452 2136 63504
rect 2188 63492 2194 63504
rect 2498 63492 2504 63504
rect 2188 63464 2504 63492
rect 2188 63452 2194 63464
rect 2498 63452 2504 63464
rect 2556 63452 2562 63504
rect 4798 63452 4804 63504
rect 4856 63492 4862 63504
rect 5166 63492 5172 63504
rect 4856 63464 5172 63492
rect 4856 63452 4862 63464
rect 5166 63452 5172 63464
rect 5224 63452 5230 63504
rect 5994 63452 6000 63504
rect 6052 63492 6058 63504
rect 6546 63492 6552 63504
rect 6052 63464 6552 63492
rect 6052 63452 6058 63464
rect 6546 63452 6552 63464
rect 6604 63452 6610 63504
rect 7650 63452 7656 63504
rect 7708 63452 7714 63504
rect 9674 63492 9680 63504
rect 8220 63464 9680 63492
rect 1210 63384 1216 63436
rect 1268 63424 1274 63436
rect 3602 63424 3608 63436
rect 1268 63396 3608 63424
rect 1268 63384 1274 63396
rect 3602 63384 3608 63396
rect 3660 63384 3666 63436
rect 5442 63384 5448 63436
rect 5500 63424 5506 63436
rect 6086 63424 6092 63436
rect 5500 63396 6092 63424
rect 5500 63384 5506 63396
rect 6086 63384 6092 63396
rect 6144 63384 6150 63436
rect 6730 63384 6736 63436
rect 6788 63424 6794 63436
rect 6917 63427 6975 63433
rect 6917 63424 6929 63427
rect 6788 63396 6929 63424
rect 6788 63384 6794 63396
rect 6917 63393 6929 63396
rect 6963 63393 6975 63427
rect 6917 63387 6975 63393
rect 7101 63427 7159 63433
rect 7101 63393 7113 63427
rect 7147 63424 7159 63427
rect 7668 63424 7696 63452
rect 8220 63424 8248 63464
rect 9674 63452 9680 63464
rect 9732 63452 9738 63504
rect 8297 63427 8355 63433
rect 8297 63424 8309 63427
rect 7147 63396 7236 63424
rect 7668 63396 8064 63424
rect 8220 63396 8309 63424
rect 7147 63393 7159 63396
rect 7101 63387 7159 63393
rect 7208 63368 7236 63396
rect 6270 63316 6276 63368
rect 6328 63356 6334 63368
rect 6825 63359 6883 63365
rect 6825 63356 6837 63359
rect 6328 63328 6837 63356
rect 6328 63316 6334 63328
rect 6825 63325 6837 63328
rect 6871 63325 6883 63359
rect 6825 63319 6883 63325
rect 7190 63316 7196 63368
rect 7248 63316 7254 63368
rect 7926 63316 7932 63368
rect 7984 63316 7990 63368
rect 8036 63365 8064 63396
rect 8297 63393 8309 63396
rect 8343 63393 8355 63427
rect 8297 63387 8355 63393
rect 8386 63384 8392 63436
rect 8444 63384 8450 63436
rect 8938 63424 8944 63436
rect 8496 63396 8944 63424
rect 8021 63359 8079 63365
rect 8021 63325 8033 63359
rect 8067 63325 8079 63359
rect 8021 63319 8079 63325
rect 8205 63359 8263 63365
rect 8205 63325 8217 63359
rect 8251 63325 8263 63359
rect 8205 63319 8263 63325
rect 7944 63288 7972 63316
rect 6840 63260 7972 63288
rect 8220 63288 8248 63319
rect 8496 63288 8524 63396
rect 8938 63384 8944 63396
rect 8996 63384 9002 63436
rect 9030 63384 9036 63436
rect 9088 63384 9094 63436
rect 8573 63359 8631 63365
rect 8573 63325 8585 63359
rect 8619 63356 8631 63359
rect 8846 63356 8852 63368
rect 8619 63328 8852 63356
rect 8619 63325 8631 63328
rect 8573 63319 8631 63325
rect 8220 63260 8524 63288
rect 6840 63232 6868 63260
rect 5534 63180 5540 63232
rect 5592 63220 5598 63232
rect 6457 63223 6515 63229
rect 6457 63220 6469 63223
rect 5592 63192 6469 63220
rect 5592 63180 5598 63192
rect 6457 63189 6469 63192
rect 6503 63189 6515 63223
rect 6457 63183 6515 63189
rect 6822 63180 6828 63232
rect 6880 63180 6886 63232
rect 7745 63223 7803 63229
rect 7745 63189 7757 63223
rect 7791 63220 7803 63223
rect 8588 63220 8616 63319
rect 8846 63316 8852 63328
rect 8904 63316 8910 63368
rect 7791 63192 8616 63220
rect 7791 63189 7803 63192
rect 7745 63183 7803 63189
rect 8754 63180 8760 63232
rect 8812 63180 8818 63232
rect 8938 63180 8944 63232
rect 8996 63220 9002 63232
rect 9048 63220 9076 63384
rect 8996 63192 9076 63220
rect 8996 63180 9002 63192
rect 1104 63130 9936 63152
rect 1104 63078 2950 63130
rect 3002 63078 3014 63130
rect 3066 63078 3078 63130
rect 3130 63078 3142 63130
rect 3194 63078 3206 63130
rect 3258 63078 4550 63130
rect 4602 63078 4614 63130
rect 4666 63078 4678 63130
rect 4730 63078 4742 63130
rect 4794 63078 4806 63130
rect 4858 63078 6150 63130
rect 6202 63078 6214 63130
rect 6266 63078 6278 63130
rect 6330 63078 6342 63130
rect 6394 63078 6406 63130
rect 6458 63078 7750 63130
rect 7802 63078 7814 63130
rect 7866 63078 7878 63130
rect 7930 63078 7942 63130
rect 7994 63078 8006 63130
rect 8058 63078 9350 63130
rect 9402 63078 9414 63130
rect 9466 63078 9478 63130
rect 9530 63078 9542 63130
rect 9594 63078 9606 63130
rect 9658 63078 9936 63130
rect 1104 63056 9936 63078
rect 4985 63019 5043 63025
rect 4985 62985 4997 63019
rect 5031 63016 5043 63019
rect 5994 63016 6000 63028
rect 5031 62988 6000 63016
rect 5031 62985 5043 62988
rect 4985 62979 5043 62985
rect 5994 62976 6000 62988
rect 6052 62976 6058 63028
rect 6730 62976 6736 63028
rect 6788 63016 6794 63028
rect 8021 63019 8079 63025
rect 8021 63016 8033 63019
rect 6788 62988 8033 63016
rect 6788 62976 6794 62988
rect 8021 62985 8033 62988
rect 8067 62985 8079 63019
rect 8021 62979 8079 62985
rect 8294 62976 8300 63028
rect 8352 63016 8358 63028
rect 8481 63019 8539 63025
rect 8481 63016 8493 63019
rect 8352 62988 8493 63016
rect 8352 62976 8358 62988
rect 8481 62985 8493 62988
rect 8527 62985 8539 63019
rect 8481 62979 8539 62985
rect 8754 62976 8760 63028
rect 8812 62976 8818 63028
rect 1026 62908 1032 62960
rect 1084 62948 1090 62960
rect 2314 62948 2320 62960
rect 1084 62920 2320 62948
rect 1084 62908 1090 62920
rect 2314 62908 2320 62920
rect 2372 62908 2378 62960
rect 8772 62948 8800 62976
rect 2746 62920 8800 62948
rect 934 62840 940 62892
rect 992 62880 998 62892
rect 1489 62883 1547 62889
rect 1489 62880 1501 62883
rect 992 62852 1501 62880
rect 992 62840 998 62852
rect 1489 62849 1501 62852
rect 1535 62849 1547 62883
rect 1489 62843 1547 62849
rect 2314 62772 2320 62824
rect 2372 62812 2378 62824
rect 2746 62812 2774 62920
rect 4798 62840 4804 62892
rect 4856 62840 4862 62892
rect 4893 62883 4951 62889
rect 4893 62849 4905 62883
rect 4939 62880 4951 62883
rect 6086 62880 6092 62892
rect 4939 62852 6092 62880
rect 4939 62849 4951 62852
rect 4893 62843 4951 62849
rect 6086 62840 6092 62852
rect 6144 62840 6150 62892
rect 6546 62884 6552 62892
rect 6472 62880 6552 62884
rect 6380 62856 6552 62880
rect 6380 62852 6500 62856
rect 2372 62784 2774 62812
rect 4816 62812 4844 62840
rect 5166 62812 5172 62824
rect 4816 62784 5172 62812
rect 2372 62772 2378 62784
rect 5166 62772 5172 62784
rect 5224 62772 5230 62824
rect 5442 62772 5448 62824
rect 5500 62812 5506 62824
rect 6380 62812 6408 62852
rect 6546 62840 6552 62856
rect 6604 62840 6610 62892
rect 6822 62889 6828 62892
rect 6816 62880 6828 62889
rect 6783 62852 6828 62880
rect 6816 62843 6828 62852
rect 6822 62840 6828 62843
rect 6880 62840 6886 62892
rect 7098 62840 7104 62892
rect 7156 62880 7162 62892
rect 7156 62852 7604 62880
rect 7156 62840 7162 62852
rect 5500 62784 6408 62812
rect 7576 62812 7604 62852
rect 7650 62840 7656 62892
rect 7708 62880 7714 62892
rect 8389 62883 8447 62889
rect 8389 62880 8401 62883
rect 7708 62852 8401 62880
rect 7708 62840 7714 62852
rect 8389 62849 8401 62852
rect 8435 62849 8447 62883
rect 8389 62843 8447 62849
rect 8662 62840 8668 62892
rect 8720 62880 8726 62892
rect 8849 62883 8907 62889
rect 8849 62880 8861 62883
rect 8720 62852 8861 62880
rect 8720 62840 8726 62852
rect 8849 62849 8861 62852
rect 8895 62849 8907 62883
rect 8849 62843 8907 62849
rect 7834 62812 7840 62824
rect 7576 62784 7840 62812
rect 5500 62772 5506 62784
rect 7834 62772 7840 62784
rect 7892 62772 7898 62824
rect 8478 62772 8484 62824
rect 8536 62812 8542 62824
rect 8573 62815 8631 62821
rect 8573 62812 8585 62815
rect 8536 62784 8585 62812
rect 8536 62772 8542 62784
rect 8573 62781 8585 62784
rect 8619 62781 8631 62815
rect 8573 62775 8631 62781
rect 8754 62772 8760 62824
rect 8812 62812 8818 62824
rect 10042 62812 10048 62824
rect 8812 62784 10048 62812
rect 8812 62772 8818 62784
rect 10042 62772 10048 62784
rect 10100 62772 10106 62824
rect 2746 62716 5120 62744
rect 1765 62679 1823 62685
rect 1765 62645 1777 62679
rect 1811 62676 1823 62679
rect 2746 62676 2774 62716
rect 1811 62648 2774 62676
rect 5092 62676 5120 62716
rect 7484 62716 10088 62744
rect 7484 62676 7512 62716
rect 10060 62688 10088 62716
rect 5092 62648 7512 62676
rect 1811 62645 1823 62648
rect 1765 62639 1823 62645
rect 7650 62636 7656 62688
rect 7708 62676 7714 62688
rect 7929 62679 7987 62685
rect 7929 62676 7941 62679
rect 7708 62648 7941 62676
rect 7708 62636 7714 62648
rect 7929 62645 7941 62648
rect 7975 62645 7987 62679
rect 7929 62639 7987 62645
rect 9033 62679 9091 62685
rect 9033 62645 9045 62679
rect 9079 62676 9091 62679
rect 9950 62676 9956 62688
rect 9079 62648 9956 62676
rect 9079 62645 9091 62648
rect 9033 62639 9091 62645
rect 9950 62636 9956 62648
rect 10008 62636 10014 62688
rect 10042 62636 10048 62688
rect 10100 62636 10106 62688
rect 1104 62586 9936 62608
rect 1104 62534 3610 62586
rect 3662 62534 3674 62586
rect 3726 62534 3738 62586
rect 3790 62534 3802 62586
rect 3854 62534 3866 62586
rect 3918 62534 5210 62586
rect 5262 62534 5274 62586
rect 5326 62534 5338 62586
rect 5390 62534 5402 62586
rect 5454 62534 5466 62586
rect 5518 62534 6810 62586
rect 6862 62534 6874 62586
rect 6926 62534 6938 62586
rect 6990 62534 7002 62586
rect 7054 62534 7066 62586
rect 7118 62534 8410 62586
rect 8462 62534 8474 62586
rect 8526 62534 8538 62586
rect 8590 62534 8602 62586
rect 8654 62534 8666 62586
rect 8718 62534 9936 62586
rect 1104 62512 9936 62534
rect 6454 62432 6460 62484
rect 6512 62472 6518 62484
rect 7469 62475 7527 62481
rect 6512 62444 7052 62472
rect 6512 62432 6518 62444
rect 4338 62404 4344 62416
rect 2332 62376 4344 62404
rect 2332 62277 2360 62376
rect 4338 62364 4344 62376
rect 4396 62364 4402 62416
rect 3804 62308 6868 62336
rect 2317 62271 2375 62277
rect 2317 62237 2329 62271
rect 2363 62237 2375 62271
rect 2317 62231 2375 62237
rect 2498 62160 2504 62212
rect 2556 62200 2562 62212
rect 3804 62200 3832 62308
rect 2556 62172 3832 62200
rect 2556 62160 2562 62172
rect 4338 62160 4344 62212
rect 4396 62200 4402 62212
rect 4706 62200 4712 62212
rect 4396 62172 4712 62200
rect 4396 62160 4402 62172
rect 4706 62160 4712 62172
rect 4764 62160 4770 62212
rect 5442 62160 5448 62212
rect 5500 62200 5506 62212
rect 6086 62200 6092 62212
rect 5500 62172 6092 62200
rect 5500 62160 5506 62172
rect 6086 62160 6092 62172
rect 6144 62200 6150 62212
rect 6840 62200 6868 62308
rect 7024 62277 7052 62444
rect 7469 62441 7481 62475
rect 7515 62472 7527 62475
rect 8846 62472 8852 62484
rect 7515 62444 8852 62472
rect 7515 62441 7527 62444
rect 7469 62435 7527 62441
rect 8846 62432 8852 62444
rect 8904 62432 8910 62484
rect 7208 62376 8064 62404
rect 7208 62348 7236 62376
rect 7190 62296 7196 62348
rect 7248 62296 7254 62348
rect 7282 62296 7288 62348
rect 7340 62296 7346 62348
rect 7558 62296 7564 62348
rect 7616 62336 7622 62348
rect 8036 62345 8064 62376
rect 7929 62339 7987 62345
rect 7929 62336 7941 62339
rect 7616 62308 7941 62336
rect 7616 62296 7622 62308
rect 7929 62305 7941 62308
rect 7975 62305 7987 62339
rect 7929 62299 7987 62305
rect 8021 62339 8079 62345
rect 8021 62305 8033 62339
rect 8067 62305 8079 62339
rect 8021 62299 8079 62305
rect 7009 62271 7067 62277
rect 7009 62237 7021 62271
rect 7055 62237 7067 62271
rect 7009 62231 7067 62237
rect 7101 62271 7159 62277
rect 7101 62237 7113 62271
rect 7147 62268 7159 62271
rect 7300 62268 7328 62296
rect 7147 62240 7328 62268
rect 7147 62237 7159 62240
rect 7101 62231 7159 62237
rect 7834 62228 7840 62280
rect 7892 62228 7898 62280
rect 8297 62271 8355 62277
rect 8297 62237 8309 62271
rect 8343 62237 8355 62271
rect 8754 62268 8760 62280
rect 8297 62231 8355 62237
rect 8404 62240 8760 62268
rect 8312 62200 8340 62231
rect 6144 62172 6767 62200
rect 6840 62172 8340 62200
rect 6144 62160 6150 62172
rect 1578 62092 1584 62144
rect 1636 62132 1642 62144
rect 2133 62135 2191 62141
rect 2133 62132 2145 62135
rect 1636 62104 2145 62132
rect 1636 62092 1642 62104
rect 2133 62101 2145 62104
rect 2179 62101 2191 62135
rect 2133 62095 2191 62101
rect 5994 62092 6000 62144
rect 6052 62132 6058 62144
rect 6641 62135 6699 62141
rect 6641 62132 6653 62135
rect 6052 62104 6653 62132
rect 6052 62092 6058 62104
rect 6641 62101 6653 62104
rect 6687 62101 6699 62135
rect 6739 62132 6767 62172
rect 8404 62132 8432 62240
rect 8754 62228 8760 62240
rect 8812 62228 8818 62280
rect 6739 62104 8432 62132
rect 8481 62135 8539 62141
rect 6641 62095 6699 62101
rect 8481 62101 8493 62135
rect 8527 62132 8539 62135
rect 11330 62132 11336 62144
rect 8527 62104 11336 62132
rect 8527 62101 8539 62104
rect 8481 62095 8539 62101
rect 11330 62092 11336 62104
rect 11388 62092 11394 62144
rect 1104 62042 9936 62064
rect 1104 61990 2950 62042
rect 3002 61990 3014 62042
rect 3066 61990 3078 62042
rect 3130 61990 3142 62042
rect 3194 61990 3206 62042
rect 3258 61990 4550 62042
rect 4602 61990 4614 62042
rect 4666 61990 4678 62042
rect 4730 61990 4742 62042
rect 4794 61990 4806 62042
rect 4858 61990 6150 62042
rect 6202 61990 6214 62042
rect 6266 61990 6278 62042
rect 6330 61990 6342 62042
rect 6394 61990 6406 62042
rect 6458 61990 7750 62042
rect 7802 61990 7814 62042
rect 7866 61990 7878 62042
rect 7930 61990 7942 62042
rect 7994 61990 8006 62042
rect 8058 61990 9350 62042
rect 9402 61990 9414 62042
rect 9466 61990 9478 62042
rect 9530 61990 9542 62042
rect 9594 61990 9606 62042
rect 9658 61990 9936 62042
rect 1104 61968 9936 61990
rect 5442 61888 5448 61940
rect 5500 61888 5506 61940
rect 8294 61888 8300 61940
rect 8352 61888 8358 61940
rect 1673 61863 1731 61869
rect 1673 61829 1685 61863
rect 1719 61860 1731 61863
rect 5460 61860 5488 61888
rect 1719 61832 5488 61860
rect 1719 61829 1731 61832
rect 1673 61823 1731 61829
rect 934 61752 940 61804
rect 992 61792 998 61804
rect 1489 61795 1547 61801
rect 1489 61792 1501 61795
rect 992 61764 1501 61792
rect 992 61752 998 61764
rect 1489 61761 1501 61764
rect 1535 61761 1547 61795
rect 1489 61755 1547 61761
rect 6546 61752 6552 61804
rect 6604 61792 6610 61804
rect 6641 61795 6699 61801
rect 6641 61792 6653 61795
rect 6604 61764 6653 61792
rect 6604 61752 6610 61764
rect 6641 61761 6653 61764
rect 6687 61761 6699 61795
rect 6641 61755 6699 61761
rect 6908 61795 6966 61801
rect 6908 61761 6920 61795
rect 6954 61792 6966 61795
rect 6954 61764 7696 61792
rect 6954 61761 6966 61764
rect 6908 61755 6966 61761
rect 7668 61656 7696 61764
rect 7742 61752 7748 61804
rect 7800 61792 7806 61804
rect 8202 61792 8208 61804
rect 7800 61764 8208 61792
rect 7800 61752 7806 61764
rect 8202 61752 8208 61764
rect 8260 61752 8266 61804
rect 8312 61792 8340 61888
rect 8386 61820 8392 61872
rect 8444 61860 8450 61872
rect 8481 61863 8539 61869
rect 8481 61860 8493 61863
rect 8444 61832 8493 61860
rect 8444 61820 8450 61832
rect 8481 61829 8493 61832
rect 8527 61829 8539 61863
rect 8481 61823 8539 61829
rect 8754 61820 8760 61872
rect 8812 61860 8818 61872
rect 8812 61832 9352 61860
rect 8812 61820 8818 61832
rect 9324 61804 9352 61832
rect 8312 61764 8708 61792
rect 8294 61684 8300 61736
rect 8352 61724 8358 61736
rect 8680 61733 8708 61764
rect 9306 61752 9312 61804
rect 9364 61752 9370 61804
rect 8573 61727 8631 61733
rect 8573 61724 8585 61727
rect 8352 61696 8585 61724
rect 8352 61684 8358 61696
rect 8573 61693 8585 61696
rect 8619 61693 8631 61727
rect 8573 61687 8631 61693
rect 8665 61727 8723 61733
rect 8665 61693 8677 61727
rect 8711 61724 8723 61727
rect 8754 61724 8760 61736
rect 8711 61696 8760 61724
rect 8711 61693 8723 61696
rect 8665 61687 8723 61693
rect 8754 61684 8760 61696
rect 8812 61684 8818 61736
rect 8938 61656 8944 61668
rect 7668 61628 8944 61656
rect 8938 61616 8944 61628
rect 8996 61616 9002 61668
rect 8018 61548 8024 61600
rect 8076 61548 8082 61600
rect 8110 61548 8116 61600
rect 8168 61548 8174 61600
rect 1104 61498 9936 61520
rect 1104 61446 3610 61498
rect 3662 61446 3674 61498
rect 3726 61446 3738 61498
rect 3790 61446 3802 61498
rect 3854 61446 3866 61498
rect 3918 61446 5210 61498
rect 5262 61446 5274 61498
rect 5326 61446 5338 61498
rect 5390 61446 5402 61498
rect 5454 61446 5466 61498
rect 5518 61446 6810 61498
rect 6862 61446 6874 61498
rect 6926 61446 6938 61498
rect 6990 61446 7002 61498
rect 7054 61446 7066 61498
rect 7118 61446 8410 61498
rect 8462 61446 8474 61498
rect 8526 61446 8538 61498
rect 8590 61446 8602 61498
rect 8654 61446 8666 61498
rect 8718 61446 9936 61498
rect 1104 61424 9936 61446
rect 7190 61344 7196 61396
rect 7248 61384 7254 61396
rect 7466 61384 7472 61396
rect 7248 61356 7472 61384
rect 7248 61344 7254 61356
rect 7466 61344 7472 61356
rect 7524 61384 7530 61396
rect 7524 61356 7880 61384
rect 7524 61344 7530 61356
rect 7650 61208 7656 61260
rect 7708 61208 7714 61260
rect 7852 61257 7880 61356
rect 8018 61344 8024 61396
rect 8076 61344 8082 61396
rect 8938 61344 8944 61396
rect 8996 61344 9002 61396
rect 7837 61251 7895 61257
rect 7837 61217 7849 61251
rect 7883 61217 7895 61251
rect 8036 61248 8064 61344
rect 8956 61316 8984 61344
rect 8588 61288 8984 61316
rect 8481 61251 8539 61257
rect 8481 61248 8493 61251
rect 8036 61220 8493 61248
rect 7837 61211 7895 61217
rect 8481 61217 8493 61220
rect 8527 61217 8539 61251
rect 8481 61211 8539 61217
rect 5258 61140 5264 61192
rect 5316 61180 5322 61192
rect 5810 61180 5816 61192
rect 5316 61152 5816 61180
rect 5316 61140 5322 61152
rect 5810 61140 5816 61152
rect 5868 61140 5874 61192
rect 7282 61140 7288 61192
rect 7340 61180 7346 61192
rect 7561 61183 7619 61189
rect 7561 61180 7573 61183
rect 7340 61152 7573 61180
rect 7340 61140 7346 61152
rect 7561 61149 7573 61152
rect 7607 61149 7619 61183
rect 7561 61143 7619 61149
rect 8389 61183 8447 61189
rect 8389 61149 8401 61183
rect 8435 61180 8447 61183
rect 8588 61180 8616 61288
rect 8665 61251 8723 61257
rect 8665 61217 8677 61251
rect 8711 61248 8723 61251
rect 8754 61248 8760 61260
rect 8711 61220 8760 61248
rect 8711 61217 8723 61220
rect 8665 61211 8723 61217
rect 8754 61208 8760 61220
rect 8812 61208 8818 61260
rect 9122 61208 9128 61260
rect 9180 61248 9186 61260
rect 9766 61248 9772 61260
rect 9180 61220 9772 61248
rect 9180 61208 9186 61220
rect 9766 61208 9772 61220
rect 9824 61208 9830 61260
rect 8435 61152 8616 61180
rect 8435 61149 8447 61152
rect 8389 61143 8447 61149
rect 8938 61140 8944 61192
rect 8996 61140 9002 61192
rect 5166 61072 5172 61124
rect 5224 61112 5230 61124
rect 5224 61084 8064 61112
rect 5224 61072 5230 61084
rect 5810 61004 5816 61056
rect 5868 61044 5874 61056
rect 8036 61053 8064 61084
rect 8754 61072 8760 61124
rect 8812 61112 8818 61124
rect 9306 61112 9312 61124
rect 8812 61084 9312 61112
rect 8812 61072 8818 61084
rect 9306 61072 9312 61084
rect 9364 61072 9370 61124
rect 7193 61047 7251 61053
rect 7193 61044 7205 61047
rect 5868 61016 7205 61044
rect 5868 61004 5874 61016
rect 7193 61013 7205 61016
rect 7239 61013 7251 61047
rect 7193 61007 7251 61013
rect 8021 61047 8079 61053
rect 8021 61013 8033 61047
rect 8067 61013 8079 61047
rect 8021 61007 8079 61013
rect 9122 61004 9128 61056
rect 9180 61004 9186 61056
rect 1104 60954 9936 60976
rect 1104 60902 2950 60954
rect 3002 60902 3014 60954
rect 3066 60902 3078 60954
rect 3130 60902 3142 60954
rect 3194 60902 3206 60954
rect 3258 60902 4550 60954
rect 4602 60902 4614 60954
rect 4666 60902 4678 60954
rect 4730 60902 4742 60954
rect 4794 60902 4806 60954
rect 4858 60902 6150 60954
rect 6202 60902 6214 60954
rect 6266 60902 6278 60954
rect 6330 60902 6342 60954
rect 6394 60902 6406 60954
rect 6458 60902 7750 60954
rect 7802 60902 7814 60954
rect 7866 60902 7878 60954
rect 7930 60902 7942 60954
rect 7994 60902 8006 60954
rect 8058 60902 9350 60954
rect 9402 60902 9414 60954
rect 9466 60902 9478 60954
rect 9530 60902 9542 60954
rect 9594 60902 9606 60954
rect 9658 60902 9936 60954
rect 1104 60880 9936 60902
rect 474 60800 480 60852
rect 532 60840 538 60852
rect 8938 60840 8944 60852
rect 532 60812 8944 60840
rect 532 60800 538 60812
rect 8938 60800 8944 60812
rect 8996 60800 9002 60852
rect 9398 60800 9404 60852
rect 9456 60840 9462 60852
rect 9858 60840 9864 60852
rect 9456 60812 9864 60840
rect 9456 60800 9462 60812
rect 9858 60800 9864 60812
rect 9916 60800 9922 60852
rect 4798 60732 4804 60784
rect 4856 60772 4862 60784
rect 5169 60775 5227 60781
rect 5169 60772 5181 60775
rect 4856 60744 5181 60772
rect 4856 60732 4862 60744
rect 5169 60741 5181 60744
rect 5215 60741 5227 60775
rect 5169 60735 5227 60741
rect 7000 60775 7058 60781
rect 7000 60741 7012 60775
rect 7046 60772 7058 60775
rect 7650 60772 7656 60784
rect 7046 60744 7656 60772
rect 7046 60741 7058 60744
rect 7000 60735 7058 60741
rect 7650 60732 7656 60744
rect 7708 60732 7714 60784
rect 934 60664 940 60716
rect 992 60704 998 60716
rect 1397 60707 1455 60713
rect 1397 60704 1409 60707
rect 992 60676 1409 60704
rect 992 60664 998 60676
rect 1397 60673 1409 60676
rect 1443 60673 1455 60707
rect 1397 60667 1455 60673
rect 2682 60664 2688 60716
rect 2740 60704 2746 60716
rect 4065 60707 4123 60713
rect 4065 60704 4077 60707
rect 2740 60676 4077 60704
rect 2740 60664 2746 60676
rect 4065 60673 4077 60676
rect 4111 60673 4123 60707
rect 4065 60667 4123 60673
rect 4430 60664 4436 60716
rect 4488 60664 4494 60716
rect 4893 60707 4951 60713
rect 4893 60673 4905 60707
rect 4939 60673 4951 60707
rect 4893 60667 4951 60673
rect 4908 60568 4936 60667
rect 6546 60664 6552 60716
rect 6604 60704 6610 60716
rect 6733 60707 6791 60713
rect 6733 60704 6745 60707
rect 6604 60676 6745 60704
rect 6604 60664 6610 60676
rect 6733 60673 6745 60676
rect 6779 60704 6791 60707
rect 7282 60704 7288 60716
rect 6779 60676 7288 60704
rect 6779 60673 6791 60676
rect 6733 60667 6791 60673
rect 7282 60664 7288 60676
rect 7340 60664 7346 60716
rect 4448 60540 4936 60568
rect 8113 60571 8171 60577
rect 4448 60512 4476 60540
rect 8113 60537 8125 60571
rect 8159 60568 8171 60571
rect 8294 60568 8300 60580
rect 8159 60540 8300 60568
rect 8159 60537 8171 60540
rect 8113 60531 8171 60537
rect 8294 60528 8300 60540
rect 8352 60528 8358 60580
rect 1581 60503 1639 60509
rect 1581 60469 1593 60503
rect 1627 60500 1639 60503
rect 2774 60500 2780 60512
rect 1627 60472 2780 60500
rect 1627 60469 1639 60472
rect 1581 60463 1639 60469
rect 2774 60460 2780 60472
rect 2832 60460 2838 60512
rect 4430 60460 4436 60512
rect 4488 60460 4494 60512
rect 4890 60460 4896 60512
rect 4948 60500 4954 60512
rect 5258 60500 5264 60512
rect 4948 60472 5264 60500
rect 4948 60460 4954 60472
rect 5258 60460 5264 60472
rect 5316 60460 5322 60512
rect 5350 60460 5356 60512
rect 5408 60500 5414 60512
rect 6546 60500 6552 60512
rect 5408 60472 6552 60500
rect 5408 60460 5414 60472
rect 6546 60460 6552 60472
rect 6604 60460 6610 60512
rect 1104 60410 9936 60432
rect 1104 60358 3610 60410
rect 3662 60358 3674 60410
rect 3726 60358 3738 60410
rect 3790 60358 3802 60410
rect 3854 60358 3866 60410
rect 3918 60358 5210 60410
rect 5262 60358 5274 60410
rect 5326 60358 5338 60410
rect 5390 60358 5402 60410
rect 5454 60358 5466 60410
rect 5518 60358 6810 60410
rect 6862 60358 6874 60410
rect 6926 60358 6938 60410
rect 6990 60358 7002 60410
rect 7054 60358 7066 60410
rect 7118 60358 8410 60410
rect 8462 60358 8474 60410
rect 8526 60358 8538 60410
rect 8590 60358 8602 60410
rect 8654 60358 8666 60410
rect 8718 60358 9936 60410
rect 1104 60336 9936 60358
rect 4798 60256 4804 60308
rect 4856 60296 4862 60308
rect 5074 60296 5080 60308
rect 4856 60268 5080 60296
rect 4856 60256 4862 60268
rect 5074 60256 5080 60268
rect 5132 60256 5138 60308
rect 7650 60256 7656 60308
rect 7708 60296 7714 60308
rect 8202 60296 8208 60308
rect 7708 60268 8208 60296
rect 7708 60256 7714 60268
rect 8202 60256 8208 60268
rect 8260 60256 8266 60308
rect 8846 60188 8852 60240
rect 8904 60228 8910 60240
rect 9214 60228 9220 60240
rect 8904 60200 9220 60228
rect 8904 60188 8910 60200
rect 9214 60188 9220 60200
rect 9272 60188 9278 60240
rect 2774 60120 2780 60172
rect 2832 60160 2838 60172
rect 3878 60160 3884 60172
rect 2832 60132 3884 60160
rect 2832 60120 2838 60132
rect 3878 60120 3884 60132
rect 3936 60120 3942 60172
rect 7282 60120 7288 60172
rect 7340 60120 7346 60172
rect 9398 60120 9404 60172
rect 9456 60120 9462 60172
rect 7552 60095 7610 60101
rect 7552 60061 7564 60095
rect 7598 60092 7610 60095
rect 9416 60092 9444 60120
rect 7598 60064 9444 60092
rect 7598 60061 7610 60064
rect 7552 60055 7610 60061
rect 8220 60036 8248 60064
rect 1486 59984 1492 60036
rect 1544 59984 1550 60036
rect 8202 59984 8208 60036
rect 8260 59984 8266 60036
rect 934 59916 940 59968
rect 992 59956 998 59968
rect 1581 59959 1639 59965
rect 1581 59956 1593 59959
rect 992 59928 1593 59956
rect 992 59916 998 59928
rect 1581 59925 1593 59928
rect 1627 59925 1639 59959
rect 1581 59919 1639 59925
rect 8294 59916 8300 59968
rect 8352 59956 8358 59968
rect 8665 59959 8723 59965
rect 8665 59956 8677 59959
rect 8352 59928 8677 59956
rect 8352 59916 8358 59928
rect 8665 59925 8677 59928
rect 8711 59925 8723 59959
rect 8665 59919 8723 59925
rect 1104 59866 9936 59888
rect 1104 59814 2950 59866
rect 3002 59814 3014 59866
rect 3066 59814 3078 59866
rect 3130 59814 3142 59866
rect 3194 59814 3206 59866
rect 3258 59814 4550 59866
rect 4602 59814 4614 59866
rect 4666 59814 4678 59866
rect 4730 59814 4742 59866
rect 4794 59814 4806 59866
rect 4858 59814 6150 59866
rect 6202 59814 6214 59866
rect 6266 59814 6278 59866
rect 6330 59814 6342 59866
rect 6394 59814 6406 59866
rect 6458 59814 7750 59866
rect 7802 59814 7814 59866
rect 7866 59814 7878 59866
rect 7930 59814 7942 59866
rect 7994 59814 8006 59866
rect 8058 59814 9350 59866
rect 9402 59814 9414 59866
rect 9466 59814 9478 59866
rect 9530 59814 9542 59866
rect 9594 59814 9606 59866
rect 9658 59814 9936 59866
rect 1104 59792 9936 59814
rect 1486 59712 1492 59764
rect 1544 59752 1550 59764
rect 4157 59755 4215 59761
rect 4157 59752 4169 59755
rect 1544 59724 4169 59752
rect 1544 59712 1550 59724
rect 4157 59721 4169 59724
rect 4203 59721 4215 59755
rect 4157 59715 4215 59721
rect 7374 59712 7380 59764
rect 7432 59752 7438 59764
rect 9125 59755 9183 59761
rect 9125 59752 9137 59755
rect 7432 59724 9137 59752
rect 7432 59712 7438 59724
rect 9125 59721 9137 59724
rect 9171 59721 9183 59755
rect 9125 59715 9183 59721
rect 1210 59644 1216 59696
rect 1268 59684 1274 59696
rect 1268 59656 5120 59684
rect 1268 59644 1274 59656
rect 3970 59576 3976 59628
rect 4028 59576 4034 59628
rect 5092 59625 5120 59656
rect 5718 59644 5724 59696
rect 5776 59684 5782 59696
rect 11606 59684 11612 59696
rect 5776 59656 11612 59684
rect 5776 59644 5782 59656
rect 11606 59644 11612 59656
rect 11664 59644 11670 59696
rect 4341 59619 4399 59625
rect 4341 59585 4353 59619
rect 4387 59616 4399 59619
rect 5077 59619 5135 59625
rect 4387 59588 5028 59616
rect 4387 59585 4399 59588
rect 4341 59579 4399 59585
rect 4890 59508 4896 59560
rect 4948 59508 4954 59560
rect 5000 59548 5028 59588
rect 5077 59585 5089 59619
rect 5123 59585 5135 59619
rect 5077 59579 5135 59585
rect 7837 59619 7895 59625
rect 7837 59585 7849 59619
rect 7883 59616 7895 59619
rect 7883 59588 11192 59616
rect 7883 59585 7895 59588
rect 7837 59579 7895 59585
rect 7282 59548 7288 59560
rect 5000 59520 7288 59548
rect 7282 59508 7288 59520
rect 7340 59508 7346 59560
rect 11164 59424 11192 59588
rect 2774 59372 2780 59424
rect 2832 59412 2838 59424
rect 3789 59415 3847 59421
rect 3789 59412 3801 59415
rect 2832 59384 3801 59412
rect 2832 59372 2838 59384
rect 3789 59381 3801 59384
rect 3835 59381 3847 59415
rect 3789 59375 3847 59381
rect 4522 59372 4528 59424
rect 4580 59412 4586 59424
rect 5261 59415 5319 59421
rect 5261 59412 5273 59415
rect 4580 59384 5273 59412
rect 4580 59372 4586 59384
rect 5261 59381 5273 59384
rect 5307 59381 5319 59415
rect 5261 59375 5319 59381
rect 11146 59372 11152 59424
rect 11204 59412 11210 59424
rect 11974 59412 11980 59424
rect 11204 59384 11980 59412
rect 11204 59372 11210 59384
rect 11974 59372 11980 59384
rect 12032 59372 12038 59424
rect 1104 59322 9936 59344
rect 1104 59270 3610 59322
rect 3662 59270 3674 59322
rect 3726 59270 3738 59322
rect 3790 59270 3802 59322
rect 3854 59270 3866 59322
rect 3918 59270 5210 59322
rect 5262 59270 5274 59322
rect 5326 59270 5338 59322
rect 5390 59270 5402 59322
rect 5454 59270 5466 59322
rect 5518 59270 6810 59322
rect 6862 59270 6874 59322
rect 6926 59270 6938 59322
rect 6990 59270 7002 59322
rect 7054 59270 7066 59322
rect 7118 59270 8410 59322
rect 8462 59270 8474 59322
rect 8526 59270 8538 59322
rect 8590 59270 8602 59322
rect 8654 59270 8666 59322
rect 8718 59270 9936 59322
rect 1104 59248 9936 59270
rect 4246 59168 4252 59220
rect 4304 59208 4310 59220
rect 6825 59211 6883 59217
rect 6825 59208 6837 59211
rect 4304 59180 6837 59208
rect 4304 59168 4310 59180
rect 6825 59177 6837 59180
rect 6871 59177 6883 59211
rect 7374 59208 7380 59220
rect 6825 59171 6883 59177
rect 7116 59180 7380 59208
rect 6546 59100 6552 59152
rect 6604 59100 6610 59152
rect 4338 59032 4344 59084
rect 4396 59072 4402 59084
rect 6564 59072 6592 59100
rect 6822 59072 6828 59084
rect 4396 59044 5212 59072
rect 6564 59044 6828 59072
rect 4396 59032 4402 59044
rect 290 58964 296 59016
rect 348 58964 354 59016
rect 1489 59007 1547 59013
rect 1489 58973 1501 59007
rect 1535 59004 1547 59007
rect 2866 59004 2872 59016
rect 1535 58976 2872 59004
rect 1535 58973 1547 58976
rect 1489 58967 1547 58973
rect 2866 58964 2872 58976
rect 2924 58964 2930 59016
rect 4246 58964 4252 59016
rect 4304 59004 4310 59016
rect 4522 59004 4528 59016
rect 4304 58976 4528 59004
rect 4304 58964 4310 58976
rect 4522 58964 4528 58976
rect 4580 58964 4586 59016
rect 4890 58964 4896 59016
rect 4948 59004 4954 59016
rect 5184 59013 5212 59044
rect 6822 59032 6828 59044
rect 6880 59032 6886 59084
rect 4985 59007 5043 59013
rect 4985 59004 4997 59007
rect 4948 58976 4997 59004
rect 4948 58964 4954 58976
rect 4985 58973 4997 58976
rect 5031 58973 5043 59007
rect 4985 58967 5043 58973
rect 5169 59007 5227 59013
rect 5169 58973 5181 59007
rect 5215 58973 5227 59007
rect 5169 58967 5227 58973
rect 5445 59007 5503 59013
rect 5445 58973 5457 59007
rect 5491 59004 5503 59007
rect 6546 59004 6552 59016
rect 5491 58976 6552 59004
rect 5491 58973 5503 58976
rect 5445 58967 5503 58973
rect 6546 58964 6552 58976
rect 6604 59004 6610 59016
rect 7116 59013 7144 59180
rect 7374 59168 7380 59180
rect 7432 59168 7438 59220
rect 7101 59007 7159 59013
rect 7101 59004 7113 59007
rect 6604 58976 7113 59004
rect 6604 58964 6610 58976
rect 7101 58973 7113 58976
rect 7147 58973 7159 59007
rect 7101 58967 7159 58973
rect 7368 59007 7426 59013
rect 7368 58973 7380 59007
rect 7414 59004 7426 59007
rect 7650 59004 7656 59016
rect 7414 58976 7656 59004
rect 7414 58973 7426 58976
rect 7368 58967 7426 58973
rect 7650 58964 7656 58976
rect 7708 59004 7714 59016
rect 9582 59004 9588 59016
rect 7708 58976 9588 59004
rect 7708 58964 7714 58976
rect 9582 58964 9588 58976
rect 9640 58964 9646 59016
rect 308 58936 336 58964
rect 5718 58945 5724 58948
rect 5690 58939 5724 58945
rect 5690 58936 5702 58939
rect 308 58908 5702 58936
rect 5690 58905 5702 58908
rect 5690 58899 5724 58905
rect 5718 58896 5724 58899
rect 5776 58896 5782 58948
rect 5902 58896 5908 58948
rect 5960 58936 5966 58948
rect 6822 58936 6828 58948
rect 5960 58908 6828 58936
rect 5960 58896 5966 58908
rect 6822 58896 6828 58908
rect 6880 58896 6886 58948
rect 934 58828 940 58880
rect 992 58868 998 58880
rect 1581 58871 1639 58877
rect 1581 58868 1593 58871
rect 992 58840 1593 58868
rect 992 58828 998 58840
rect 1581 58837 1593 58840
rect 1627 58837 1639 58871
rect 1581 58831 1639 58837
rect 5074 58828 5080 58880
rect 5132 58868 5138 58880
rect 5353 58871 5411 58877
rect 5353 58868 5365 58871
rect 5132 58840 5365 58868
rect 5132 58828 5138 58840
rect 5353 58837 5365 58840
rect 5399 58837 5411 58871
rect 5353 58831 5411 58837
rect 7374 58828 7380 58880
rect 7432 58868 7438 58880
rect 7742 58868 7748 58880
rect 7432 58840 7748 58868
rect 7432 58828 7438 58840
rect 7742 58828 7748 58840
rect 7800 58828 7806 58880
rect 8386 58828 8392 58880
rect 8444 58868 8450 58880
rect 8481 58871 8539 58877
rect 8481 58868 8493 58871
rect 8444 58840 8493 58868
rect 8444 58828 8450 58840
rect 8481 58837 8493 58840
rect 8527 58837 8539 58871
rect 8481 58831 8539 58837
rect 1104 58778 9936 58800
rect 1104 58726 2950 58778
rect 3002 58726 3014 58778
rect 3066 58726 3078 58778
rect 3130 58726 3142 58778
rect 3194 58726 3206 58778
rect 3258 58726 4550 58778
rect 4602 58726 4614 58778
rect 4666 58726 4678 58778
rect 4730 58726 4742 58778
rect 4794 58726 4806 58778
rect 4858 58726 6150 58778
rect 6202 58726 6214 58778
rect 6266 58726 6278 58778
rect 6330 58726 6342 58778
rect 6394 58726 6406 58778
rect 6458 58726 7750 58778
rect 7802 58726 7814 58778
rect 7866 58726 7878 58778
rect 7930 58726 7942 58778
rect 7994 58726 8006 58778
rect 8058 58726 9350 58778
rect 9402 58726 9414 58778
rect 9466 58726 9478 58778
rect 9530 58726 9542 58778
rect 9594 58726 9606 58778
rect 9658 58726 9936 58778
rect 1104 58704 9936 58726
rect 5718 58624 5724 58676
rect 5776 58664 5782 58676
rect 6086 58664 6092 58676
rect 5776 58636 6092 58664
rect 5776 58624 5782 58636
rect 6086 58624 6092 58636
rect 6144 58624 6150 58676
rect 6362 58624 6368 58676
rect 6420 58664 6426 58676
rect 6914 58664 6920 58676
rect 6420 58636 6920 58664
rect 6420 58624 6426 58636
rect 6914 58624 6920 58636
rect 6972 58624 6978 58676
rect 8205 58667 8263 58673
rect 8205 58633 8217 58667
rect 8251 58664 8263 58667
rect 8294 58664 8300 58676
rect 8251 58636 8300 58664
rect 8251 58633 8263 58636
rect 8205 58627 8263 58633
rect 8294 58624 8300 58636
rect 8352 58624 8358 58676
rect 9030 58624 9036 58676
rect 9088 58664 9094 58676
rect 9306 58664 9312 58676
rect 9088 58636 9312 58664
rect 9088 58624 9094 58636
rect 9306 58624 9312 58636
rect 9364 58624 9370 58676
rect 10318 58596 10324 58608
rect 5992 58568 10324 58596
rect 4890 58488 4896 58540
rect 4948 58488 4954 58540
rect 5992 58537 6020 58568
rect 10318 58556 10324 58568
rect 10376 58556 10382 58608
rect 5992 58531 6055 58537
rect 5992 58498 6009 58531
rect 5997 58497 6009 58498
rect 6043 58497 6055 58531
rect 5997 58491 6055 58497
rect 6733 58531 6791 58537
rect 6733 58497 6745 58531
rect 6779 58528 6791 58531
rect 6822 58528 6828 58540
rect 6779 58500 6828 58528
rect 6779 58497 6791 58500
rect 6733 58491 6791 58497
rect 6822 58488 6828 58500
rect 6880 58488 6886 58540
rect 7190 58488 7196 58540
rect 7248 58488 7254 58540
rect 8113 58531 8171 58537
rect 8113 58497 8125 58531
rect 8159 58528 8171 58531
rect 8202 58528 8208 58540
rect 8159 58500 8208 58528
rect 8159 58497 8171 58500
rect 8113 58491 8171 58497
rect 8202 58488 8208 58500
rect 8260 58488 8266 58540
rect 8573 58531 8631 58537
rect 8573 58497 8585 58531
rect 8619 58528 8631 58531
rect 10870 58528 10876 58540
rect 8619 58500 10876 58528
rect 8619 58497 8631 58500
rect 8573 58491 8631 58497
rect 10870 58488 10876 58500
rect 10928 58488 10934 58540
rect 4908 58460 4936 58488
rect 6549 58463 6607 58469
rect 6549 58460 6561 58463
rect 4908 58432 6561 58460
rect 6549 58429 6561 58432
rect 6595 58460 6607 58463
rect 7009 58463 7067 58469
rect 7009 58460 7021 58463
rect 6595 58432 7021 58460
rect 6595 58429 6607 58432
rect 6549 58423 6607 58429
rect 7009 58429 7021 58432
rect 7055 58429 7067 58463
rect 7009 58423 7067 58429
rect 4890 58352 4896 58404
rect 4948 58392 4954 58404
rect 5166 58392 5172 58404
rect 4948 58364 5172 58392
rect 4948 58352 4954 58364
rect 5166 58352 5172 58364
rect 5224 58352 5230 58404
rect 5718 58352 5724 58404
rect 5776 58392 5782 58404
rect 6917 58395 6975 58401
rect 6917 58392 6929 58395
rect 5776 58364 6929 58392
rect 5776 58352 5782 58364
rect 6917 58361 6929 58364
rect 6963 58361 6975 58395
rect 7024 58392 7052 58423
rect 7466 58420 7472 58472
rect 7524 58460 7530 58472
rect 7650 58460 7656 58472
rect 7524 58432 7656 58460
rect 7524 58420 7530 58432
rect 7650 58420 7656 58432
rect 7708 58460 7714 58472
rect 8297 58463 8355 58469
rect 8297 58460 8309 58463
rect 7708 58432 8309 58460
rect 7708 58420 7714 58432
rect 8297 58429 8309 58432
rect 8343 58429 8355 58463
rect 8297 58423 8355 58429
rect 8754 58420 8760 58472
rect 8812 58420 8818 58472
rect 7190 58392 7196 58404
rect 7024 58364 7196 58392
rect 6917 58355 6975 58361
rect 7190 58352 7196 58364
rect 7248 58352 7254 58404
rect 7300 58364 7788 58392
rect 5902 58284 5908 58336
rect 5960 58324 5966 58336
rect 6181 58327 6239 58333
rect 6181 58324 6193 58327
rect 5960 58296 6193 58324
rect 5960 58284 5966 58296
rect 6181 58293 6193 58296
rect 6227 58293 6239 58327
rect 6181 58287 6239 58293
rect 6454 58284 6460 58336
rect 6512 58324 6518 58336
rect 7300 58324 7328 58364
rect 6512 58296 7328 58324
rect 7377 58327 7435 58333
rect 6512 58284 6518 58296
rect 7377 58293 7389 58327
rect 7423 58324 7435 58327
rect 7466 58324 7472 58336
rect 7423 58296 7472 58324
rect 7423 58293 7435 58296
rect 7377 58287 7435 58293
rect 7466 58284 7472 58296
rect 7524 58284 7530 58336
rect 7760 58333 7788 58364
rect 8202 58352 8208 58404
rect 8260 58392 8266 58404
rect 8772 58392 8800 58420
rect 8260 58364 8800 58392
rect 8260 58352 8266 58364
rect 7745 58327 7803 58333
rect 7745 58293 7757 58327
rect 7791 58293 7803 58327
rect 7745 58287 7803 58293
rect 8754 58284 8760 58336
rect 8812 58284 8818 58336
rect 1104 58234 9936 58256
rect 1104 58182 3610 58234
rect 3662 58182 3674 58234
rect 3726 58182 3738 58234
rect 3790 58182 3802 58234
rect 3854 58182 3866 58234
rect 3918 58182 5210 58234
rect 5262 58182 5274 58234
rect 5326 58182 5338 58234
rect 5390 58182 5402 58234
rect 5454 58182 5466 58234
rect 5518 58182 6810 58234
rect 6862 58182 6874 58234
rect 6926 58182 6938 58234
rect 6990 58182 7002 58234
rect 7054 58182 7066 58234
rect 7118 58182 8410 58234
rect 8462 58182 8474 58234
rect 8526 58182 8538 58234
rect 8590 58182 8602 58234
rect 8654 58182 8666 58234
rect 8718 58182 9936 58234
rect 1104 58160 9936 58182
rect 4890 58080 4896 58132
rect 4948 58120 4954 58132
rect 5166 58120 5172 58132
rect 4948 58092 5172 58120
rect 4948 58080 4954 58092
rect 5166 58080 5172 58092
rect 5224 58080 5230 58132
rect 7101 58123 7159 58129
rect 7101 58089 7113 58123
rect 7147 58120 7159 58123
rect 7190 58120 7196 58132
rect 7147 58092 7196 58120
rect 7147 58089 7159 58092
rect 7101 58083 7159 58089
rect 7190 58080 7196 58092
rect 7248 58080 7254 58132
rect 7282 58080 7288 58132
rect 7340 58120 7346 58132
rect 7653 58123 7711 58129
rect 7653 58120 7665 58123
rect 7340 58092 7665 58120
rect 7340 58080 7346 58092
rect 7653 58089 7665 58092
rect 7699 58089 7711 58123
rect 7653 58083 7711 58089
rect 7208 57993 7236 58080
rect 8220 58024 8432 58052
rect 8220 57993 8248 58024
rect 7193 57987 7251 57993
rect 7193 57953 7205 57987
rect 7239 57953 7251 57987
rect 7193 57947 7251 57953
rect 8205 57987 8263 57993
rect 8205 57953 8217 57987
rect 8251 57953 8263 57987
rect 8205 57947 8263 57953
rect 8294 57944 8300 57996
rect 8352 57944 8358 57996
rect 8404 57984 8432 58024
rect 8404 57956 8708 57984
rect 1489 57919 1547 57925
rect 1489 57885 1501 57919
rect 1535 57916 1547 57919
rect 2682 57916 2688 57928
rect 1535 57888 2688 57916
rect 1535 57885 1547 57888
rect 1489 57879 1547 57885
rect 2682 57876 2688 57888
rect 2740 57876 2746 57928
rect 6362 57876 6368 57928
rect 6420 57916 6426 57928
rect 6917 57919 6975 57925
rect 6917 57916 6929 57919
rect 6420 57888 6929 57916
rect 6420 57876 6426 57888
rect 6917 57885 6929 57888
rect 6963 57916 6975 57919
rect 7377 57919 7435 57925
rect 6963 57888 7236 57916
rect 6963 57885 6975 57888
rect 6917 57879 6975 57885
rect 7208 57792 7236 57888
rect 7377 57885 7389 57919
rect 7423 57916 7435 57919
rect 7558 57916 7564 57928
rect 7423 57888 7564 57916
rect 7423 57885 7435 57888
rect 7377 57879 7435 57885
rect 7558 57876 7564 57888
rect 7616 57876 7622 57928
rect 7742 57876 7748 57928
rect 7800 57916 7806 57928
rect 8021 57919 8079 57925
rect 8021 57916 8033 57919
rect 7800 57888 8033 57916
rect 7800 57876 7806 57888
rect 8021 57885 8033 57888
rect 8067 57885 8079 57919
rect 8021 57879 8079 57885
rect 8113 57919 8171 57925
rect 8113 57885 8125 57919
rect 8159 57916 8171 57919
rect 8312 57916 8340 57944
rect 8159 57888 8340 57916
rect 8573 57919 8631 57925
rect 8159 57885 8171 57888
rect 8113 57879 8171 57885
rect 8573 57885 8585 57919
rect 8619 57885 8631 57919
rect 8573 57879 8631 57885
rect 8202 57808 8208 57860
rect 8260 57848 8266 57860
rect 8588 57848 8616 57879
rect 8260 57820 8616 57848
rect 8260 57808 8266 57820
rect 8588 57792 8616 57820
rect 1578 57740 1584 57792
rect 1636 57740 1642 57792
rect 5442 57740 5448 57792
rect 5500 57780 5506 57792
rect 6086 57780 6092 57792
rect 5500 57752 6092 57780
rect 5500 57740 5506 57752
rect 6086 57740 6092 57752
rect 6144 57740 6150 57792
rect 7190 57740 7196 57792
rect 7248 57740 7254 57792
rect 7282 57740 7288 57792
rect 7340 57780 7346 57792
rect 7561 57783 7619 57789
rect 7561 57780 7573 57783
rect 7340 57752 7573 57780
rect 7340 57740 7346 57752
rect 7561 57749 7573 57752
rect 7607 57749 7619 57783
rect 7561 57743 7619 57749
rect 8570 57740 8576 57792
rect 8628 57740 8634 57792
rect 8680 57789 8708 57956
rect 8941 57919 8999 57925
rect 8941 57885 8953 57919
rect 8987 57916 8999 57919
rect 11238 57916 11244 57928
rect 8987 57888 11244 57916
rect 8987 57885 8999 57888
rect 8941 57879 8999 57885
rect 11238 57876 11244 57888
rect 11296 57876 11302 57928
rect 8665 57783 8723 57789
rect 8665 57749 8677 57783
rect 8711 57780 8723 57783
rect 8846 57780 8852 57792
rect 8711 57752 8852 57780
rect 8711 57749 8723 57752
rect 8665 57743 8723 57749
rect 8846 57740 8852 57752
rect 8904 57740 8910 57792
rect 9122 57740 9128 57792
rect 9180 57740 9186 57792
rect 1104 57690 9936 57712
rect 1104 57638 2950 57690
rect 3002 57638 3014 57690
rect 3066 57638 3078 57690
rect 3130 57638 3142 57690
rect 3194 57638 3206 57690
rect 3258 57638 4550 57690
rect 4602 57638 4614 57690
rect 4666 57638 4678 57690
rect 4730 57638 4742 57690
rect 4794 57638 4806 57690
rect 4858 57638 6150 57690
rect 6202 57638 6214 57690
rect 6266 57638 6278 57690
rect 6330 57638 6342 57690
rect 6394 57638 6406 57690
rect 6458 57638 7750 57690
rect 7802 57638 7814 57690
rect 7866 57638 7878 57690
rect 7930 57638 7942 57690
rect 7994 57638 8006 57690
rect 8058 57638 9350 57690
rect 9402 57638 9414 57690
rect 9466 57638 9478 57690
rect 9530 57638 9542 57690
rect 9594 57638 9606 57690
rect 9658 57638 9936 57690
rect 1104 57616 9936 57638
rect 2590 57536 2596 57588
rect 2648 57576 2654 57588
rect 2648 57548 2774 57576
rect 2648 57536 2654 57548
rect 2746 57372 2774 57548
rect 4154 57536 4160 57588
rect 4212 57576 4218 57588
rect 4341 57579 4399 57585
rect 4341 57576 4353 57579
rect 4212 57548 4353 57576
rect 4212 57536 4218 57548
rect 4341 57545 4353 57548
rect 4387 57545 4399 57579
rect 4341 57539 4399 57545
rect 5166 57536 5172 57588
rect 5224 57576 5230 57588
rect 6270 57576 6276 57588
rect 5224 57548 6276 57576
rect 5224 57536 5230 57548
rect 6270 57536 6276 57548
rect 6328 57536 6334 57588
rect 6362 57536 6368 57588
rect 6420 57576 6426 57588
rect 6546 57576 6552 57588
rect 6420 57548 6552 57576
rect 6420 57536 6426 57548
rect 6546 57536 6552 57548
rect 6604 57536 6610 57588
rect 4430 57468 4436 57520
rect 4488 57508 4494 57520
rect 4890 57508 4896 57520
rect 4488 57480 4896 57508
rect 4488 57468 4494 57480
rect 4890 57468 4896 57480
rect 4948 57468 4954 57520
rect 7098 57508 7104 57520
rect 6288 57480 7104 57508
rect 3881 57443 3939 57449
rect 3881 57409 3893 57443
rect 3927 57440 3939 57443
rect 4448 57440 4476 57468
rect 3927 57412 4476 57440
rect 4709 57443 4767 57449
rect 3927 57409 3939 57412
rect 3881 57403 3939 57409
rect 4709 57409 4721 57443
rect 4755 57440 4767 57443
rect 6288 57440 6316 57480
rect 7098 57468 7104 57480
rect 7156 57468 7162 57520
rect 4755 57412 6316 57440
rect 4755 57409 4767 57412
rect 4709 57403 4767 57409
rect 6362 57400 6368 57452
rect 6420 57400 6426 57452
rect 6621 57443 6679 57449
rect 6621 57440 6633 57443
rect 6472 57412 6633 57440
rect 6472 57372 6500 57412
rect 6621 57409 6633 57412
rect 6667 57409 6679 57443
rect 6621 57403 6679 57409
rect 7190 57400 7196 57452
rect 7248 57440 7254 57452
rect 8021 57443 8079 57449
rect 7248 57412 7604 57440
rect 7248 57400 7254 57412
rect 7576 57384 7604 57412
rect 8021 57409 8033 57443
rect 8067 57440 8079 57443
rect 8938 57440 8944 57452
rect 8067 57412 8944 57440
rect 8067 57409 8079 57412
rect 8021 57403 8079 57409
rect 8938 57400 8944 57412
rect 8996 57400 9002 57452
rect 2746 57344 6500 57372
rect 6380 57316 6408 57344
rect 7558 57332 7564 57384
rect 7616 57372 7622 57384
rect 7837 57375 7895 57381
rect 7837 57372 7849 57375
rect 7616 57344 7849 57372
rect 7616 57332 7622 57344
rect 7837 57341 7849 57344
rect 7883 57341 7895 57375
rect 7837 57335 7895 57341
rect 4338 57304 4344 57316
rect 4080 57276 4344 57304
rect 4080 57245 4108 57276
rect 4338 57264 4344 57276
rect 4396 57264 4402 57316
rect 4430 57264 4436 57316
rect 4488 57304 4494 57316
rect 5350 57304 5356 57316
rect 4488 57276 5356 57304
rect 4488 57264 4494 57276
rect 5350 57264 5356 57276
rect 5408 57264 5414 57316
rect 5626 57264 5632 57316
rect 5684 57264 5690 57316
rect 6362 57264 6368 57316
rect 6420 57264 6426 57316
rect 7374 57264 7380 57316
rect 7432 57304 7438 57316
rect 8205 57307 8263 57313
rect 8205 57304 8217 57307
rect 7432 57276 8217 57304
rect 7432 57264 7438 57276
rect 8205 57273 8217 57276
rect 8251 57273 8263 57307
rect 8205 57267 8263 57273
rect 8570 57264 8576 57316
rect 8628 57304 8634 57316
rect 8938 57304 8944 57316
rect 8628 57276 8944 57304
rect 8628 57264 8634 57276
rect 8938 57264 8944 57276
rect 8996 57264 9002 57316
rect 4065 57239 4123 57245
rect 4065 57205 4077 57239
rect 4111 57205 4123 57239
rect 4065 57199 4123 57205
rect 4246 57196 4252 57248
rect 4304 57236 4310 57248
rect 4525 57239 4583 57245
rect 4525 57236 4537 57239
rect 4304 57208 4537 57236
rect 4304 57196 4310 57208
rect 4525 57205 4537 57208
rect 4571 57205 4583 57239
rect 5644 57236 5672 57264
rect 7745 57239 7803 57245
rect 7745 57236 7757 57239
rect 5644 57208 7757 57236
rect 4525 57199 4583 57205
rect 7745 57205 7757 57208
rect 7791 57205 7803 57239
rect 7745 57199 7803 57205
rect 1104 57146 9936 57168
rect 1104 57094 3610 57146
rect 3662 57094 3674 57146
rect 3726 57094 3738 57146
rect 3790 57094 3802 57146
rect 3854 57094 3866 57146
rect 3918 57094 5210 57146
rect 5262 57094 5274 57146
rect 5326 57094 5338 57146
rect 5390 57094 5402 57146
rect 5454 57094 5466 57146
rect 5518 57094 6810 57146
rect 6862 57094 6874 57146
rect 6926 57094 6938 57146
rect 6990 57094 7002 57146
rect 7054 57094 7066 57146
rect 7118 57094 8410 57146
rect 8462 57094 8474 57146
rect 8526 57094 8538 57146
rect 8590 57094 8602 57146
rect 8654 57094 8666 57146
rect 8718 57094 9936 57146
rect 1104 57072 9936 57094
rect 6270 56856 6276 56908
rect 6328 56896 6334 56908
rect 6822 56896 6828 56908
rect 6328 56868 6828 56896
rect 6328 56856 6334 56868
rect 6822 56856 6828 56868
rect 6880 56856 6886 56908
rect 1489 56831 1547 56837
rect 1489 56797 1501 56831
rect 1535 56828 1547 56831
rect 3510 56828 3516 56840
rect 1535 56800 3516 56828
rect 1535 56797 1547 56800
rect 1489 56791 1547 56797
rect 3510 56788 3516 56800
rect 3568 56788 3574 56840
rect 4157 56831 4215 56837
rect 4157 56797 4169 56831
rect 4203 56828 4215 56831
rect 6730 56828 6736 56840
rect 4203 56800 6736 56828
rect 4203 56797 4215 56800
rect 4157 56791 4215 56797
rect 6730 56788 6736 56800
rect 6788 56788 6794 56840
rect 7561 56831 7619 56837
rect 7561 56797 7573 56831
rect 7607 56828 7619 56831
rect 9214 56828 9220 56840
rect 7607 56800 9220 56828
rect 7607 56797 7619 56800
rect 7561 56791 7619 56797
rect 9214 56788 9220 56800
rect 9272 56788 9278 56840
rect 6638 56720 6644 56772
rect 6696 56760 6702 56772
rect 11054 56760 11060 56772
rect 6696 56732 11060 56760
rect 6696 56720 6702 56732
rect 11054 56720 11060 56732
rect 11112 56720 11118 56772
rect 934 56652 940 56704
rect 992 56692 998 56704
rect 1581 56695 1639 56701
rect 1581 56692 1593 56695
rect 992 56664 1593 56692
rect 992 56652 998 56664
rect 1581 56661 1593 56664
rect 1627 56661 1639 56695
rect 1581 56655 1639 56661
rect 3510 56652 3516 56704
rect 3568 56692 3574 56704
rect 4341 56695 4399 56701
rect 4341 56692 4353 56695
rect 3568 56664 4353 56692
rect 3568 56652 3574 56664
rect 4341 56661 4353 56664
rect 4387 56661 4399 56695
rect 4341 56655 4399 56661
rect 6362 56652 6368 56704
rect 6420 56692 6426 56704
rect 6730 56692 6736 56704
rect 6420 56664 6736 56692
rect 6420 56652 6426 56664
rect 6730 56652 6736 56664
rect 6788 56652 6794 56704
rect 7190 56652 7196 56704
rect 7248 56692 7254 56704
rect 7745 56695 7803 56701
rect 7745 56692 7757 56695
rect 7248 56664 7757 56692
rect 7248 56652 7254 56664
rect 7745 56661 7757 56664
rect 7791 56661 7803 56695
rect 7745 56655 7803 56661
rect 1104 56602 9936 56624
rect 1104 56550 2950 56602
rect 3002 56550 3014 56602
rect 3066 56550 3078 56602
rect 3130 56550 3142 56602
rect 3194 56550 3206 56602
rect 3258 56550 4550 56602
rect 4602 56550 4614 56602
rect 4666 56550 4678 56602
rect 4730 56550 4742 56602
rect 4794 56550 4806 56602
rect 4858 56550 6150 56602
rect 6202 56550 6214 56602
rect 6266 56550 6278 56602
rect 6330 56550 6342 56602
rect 6394 56550 6406 56602
rect 6458 56550 7750 56602
rect 7802 56550 7814 56602
rect 7866 56550 7878 56602
rect 7930 56550 7942 56602
rect 7994 56550 8006 56602
rect 8058 56550 9350 56602
rect 9402 56550 9414 56602
rect 9466 56550 9478 56602
rect 9530 56550 9542 56602
rect 9594 56550 9606 56602
rect 9658 56550 9936 56602
rect 1104 56528 9936 56550
rect 7561 56491 7619 56497
rect 7561 56457 7573 56491
rect 7607 56488 7619 56491
rect 7650 56488 7656 56500
rect 7607 56460 7656 56488
rect 7607 56457 7619 56460
rect 7561 56451 7619 56457
rect 7650 56448 7656 56460
rect 7708 56448 7714 56500
rect 1489 56423 1547 56429
rect 1489 56389 1501 56423
rect 1535 56420 1547 56423
rect 3326 56420 3332 56432
rect 1535 56392 3332 56420
rect 1535 56389 1547 56392
rect 1489 56383 1547 56389
rect 3326 56380 3332 56392
rect 3384 56380 3390 56432
rect 4249 56355 4307 56361
rect 4249 56321 4261 56355
rect 4295 56352 4307 56355
rect 4430 56352 4436 56364
rect 4295 56324 4436 56352
rect 4295 56321 4307 56324
rect 4249 56315 4307 56321
rect 4430 56312 4436 56324
rect 4488 56312 4494 56364
rect 4709 56355 4767 56361
rect 4709 56321 4721 56355
rect 4755 56352 4767 56355
rect 4982 56352 4988 56364
rect 4755 56324 4988 56352
rect 4755 56321 4767 56324
rect 4709 56315 4767 56321
rect 4982 56312 4988 56324
rect 5040 56312 5046 56364
rect 5074 56312 5080 56364
rect 5132 56312 5138 56364
rect 7469 56355 7527 56361
rect 7469 56321 7481 56355
rect 7515 56352 7527 56355
rect 8846 56352 8852 56364
rect 7515 56324 8852 56352
rect 7515 56321 7527 56324
rect 7469 56315 7527 56321
rect 8846 56312 8852 56324
rect 8904 56312 8910 56364
rect 3326 56244 3332 56296
rect 3384 56284 3390 56296
rect 3510 56284 3516 56296
rect 3384 56256 3516 56284
rect 3384 56244 3390 56256
rect 3510 56244 3516 56256
rect 3568 56244 3574 56296
rect 1486 56176 1492 56228
rect 1544 56216 1550 56228
rect 4525 56219 4583 56225
rect 4525 56216 4537 56219
rect 1544 56188 4537 56216
rect 1544 56176 1550 56188
rect 4525 56185 4537 56188
rect 4571 56185 4583 56219
rect 4525 56179 4583 56185
rect 5092 56160 5120 56312
rect 6638 56244 6644 56296
rect 6696 56284 6702 56296
rect 8202 56284 8208 56296
rect 6696 56256 8208 56284
rect 6696 56244 6702 56256
rect 8202 56244 8208 56256
rect 8260 56244 8266 56296
rect 934 56108 940 56160
rect 992 56148 998 56160
rect 1581 56151 1639 56157
rect 1581 56148 1593 56151
rect 992 56120 1593 56148
rect 992 56108 998 56120
rect 1581 56117 1593 56120
rect 1627 56117 1639 56151
rect 1581 56111 1639 56117
rect 2682 56108 2688 56160
rect 2740 56148 2746 56160
rect 4433 56151 4491 56157
rect 4433 56148 4445 56151
rect 2740 56120 4445 56148
rect 2740 56108 2746 56120
rect 4433 56117 4445 56120
rect 4479 56117 4491 56151
rect 4433 56111 4491 56117
rect 5074 56108 5080 56160
rect 5132 56108 5138 56160
rect 6822 56108 6828 56160
rect 6880 56148 6886 56160
rect 7650 56148 7656 56160
rect 6880 56120 7656 56148
rect 6880 56108 6886 56120
rect 7650 56108 7656 56120
rect 7708 56108 7714 56160
rect 1104 56058 9936 56080
rect 1104 56006 3610 56058
rect 3662 56006 3674 56058
rect 3726 56006 3738 56058
rect 3790 56006 3802 56058
rect 3854 56006 3866 56058
rect 3918 56006 5210 56058
rect 5262 56006 5274 56058
rect 5326 56006 5338 56058
rect 5390 56006 5402 56058
rect 5454 56006 5466 56058
rect 5518 56006 6810 56058
rect 6862 56006 6874 56058
rect 6926 56006 6938 56058
rect 6990 56006 7002 56058
rect 7054 56006 7066 56058
rect 7118 56006 8410 56058
rect 8462 56006 8474 56058
rect 8526 56006 8538 56058
rect 8590 56006 8602 56058
rect 8654 56006 8666 56058
rect 8718 56006 9936 56058
rect 1104 55984 9936 56006
rect 1210 55904 1216 55956
rect 1268 55944 1274 55956
rect 4157 55947 4215 55953
rect 4157 55944 4169 55947
rect 1268 55916 4169 55944
rect 1268 55904 1274 55916
rect 4157 55913 4169 55916
rect 4203 55913 4215 55947
rect 4157 55907 4215 55913
rect 2130 55836 2136 55888
rect 2188 55876 2194 55888
rect 9674 55876 9680 55888
rect 2188 55848 9680 55876
rect 2188 55836 2194 55848
rect 9674 55836 9680 55848
rect 9732 55836 9738 55888
rect 8202 55808 8208 55820
rect 7208 55780 8208 55808
rect 7208 55749 7236 55780
rect 8202 55768 8208 55780
rect 8260 55768 8266 55820
rect 7101 55743 7159 55749
rect 7101 55709 7113 55743
rect 7147 55709 7159 55743
rect 7101 55703 7159 55709
rect 7193 55743 7251 55749
rect 7193 55709 7205 55743
rect 7239 55709 7251 55743
rect 7193 55703 7251 55709
rect 4065 55675 4123 55681
rect 4065 55641 4077 55675
rect 4111 55672 4123 55675
rect 4430 55672 4436 55684
rect 4111 55644 4436 55672
rect 4111 55641 4123 55644
rect 4065 55635 4123 55641
rect 4430 55632 4436 55644
rect 4488 55632 4494 55684
rect 7116 55672 7144 55703
rect 7558 55700 7564 55752
rect 7616 55700 7622 55752
rect 7653 55743 7711 55749
rect 7653 55709 7665 55743
rect 7699 55740 7711 55743
rect 8110 55740 8116 55752
rect 7699 55712 8116 55740
rect 7699 55709 7711 55712
rect 7653 55703 7711 55709
rect 8110 55700 8116 55712
rect 8168 55700 8174 55752
rect 7576 55672 7604 55700
rect 7116 55644 7604 55672
rect 5534 55564 5540 55616
rect 5592 55604 5598 55616
rect 7377 55607 7435 55613
rect 7377 55604 7389 55607
rect 5592 55576 7389 55604
rect 5592 55564 5598 55576
rect 7377 55573 7389 55576
rect 7423 55573 7435 55607
rect 7377 55567 7435 55573
rect 7837 55607 7895 55613
rect 7837 55573 7849 55607
rect 7883 55604 7895 55607
rect 8202 55604 8208 55616
rect 7883 55576 8208 55604
rect 7883 55573 7895 55576
rect 7837 55567 7895 55573
rect 8202 55564 8208 55576
rect 8260 55564 8266 55616
rect 1104 55514 9936 55536
rect 1104 55462 2950 55514
rect 3002 55462 3014 55514
rect 3066 55462 3078 55514
rect 3130 55462 3142 55514
rect 3194 55462 3206 55514
rect 3258 55462 4550 55514
rect 4602 55462 4614 55514
rect 4666 55462 4678 55514
rect 4730 55462 4742 55514
rect 4794 55462 4806 55514
rect 4858 55462 6150 55514
rect 6202 55462 6214 55514
rect 6266 55462 6278 55514
rect 6330 55462 6342 55514
rect 6394 55462 6406 55514
rect 6458 55462 7750 55514
rect 7802 55462 7814 55514
rect 7866 55462 7878 55514
rect 7930 55462 7942 55514
rect 7994 55462 8006 55514
rect 8058 55462 9350 55514
rect 9402 55462 9414 55514
rect 9466 55462 9478 55514
rect 9530 55462 9542 55514
rect 9594 55462 9606 55514
rect 9658 55462 9936 55514
rect 1104 55440 9936 55462
rect 7558 55360 7564 55412
rect 7616 55400 7622 55412
rect 8110 55400 8116 55412
rect 7616 55372 8116 55400
rect 7616 55360 7622 55372
rect 8110 55360 8116 55372
rect 8168 55360 8174 55412
rect 1489 55335 1547 55341
rect 1489 55301 1501 55335
rect 1535 55332 1547 55335
rect 2406 55332 2412 55344
rect 1535 55304 2412 55332
rect 1535 55301 1547 55304
rect 1489 55295 1547 55301
rect 2406 55292 2412 55304
rect 2464 55292 2470 55344
rect 9674 55224 9680 55276
rect 9732 55264 9738 55276
rect 9858 55264 9864 55276
rect 9732 55236 9864 55264
rect 9732 55224 9738 55236
rect 9858 55224 9864 55236
rect 9916 55224 9922 55276
rect 934 55020 940 55072
rect 992 55060 998 55072
rect 1581 55063 1639 55069
rect 1581 55060 1593 55063
rect 992 55032 1593 55060
rect 992 55020 998 55032
rect 1581 55029 1593 55032
rect 1627 55029 1639 55063
rect 1581 55023 1639 55029
rect 1104 54970 9936 54992
rect 1104 54918 3610 54970
rect 3662 54918 3674 54970
rect 3726 54918 3738 54970
rect 3790 54918 3802 54970
rect 3854 54918 3866 54970
rect 3918 54918 5210 54970
rect 5262 54918 5274 54970
rect 5326 54918 5338 54970
rect 5390 54918 5402 54970
rect 5454 54918 5466 54970
rect 5518 54918 6810 54970
rect 6862 54918 6874 54970
rect 6926 54918 6938 54970
rect 6990 54918 7002 54970
rect 7054 54918 7066 54970
rect 7118 54918 8410 54970
rect 8462 54918 8474 54970
rect 8526 54918 8538 54970
rect 8590 54918 8602 54970
rect 8654 54918 8666 54970
rect 8718 54918 9936 54970
rect 1104 54896 9936 54918
rect 4433 54655 4491 54661
rect 4433 54621 4445 54655
rect 4479 54652 4491 54655
rect 6638 54652 6644 54664
rect 4479 54624 6644 54652
rect 4479 54621 4491 54624
rect 4433 54615 4491 54621
rect 6638 54612 6644 54624
rect 6696 54612 6702 54664
rect 6733 54655 6791 54661
rect 6733 54621 6745 54655
rect 6779 54652 6791 54655
rect 8938 54652 8944 54664
rect 6779 54624 8944 54652
rect 6779 54621 6791 54624
rect 6733 54615 6791 54621
rect 8938 54612 8944 54624
rect 8996 54612 9002 54664
rect 6917 54587 6975 54593
rect 6917 54553 6929 54587
rect 6963 54584 6975 54587
rect 9214 54584 9220 54596
rect 6963 54556 9220 54584
rect 6963 54553 6975 54556
rect 6917 54547 6975 54553
rect 9214 54544 9220 54556
rect 9272 54544 9278 54596
rect 2866 54476 2872 54528
rect 2924 54516 2930 54528
rect 4249 54519 4307 54525
rect 4249 54516 4261 54519
rect 2924 54488 4261 54516
rect 2924 54476 2930 54488
rect 4249 54485 4261 54488
rect 4295 54485 4307 54519
rect 4249 54479 4307 54485
rect 1104 54426 9936 54448
rect 1104 54374 2950 54426
rect 3002 54374 3014 54426
rect 3066 54374 3078 54426
rect 3130 54374 3142 54426
rect 3194 54374 3206 54426
rect 3258 54374 4550 54426
rect 4602 54374 4614 54426
rect 4666 54374 4678 54426
rect 4730 54374 4742 54426
rect 4794 54374 4806 54426
rect 4858 54374 6150 54426
rect 6202 54374 6214 54426
rect 6266 54374 6278 54426
rect 6330 54374 6342 54426
rect 6394 54374 6406 54426
rect 6458 54374 7750 54426
rect 7802 54374 7814 54426
rect 7866 54374 7878 54426
rect 7930 54374 7942 54426
rect 7994 54374 8006 54426
rect 8058 54374 9350 54426
rect 9402 54374 9414 54426
rect 9466 54374 9478 54426
rect 9530 54374 9542 54426
rect 9594 54374 9606 54426
rect 9658 54374 9936 54426
rect 1104 54352 9936 54374
rect 9674 54312 9680 54324
rect 7300 54284 9680 54312
rect 1394 54204 1400 54256
rect 1452 54244 1458 54256
rect 1489 54247 1547 54253
rect 1489 54244 1501 54247
rect 1452 54216 1501 54244
rect 1452 54204 1458 54216
rect 1489 54213 1501 54216
rect 1535 54213 1547 54247
rect 5810 54244 5816 54256
rect 1489 54207 1547 54213
rect 4448 54216 5816 54244
rect 4448 54185 4476 54216
rect 5810 54204 5816 54216
rect 5868 54204 5874 54256
rect 4433 54179 4491 54185
rect 4433 54145 4445 54179
rect 4479 54145 4491 54179
rect 4433 54139 4491 54145
rect 4525 54179 4583 54185
rect 4525 54145 4537 54179
rect 4571 54176 4583 54179
rect 5994 54176 6000 54188
rect 4571 54148 6000 54176
rect 4571 54145 4583 54148
rect 4525 54139 4583 54145
rect 5994 54136 6000 54148
rect 6052 54136 6058 54188
rect 6638 54136 6644 54188
rect 6696 54176 6702 54188
rect 7193 54179 7251 54185
rect 7193 54176 7205 54179
rect 6696 54148 7205 54176
rect 6696 54136 6702 54148
rect 2590 54000 2596 54052
rect 2648 54040 2654 54052
rect 4709 54043 4767 54049
rect 4709 54040 4721 54043
rect 2648 54012 4721 54040
rect 2648 54000 2654 54012
rect 4709 54009 4721 54012
rect 4755 54009 4767 54043
rect 7024 54040 7052 54148
rect 7193 54145 7205 54148
rect 7239 54145 7251 54179
rect 7300 54176 7328 54284
rect 9674 54272 9680 54284
rect 9732 54312 9738 54324
rect 9732 54284 10824 54312
rect 9732 54272 9738 54284
rect 10796 54256 10824 54284
rect 7377 54247 7435 54253
rect 7377 54213 7389 54247
rect 7423 54244 7435 54247
rect 7466 54244 7472 54256
rect 7423 54216 7472 54244
rect 7423 54213 7435 54216
rect 7377 54207 7435 54213
rect 7466 54204 7472 54216
rect 7524 54244 7530 54256
rect 7524 54216 8984 54244
rect 7524 54204 7530 54216
rect 8956 54188 8984 54216
rect 10778 54204 10784 54256
rect 10836 54204 10842 54256
rect 7653 54179 7711 54185
rect 7653 54176 7665 54179
rect 7300 54148 7665 54176
rect 7193 54139 7251 54145
rect 7653 54145 7665 54148
rect 7699 54145 7711 54179
rect 7834 54176 7840 54188
rect 7795 54148 7840 54176
rect 7653 54139 7711 54145
rect 7834 54136 7840 54148
rect 7892 54136 7898 54188
rect 8938 54136 8944 54188
rect 8996 54136 9002 54188
rect 11514 54040 11520 54052
rect 7024 54012 11520 54040
rect 4709 54003 4767 54009
rect 11514 54000 11520 54012
rect 11572 54000 11578 54052
rect 934 53932 940 53984
rect 992 53972 998 53984
rect 1581 53975 1639 53981
rect 1581 53972 1593 53975
rect 992 53944 1593 53972
rect 992 53932 998 53944
rect 1581 53941 1593 53944
rect 1627 53941 1639 53975
rect 1581 53935 1639 53941
rect 2682 53932 2688 53984
rect 2740 53972 2746 53984
rect 4249 53975 4307 53981
rect 4249 53972 4261 53975
rect 2740 53944 4261 53972
rect 2740 53932 2746 53944
rect 4249 53941 4261 53944
rect 4295 53941 4307 53975
rect 4249 53935 4307 53941
rect 7558 53932 7564 53984
rect 7616 53932 7622 53984
rect 7650 53932 7656 53984
rect 7708 53972 7714 53984
rect 8021 53975 8079 53981
rect 8021 53972 8033 53975
rect 7708 53944 8033 53972
rect 7708 53932 7714 53944
rect 8021 53941 8033 53944
rect 8067 53941 8079 53975
rect 8021 53935 8079 53941
rect 1104 53882 9936 53904
rect 1104 53830 3610 53882
rect 3662 53830 3674 53882
rect 3726 53830 3738 53882
rect 3790 53830 3802 53882
rect 3854 53830 3866 53882
rect 3918 53830 5210 53882
rect 5262 53830 5274 53882
rect 5326 53830 5338 53882
rect 5390 53830 5402 53882
rect 5454 53830 5466 53882
rect 5518 53830 6810 53882
rect 6862 53830 6874 53882
rect 6926 53830 6938 53882
rect 6990 53830 7002 53882
rect 7054 53830 7066 53882
rect 7118 53830 8410 53882
rect 8462 53830 8474 53882
rect 8526 53830 8538 53882
rect 8590 53830 8602 53882
rect 8654 53830 8666 53882
rect 8718 53830 9936 53882
rect 1104 53808 9936 53830
rect 4890 53728 4896 53780
rect 4948 53768 4954 53780
rect 4985 53771 5043 53777
rect 4985 53768 4997 53771
rect 4948 53740 4997 53768
rect 4948 53728 4954 53740
rect 4985 53737 4997 53740
rect 5031 53737 5043 53771
rect 4985 53731 5043 53737
rect 7006 53728 7012 53780
rect 7064 53768 7070 53780
rect 10226 53768 10232 53780
rect 7064 53740 10232 53768
rect 7064 53728 7070 53740
rect 10226 53728 10232 53740
rect 10284 53728 10290 53780
rect 11422 53728 11428 53780
rect 11480 53728 11486 53780
rect 4798 53660 4804 53712
rect 4856 53700 4862 53712
rect 7024 53700 7052 53728
rect 11440 53700 11468 53728
rect 4856 53672 7052 53700
rect 9646 53672 11468 53700
rect 4856 53660 4862 53672
rect 9646 53632 9674 53672
rect 6932 53604 9674 53632
rect 2130 53524 2136 53576
rect 2188 53564 2194 53576
rect 4154 53564 4160 53576
rect 2188 53536 4160 53564
rect 2188 53524 2194 53536
rect 4154 53524 4160 53536
rect 4212 53524 4218 53576
rect 4430 53524 4436 53576
rect 4488 53564 4494 53576
rect 4893 53567 4951 53573
rect 4893 53564 4905 53567
rect 4488 53536 4905 53564
rect 4488 53524 4494 53536
rect 4893 53533 4905 53536
rect 4939 53533 4951 53567
rect 4893 53527 4951 53533
rect 3970 53456 3976 53508
rect 4028 53496 4034 53508
rect 6932 53496 6960 53604
rect 7098 53524 7104 53576
rect 7156 53564 7162 53576
rect 7193 53567 7251 53573
rect 7193 53564 7205 53567
rect 7156 53536 7205 53564
rect 7156 53524 7162 53536
rect 7193 53533 7205 53536
rect 7239 53564 7251 53567
rect 7282 53564 7288 53576
rect 7239 53536 7288 53564
rect 7239 53533 7251 53536
rect 7193 53527 7251 53533
rect 7282 53524 7288 53536
rect 7340 53524 7346 53576
rect 7374 53524 7380 53576
rect 7432 53524 7438 53576
rect 7742 53524 7748 53576
rect 7800 53524 7806 53576
rect 7009 53499 7067 53505
rect 7009 53496 7021 53499
rect 4028 53468 7021 53496
rect 4028 53456 4034 53468
rect 7009 53465 7021 53468
rect 7055 53465 7067 53499
rect 7392 53496 7420 53524
rect 7009 53459 7067 53465
rect 7300 53468 7420 53496
rect 3510 53388 3516 53440
rect 3568 53428 3574 53440
rect 7098 53428 7104 53440
rect 3568 53400 7104 53428
rect 3568 53388 3574 53400
rect 7098 53388 7104 53400
rect 7156 53428 7162 53440
rect 7300 53428 7328 53468
rect 7156 53400 7328 53428
rect 7156 53388 7162 53400
rect 7374 53388 7380 53440
rect 7432 53388 7438 53440
rect 7466 53388 7472 53440
rect 7524 53428 7530 53440
rect 7929 53431 7987 53437
rect 7929 53428 7941 53431
rect 7524 53400 7941 53428
rect 7524 53388 7530 53400
rect 7929 53397 7941 53400
rect 7975 53397 7987 53431
rect 7929 53391 7987 53397
rect 1104 53338 9936 53360
rect 1104 53286 2950 53338
rect 3002 53286 3014 53338
rect 3066 53286 3078 53338
rect 3130 53286 3142 53338
rect 3194 53286 3206 53338
rect 3258 53286 4550 53338
rect 4602 53286 4614 53338
rect 4666 53286 4678 53338
rect 4730 53286 4742 53338
rect 4794 53286 4806 53338
rect 4858 53286 6150 53338
rect 6202 53286 6214 53338
rect 6266 53286 6278 53338
rect 6330 53286 6342 53338
rect 6394 53286 6406 53338
rect 6458 53286 7750 53338
rect 7802 53286 7814 53338
rect 7866 53286 7878 53338
rect 7930 53286 7942 53338
rect 7994 53286 8006 53338
rect 8058 53286 9350 53338
rect 9402 53286 9414 53338
rect 9466 53286 9478 53338
rect 9530 53286 9542 53338
rect 9594 53286 9606 53338
rect 9658 53286 9936 53338
rect 1104 53264 9936 53286
rect 5718 53184 5724 53236
rect 5776 53184 5782 53236
rect 7006 53184 7012 53236
rect 7064 53184 7070 53236
rect 7190 53184 7196 53236
rect 7248 53224 7254 53236
rect 7248 53196 7328 53224
rect 7248 53184 7254 53196
rect 1489 53159 1547 53165
rect 1489 53125 1501 53159
rect 1535 53156 1547 53159
rect 2774 53156 2780 53168
rect 1535 53128 2780 53156
rect 1535 53125 1547 53128
rect 1489 53119 1547 53125
rect 2774 53116 2780 53128
rect 2832 53116 2838 53168
rect 4525 53159 4583 53165
rect 4525 53125 4537 53159
rect 4571 53156 4583 53159
rect 5074 53156 5080 53168
rect 4571 53128 5080 53156
rect 4571 53125 4583 53128
rect 4525 53119 4583 53125
rect 5074 53116 5080 53128
rect 5132 53116 5138 53168
rect 750 53048 756 53100
rect 808 53088 814 53100
rect 4154 53088 4160 53100
rect 808 53060 4160 53088
rect 808 53048 814 53060
rect 4154 53048 4160 53060
rect 4212 53088 4218 53100
rect 4341 53091 4399 53097
rect 4341 53088 4353 53091
rect 4212 53060 4353 53088
rect 4212 53048 4218 53060
rect 4341 53057 4353 53060
rect 4387 53057 4399 53091
rect 4798 53088 4804 53100
rect 4341 53051 4399 53057
rect 4448 53060 4804 53088
rect 1118 52980 1124 53032
rect 1176 53020 1182 53032
rect 4448 53020 4476 53060
rect 4798 53048 4804 53060
rect 4856 53048 4862 53100
rect 4985 53091 5043 53097
rect 4985 53057 4997 53091
rect 5031 53088 5043 53091
rect 5736 53088 5764 53184
rect 5031 53060 5764 53088
rect 5031 53057 5043 53060
rect 4985 53051 5043 53057
rect 1176 52992 4476 53020
rect 4709 53023 4767 53029
rect 1176 52980 1182 52992
rect 4709 52989 4721 53023
rect 4755 53020 4767 53023
rect 5626 53020 5632 53032
rect 4755 52992 5632 53020
rect 4755 52989 4767 52992
rect 4709 52983 4767 52989
rect 5626 52980 5632 52992
rect 5684 52980 5690 53032
rect 2774 52912 2780 52964
rect 2832 52952 2838 52964
rect 3786 52952 3792 52964
rect 2832 52924 3792 52952
rect 2832 52912 2838 52924
rect 3786 52912 3792 52924
rect 3844 52912 3850 52964
rect 5736 52952 5764 53060
rect 6454 53048 6460 53100
rect 6512 53088 6518 53100
rect 6638 53088 6644 53100
rect 6512 53060 6644 53088
rect 6512 53048 6518 53060
rect 6638 53048 6644 53060
rect 6696 53048 6702 53100
rect 7024 53097 7052 53184
rect 7098 53116 7104 53168
rect 7156 53116 7162 53168
rect 7009 53091 7067 53097
rect 7009 53057 7021 53091
rect 7055 53057 7067 53091
rect 7116 53088 7144 53116
rect 7193 53091 7251 53097
rect 7193 53088 7205 53091
rect 7116 53060 7205 53088
rect 7009 53051 7067 53057
rect 7193 53057 7205 53060
rect 7239 53057 7251 53091
rect 7193 53051 7251 53057
rect 7300 52964 7328 53196
rect 7374 53184 7380 53236
rect 7432 53184 7438 53236
rect 7558 53184 7564 53236
rect 7616 53224 7622 53236
rect 7616 53196 8248 53224
rect 7616 53184 7622 53196
rect 7392 53156 7420 53184
rect 7392 53128 7972 53156
rect 7650 53048 7656 53100
rect 7708 53048 7714 53100
rect 7944 53097 7972 53128
rect 8220 53097 8248 53196
rect 9766 53116 9772 53168
rect 9824 53156 9830 53168
rect 10042 53156 10048 53168
rect 9824 53128 10048 53156
rect 9824 53116 9830 53128
rect 10042 53116 10048 53128
rect 10100 53116 10106 53168
rect 7929 53091 7987 53097
rect 7929 53057 7941 53091
rect 7975 53057 7987 53091
rect 7929 53051 7987 53057
rect 8205 53091 8263 53097
rect 8205 53057 8217 53091
rect 8251 53057 8263 53091
rect 8205 53051 8263 53057
rect 7377 53023 7435 53029
rect 7377 52989 7389 53023
rect 7423 53020 7435 53023
rect 8294 53020 8300 53032
rect 7423 52992 8300 53020
rect 7423 52989 7435 52992
rect 7377 52983 7435 52989
rect 8294 52980 8300 52992
rect 8352 52980 8358 53032
rect 4540 52924 5764 52952
rect 934 52844 940 52896
rect 992 52884 998 52896
rect 1581 52887 1639 52893
rect 1581 52884 1593 52887
rect 992 52856 1593 52884
rect 992 52844 998 52856
rect 1581 52853 1593 52856
rect 1627 52853 1639 52887
rect 1581 52847 1639 52853
rect 2406 52844 2412 52896
rect 2464 52884 2470 52896
rect 4540 52884 4568 52924
rect 7282 52912 7288 52964
rect 7340 52912 7346 52964
rect 7558 52912 7564 52964
rect 7616 52952 7622 52964
rect 8021 52955 8079 52961
rect 8021 52952 8033 52955
rect 7616 52924 8033 52952
rect 7616 52912 7622 52924
rect 8021 52921 8033 52924
rect 8067 52921 8079 52955
rect 8021 52915 8079 52921
rect 2464 52856 4568 52884
rect 2464 52844 2470 52856
rect 4798 52844 4804 52896
rect 4856 52884 4862 52896
rect 5074 52884 5080 52896
rect 4856 52856 5080 52884
rect 4856 52844 4862 52856
rect 5074 52844 5080 52856
rect 5132 52844 5138 52896
rect 5169 52887 5227 52893
rect 5169 52853 5181 52887
rect 5215 52884 5227 52887
rect 6178 52884 6184 52896
rect 5215 52856 6184 52884
rect 5215 52853 5227 52856
rect 5169 52847 5227 52853
rect 6178 52844 6184 52856
rect 6236 52844 6242 52896
rect 7466 52844 7472 52896
rect 7524 52844 7530 52896
rect 7742 52844 7748 52896
rect 7800 52844 7806 52896
rect 1104 52794 9936 52816
rect 1104 52742 3610 52794
rect 3662 52742 3674 52794
rect 3726 52742 3738 52794
rect 3790 52742 3802 52794
rect 3854 52742 3866 52794
rect 3918 52742 5210 52794
rect 5262 52742 5274 52794
rect 5326 52742 5338 52794
rect 5390 52742 5402 52794
rect 5454 52742 5466 52794
rect 5518 52742 6810 52794
rect 6862 52742 6874 52794
rect 6926 52742 6938 52794
rect 6990 52742 7002 52794
rect 7054 52742 7066 52794
rect 7118 52742 8410 52794
rect 8462 52742 8474 52794
rect 8526 52742 8538 52794
rect 8590 52742 8602 52794
rect 8654 52742 8666 52794
rect 8718 52742 9936 52794
rect 1104 52720 9936 52742
rect 5718 52640 5724 52692
rect 5776 52680 5782 52692
rect 5902 52680 5908 52692
rect 5776 52652 5908 52680
rect 5776 52640 5782 52652
rect 5902 52640 5908 52652
rect 5960 52640 5966 52692
rect 6638 52640 6644 52692
rect 6696 52680 6702 52692
rect 6696 52652 8156 52680
rect 6696 52640 6702 52652
rect 8128 52621 8156 52652
rect 5997 52615 6055 52621
rect 5997 52581 6009 52615
rect 6043 52581 6055 52615
rect 5997 52575 6055 52581
rect 8113 52615 8171 52621
rect 8113 52581 8125 52615
rect 8159 52581 8171 52615
rect 8113 52575 8171 52581
rect 6012 52544 6040 52575
rect 6012 52516 6868 52544
rect 6178 52436 6184 52488
rect 6236 52436 6242 52488
rect 6730 52436 6736 52488
rect 6788 52436 6794 52488
rect 6840 52476 6868 52516
rect 6989 52479 7047 52485
rect 6989 52476 7001 52479
rect 6840 52448 7001 52476
rect 6989 52445 7001 52448
rect 7035 52445 7047 52479
rect 6989 52439 7047 52445
rect 1489 52411 1547 52417
rect 1489 52377 1501 52411
rect 1535 52408 1547 52411
rect 4246 52408 4252 52420
rect 1535 52380 4252 52408
rect 1535 52377 1547 52380
rect 1489 52371 1547 52377
rect 4246 52368 4252 52380
rect 4304 52368 4310 52420
rect 1578 52300 1584 52352
rect 1636 52300 1642 52352
rect 5902 52300 5908 52352
rect 5960 52340 5966 52352
rect 6454 52340 6460 52352
rect 5960 52312 6460 52340
rect 5960 52300 5966 52312
rect 6454 52300 6460 52312
rect 6512 52300 6518 52352
rect 7282 52300 7288 52352
rect 7340 52340 7346 52352
rect 7742 52340 7748 52352
rect 7340 52312 7748 52340
rect 7340 52300 7346 52312
rect 7742 52300 7748 52312
rect 7800 52300 7806 52352
rect 1104 52250 9936 52272
rect 1104 52198 2950 52250
rect 3002 52198 3014 52250
rect 3066 52198 3078 52250
rect 3130 52198 3142 52250
rect 3194 52198 3206 52250
rect 3258 52198 4550 52250
rect 4602 52198 4614 52250
rect 4666 52198 4678 52250
rect 4730 52198 4742 52250
rect 4794 52198 4806 52250
rect 4858 52198 6150 52250
rect 6202 52198 6214 52250
rect 6266 52198 6278 52250
rect 6330 52198 6342 52250
rect 6394 52198 6406 52250
rect 6458 52198 7750 52250
rect 7802 52198 7814 52250
rect 7866 52198 7878 52250
rect 7930 52198 7942 52250
rect 7994 52198 8006 52250
rect 8058 52198 9350 52250
rect 9402 52198 9414 52250
rect 9466 52198 9478 52250
rect 9530 52198 9542 52250
rect 9594 52198 9606 52250
rect 9658 52198 9936 52250
rect 1104 52176 9936 52198
rect 4798 52096 4804 52148
rect 4856 52136 4862 52148
rect 5902 52136 5908 52148
rect 4856 52108 5908 52136
rect 4856 52096 4862 52108
rect 5902 52096 5908 52108
rect 5960 52096 5966 52148
rect 7000 52071 7058 52077
rect 7000 52037 7012 52071
rect 7046 52068 7058 52071
rect 7558 52068 7564 52080
rect 7046 52040 7564 52068
rect 7046 52037 7058 52040
rect 7000 52031 7058 52037
rect 7558 52028 7564 52040
rect 7616 52028 7622 52080
rect 4341 52003 4399 52009
rect 4341 51969 4353 52003
rect 4387 52000 4399 52003
rect 6454 52000 6460 52012
rect 4387 51972 6460 52000
rect 4387 51969 4399 51972
rect 4341 51963 4399 51969
rect 6454 51960 6460 51972
rect 6512 51960 6518 52012
rect 6822 52000 6828 52012
rect 6656 51972 6828 52000
rect 6546 51892 6552 51944
rect 6604 51932 6610 51944
rect 6656 51932 6684 51972
rect 6822 51960 6828 51972
rect 6880 51960 6886 52012
rect 7466 51960 7472 52012
rect 7524 52000 7530 52012
rect 7742 52000 7748 52012
rect 7524 51972 7748 52000
rect 7524 51960 7530 51972
rect 7742 51960 7748 51972
rect 7800 51960 7806 52012
rect 10134 51960 10140 52012
rect 10192 51960 10198 52012
rect 6604 51904 6684 51932
rect 6604 51892 6610 51904
rect 6730 51892 6736 51944
rect 6788 51892 6794 51944
rect 10152 51864 10180 51960
rect 7668 51836 10180 51864
rect 1578 51756 1584 51808
rect 1636 51796 1642 51808
rect 4525 51799 4583 51805
rect 4525 51796 4537 51799
rect 1636 51768 4537 51796
rect 1636 51756 1642 51768
rect 4525 51765 4537 51768
rect 4571 51765 4583 51799
rect 4525 51759 4583 51765
rect 6362 51756 6368 51808
rect 6420 51796 6426 51808
rect 7668 51796 7696 51836
rect 6420 51768 7696 51796
rect 6420 51756 6426 51768
rect 8110 51756 8116 51808
rect 8168 51756 8174 51808
rect 1104 51706 9936 51728
rect 1104 51654 3610 51706
rect 3662 51654 3674 51706
rect 3726 51654 3738 51706
rect 3790 51654 3802 51706
rect 3854 51654 3866 51706
rect 3918 51654 5210 51706
rect 5262 51654 5274 51706
rect 5326 51654 5338 51706
rect 5390 51654 5402 51706
rect 5454 51654 5466 51706
rect 5518 51654 6810 51706
rect 6862 51654 6874 51706
rect 6926 51654 6938 51706
rect 6990 51654 7002 51706
rect 7054 51654 7066 51706
rect 7118 51654 8410 51706
rect 8462 51654 8474 51706
rect 8526 51654 8538 51706
rect 8590 51654 8602 51706
rect 8654 51654 8666 51706
rect 8718 51654 9936 51706
rect 1104 51632 9936 51654
rect 7006 51552 7012 51604
rect 7064 51592 7070 51604
rect 7064 51564 8156 51592
rect 7064 51552 7070 51564
rect 8128 51533 8156 51564
rect 8662 51552 8668 51604
rect 8720 51592 8726 51604
rect 9582 51592 9588 51604
rect 8720 51564 9588 51592
rect 8720 51552 8726 51564
rect 9582 51552 9588 51564
rect 9640 51552 9646 51604
rect 8113 51527 8171 51533
rect 8113 51493 8125 51527
rect 8159 51493 8171 51527
rect 8113 51487 8171 51493
rect 4890 51416 4896 51468
rect 4948 51416 4954 51468
rect 1486 51348 1492 51400
rect 1544 51348 1550 51400
rect 4908 51388 4936 51416
rect 5074 51388 5080 51400
rect 4908 51360 5080 51388
rect 5074 51348 5080 51360
rect 5132 51348 5138 51400
rect 5902 51348 5908 51400
rect 5960 51388 5966 51400
rect 6273 51391 6331 51397
rect 6273 51388 6285 51391
rect 5960 51360 6285 51388
rect 5960 51348 5966 51360
rect 6273 51357 6285 51360
rect 6319 51388 6331 51391
rect 6362 51388 6368 51400
rect 6319 51360 6368 51388
rect 6319 51357 6331 51360
rect 6273 51351 6331 51357
rect 6362 51348 6368 51360
rect 6420 51348 6426 51400
rect 6730 51348 6736 51400
rect 6788 51348 6794 51400
rect 8202 51388 8208 51400
rect 6840 51360 8208 51388
rect 6457 51323 6515 51329
rect 6457 51289 6469 51323
rect 6503 51320 6515 51323
rect 6840 51320 6868 51360
rect 8202 51348 8208 51360
rect 8260 51348 8266 51400
rect 8294 51348 8300 51400
rect 8352 51388 8358 51400
rect 8389 51391 8447 51397
rect 8389 51388 8401 51391
rect 8352 51360 8401 51388
rect 8352 51348 8358 51360
rect 8389 51357 8401 51360
rect 8435 51357 8447 51391
rect 8389 51351 8447 51357
rect 8481 51391 8539 51397
rect 8481 51357 8493 51391
rect 8527 51388 8539 51391
rect 8846 51388 8852 51400
rect 8527 51360 8852 51388
rect 8527 51357 8539 51360
rect 8481 51351 8539 51357
rect 8588 51332 8616 51360
rect 8846 51348 8852 51360
rect 8904 51348 8910 51400
rect 6503 51292 6868 51320
rect 7000 51323 7058 51329
rect 6503 51289 6515 51292
rect 6457 51283 6515 51289
rect 7000 51289 7012 51323
rect 7046 51320 7058 51323
rect 7282 51320 7288 51332
rect 7046 51292 7288 51320
rect 7046 51289 7058 51292
rect 7000 51283 7058 51289
rect 934 51212 940 51264
rect 992 51252 998 51264
rect 1581 51255 1639 51261
rect 1581 51252 1593 51255
rect 992 51224 1593 51252
rect 992 51212 998 51224
rect 1581 51221 1593 51224
rect 1627 51221 1639 51255
rect 1581 51215 1639 51221
rect 4246 51212 4252 51264
rect 4304 51252 4310 51264
rect 6472 51252 6500 51283
rect 7282 51280 7288 51292
rect 7340 51280 7346 51332
rect 7466 51280 7472 51332
rect 7524 51320 7530 51332
rect 7742 51320 7748 51332
rect 7524 51292 7748 51320
rect 7524 51280 7530 51292
rect 7742 51280 7748 51292
rect 7800 51280 7806 51332
rect 8036 51292 8340 51320
rect 4304 51224 6500 51252
rect 6641 51255 6699 51261
rect 4304 51212 4310 51224
rect 6641 51221 6653 51255
rect 6687 51252 6699 51255
rect 8036 51252 8064 51292
rect 8312 51264 8340 51292
rect 8570 51280 8576 51332
rect 8628 51280 8634 51332
rect 6687 51224 8064 51252
rect 6687 51221 6699 51224
rect 6641 51215 6699 51221
rect 8202 51212 8208 51264
rect 8260 51212 8266 51264
rect 8294 51212 8300 51264
rect 8352 51212 8358 51264
rect 8665 51255 8723 51261
rect 8665 51221 8677 51255
rect 8711 51252 8723 51255
rect 9214 51252 9220 51264
rect 8711 51224 9220 51252
rect 8711 51221 8723 51224
rect 8665 51215 8723 51221
rect 9214 51212 9220 51224
rect 9272 51212 9278 51264
rect 1104 51162 9936 51184
rect 1104 51110 2950 51162
rect 3002 51110 3014 51162
rect 3066 51110 3078 51162
rect 3130 51110 3142 51162
rect 3194 51110 3206 51162
rect 3258 51110 4550 51162
rect 4602 51110 4614 51162
rect 4666 51110 4678 51162
rect 4730 51110 4742 51162
rect 4794 51110 4806 51162
rect 4858 51110 6150 51162
rect 6202 51110 6214 51162
rect 6266 51110 6278 51162
rect 6330 51110 6342 51162
rect 6394 51110 6406 51162
rect 6458 51110 7750 51162
rect 7802 51110 7814 51162
rect 7866 51110 7878 51162
rect 7930 51110 7942 51162
rect 7994 51110 8006 51162
rect 8058 51110 9350 51162
rect 9402 51110 9414 51162
rect 9466 51110 9478 51162
rect 9530 51110 9542 51162
rect 9594 51110 9606 51162
rect 9658 51110 9936 51162
rect 1104 51088 9936 51110
rect 2222 51008 2228 51060
rect 2280 51048 2286 51060
rect 2498 51048 2504 51060
rect 2280 51020 2504 51048
rect 2280 51008 2286 51020
rect 2498 51008 2504 51020
rect 2556 51008 2562 51060
rect 2590 51008 2596 51060
rect 2648 51008 2654 51060
rect 7006 51048 7012 51060
rect 6104 51020 7012 51048
rect 2406 50980 2412 50992
rect 2332 50952 2412 50980
rect 2332 50708 2360 50952
rect 2406 50940 2412 50952
rect 2464 50940 2470 50992
rect 2406 50736 2412 50788
rect 2464 50776 2470 50788
rect 2608 50776 2636 51008
rect 5994 50940 6000 50992
rect 6052 50980 6058 50992
rect 6104 50980 6132 51020
rect 7006 51008 7012 51020
rect 7064 51008 7070 51060
rect 6052 50952 6132 50980
rect 6908 50983 6966 50989
rect 6052 50940 6058 50952
rect 6908 50949 6920 50983
rect 6954 50980 6966 50983
rect 7466 50980 7472 50992
rect 6954 50952 7472 50980
rect 6954 50949 6966 50952
rect 6908 50943 6966 50949
rect 7466 50940 7472 50952
rect 7524 50940 7530 50992
rect 5626 50872 5632 50924
rect 5684 50912 5690 50924
rect 6549 50915 6607 50921
rect 6549 50912 6561 50915
rect 5684 50884 6561 50912
rect 5684 50872 5690 50884
rect 6549 50881 6561 50884
rect 6595 50881 6607 50915
rect 6549 50875 6607 50881
rect 6641 50915 6699 50921
rect 6641 50881 6653 50915
rect 6687 50912 6699 50915
rect 6730 50912 6736 50924
rect 6687 50884 6736 50912
rect 6687 50881 6699 50884
rect 6641 50875 6699 50881
rect 6730 50872 6736 50884
rect 6788 50872 6794 50924
rect 8662 50804 8668 50856
rect 8720 50844 8726 50856
rect 9582 50844 9588 50856
rect 8720 50816 9588 50844
rect 8720 50804 8726 50816
rect 9582 50804 9588 50816
rect 9640 50804 9646 50856
rect 2464 50748 2636 50776
rect 2464 50736 2470 50748
rect 2498 50708 2504 50720
rect 2332 50680 2504 50708
rect 2498 50668 2504 50680
rect 2556 50668 2562 50720
rect 6365 50711 6423 50717
rect 6365 50677 6377 50711
rect 6411 50708 6423 50711
rect 7006 50708 7012 50720
rect 6411 50680 7012 50708
rect 6411 50677 6423 50680
rect 6365 50671 6423 50677
rect 7006 50668 7012 50680
rect 7064 50668 7070 50720
rect 7282 50668 7288 50720
rect 7340 50708 7346 50720
rect 8021 50711 8079 50717
rect 8021 50708 8033 50711
rect 7340 50680 8033 50708
rect 7340 50668 7346 50680
rect 8021 50677 8033 50680
rect 8067 50677 8079 50711
rect 8021 50671 8079 50677
rect 1104 50618 9936 50640
rect 1104 50566 3610 50618
rect 3662 50566 3674 50618
rect 3726 50566 3738 50618
rect 3790 50566 3802 50618
rect 3854 50566 3866 50618
rect 3918 50566 5210 50618
rect 5262 50566 5274 50618
rect 5326 50566 5338 50618
rect 5390 50566 5402 50618
rect 5454 50566 5466 50618
rect 5518 50566 6810 50618
rect 6862 50566 6874 50618
rect 6926 50566 6938 50618
rect 6990 50566 7002 50618
rect 7054 50566 7066 50618
rect 7118 50566 8410 50618
rect 8462 50566 8474 50618
rect 8526 50566 8538 50618
rect 8590 50566 8602 50618
rect 8654 50566 8666 50618
rect 8718 50566 9936 50618
rect 1104 50544 9936 50566
rect 1489 50303 1547 50309
rect 1489 50269 1501 50303
rect 1535 50300 1547 50303
rect 3326 50300 3332 50312
rect 1535 50272 3332 50300
rect 1535 50269 1547 50272
rect 1489 50263 1547 50269
rect 3326 50260 3332 50272
rect 3384 50260 3390 50312
rect 3786 50192 3792 50244
rect 3844 50232 3850 50244
rect 4338 50232 4344 50244
rect 3844 50204 4344 50232
rect 3844 50192 3850 50204
rect 4338 50192 4344 50204
rect 4396 50192 4402 50244
rect 934 50124 940 50176
rect 992 50164 998 50176
rect 1581 50167 1639 50173
rect 1581 50164 1593 50167
rect 992 50136 1593 50164
rect 992 50124 998 50136
rect 1581 50133 1593 50136
rect 1627 50133 1639 50167
rect 1581 50127 1639 50133
rect 5626 50124 5632 50176
rect 5684 50164 5690 50176
rect 6086 50164 6092 50176
rect 5684 50136 6092 50164
rect 5684 50124 5690 50136
rect 6086 50124 6092 50136
rect 6144 50124 6150 50176
rect 1104 50074 9936 50096
rect 1104 50022 2950 50074
rect 3002 50022 3014 50074
rect 3066 50022 3078 50074
rect 3130 50022 3142 50074
rect 3194 50022 3206 50074
rect 3258 50022 4550 50074
rect 4602 50022 4614 50074
rect 4666 50022 4678 50074
rect 4730 50022 4742 50074
rect 4794 50022 4806 50074
rect 4858 50022 6150 50074
rect 6202 50022 6214 50074
rect 6266 50022 6278 50074
rect 6330 50022 6342 50074
rect 6394 50022 6406 50074
rect 6458 50022 7750 50074
rect 7802 50022 7814 50074
rect 7866 50022 7878 50074
rect 7930 50022 7942 50074
rect 7994 50022 8006 50074
rect 8058 50022 9350 50074
rect 9402 50022 9414 50074
rect 9466 50022 9478 50074
rect 9530 50022 9542 50074
rect 9594 50022 9606 50074
rect 9658 50022 9936 50074
rect 1104 50000 9936 50022
rect 2746 49932 4384 49960
rect 2314 49852 2320 49904
rect 2372 49892 2378 49904
rect 2746 49892 2774 49932
rect 2372 49864 2774 49892
rect 2372 49852 2378 49864
rect 3786 49852 3792 49904
rect 3844 49892 3850 49904
rect 4249 49895 4307 49901
rect 4249 49892 4261 49895
rect 3844 49864 4261 49892
rect 3844 49852 3850 49864
rect 4249 49861 4261 49864
rect 4295 49861 4307 49895
rect 4249 49855 4307 49861
rect 1026 49784 1032 49836
rect 1084 49824 1090 49836
rect 3804 49824 3832 49852
rect 1084 49796 3832 49824
rect 4356 49824 4384 49932
rect 4430 49920 4436 49972
rect 4488 49960 4494 49972
rect 5074 49960 5080 49972
rect 4488 49932 5080 49960
rect 4488 49920 4494 49932
rect 5074 49920 5080 49932
rect 5132 49920 5138 49972
rect 7650 49960 7656 49972
rect 6196 49932 7656 49960
rect 4706 49852 4712 49904
rect 4764 49892 4770 49904
rect 4985 49895 5043 49901
rect 4985 49892 4997 49895
rect 4764 49864 4997 49892
rect 4764 49852 4770 49864
rect 4985 49861 4997 49864
rect 5031 49892 5043 49895
rect 5534 49892 5540 49904
rect 5031 49864 5540 49892
rect 5031 49861 5043 49864
rect 4985 49855 5043 49861
rect 5534 49852 5540 49864
rect 5592 49852 5598 49904
rect 4801 49827 4859 49833
rect 4801 49824 4813 49827
rect 4356 49796 4813 49824
rect 1084 49784 1090 49796
rect 3326 49716 3332 49768
rect 3384 49756 3390 49768
rect 4338 49756 4344 49768
rect 3384 49728 4344 49756
rect 3384 49716 3390 49728
rect 4338 49716 4344 49728
rect 4396 49756 4402 49768
rect 4396 49728 4568 49756
rect 4396 49716 4402 49728
rect 4540 49697 4568 49728
rect 4525 49691 4583 49697
rect 4525 49657 4537 49691
rect 4571 49657 4583 49691
rect 4525 49651 4583 49657
rect 4338 49580 4344 49632
rect 4396 49620 4402 49632
rect 4632 49620 4660 49796
rect 4801 49793 4813 49796
rect 4847 49793 4859 49827
rect 4801 49787 4859 49793
rect 4709 49759 4767 49765
rect 4709 49725 4721 49759
rect 4755 49756 4767 49759
rect 6196 49756 6224 49932
rect 7650 49920 7656 49932
rect 7708 49920 7714 49972
rect 8113 49963 8171 49969
rect 8113 49929 8125 49963
rect 8159 49929 8171 49963
rect 8113 49923 8171 49929
rect 6908 49895 6966 49901
rect 6908 49861 6920 49895
rect 6954 49892 6966 49895
rect 8128 49892 8156 49923
rect 6954 49864 8156 49892
rect 6954 49861 6966 49864
rect 6908 49855 6966 49861
rect 6641 49827 6699 49833
rect 6641 49793 6653 49827
rect 6687 49824 6699 49827
rect 6730 49824 6736 49836
rect 6687 49796 6736 49824
rect 6687 49793 6699 49796
rect 6641 49787 6699 49793
rect 6730 49784 6736 49796
rect 6788 49784 6794 49836
rect 8294 49784 8300 49836
rect 8352 49784 8358 49836
rect 4755 49728 6224 49756
rect 4755 49725 4767 49728
rect 4709 49719 4767 49725
rect 4396 49592 4660 49620
rect 4396 49580 4402 49592
rect 4890 49580 4896 49632
rect 4948 49620 4954 49632
rect 5169 49623 5227 49629
rect 5169 49620 5181 49623
rect 4948 49592 5181 49620
rect 4948 49580 4954 49592
rect 5169 49589 5181 49592
rect 5215 49589 5227 49623
rect 5169 49583 5227 49589
rect 8021 49623 8079 49629
rect 8021 49589 8033 49623
rect 8067 49620 8079 49623
rect 8294 49620 8300 49632
rect 8067 49592 8300 49620
rect 8067 49589 8079 49592
rect 8021 49583 8079 49589
rect 8294 49580 8300 49592
rect 8352 49580 8358 49632
rect 1104 49530 9936 49552
rect 1104 49478 3610 49530
rect 3662 49478 3674 49530
rect 3726 49478 3738 49530
rect 3790 49478 3802 49530
rect 3854 49478 3866 49530
rect 3918 49478 5210 49530
rect 5262 49478 5274 49530
rect 5326 49478 5338 49530
rect 5390 49478 5402 49530
rect 5454 49478 5466 49530
rect 5518 49478 6810 49530
rect 6862 49478 6874 49530
rect 6926 49478 6938 49530
rect 6990 49478 7002 49530
rect 7054 49478 7066 49530
rect 7118 49478 8410 49530
rect 8462 49478 8474 49530
rect 8526 49478 8538 49530
rect 8590 49478 8602 49530
rect 8654 49478 8666 49530
rect 8718 49478 9936 49530
rect 1104 49456 9936 49478
rect 2222 49416 2228 49428
rect 1504 49388 2228 49416
rect 1504 49221 1532 49388
rect 2222 49376 2228 49388
rect 2280 49376 2286 49428
rect 4706 49376 4712 49428
rect 4764 49416 4770 49428
rect 5166 49416 5172 49428
rect 4764 49388 5172 49416
rect 4764 49376 4770 49388
rect 5166 49376 5172 49388
rect 5224 49376 5230 49428
rect 6457 49419 6515 49425
rect 6457 49385 6469 49419
rect 6503 49416 6515 49419
rect 6638 49416 6644 49428
rect 6503 49388 6644 49416
rect 6503 49385 6515 49388
rect 6457 49379 6515 49385
rect 6638 49376 6644 49388
rect 6696 49376 6702 49428
rect 8110 49376 8116 49428
rect 8168 49416 8174 49428
rect 8297 49419 8355 49425
rect 8297 49416 8309 49419
rect 8168 49388 8309 49416
rect 8168 49376 8174 49388
rect 8297 49385 8309 49388
rect 8343 49385 8355 49419
rect 8297 49379 8355 49385
rect 9214 49376 9220 49428
rect 9272 49376 9278 49428
rect 9232 49348 9260 49376
rect 8220 49320 9260 49348
rect 6196 49252 6868 49280
rect 6196 49221 6224 49252
rect 1489 49215 1547 49221
rect 1489 49181 1501 49215
rect 1535 49181 1547 49215
rect 1489 49175 1547 49181
rect 6181 49215 6239 49221
rect 6181 49181 6193 49215
rect 6227 49181 6239 49215
rect 6181 49175 6239 49181
rect 6730 49172 6736 49224
rect 6788 49172 6794 49224
rect 6840 49212 6868 49252
rect 7466 49212 7472 49224
rect 6840 49184 7472 49212
rect 7466 49172 7472 49184
rect 7524 49212 7530 49224
rect 8220 49221 8248 49320
rect 8570 49240 8576 49292
rect 8628 49280 8634 49292
rect 9122 49280 9128 49292
rect 8628 49252 9128 49280
rect 8628 49240 8634 49252
rect 9122 49240 9128 49252
rect 9180 49240 9186 49292
rect 8205 49215 8263 49221
rect 8205 49212 8217 49215
rect 7524 49184 8217 49212
rect 7524 49172 7530 49184
rect 8205 49181 8217 49184
rect 8251 49181 8263 49215
rect 8205 49175 8263 49181
rect 11330 49172 11336 49224
rect 11388 49172 11394 49224
rect 7000 49147 7058 49153
rect 7000 49113 7012 49147
rect 7046 49144 7058 49147
rect 7650 49144 7656 49156
rect 7046 49116 7656 49144
rect 7046 49113 7058 49116
rect 7000 49107 7058 49113
rect 7650 49104 7656 49116
rect 7708 49144 7714 49156
rect 11348 49144 11376 49172
rect 7708 49116 11376 49144
rect 7708 49104 7714 49116
rect 934 49036 940 49088
rect 992 49076 998 49088
rect 1581 49079 1639 49085
rect 1581 49076 1593 49079
rect 992 49048 1593 49076
rect 992 49036 998 49048
rect 1581 49045 1593 49048
rect 1627 49045 1639 49079
rect 1581 49039 1639 49045
rect 6638 49036 6644 49088
rect 6696 49036 6702 49088
rect 8110 49036 8116 49088
rect 8168 49036 8174 49088
rect 8665 49079 8723 49085
rect 8665 49045 8677 49079
rect 8711 49076 8723 49079
rect 8754 49076 8760 49088
rect 8711 49048 8760 49076
rect 8711 49045 8723 49048
rect 8665 49039 8723 49045
rect 8754 49036 8760 49048
rect 8812 49036 8818 49088
rect 1104 48986 9936 49008
rect 1104 48934 2950 48986
rect 3002 48934 3014 48986
rect 3066 48934 3078 48986
rect 3130 48934 3142 48986
rect 3194 48934 3206 48986
rect 3258 48934 4550 48986
rect 4602 48934 4614 48986
rect 4666 48934 4678 48986
rect 4730 48934 4742 48986
rect 4794 48934 4806 48986
rect 4858 48934 6150 48986
rect 6202 48934 6214 48986
rect 6266 48934 6278 48986
rect 6330 48934 6342 48986
rect 6394 48934 6406 48986
rect 6458 48934 7750 48986
rect 7802 48934 7814 48986
rect 7866 48934 7878 48986
rect 7930 48934 7942 48986
rect 7994 48934 8006 48986
rect 8058 48934 9350 48986
rect 9402 48934 9414 48986
rect 9466 48934 9478 48986
rect 9530 48934 9542 48986
rect 9594 48934 9606 48986
rect 9658 48934 9936 48986
rect 1104 48912 9936 48934
rect 4154 48832 4160 48884
rect 4212 48872 4218 48884
rect 4798 48872 4804 48884
rect 4212 48844 4804 48872
rect 4212 48832 4218 48844
rect 4798 48832 4804 48844
rect 4856 48832 4862 48884
rect 4890 48832 4896 48884
rect 4948 48832 4954 48884
rect 1489 48807 1547 48813
rect 1489 48773 1501 48807
rect 1535 48804 1547 48807
rect 2866 48804 2872 48816
rect 1535 48776 2872 48804
rect 1535 48773 1547 48776
rect 1489 48767 1547 48773
rect 2866 48764 2872 48776
rect 2924 48764 2930 48816
rect 4709 48739 4767 48745
rect 4709 48705 4721 48739
rect 4755 48736 4767 48739
rect 4908 48736 4936 48832
rect 6908 48807 6966 48813
rect 5368 48776 6868 48804
rect 5368 48745 5396 48776
rect 4755 48708 4936 48736
rect 5353 48739 5411 48745
rect 4755 48705 4767 48708
rect 4709 48699 4767 48705
rect 5353 48705 5365 48739
rect 5399 48705 5411 48739
rect 5353 48699 5411 48705
rect 5629 48739 5687 48745
rect 5629 48705 5641 48739
rect 5675 48736 5687 48739
rect 6086 48736 6092 48748
rect 5675 48708 6092 48736
rect 5675 48705 5687 48708
rect 5629 48699 5687 48705
rect 6086 48696 6092 48708
rect 6144 48696 6150 48748
rect 6641 48739 6699 48745
rect 6641 48705 6653 48739
rect 6687 48736 6699 48739
rect 6730 48736 6736 48748
rect 6687 48708 6736 48736
rect 6687 48705 6699 48708
rect 6641 48699 6699 48705
rect 6730 48696 6736 48708
rect 6788 48696 6794 48748
rect 6840 48736 6868 48776
rect 6908 48773 6920 48807
rect 6954 48804 6966 48807
rect 8202 48804 8208 48816
rect 6954 48776 8208 48804
rect 6954 48773 6966 48776
rect 6908 48767 6966 48773
rect 8202 48764 8208 48776
rect 8260 48764 8266 48816
rect 8662 48736 8668 48748
rect 6840 48708 8668 48736
rect 8662 48696 8668 48708
rect 8720 48736 8726 48748
rect 9122 48736 9128 48748
rect 8720 48708 9128 48736
rect 8720 48696 8726 48708
rect 9122 48696 9128 48708
rect 9180 48696 9186 48748
rect 4706 48560 4712 48612
rect 4764 48600 4770 48612
rect 5166 48600 5172 48612
rect 4764 48572 5172 48600
rect 4764 48560 4770 48572
rect 5166 48560 5172 48572
rect 5224 48560 5230 48612
rect 1578 48492 1584 48544
rect 1636 48492 1642 48544
rect 4246 48492 4252 48544
rect 4304 48532 4310 48544
rect 4525 48535 4583 48541
rect 4525 48532 4537 48535
rect 4304 48504 4537 48532
rect 4304 48492 4310 48504
rect 4525 48501 4537 48504
rect 4571 48501 4583 48535
rect 4525 48495 4583 48501
rect 8021 48535 8079 48541
rect 8021 48501 8033 48535
rect 8067 48532 8079 48535
rect 8202 48532 8208 48544
rect 8067 48504 8208 48532
rect 8067 48501 8079 48504
rect 8021 48495 8079 48501
rect 8202 48492 8208 48504
rect 8260 48492 8266 48544
rect 8570 48492 8576 48544
rect 8628 48532 8634 48544
rect 8938 48532 8944 48544
rect 8628 48504 8944 48532
rect 8628 48492 8634 48504
rect 8938 48492 8944 48504
rect 8996 48492 9002 48544
rect 1104 48442 9936 48464
rect 1104 48390 3610 48442
rect 3662 48390 3674 48442
rect 3726 48390 3738 48442
rect 3790 48390 3802 48442
rect 3854 48390 3866 48442
rect 3918 48390 5210 48442
rect 5262 48390 5274 48442
rect 5326 48390 5338 48442
rect 5390 48390 5402 48442
rect 5454 48390 5466 48442
rect 5518 48390 6810 48442
rect 6862 48390 6874 48442
rect 6926 48390 6938 48442
rect 6990 48390 7002 48442
rect 7054 48390 7066 48442
rect 7118 48390 8410 48442
rect 8462 48390 8474 48442
rect 8526 48390 8538 48442
rect 8590 48390 8602 48442
rect 8654 48390 8666 48442
rect 8718 48390 9936 48442
rect 1104 48368 9936 48390
rect 4706 48288 4712 48340
rect 4764 48328 4770 48340
rect 5166 48328 5172 48340
rect 4764 48300 5172 48328
rect 4764 48288 4770 48300
rect 5166 48288 5172 48300
rect 5224 48288 5230 48340
rect 6641 48127 6699 48133
rect 6641 48093 6653 48127
rect 6687 48124 6699 48127
rect 6730 48124 6736 48136
rect 6687 48096 6736 48124
rect 6687 48093 6699 48096
rect 6641 48087 6699 48093
rect 6730 48084 6736 48096
rect 6788 48084 6794 48136
rect 6908 48127 6966 48133
rect 6908 48093 6920 48127
rect 6954 48124 6966 48127
rect 7190 48124 7196 48136
rect 6954 48096 7196 48124
rect 6954 48093 6966 48096
rect 6908 48087 6966 48093
rect 7190 48084 7196 48096
rect 7248 48084 7254 48136
rect 7466 48084 7472 48136
rect 7524 48084 7530 48136
rect 7484 48056 7512 48084
rect 7208 48028 7512 48056
rect 7208 48000 7236 48028
rect 6086 47948 6092 48000
rect 6144 47988 6150 48000
rect 6822 47988 6828 48000
rect 6144 47960 6828 47988
rect 6144 47948 6150 47960
rect 6822 47948 6828 47960
rect 6880 47948 6886 48000
rect 7190 47948 7196 48000
rect 7248 47948 7254 48000
rect 7466 47948 7472 48000
rect 7524 47988 7530 48000
rect 8021 47991 8079 47997
rect 8021 47988 8033 47991
rect 7524 47960 8033 47988
rect 7524 47948 7530 47960
rect 8021 47957 8033 47960
rect 8067 47957 8079 47991
rect 8021 47951 8079 47957
rect 1104 47898 9936 47920
rect 1104 47846 2950 47898
rect 3002 47846 3014 47898
rect 3066 47846 3078 47898
rect 3130 47846 3142 47898
rect 3194 47846 3206 47898
rect 3258 47846 4550 47898
rect 4602 47846 4614 47898
rect 4666 47846 4678 47898
rect 4730 47846 4742 47898
rect 4794 47846 4806 47898
rect 4858 47846 6150 47898
rect 6202 47846 6214 47898
rect 6266 47846 6278 47898
rect 6330 47846 6342 47898
rect 6394 47846 6406 47898
rect 6458 47846 7750 47898
rect 7802 47846 7814 47898
rect 7866 47846 7878 47898
rect 7930 47846 7942 47898
rect 7994 47846 8006 47898
rect 8058 47846 9350 47898
rect 9402 47846 9414 47898
rect 9466 47846 9478 47898
rect 9530 47846 9542 47898
rect 9594 47846 9606 47898
rect 9658 47846 9936 47898
rect 1104 47824 9936 47846
rect 1489 47719 1547 47725
rect 1489 47685 1501 47719
rect 1535 47716 1547 47719
rect 2682 47716 2688 47728
rect 1535 47688 2688 47716
rect 1535 47685 1547 47688
rect 1489 47679 1547 47685
rect 2682 47676 2688 47688
rect 2740 47676 2746 47728
rect 6454 47608 6460 47660
rect 6512 47648 6518 47660
rect 6822 47648 6828 47660
rect 6512 47620 6828 47648
rect 6512 47608 6518 47620
rect 6822 47608 6828 47620
rect 6880 47648 6886 47660
rect 6917 47651 6975 47657
rect 6917 47648 6929 47651
rect 6880 47620 6929 47648
rect 6880 47608 6886 47620
rect 6917 47617 6929 47620
rect 6963 47617 6975 47651
rect 6917 47611 6975 47617
rect 4890 47472 4896 47524
rect 4948 47512 4954 47524
rect 7377 47515 7435 47521
rect 7377 47512 7389 47515
rect 4948 47484 7389 47512
rect 4948 47472 4954 47484
rect 7377 47481 7389 47484
rect 7423 47481 7435 47515
rect 7377 47475 7435 47481
rect 9030 47472 9036 47524
rect 9088 47512 9094 47524
rect 9306 47512 9312 47524
rect 9088 47484 9312 47512
rect 9088 47472 9094 47484
rect 9306 47472 9312 47484
rect 9364 47472 9370 47524
rect 934 47404 940 47456
rect 992 47444 998 47456
rect 1581 47447 1639 47453
rect 1581 47444 1593 47447
rect 992 47416 1593 47444
rect 992 47404 998 47416
rect 1581 47413 1593 47416
rect 1627 47413 1639 47447
rect 1581 47407 1639 47413
rect 2866 47404 2872 47456
rect 2924 47444 2930 47456
rect 5166 47444 5172 47456
rect 2924 47416 5172 47444
rect 2924 47404 2930 47416
rect 5166 47404 5172 47416
rect 5224 47404 5230 47456
rect 7193 47447 7251 47453
rect 7193 47413 7205 47447
rect 7239 47444 7251 47447
rect 7282 47444 7288 47456
rect 7239 47416 7288 47444
rect 7239 47413 7251 47416
rect 7193 47407 7251 47413
rect 7282 47404 7288 47416
rect 7340 47404 7346 47456
rect 1104 47354 9936 47376
rect 1104 47302 3610 47354
rect 3662 47302 3674 47354
rect 3726 47302 3738 47354
rect 3790 47302 3802 47354
rect 3854 47302 3866 47354
rect 3918 47302 5210 47354
rect 5262 47302 5274 47354
rect 5326 47302 5338 47354
rect 5390 47302 5402 47354
rect 5454 47302 5466 47354
rect 5518 47302 6810 47354
rect 6862 47302 6874 47354
rect 6926 47302 6938 47354
rect 6990 47302 7002 47354
rect 7054 47302 7066 47354
rect 7118 47302 8410 47354
rect 8462 47302 8474 47354
rect 8526 47302 8538 47354
rect 8590 47302 8602 47354
rect 8654 47302 8666 47354
rect 8718 47302 9936 47354
rect 1104 47280 9936 47302
rect 1578 47064 1584 47116
rect 1636 47104 1642 47116
rect 3326 47104 3332 47116
rect 1636 47076 3332 47104
rect 1636 47064 1642 47076
rect 3326 47064 3332 47076
rect 3384 47064 3390 47116
rect 8846 47064 8852 47116
rect 8904 47104 8910 47116
rect 9030 47104 9036 47116
rect 8904 47076 9036 47104
rect 8904 47064 8910 47076
rect 9030 47064 9036 47076
rect 9088 47064 9094 47116
rect 9214 47064 9220 47116
rect 9272 47064 9278 47116
rect 3789 47039 3847 47045
rect 3789 47005 3801 47039
rect 3835 47036 3847 47039
rect 6733 47039 6791 47045
rect 6733 47036 6745 47039
rect 3835 47008 6745 47036
rect 3835 47005 3847 47008
rect 3789 46999 3847 47005
rect 6733 47005 6745 47008
rect 6779 47036 6791 47039
rect 6822 47036 6828 47048
rect 6779 47008 6828 47036
rect 6779 47005 6791 47008
rect 6733 46999 6791 47005
rect 6822 46996 6828 47008
rect 6880 46996 6886 47048
rect 9232 47036 9260 47064
rect 7116 47008 9260 47036
rect 7116 46980 7144 47008
rect 2774 46928 2780 46980
rect 2832 46968 2838 46980
rect 3326 46968 3332 46980
rect 2832 46940 3332 46968
rect 2832 46928 2838 46940
rect 3326 46928 3332 46940
rect 3384 46928 3390 46980
rect 4056 46971 4114 46977
rect 4056 46937 4068 46971
rect 4102 46968 4114 46971
rect 4246 46968 4252 46980
rect 4102 46940 4252 46968
rect 4102 46937 4114 46940
rect 4056 46931 4114 46937
rect 4246 46928 4252 46940
rect 4304 46928 4310 46980
rect 5534 46928 5540 46980
rect 5592 46968 5598 46980
rect 6454 46968 6460 46980
rect 5592 46940 6460 46968
rect 5592 46928 5598 46940
rect 6454 46928 6460 46940
rect 6512 46928 6518 46980
rect 7000 46971 7058 46977
rect 7000 46937 7012 46971
rect 7046 46968 7058 46971
rect 7098 46968 7104 46980
rect 7046 46940 7104 46968
rect 7046 46937 7058 46940
rect 7000 46931 7058 46937
rect 7098 46928 7104 46940
rect 7156 46928 7162 46980
rect 5166 46860 5172 46912
rect 5224 46860 5230 46912
rect 5718 46860 5724 46912
rect 5776 46900 5782 46912
rect 6730 46900 6736 46912
rect 5776 46872 6736 46900
rect 5776 46860 5782 46872
rect 6730 46860 6736 46872
rect 6788 46860 6794 46912
rect 8113 46903 8171 46909
rect 8113 46869 8125 46903
rect 8159 46900 8171 46903
rect 8846 46900 8852 46912
rect 8159 46872 8852 46900
rect 8159 46869 8171 46872
rect 8113 46863 8171 46869
rect 8846 46860 8852 46872
rect 8904 46860 8910 46912
rect 1104 46810 9936 46832
rect 1104 46758 2950 46810
rect 3002 46758 3014 46810
rect 3066 46758 3078 46810
rect 3130 46758 3142 46810
rect 3194 46758 3206 46810
rect 3258 46758 4550 46810
rect 4602 46758 4614 46810
rect 4666 46758 4678 46810
rect 4730 46758 4742 46810
rect 4794 46758 4806 46810
rect 4858 46758 6150 46810
rect 6202 46758 6214 46810
rect 6266 46758 6278 46810
rect 6330 46758 6342 46810
rect 6394 46758 6406 46810
rect 6458 46758 7750 46810
rect 7802 46758 7814 46810
rect 7866 46758 7878 46810
rect 7930 46758 7942 46810
rect 7994 46758 8006 46810
rect 8058 46758 9350 46810
rect 9402 46758 9414 46810
rect 9466 46758 9478 46810
rect 9530 46758 9542 46810
rect 9594 46758 9606 46810
rect 9658 46758 9936 46810
rect 1104 46736 9936 46758
rect 5718 46656 5724 46708
rect 5776 46696 5782 46708
rect 5902 46696 5908 46708
rect 5776 46668 5908 46696
rect 5776 46656 5782 46668
rect 5902 46656 5908 46668
rect 5960 46656 5966 46708
rect 6822 46656 6828 46708
rect 6880 46696 6886 46708
rect 9125 46699 9183 46705
rect 9125 46696 9137 46699
rect 6880 46668 9137 46696
rect 6880 46656 6886 46668
rect 9125 46665 9137 46668
rect 9171 46665 9183 46699
rect 9125 46659 9183 46665
rect 1489 46631 1547 46637
rect 1489 46597 1501 46631
rect 1535 46628 1547 46631
rect 2406 46628 2412 46640
rect 1535 46600 2412 46628
rect 1535 46597 1547 46600
rect 1489 46591 1547 46597
rect 2406 46588 2412 46600
rect 2464 46588 2470 46640
rect 6454 46588 6460 46640
rect 6512 46628 6518 46640
rect 6730 46628 6736 46640
rect 6512 46600 6736 46628
rect 6512 46588 6518 46600
rect 6730 46588 6736 46600
rect 6788 46588 6794 46640
rect 7190 46588 7196 46640
rect 7248 46628 7254 46640
rect 7837 46631 7895 46637
rect 7837 46628 7849 46631
rect 7248 46600 7849 46628
rect 7248 46588 7254 46600
rect 7837 46597 7849 46600
rect 7883 46628 7895 46631
rect 11146 46628 11152 46640
rect 7883 46600 11152 46628
rect 7883 46597 7895 46600
rect 7837 46591 7895 46597
rect 11146 46588 11152 46600
rect 11204 46588 11210 46640
rect 5534 46520 5540 46572
rect 5592 46560 5598 46572
rect 5721 46563 5779 46569
rect 5721 46560 5733 46563
rect 5592 46532 5733 46560
rect 5592 46520 5598 46532
rect 5721 46529 5733 46532
rect 5767 46560 5779 46563
rect 6632 46563 6690 46569
rect 5767 46532 6132 46560
rect 5767 46529 5779 46532
rect 5721 46523 5779 46529
rect 5994 46452 6000 46504
rect 6052 46452 6058 46504
rect 6012 46424 6040 46452
rect 6104 46436 6132 46532
rect 6632 46529 6644 46563
rect 6678 46560 6690 46563
rect 6678 46532 9674 46560
rect 6678 46529 6690 46532
rect 6632 46523 6690 46529
rect 6362 46452 6368 46504
rect 6420 46452 6426 46504
rect 9646 46492 9674 46532
rect 9950 46520 9956 46572
rect 10008 46520 10014 46572
rect 9968 46492 9996 46520
rect 9646 46464 9996 46492
rect 5828 46396 6040 46424
rect 934 46316 940 46368
rect 992 46356 998 46368
rect 1581 46359 1639 46365
rect 1581 46356 1593 46359
rect 992 46328 1593 46356
rect 992 46316 998 46328
rect 1581 46325 1593 46328
rect 1627 46325 1639 46359
rect 1581 46319 1639 46325
rect 4338 46316 4344 46368
rect 4396 46356 4402 46368
rect 5166 46356 5172 46368
rect 4396 46328 5172 46356
rect 4396 46316 4402 46328
rect 5166 46316 5172 46328
rect 5224 46316 5230 46368
rect 5828 46365 5856 46396
rect 6086 46384 6092 46436
rect 6144 46384 6150 46436
rect 5813 46359 5871 46365
rect 5813 46325 5825 46359
rect 5859 46325 5871 46359
rect 5813 46319 5871 46325
rect 5902 46316 5908 46368
rect 5960 46356 5966 46368
rect 6181 46359 6239 46365
rect 6181 46356 6193 46359
rect 5960 46328 6193 46356
rect 5960 46316 5966 46328
rect 6181 46325 6193 46328
rect 6227 46325 6239 46359
rect 6181 46319 6239 46325
rect 6270 46316 6276 46368
rect 6328 46356 6334 46368
rect 7745 46359 7803 46365
rect 7745 46356 7757 46359
rect 6328 46328 7757 46356
rect 6328 46316 6334 46328
rect 7745 46325 7757 46328
rect 7791 46325 7803 46359
rect 7745 46319 7803 46325
rect 1104 46266 9936 46288
rect 1104 46214 3610 46266
rect 3662 46214 3674 46266
rect 3726 46214 3738 46266
rect 3790 46214 3802 46266
rect 3854 46214 3866 46266
rect 3918 46214 5210 46266
rect 5262 46214 5274 46266
rect 5326 46214 5338 46266
rect 5390 46214 5402 46266
rect 5454 46214 5466 46266
rect 5518 46214 6810 46266
rect 6862 46214 6874 46266
rect 6926 46214 6938 46266
rect 6990 46214 7002 46266
rect 7054 46214 7066 46266
rect 7118 46214 8410 46266
rect 8462 46214 8474 46266
rect 8526 46214 8538 46266
rect 8590 46214 8602 46266
rect 8654 46214 8666 46266
rect 8718 46214 9936 46266
rect 1104 46192 9936 46214
rect 2498 46112 2504 46164
rect 2556 46152 2562 46164
rect 2866 46152 2872 46164
rect 2556 46124 2872 46152
rect 2556 46112 2562 46124
rect 2866 46112 2872 46124
rect 2924 46112 2930 46164
rect 7006 46112 7012 46164
rect 7064 46152 7070 46164
rect 7282 46152 7288 46164
rect 7064 46124 7288 46152
rect 7064 46112 7070 46124
rect 7282 46112 7288 46124
rect 7340 46152 7346 46164
rect 7340 46124 8064 46152
rect 7340 46112 7346 46124
rect 6362 45976 6368 46028
rect 6420 46016 6426 46028
rect 6638 46016 6644 46028
rect 6420 45988 6644 46016
rect 6420 45976 6426 45988
rect 6638 45976 6644 45988
rect 6696 45976 6702 46028
rect 4522 45908 4528 45960
rect 4580 45948 4586 45960
rect 5166 45948 5172 45960
rect 4580 45920 5172 45948
rect 4580 45908 4586 45920
rect 5166 45908 5172 45920
rect 5224 45908 5230 45960
rect 6454 45908 6460 45960
rect 6512 45908 6518 45960
rect 8036 45948 8064 46124
rect 8202 46112 8208 46164
rect 8260 46112 8266 46164
rect 8294 46112 8300 46164
rect 8352 46112 8358 46164
rect 8662 46112 8668 46164
rect 8720 46152 8726 46164
rect 8938 46152 8944 46164
rect 8720 46124 8944 46152
rect 8720 46112 8726 46124
rect 8938 46112 8944 46124
rect 8996 46112 9002 46164
rect 9033 46155 9091 46161
rect 9033 46121 9045 46155
rect 9079 46121 9091 46155
rect 9033 46115 9091 46121
rect 8220 46084 8248 46112
rect 9048 46084 9076 46115
rect 8220 46056 9076 46084
rect 8205 45951 8263 45957
rect 8205 45948 8217 45951
rect 8036 45920 8217 45948
rect 8205 45917 8217 45920
rect 8251 45948 8263 45951
rect 8941 45951 8999 45957
rect 8941 45948 8953 45951
rect 8251 45920 8953 45948
rect 8251 45917 8263 45920
rect 8205 45911 8263 45917
rect 8941 45917 8953 45920
rect 8987 45917 8999 45951
rect 8941 45911 8999 45917
rect 5534 45840 5540 45892
rect 5592 45880 5598 45892
rect 6472 45880 6500 45908
rect 6897 45883 6955 45889
rect 6897 45880 6909 45883
rect 5592 45852 6909 45880
rect 5592 45840 5598 45852
rect 6897 45849 6909 45852
rect 6943 45849 6955 45883
rect 6897 45843 6955 45849
rect 8386 45840 8392 45892
rect 8444 45880 8450 45892
rect 9306 45880 9312 45892
rect 8444 45852 9312 45880
rect 8444 45840 8450 45852
rect 9306 45840 9312 45852
rect 9364 45840 9370 45892
rect 2498 45772 2504 45824
rect 2556 45812 2562 45824
rect 4154 45812 4160 45824
rect 2556 45784 4160 45812
rect 2556 45772 2562 45784
rect 4154 45772 4160 45784
rect 4212 45772 4218 45824
rect 7374 45772 7380 45824
rect 7432 45812 7438 45824
rect 8021 45815 8079 45821
rect 8021 45812 8033 45815
rect 7432 45784 8033 45812
rect 7432 45772 7438 45784
rect 8021 45781 8033 45784
rect 8067 45781 8079 45815
rect 8021 45775 8079 45781
rect 8294 45772 8300 45824
rect 8352 45812 8358 45824
rect 8665 45815 8723 45821
rect 8665 45812 8677 45815
rect 8352 45784 8677 45812
rect 8352 45772 8358 45784
rect 8665 45781 8677 45784
rect 8711 45781 8723 45815
rect 8665 45775 8723 45781
rect 8938 45772 8944 45824
rect 8996 45812 9002 45824
rect 9401 45815 9459 45821
rect 9401 45812 9413 45815
rect 8996 45784 9413 45812
rect 8996 45772 9002 45784
rect 9401 45781 9413 45784
rect 9447 45781 9459 45815
rect 9401 45775 9459 45781
rect 1104 45722 9936 45744
rect 1104 45670 2950 45722
rect 3002 45670 3014 45722
rect 3066 45670 3078 45722
rect 3130 45670 3142 45722
rect 3194 45670 3206 45722
rect 3258 45670 4550 45722
rect 4602 45670 4614 45722
rect 4666 45670 4678 45722
rect 4730 45670 4742 45722
rect 4794 45670 4806 45722
rect 4858 45670 6150 45722
rect 6202 45670 6214 45722
rect 6266 45670 6278 45722
rect 6330 45670 6342 45722
rect 6394 45670 6406 45722
rect 6458 45670 7750 45722
rect 7802 45670 7814 45722
rect 7866 45670 7878 45722
rect 7930 45670 7942 45722
rect 7994 45670 8006 45722
rect 8058 45670 9350 45722
rect 9402 45670 9414 45722
rect 9466 45670 9478 45722
rect 9530 45670 9542 45722
rect 9594 45670 9606 45722
rect 9658 45670 9936 45722
rect 1104 45648 9936 45670
rect 7834 45568 7840 45620
rect 7892 45608 7898 45620
rect 8386 45608 8392 45620
rect 7892 45580 8392 45608
rect 7892 45568 7898 45580
rect 8386 45568 8392 45580
rect 8444 45568 8450 45620
rect 1486 45500 1492 45552
rect 1544 45500 1550 45552
rect 4908 45512 8800 45540
rect 4246 45432 4252 45484
rect 4304 45432 4310 45484
rect 4614 45432 4620 45484
rect 4672 45432 4678 45484
rect 4908 45481 4936 45512
rect 8772 45484 8800 45512
rect 9122 45500 9128 45552
rect 9180 45500 9186 45552
rect 4893 45475 4951 45481
rect 4893 45441 4905 45475
rect 4939 45441 4951 45475
rect 4893 45435 4951 45441
rect 4982 45432 4988 45484
rect 5040 45432 5046 45484
rect 5442 45432 5448 45484
rect 5500 45432 5506 45484
rect 7006 45432 7012 45484
rect 7064 45472 7070 45484
rect 7193 45475 7251 45481
rect 7193 45472 7205 45475
rect 7064 45444 7205 45472
rect 7064 45432 7070 45444
rect 7193 45441 7205 45444
rect 7239 45441 7251 45475
rect 7193 45435 7251 45441
rect 8205 45475 8263 45481
rect 8205 45441 8217 45475
rect 8251 45441 8263 45475
rect 8205 45435 8263 45441
rect 4264 45336 4292 45432
rect 4801 45407 4859 45413
rect 4801 45373 4813 45407
rect 4847 45404 4859 45407
rect 5000 45404 5028 45432
rect 4847 45376 5028 45404
rect 4847 45373 4859 45376
rect 4801 45367 4859 45373
rect 4172 45308 4292 45336
rect 4709 45339 4767 45345
rect 4172 45280 4200 45308
rect 4709 45305 4721 45339
rect 4755 45305 4767 45339
rect 4709 45299 4767 45305
rect 934 45228 940 45280
rect 992 45268 998 45280
rect 1581 45271 1639 45277
rect 1581 45268 1593 45271
rect 992 45240 1593 45268
rect 992 45228 998 45240
rect 1581 45237 1593 45240
rect 1627 45237 1639 45271
rect 1581 45231 1639 45237
rect 4154 45228 4160 45280
rect 4212 45228 4218 45280
rect 4246 45228 4252 45280
rect 4304 45268 4310 45280
rect 4433 45271 4491 45277
rect 4433 45268 4445 45271
rect 4304 45240 4445 45268
rect 4304 45228 4310 45240
rect 4433 45237 4445 45240
rect 4479 45237 4491 45271
rect 4724 45268 4752 45299
rect 4982 45296 4988 45348
rect 5040 45336 5046 45348
rect 5460 45336 5488 45432
rect 8220 45404 8248 45435
rect 8754 45432 8760 45484
rect 8812 45432 8818 45484
rect 9140 45404 9168 45500
rect 8220 45376 9168 45404
rect 8389 45339 8447 45345
rect 5040 45308 5488 45336
rect 5552 45308 7788 45336
rect 5040 45296 5046 45308
rect 5552 45268 5580 45308
rect 4724 45240 5580 45268
rect 4433 45231 4491 45237
rect 7466 45228 7472 45280
rect 7524 45228 7530 45280
rect 7650 45228 7656 45280
rect 7708 45228 7714 45280
rect 7760 45268 7788 45308
rect 8389 45305 8401 45339
rect 8435 45336 8447 45339
rect 9122 45336 9128 45348
rect 8435 45308 9128 45336
rect 8435 45305 8447 45308
rect 8389 45299 8447 45305
rect 9122 45296 9128 45308
rect 9180 45296 9186 45348
rect 9214 45268 9220 45280
rect 7760 45240 9220 45268
rect 9214 45228 9220 45240
rect 9272 45228 9278 45280
rect 1104 45178 9936 45200
rect 1104 45126 3610 45178
rect 3662 45126 3674 45178
rect 3726 45126 3738 45178
rect 3790 45126 3802 45178
rect 3854 45126 3866 45178
rect 3918 45126 5210 45178
rect 5262 45126 5274 45178
rect 5326 45126 5338 45178
rect 5390 45126 5402 45178
rect 5454 45126 5466 45178
rect 5518 45126 6810 45178
rect 6862 45126 6874 45178
rect 6926 45126 6938 45178
rect 6990 45126 7002 45178
rect 7054 45126 7066 45178
rect 7118 45126 8410 45178
rect 8462 45126 8474 45178
rect 8526 45126 8538 45178
rect 8590 45126 8602 45178
rect 8654 45126 8666 45178
rect 8718 45126 9936 45178
rect 1104 45104 9936 45126
rect 4338 45024 4344 45076
rect 4396 45064 4402 45076
rect 4614 45064 4620 45076
rect 4396 45036 4620 45064
rect 4396 45024 4402 45036
rect 4614 45024 4620 45036
rect 4672 45024 4678 45076
rect 4816 45036 9628 45064
rect 2314 44956 2320 45008
rect 2372 44996 2378 45008
rect 4816 45005 4844 45036
rect 9600 45008 9628 45036
rect 4709 44999 4767 45005
rect 4709 44996 4721 44999
rect 2372 44968 4721 44996
rect 2372 44956 2378 44968
rect 4709 44965 4721 44968
rect 4755 44965 4767 44999
rect 4709 44959 4767 44965
rect 4801 44999 4859 45005
rect 4801 44965 4813 44999
rect 4847 44965 4859 44999
rect 4801 44959 4859 44965
rect 5353 44999 5411 45005
rect 5353 44965 5365 44999
rect 5399 44996 5411 44999
rect 5626 44996 5632 45008
rect 5399 44968 5632 44996
rect 5399 44965 5411 44968
rect 5353 44959 5411 44965
rect 5626 44956 5632 44968
rect 5684 44956 5690 45008
rect 6733 44999 6791 45005
rect 6733 44965 6745 44999
rect 6779 44996 6791 44999
rect 9214 44996 9220 45008
rect 6779 44968 9220 44996
rect 6779 44965 6791 44968
rect 6733 44959 6791 44965
rect 9214 44956 9220 44968
rect 9272 44956 9278 45008
rect 9582 44956 9588 45008
rect 9640 44956 9646 45008
rect 2038 44888 2044 44940
rect 2096 44928 2102 44940
rect 4433 44931 4491 44937
rect 4433 44928 4445 44931
rect 2096 44900 4445 44928
rect 2096 44888 2102 44900
rect 4433 44897 4445 44900
rect 4479 44897 4491 44931
rect 4433 44891 4491 44897
rect 4522 44888 4528 44940
rect 4580 44928 4586 44940
rect 7377 44931 7435 44937
rect 7377 44928 7389 44931
rect 4580 44900 4844 44928
rect 4580 44888 4586 44900
rect 934 44820 940 44872
rect 992 44860 998 44872
rect 1397 44863 1455 44869
rect 1397 44860 1409 44863
rect 992 44832 1409 44860
rect 992 44820 998 44832
rect 1397 44829 1409 44832
rect 1443 44829 1455 44863
rect 1397 44823 1455 44829
rect 4183 44863 4241 44869
rect 4183 44829 4195 44863
rect 4229 44860 4241 44863
rect 4229 44832 4568 44860
rect 4229 44829 4241 44832
rect 4183 44823 4241 44829
rect 4540 44792 4568 44832
rect 4614 44820 4620 44872
rect 4672 44820 4678 44872
rect 4816 44860 4844 44900
rect 5368 44900 7389 44928
rect 4905 44863 4963 44869
rect 4905 44860 4917 44863
rect 4816 44832 4917 44860
rect 4905 44829 4917 44832
rect 4951 44829 4963 44863
rect 4905 44823 4963 44829
rect 5258 44820 5264 44872
rect 5316 44820 5322 44872
rect 5368 44792 5396 44900
rect 7377 44897 7389 44900
rect 7423 44928 7435 44931
rect 7834 44928 7840 44940
rect 7423 44900 7840 44928
rect 7423 44897 7435 44900
rect 7377 44891 7435 44897
rect 7834 44888 7840 44900
rect 7892 44888 7898 44940
rect 8110 44888 8116 44940
rect 8168 44888 8174 44940
rect 5442 44820 5448 44872
rect 5500 44820 5506 44872
rect 5537 44863 5595 44869
rect 5537 44829 5549 44863
rect 5583 44860 5595 44863
rect 5902 44860 5908 44872
rect 5583 44832 5908 44860
rect 5583 44829 5595 44832
rect 5537 44823 5595 44829
rect 5902 44820 5908 44832
rect 5960 44820 5966 44872
rect 7193 44863 7251 44869
rect 7193 44829 7205 44863
rect 7239 44860 7251 44863
rect 8128 44860 8156 44888
rect 7239 44832 8156 44860
rect 7239 44829 7251 44832
rect 7193 44823 7251 44829
rect 3528 44764 4476 44792
rect 4540 44764 5396 44792
rect 7101 44795 7159 44801
rect 3528 44736 3556 44764
rect 1581 44727 1639 44733
rect 1581 44693 1593 44727
rect 1627 44724 1639 44727
rect 2682 44724 2688 44736
rect 1627 44696 2688 44724
rect 1627 44693 1639 44696
rect 1581 44687 1639 44693
rect 2682 44684 2688 44696
rect 2740 44684 2746 44736
rect 3510 44684 3516 44736
rect 3568 44684 3574 44736
rect 4448 44724 4476 44764
rect 7101 44761 7113 44795
rect 7147 44792 7159 44795
rect 7742 44792 7748 44804
rect 7147 44764 7748 44792
rect 7147 44761 7159 44764
rect 7101 44755 7159 44761
rect 7742 44752 7748 44764
rect 7800 44752 7806 44804
rect 5077 44727 5135 44733
rect 5077 44724 5089 44727
rect 4448 44696 5089 44724
rect 5077 44693 5089 44696
rect 5123 44693 5135 44727
rect 5077 44687 5135 44693
rect 5902 44684 5908 44736
rect 5960 44724 5966 44736
rect 6086 44724 6092 44736
rect 5960 44696 6092 44724
rect 5960 44684 5966 44696
rect 6086 44684 6092 44696
rect 6144 44684 6150 44736
rect 1104 44634 9936 44656
rect 1104 44582 2950 44634
rect 3002 44582 3014 44634
rect 3066 44582 3078 44634
rect 3130 44582 3142 44634
rect 3194 44582 3206 44634
rect 3258 44582 4550 44634
rect 4602 44582 4614 44634
rect 4666 44582 4678 44634
rect 4730 44582 4742 44634
rect 4794 44582 4806 44634
rect 4858 44582 6150 44634
rect 6202 44582 6214 44634
rect 6266 44582 6278 44634
rect 6330 44582 6342 44634
rect 6394 44582 6406 44634
rect 6458 44582 7750 44634
rect 7802 44582 7814 44634
rect 7866 44582 7878 44634
rect 7930 44582 7942 44634
rect 7994 44582 8006 44634
rect 8058 44582 9350 44634
rect 9402 44582 9414 44634
rect 9466 44582 9478 44634
rect 9530 44582 9542 44634
rect 9594 44582 9606 44634
rect 9658 44582 9936 44634
rect 1104 44560 9936 44582
rect 4157 44523 4215 44529
rect 4157 44489 4169 44523
rect 4203 44520 4215 44523
rect 4706 44520 4712 44532
rect 4203 44492 4712 44520
rect 4203 44489 4215 44492
rect 4157 44483 4215 44489
rect 4706 44480 4712 44492
rect 4764 44480 4770 44532
rect 5258 44520 5264 44532
rect 5184 44492 5264 44520
rect 5184 44452 5212 44492
rect 5258 44480 5264 44492
rect 5316 44480 5322 44532
rect 7650 44480 7656 44532
rect 7708 44480 7714 44532
rect 7742 44480 7748 44532
rect 7800 44520 7806 44532
rect 8202 44520 8208 44532
rect 7800 44492 8208 44520
rect 7800 44480 7806 44492
rect 8202 44480 8208 44492
rect 8260 44480 8266 44532
rect 7668 44452 7696 44480
rect 4356 44424 5212 44452
rect 5276 44424 7696 44452
rect 4356 44396 4384 44424
rect 2866 44344 2872 44396
rect 2924 44344 2930 44396
rect 4338 44393 4344 44396
rect 4331 44387 4344 44393
rect 4331 44384 4343 44387
rect 4299 44356 4343 44384
rect 4331 44353 4343 44356
rect 4331 44347 4344 44353
rect 4338 44344 4344 44347
rect 4396 44344 4402 44396
rect 4617 44387 4675 44393
rect 4617 44353 4629 44387
rect 4663 44384 4675 44387
rect 4706 44384 4712 44396
rect 4663 44356 4712 44384
rect 4663 44353 4675 44356
rect 4617 44347 4675 44353
rect 4706 44344 4712 44356
rect 4764 44344 4770 44396
rect 5000 44393 5028 44424
rect 4985 44387 5043 44393
rect 4985 44353 4997 44387
rect 5031 44353 5043 44387
rect 4985 44347 5043 44353
rect 5074 44344 5080 44396
rect 5132 44344 5138 44396
rect 5166 44344 5172 44396
rect 5224 44344 5230 44396
rect 5276 44393 5304 44424
rect 5261 44387 5319 44393
rect 5261 44353 5273 44387
rect 5307 44353 5319 44387
rect 5261 44347 5319 44353
rect 6638 44344 6644 44396
rect 6696 44384 6702 44396
rect 6733 44387 6791 44393
rect 6733 44384 6745 44387
rect 6696 44356 6745 44384
rect 6696 44344 6702 44356
rect 6733 44353 6745 44356
rect 6779 44353 6791 44387
rect 6733 44347 6791 44353
rect 7000 44387 7058 44393
rect 7000 44353 7012 44387
rect 7046 44384 7058 44387
rect 7558 44384 7564 44396
rect 7046 44356 7564 44384
rect 7046 44353 7058 44356
rect 7000 44347 7058 44353
rect 7558 44344 7564 44356
rect 7616 44344 7622 44396
rect 8110 44344 8116 44396
rect 8168 44344 8174 44396
rect 2884 44316 2912 44344
rect 4433 44319 4491 44325
rect 4433 44316 4445 44319
rect 2884 44288 4445 44316
rect 4433 44285 4445 44288
rect 4479 44285 4491 44319
rect 4433 44279 4491 44285
rect 4525 44319 4583 44325
rect 4525 44285 4537 44319
rect 4571 44316 4583 44319
rect 4890 44316 4896 44328
rect 4571 44288 4896 44316
rect 4571 44285 4583 44288
rect 4525 44279 4583 44285
rect 4890 44276 4896 44288
rect 4948 44276 4954 44328
rect 4706 44208 4712 44260
rect 4764 44248 4770 44260
rect 6730 44248 6736 44260
rect 4764 44220 6736 44248
rect 4764 44208 4770 44220
rect 6730 44208 6736 44220
rect 6788 44208 6794 44260
rect 8128 44248 8156 44344
rect 8128 44220 8248 44248
rect 8220 44192 8248 44220
rect 4338 44140 4344 44192
rect 4396 44180 4402 44192
rect 4801 44183 4859 44189
rect 4801 44180 4813 44183
rect 4396 44152 4813 44180
rect 4396 44140 4402 44152
rect 4801 44149 4813 44152
rect 4847 44149 4859 44183
rect 4801 44143 4859 44149
rect 8110 44140 8116 44192
rect 8168 44140 8174 44192
rect 8202 44140 8208 44192
rect 8260 44140 8266 44192
rect 1104 44090 9936 44112
rect 1104 44038 3610 44090
rect 3662 44038 3674 44090
rect 3726 44038 3738 44090
rect 3790 44038 3802 44090
rect 3854 44038 3866 44090
rect 3918 44038 5210 44090
rect 5262 44038 5274 44090
rect 5326 44038 5338 44090
rect 5390 44038 5402 44090
rect 5454 44038 5466 44090
rect 5518 44038 6810 44090
rect 6862 44038 6874 44090
rect 6926 44038 6938 44090
rect 6990 44038 7002 44090
rect 7054 44038 7066 44090
rect 7118 44038 8410 44090
rect 8462 44038 8474 44090
rect 8526 44038 8538 44090
rect 8590 44038 8602 44090
rect 8654 44038 8666 44090
rect 8718 44038 9936 44090
rect 1104 44016 9936 44038
rect 4062 43936 4068 43988
rect 4120 43976 4126 43988
rect 4341 43979 4399 43985
rect 4341 43976 4353 43979
rect 4120 43948 4353 43976
rect 4120 43936 4126 43948
rect 4341 43945 4353 43948
rect 4387 43945 4399 43979
rect 8202 43976 8208 43988
rect 4341 43939 4399 43945
rect 6564 43948 8208 43976
rect 934 43732 940 43784
rect 992 43772 998 43784
rect 1397 43775 1455 43781
rect 1397 43772 1409 43775
rect 992 43744 1409 43772
rect 992 43732 998 43744
rect 1397 43741 1409 43744
rect 1443 43741 1455 43775
rect 1397 43735 1455 43741
rect 4249 43775 4307 43781
rect 4249 43741 4261 43775
rect 4295 43772 4307 43775
rect 6564 43772 6592 43948
rect 8202 43936 8208 43948
rect 8260 43936 8266 43988
rect 6638 43800 6644 43852
rect 6696 43840 6702 43852
rect 6733 43843 6791 43849
rect 6733 43840 6745 43843
rect 6696 43812 6745 43840
rect 6696 43800 6702 43812
rect 6733 43809 6745 43812
rect 6779 43809 6791 43843
rect 6733 43803 6791 43809
rect 4295 43744 6592 43772
rect 7000 43775 7058 43781
rect 4295 43741 4307 43744
rect 4249 43735 4307 43741
rect 7000 43741 7012 43775
rect 7046 43772 7058 43775
rect 8754 43772 8760 43784
rect 7046 43744 8760 43772
rect 7046 43741 7058 43744
rect 7000 43735 7058 43741
rect 8754 43732 8760 43744
rect 8812 43772 8818 43784
rect 9030 43772 9036 43784
rect 8812 43744 9036 43772
rect 8812 43732 8818 43744
rect 9030 43732 9036 43744
rect 9088 43732 9094 43784
rect 2746 43676 7236 43704
rect 1581 43639 1639 43645
rect 1581 43605 1593 43639
rect 1627 43636 1639 43639
rect 2746 43636 2774 43676
rect 7208 43648 7236 43676
rect 1627 43608 2774 43636
rect 4709 43639 4767 43645
rect 1627 43605 1639 43608
rect 1581 43599 1639 43605
rect 4709 43605 4721 43639
rect 4755 43636 4767 43639
rect 4890 43636 4896 43648
rect 4755 43608 4896 43636
rect 4755 43605 4767 43608
rect 4709 43599 4767 43605
rect 4890 43596 4896 43608
rect 4948 43596 4954 43648
rect 7190 43596 7196 43648
rect 7248 43596 7254 43648
rect 8113 43639 8171 43645
rect 8113 43605 8125 43639
rect 8159 43636 8171 43639
rect 9030 43636 9036 43648
rect 8159 43608 9036 43636
rect 8159 43605 8171 43608
rect 8113 43599 8171 43605
rect 9030 43596 9036 43608
rect 9088 43596 9094 43648
rect 1104 43546 9936 43568
rect 1104 43494 2950 43546
rect 3002 43494 3014 43546
rect 3066 43494 3078 43546
rect 3130 43494 3142 43546
rect 3194 43494 3206 43546
rect 3258 43494 4550 43546
rect 4602 43494 4614 43546
rect 4666 43494 4678 43546
rect 4730 43494 4742 43546
rect 4794 43494 4806 43546
rect 4858 43494 6150 43546
rect 6202 43494 6214 43546
rect 6266 43494 6278 43546
rect 6330 43494 6342 43546
rect 6394 43494 6406 43546
rect 6458 43494 7750 43546
rect 7802 43494 7814 43546
rect 7866 43494 7878 43546
rect 7930 43494 7942 43546
rect 7994 43494 8006 43546
rect 8058 43494 9350 43546
rect 9402 43494 9414 43546
rect 9466 43494 9478 43546
rect 9530 43494 9542 43546
rect 9594 43494 9606 43546
rect 9658 43494 9936 43546
rect 1104 43472 9936 43494
rect 7742 43392 7748 43444
rect 7800 43432 7806 43444
rect 8202 43432 8208 43444
rect 7800 43404 8208 43432
rect 7800 43392 7806 43404
rect 8202 43392 8208 43404
rect 8260 43392 8266 43444
rect 7000 43367 7058 43373
rect 7000 43333 7012 43367
rect 7046 43364 7058 43367
rect 7650 43364 7656 43376
rect 7046 43336 7656 43364
rect 7046 43333 7058 43336
rect 7000 43327 7058 43333
rect 7650 43324 7656 43336
rect 7708 43364 7714 43376
rect 8662 43364 8668 43376
rect 7708 43336 8668 43364
rect 7708 43324 7714 43336
rect 8662 43324 8668 43336
rect 8720 43324 8726 43376
rect 6638 43256 6644 43308
rect 6696 43296 6702 43308
rect 6733 43299 6791 43305
rect 6733 43296 6745 43299
rect 6696 43268 6745 43296
rect 6696 43256 6702 43268
rect 6733 43265 6745 43268
rect 6779 43265 6791 43299
rect 6733 43259 6791 43265
rect 8110 43052 8116 43104
rect 8168 43052 8174 43104
rect 1104 43002 9936 43024
rect 1104 42950 3610 43002
rect 3662 42950 3674 43002
rect 3726 42950 3738 43002
rect 3790 42950 3802 43002
rect 3854 42950 3866 43002
rect 3918 42950 5210 43002
rect 5262 42950 5274 43002
rect 5326 42950 5338 43002
rect 5390 42950 5402 43002
rect 5454 42950 5466 43002
rect 5518 42950 6810 43002
rect 6862 42950 6874 43002
rect 6926 42950 6938 43002
rect 6990 42950 7002 43002
rect 7054 42950 7066 43002
rect 7118 42950 8410 43002
rect 8462 42950 8474 43002
rect 8526 42950 8538 43002
rect 8590 42950 8602 43002
rect 8654 42950 8666 43002
rect 8718 42950 9936 43002
rect 1104 42928 9936 42950
rect 5902 42888 5908 42900
rect 5368 42860 5908 42888
rect 3970 42780 3976 42832
rect 4028 42820 4034 42832
rect 4801 42823 4859 42829
rect 4801 42820 4813 42823
rect 4028 42792 4813 42820
rect 4028 42780 4034 42792
rect 4801 42789 4813 42792
rect 4847 42789 4859 42823
rect 4801 42783 4859 42789
rect 3326 42712 3332 42764
rect 3384 42752 3390 42764
rect 3384 42724 4292 42752
rect 3384 42712 3390 42724
rect 1946 42644 1952 42696
rect 2004 42684 2010 42696
rect 2590 42684 2596 42696
rect 2004 42656 2596 42684
rect 2004 42644 2010 42656
rect 2590 42644 2596 42656
rect 2648 42684 2654 42696
rect 4264 42693 4292 42724
rect 4522 42712 4528 42764
rect 4580 42752 4586 42764
rect 4893 42755 4951 42761
rect 4893 42752 4905 42755
rect 4580 42724 4905 42752
rect 4580 42712 4586 42724
rect 4893 42721 4905 42724
rect 4939 42721 4951 42755
rect 4893 42715 4951 42721
rect 4065 42687 4123 42693
rect 4065 42684 4077 42687
rect 2648 42656 4077 42684
rect 2648 42644 2654 42656
rect 4065 42653 4077 42656
rect 4111 42653 4123 42687
rect 4065 42647 4123 42653
rect 4249 42687 4307 42693
rect 4249 42653 4261 42687
rect 4295 42653 4307 42687
rect 4709 42687 4767 42693
rect 4709 42684 4721 42687
rect 4249 42647 4307 42653
rect 4356 42656 4721 42684
rect 934 42576 940 42628
rect 992 42616 998 42628
rect 1489 42619 1547 42625
rect 1489 42616 1501 42619
rect 992 42588 1501 42616
rect 992 42576 998 42588
rect 1489 42585 1501 42588
rect 1535 42585 1547 42619
rect 1489 42579 1547 42585
rect 1857 42619 1915 42625
rect 1857 42585 1869 42619
rect 1903 42616 1915 42619
rect 4356 42616 4384 42656
rect 4709 42653 4721 42656
rect 4755 42653 4767 42687
rect 4709 42647 4767 42653
rect 4985 42687 5043 42693
rect 4985 42653 4997 42687
rect 5031 42684 5043 42687
rect 5258 42684 5264 42696
rect 5031 42656 5264 42684
rect 5031 42653 5043 42656
rect 4985 42647 5043 42653
rect 1903 42588 2774 42616
rect 1903 42585 1915 42588
rect 1857 42579 1915 42585
rect 2746 42548 2774 42588
rect 4080 42588 4384 42616
rect 4433 42619 4491 42625
rect 4080 42560 4108 42588
rect 4433 42585 4445 42619
rect 4479 42616 4491 42619
rect 4724 42616 4752 42647
rect 5258 42644 5264 42656
rect 5316 42644 5322 42696
rect 5368 42693 5396 42860
rect 5902 42848 5908 42860
rect 5960 42848 5966 42900
rect 7190 42780 7196 42832
rect 7248 42820 7254 42832
rect 8662 42820 8668 42832
rect 7248 42792 8668 42820
rect 7248 42780 7254 42792
rect 8662 42780 8668 42792
rect 8720 42780 8726 42832
rect 5537 42755 5595 42761
rect 5537 42721 5549 42755
rect 5583 42752 5595 42755
rect 5718 42752 5724 42764
rect 5583 42724 5724 42752
rect 5583 42721 5595 42724
rect 5537 42715 5595 42721
rect 5718 42712 5724 42724
rect 5776 42712 5782 42764
rect 7101 42755 7159 42761
rect 7101 42721 7113 42755
rect 7147 42752 7159 42755
rect 7742 42752 7748 42764
rect 7147 42724 7748 42752
rect 7147 42721 7159 42724
rect 7101 42715 7159 42721
rect 7742 42712 7748 42724
rect 7800 42712 7806 42764
rect 5353 42687 5411 42693
rect 5353 42653 5365 42687
rect 5399 42653 5411 42687
rect 5353 42647 5411 42653
rect 5368 42616 5396 42647
rect 5442 42644 5448 42696
rect 5500 42644 5506 42696
rect 5629 42687 5687 42693
rect 5629 42653 5641 42687
rect 5675 42684 5687 42687
rect 8294 42684 8300 42696
rect 5675 42656 8300 42684
rect 5675 42653 5687 42656
rect 5629 42647 5687 42653
rect 8294 42644 8300 42656
rect 8352 42644 8358 42696
rect 8570 42644 8576 42696
rect 8628 42684 8634 42696
rect 8846 42684 8852 42696
rect 8628 42656 8852 42684
rect 8628 42644 8634 42656
rect 8846 42644 8852 42656
rect 8904 42644 8910 42696
rect 4479 42588 4672 42616
rect 4724 42588 5396 42616
rect 4479 42585 4491 42588
rect 4433 42579 4491 42585
rect 3878 42548 3884 42560
rect 2746 42520 3884 42548
rect 3878 42508 3884 42520
rect 3936 42508 3942 42560
rect 4062 42508 4068 42560
rect 4120 42508 4126 42560
rect 4338 42508 4344 42560
rect 4396 42548 4402 42560
rect 4525 42551 4583 42557
rect 4525 42548 4537 42551
rect 4396 42520 4537 42548
rect 4396 42508 4402 42520
rect 4525 42517 4537 42520
rect 4571 42517 4583 42551
rect 4644 42548 4672 42588
rect 5534 42576 5540 42628
rect 5592 42616 5598 42628
rect 6825 42619 6883 42625
rect 6825 42616 6837 42619
rect 5592 42588 6837 42616
rect 5592 42576 5598 42588
rect 6825 42585 6837 42588
rect 6871 42585 6883 42619
rect 6825 42579 6883 42585
rect 5074 42548 5080 42560
rect 4644 42520 5080 42548
rect 4525 42511 4583 42517
rect 5074 42508 5080 42520
rect 5132 42508 5138 42560
rect 5166 42508 5172 42560
rect 5224 42508 5230 42560
rect 5258 42508 5264 42560
rect 5316 42548 5322 42560
rect 6457 42551 6515 42557
rect 6457 42548 6469 42551
rect 5316 42520 6469 42548
rect 5316 42508 5322 42520
rect 6457 42517 6469 42520
rect 6503 42517 6515 42551
rect 6457 42511 6515 42517
rect 6917 42551 6975 42557
rect 6917 42517 6929 42551
rect 6963 42548 6975 42551
rect 7374 42548 7380 42560
rect 6963 42520 7380 42548
rect 6963 42517 6975 42520
rect 6917 42511 6975 42517
rect 7374 42508 7380 42520
rect 7432 42508 7438 42560
rect 7742 42508 7748 42560
rect 7800 42548 7806 42560
rect 8294 42548 8300 42560
rect 7800 42520 8300 42548
rect 7800 42508 7806 42520
rect 8294 42508 8300 42520
rect 8352 42508 8358 42560
rect 1104 42458 9936 42480
rect 1104 42406 2950 42458
rect 3002 42406 3014 42458
rect 3066 42406 3078 42458
rect 3130 42406 3142 42458
rect 3194 42406 3206 42458
rect 3258 42406 4550 42458
rect 4602 42406 4614 42458
rect 4666 42406 4678 42458
rect 4730 42406 4742 42458
rect 4794 42406 4806 42458
rect 4858 42406 6150 42458
rect 6202 42406 6214 42458
rect 6266 42406 6278 42458
rect 6330 42406 6342 42458
rect 6394 42406 6406 42458
rect 6458 42406 7750 42458
rect 7802 42406 7814 42458
rect 7866 42406 7878 42458
rect 7930 42406 7942 42458
rect 7994 42406 8006 42458
rect 8058 42406 9350 42458
rect 9402 42406 9414 42458
rect 9466 42406 9478 42458
rect 9530 42406 9542 42458
rect 9594 42406 9606 42458
rect 9658 42406 9936 42458
rect 1104 42384 9936 42406
rect 2498 42304 2504 42356
rect 2556 42304 2562 42356
rect 3970 42304 3976 42356
rect 4028 42344 4034 42356
rect 5258 42344 5264 42356
rect 4028 42316 5264 42344
rect 4028 42304 4034 42316
rect 5258 42304 5264 42316
rect 5316 42304 5322 42356
rect 7742 42304 7748 42356
rect 7800 42344 7806 42356
rect 9950 42344 9956 42356
rect 7800 42316 9956 42344
rect 7800 42304 7806 42316
rect 9950 42304 9956 42316
rect 10008 42304 10014 42356
rect 2516 42276 2544 42304
rect 5442 42276 5448 42288
rect 2516 42248 5448 42276
rect 5442 42236 5448 42248
rect 5500 42236 5506 42288
rect 7000 42279 7058 42285
rect 7000 42245 7012 42279
rect 7046 42276 7058 42279
rect 7282 42276 7288 42288
rect 7046 42248 7288 42276
rect 7046 42245 7058 42248
rect 7000 42239 7058 42245
rect 7282 42236 7288 42248
rect 7340 42236 7346 42288
rect 2590 42168 2596 42220
rect 2648 42208 2654 42220
rect 2648 42180 2774 42208
rect 2648 42168 2654 42180
rect 2746 42140 2774 42180
rect 6638 42168 6644 42220
rect 6696 42208 6702 42220
rect 6733 42211 6791 42217
rect 6733 42208 6745 42211
rect 6696 42180 6745 42208
rect 6696 42168 6702 42180
rect 6733 42177 6745 42180
rect 6779 42177 6791 42211
rect 10042 42208 10048 42220
rect 6733 42171 6791 42177
rect 6840 42180 10048 42208
rect 6840 42140 6868 42180
rect 10042 42168 10048 42180
rect 10100 42168 10106 42220
rect 2746 42112 6868 42140
rect 1578 42032 1584 42084
rect 1636 42072 1642 42084
rect 3326 42072 3332 42084
rect 1636 42044 3332 42072
rect 1636 42032 1642 42044
rect 3326 42032 3332 42044
rect 3384 42032 3390 42084
rect 3878 42032 3884 42084
rect 3936 42072 3942 42084
rect 3936 42044 5580 42072
rect 3936 42032 3942 42044
rect 5552 42016 5580 42044
rect 1946 41964 1952 42016
rect 2004 42004 2010 42016
rect 5166 42004 5172 42016
rect 2004 41976 5172 42004
rect 2004 41964 2010 41976
rect 5166 41964 5172 41976
rect 5224 41964 5230 42016
rect 5534 41964 5540 42016
rect 5592 41964 5598 42016
rect 7374 41964 7380 42016
rect 7432 42004 7438 42016
rect 8113 42007 8171 42013
rect 8113 42004 8125 42007
rect 7432 41976 8125 42004
rect 7432 41964 7438 41976
rect 8113 41973 8125 41976
rect 8159 41973 8171 42007
rect 8113 41967 8171 41973
rect 8570 41964 8576 42016
rect 8628 42004 8634 42016
rect 8846 42004 8852 42016
rect 8628 41976 8852 42004
rect 8628 41964 8634 41976
rect 8846 41964 8852 41976
rect 8904 41964 8910 42016
rect 1104 41914 9936 41936
rect 1104 41862 3610 41914
rect 3662 41862 3674 41914
rect 3726 41862 3738 41914
rect 3790 41862 3802 41914
rect 3854 41862 3866 41914
rect 3918 41862 5210 41914
rect 5262 41862 5274 41914
rect 5326 41862 5338 41914
rect 5390 41862 5402 41914
rect 5454 41862 5466 41914
rect 5518 41862 6810 41914
rect 6862 41862 6874 41914
rect 6926 41862 6938 41914
rect 6990 41862 7002 41914
rect 7054 41862 7066 41914
rect 7118 41862 8410 41914
rect 8462 41862 8474 41914
rect 8526 41862 8538 41914
rect 8590 41862 8602 41914
rect 8654 41862 8666 41914
rect 8718 41862 9936 41914
rect 1104 41840 9936 41862
rect 4154 41760 4160 41812
rect 4212 41800 4218 41812
rect 4212 41772 4568 41800
rect 4212 41760 4218 41772
rect 2774 41692 2780 41744
rect 2832 41732 2838 41744
rect 4540 41741 4568 41772
rect 4433 41735 4491 41741
rect 4433 41732 4445 41735
rect 2832 41704 4445 41732
rect 2832 41692 2838 41704
rect 4433 41701 4445 41704
rect 4479 41701 4491 41735
rect 4433 41695 4491 41701
rect 4525 41735 4583 41741
rect 4525 41701 4537 41735
rect 4571 41701 4583 41735
rect 4525 41695 4583 41701
rect 4341 41599 4399 41605
rect 4341 41565 4353 41599
rect 4387 41596 4399 41599
rect 4522 41596 4528 41608
rect 4387 41568 4528 41596
rect 4387 41565 4399 41568
rect 4341 41559 4399 41565
rect 4522 41556 4528 41568
rect 4580 41556 4586 41608
rect 4617 41599 4675 41605
rect 4617 41565 4629 41599
rect 4663 41596 4675 41599
rect 4890 41596 4896 41608
rect 4663 41568 4896 41596
rect 4663 41565 4675 41568
rect 4617 41559 4675 41565
rect 4890 41556 4896 41568
rect 4948 41556 4954 41608
rect 7282 41556 7288 41608
rect 7340 41596 7346 41608
rect 7650 41596 7656 41608
rect 7340 41568 7656 41596
rect 7340 41556 7346 41568
rect 7650 41556 7656 41568
rect 7708 41556 7714 41608
rect 934 41488 940 41540
rect 992 41528 998 41540
rect 1489 41531 1547 41537
rect 1489 41528 1501 41531
rect 992 41500 1501 41528
rect 992 41488 998 41500
rect 1489 41497 1501 41500
rect 1535 41497 1547 41531
rect 1489 41491 1547 41497
rect 1857 41531 1915 41537
rect 1857 41497 1869 41531
rect 1903 41528 1915 41531
rect 2130 41528 2136 41540
rect 1903 41500 2136 41528
rect 1903 41497 1915 41500
rect 1857 41491 1915 41497
rect 2130 41488 2136 41500
rect 2188 41488 2194 41540
rect 2498 41420 2504 41472
rect 2556 41460 2562 41472
rect 4157 41463 4215 41469
rect 4157 41460 4169 41463
rect 2556 41432 4169 41460
rect 2556 41420 2562 41432
rect 4157 41429 4169 41432
rect 4203 41429 4215 41463
rect 4157 41423 4215 41429
rect 1104 41370 9936 41392
rect 1104 41318 2950 41370
rect 3002 41318 3014 41370
rect 3066 41318 3078 41370
rect 3130 41318 3142 41370
rect 3194 41318 3206 41370
rect 3258 41318 4550 41370
rect 4602 41318 4614 41370
rect 4666 41318 4678 41370
rect 4730 41318 4742 41370
rect 4794 41318 4806 41370
rect 4858 41318 6150 41370
rect 6202 41318 6214 41370
rect 6266 41318 6278 41370
rect 6330 41318 6342 41370
rect 6394 41318 6406 41370
rect 6458 41318 7750 41370
rect 7802 41318 7814 41370
rect 7866 41318 7878 41370
rect 7930 41318 7942 41370
rect 7994 41318 8006 41370
rect 8058 41318 9350 41370
rect 9402 41318 9414 41370
rect 9466 41318 9478 41370
rect 9530 41318 9542 41370
rect 9594 41318 9606 41370
rect 9658 41318 9936 41370
rect 1104 41296 9936 41318
rect 1026 41080 1032 41132
rect 1084 41120 1090 41132
rect 1489 41123 1547 41129
rect 1489 41120 1501 41123
rect 1084 41092 1501 41120
rect 1084 41080 1090 41092
rect 1489 41089 1501 41092
rect 1535 41089 1547 41123
rect 1489 41083 1547 41089
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 4062 40916 4068 40928
rect 1811 40888 4068 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 4062 40876 4068 40888
rect 4120 40876 4126 40928
rect 1104 40826 9936 40848
rect 1104 40774 3610 40826
rect 3662 40774 3674 40826
rect 3726 40774 3738 40826
rect 3790 40774 3802 40826
rect 3854 40774 3866 40826
rect 3918 40774 5210 40826
rect 5262 40774 5274 40826
rect 5326 40774 5338 40826
rect 5390 40774 5402 40826
rect 5454 40774 5466 40826
rect 5518 40774 6810 40826
rect 6862 40774 6874 40826
rect 6926 40774 6938 40826
rect 6990 40774 7002 40826
rect 7054 40774 7066 40826
rect 7118 40774 8410 40826
rect 8462 40774 8474 40826
rect 8526 40774 8538 40826
rect 8590 40774 8602 40826
rect 8654 40774 8666 40826
rect 8718 40774 9936 40826
rect 1104 40752 9936 40774
rect 5626 40672 5632 40724
rect 5684 40712 5690 40724
rect 6822 40712 6828 40724
rect 5684 40684 6828 40712
rect 5684 40672 5690 40684
rect 6822 40672 6828 40684
rect 6880 40672 6886 40724
rect 9122 40712 9128 40724
rect 7668 40684 9128 40712
rect 7558 40644 7564 40656
rect 7392 40616 7564 40644
rect 4338 40536 4344 40588
rect 4396 40576 4402 40588
rect 4798 40576 4804 40588
rect 4396 40548 4804 40576
rect 4396 40536 4402 40548
rect 4798 40536 4804 40548
rect 4856 40536 4862 40588
rect 566 40468 572 40520
rect 624 40468 630 40520
rect 2590 40468 2596 40520
rect 2648 40508 2654 40520
rect 7392 40517 7420 40616
rect 7558 40604 7564 40616
rect 7616 40604 7622 40656
rect 7668 40585 7696 40684
rect 9122 40672 9128 40684
rect 9180 40672 9186 40724
rect 8018 40604 8024 40656
rect 8076 40604 8082 40656
rect 7653 40579 7711 40585
rect 7653 40545 7665 40579
rect 7699 40545 7711 40579
rect 7653 40539 7711 40545
rect 7377 40511 7435 40517
rect 2648 40480 7328 40508
rect 2648 40468 2654 40480
rect 584 40440 612 40468
rect 4338 40440 4344 40452
rect 584 40412 4344 40440
rect 4338 40400 4344 40412
rect 4396 40440 4402 40452
rect 4525 40443 4583 40449
rect 4525 40440 4537 40443
rect 4396 40412 4537 40440
rect 4396 40400 4402 40412
rect 4525 40409 4537 40412
rect 4571 40409 4583 40443
rect 4525 40403 4583 40409
rect 4709 40443 4767 40449
rect 4709 40409 4721 40443
rect 4755 40440 4767 40443
rect 5902 40440 5908 40452
rect 4755 40412 5908 40440
rect 4755 40409 4767 40412
rect 4709 40403 4767 40409
rect 5902 40400 5908 40412
rect 5960 40400 5966 40452
rect 5994 40400 6000 40452
rect 6052 40440 6058 40452
rect 7098 40440 7104 40452
rect 6052 40412 7104 40440
rect 6052 40400 6058 40412
rect 7098 40400 7104 40412
rect 7156 40400 7162 40452
rect 4798 40332 4804 40384
rect 4856 40372 4862 40384
rect 4982 40372 4988 40384
rect 4856 40344 4988 40372
rect 4856 40332 4862 40344
rect 4982 40332 4988 40344
rect 5040 40332 5046 40384
rect 5626 40332 5632 40384
rect 5684 40372 5690 40384
rect 7009 40375 7067 40381
rect 7009 40372 7021 40375
rect 5684 40344 7021 40372
rect 5684 40332 5690 40344
rect 7009 40341 7021 40344
rect 7055 40341 7067 40375
rect 7300 40372 7328 40480
rect 7377 40477 7389 40511
rect 7423 40477 7435 40511
rect 7377 40471 7435 40477
rect 7558 40468 7564 40520
rect 7616 40508 7622 40520
rect 8036 40508 8064 40604
rect 8846 40536 8852 40588
rect 8904 40536 8910 40588
rect 7616 40480 8064 40508
rect 7616 40468 7622 40480
rect 7469 40443 7527 40449
rect 7469 40409 7481 40443
rect 7515 40440 7527 40443
rect 8864 40440 8892 40536
rect 7515 40412 8892 40440
rect 7515 40409 7527 40412
rect 7469 40403 7527 40409
rect 8386 40372 8392 40384
rect 7300 40344 8392 40372
rect 7009 40335 7067 40341
rect 8386 40332 8392 40344
rect 8444 40332 8450 40384
rect 1104 40282 9936 40304
rect 1104 40230 2950 40282
rect 3002 40230 3014 40282
rect 3066 40230 3078 40282
rect 3130 40230 3142 40282
rect 3194 40230 3206 40282
rect 3258 40230 4550 40282
rect 4602 40230 4614 40282
rect 4666 40230 4678 40282
rect 4730 40230 4742 40282
rect 4794 40230 4806 40282
rect 4858 40230 6150 40282
rect 6202 40230 6214 40282
rect 6266 40230 6278 40282
rect 6330 40230 6342 40282
rect 6394 40230 6406 40282
rect 6458 40230 7750 40282
rect 7802 40230 7814 40282
rect 7866 40230 7878 40282
rect 7930 40230 7942 40282
rect 7994 40230 8006 40282
rect 8058 40230 9350 40282
rect 9402 40230 9414 40282
rect 9466 40230 9478 40282
rect 9530 40230 9542 40282
rect 9594 40230 9606 40282
rect 9658 40230 9936 40282
rect 1104 40208 9936 40230
rect 4798 40128 4804 40180
rect 4856 40168 4862 40180
rect 5166 40168 5172 40180
rect 4856 40140 5172 40168
rect 4856 40128 4862 40140
rect 5166 40128 5172 40140
rect 5224 40128 5230 40180
rect 5810 40128 5816 40180
rect 5868 40168 5874 40180
rect 6917 40171 6975 40177
rect 6917 40168 6929 40171
rect 5868 40140 6929 40168
rect 5868 40128 5874 40140
rect 6917 40137 6929 40140
rect 6963 40137 6975 40171
rect 6917 40131 6975 40137
rect 7098 40128 7104 40180
rect 7156 40168 7162 40180
rect 7377 40171 7435 40177
rect 7377 40168 7389 40171
rect 7156 40140 7389 40168
rect 7156 40128 7162 40140
rect 7377 40137 7389 40140
rect 7423 40137 7435 40171
rect 7377 40131 7435 40137
rect 7466 40128 7472 40180
rect 7524 40168 7530 40180
rect 8113 40171 8171 40177
rect 8113 40168 8125 40171
rect 7524 40140 8125 40168
rect 7524 40128 7530 40140
rect 8113 40137 8125 40140
rect 8159 40137 8171 40171
rect 8113 40131 8171 40137
rect 8573 40171 8631 40177
rect 8573 40137 8585 40171
rect 8619 40137 8631 40171
rect 8573 40131 8631 40137
rect 1486 40060 1492 40112
rect 1544 40060 1550 40112
rect 7285 40103 7343 40109
rect 7285 40069 7297 40103
rect 7331 40100 7343 40103
rect 7650 40100 7656 40112
rect 7331 40072 7656 40100
rect 7331 40069 7343 40072
rect 7285 40063 7343 40069
rect 7650 40060 7656 40072
rect 7708 40060 7714 40112
rect 8588 40100 8616 40131
rect 8938 40128 8944 40180
rect 8996 40128 9002 40180
rect 9950 40100 9956 40112
rect 8588 40072 9956 40100
rect 9950 40060 9956 40072
rect 10008 40060 10014 40112
rect 7576 40004 8432 40032
rect 7466 39924 7472 39976
rect 7524 39964 7530 39976
rect 7576 39973 7604 40004
rect 7561 39967 7619 39973
rect 7561 39964 7573 39967
rect 7524 39936 7573 39964
rect 7524 39924 7530 39936
rect 7561 39933 7573 39936
rect 7607 39933 7619 39967
rect 7561 39927 7619 39933
rect 8018 39924 8024 39976
rect 8076 39924 8082 39976
rect 8110 39924 8116 39976
rect 8168 39964 8174 39976
rect 8205 39967 8263 39973
rect 8205 39964 8217 39967
rect 8168 39936 8217 39964
rect 8168 39924 8174 39936
rect 8205 39933 8217 39936
rect 8251 39933 8263 39967
rect 8205 39927 8263 39933
rect 8294 39924 8300 39976
rect 8352 39924 8358 39976
rect 8404 39964 8432 40004
rect 9030 39992 9036 40044
rect 9088 39992 9094 40044
rect 9122 39992 9128 40044
rect 9180 40032 9186 40044
rect 9180 40004 9260 40032
rect 9180 39992 9186 40004
rect 9232 39973 9260 40004
rect 9217 39967 9275 39973
rect 9217 39964 9229 39967
rect 8404 39936 9229 39964
rect 9217 39933 9229 39936
rect 9263 39933 9275 39967
rect 9217 39927 9275 39933
rect 6822 39856 6828 39908
rect 6880 39896 6886 39908
rect 8036 39896 8064 39924
rect 6880 39868 8064 39896
rect 6880 39856 6886 39868
rect 1765 39831 1823 39837
rect 1765 39797 1777 39831
rect 1811 39828 1823 39831
rect 2682 39828 2688 39840
rect 1811 39800 2688 39828
rect 1811 39797 1823 39800
rect 1765 39791 1823 39797
rect 2682 39788 2688 39800
rect 2740 39788 2746 39840
rect 7745 39831 7803 39837
rect 7745 39797 7757 39831
rect 7791 39828 7803 39831
rect 8846 39828 8852 39840
rect 7791 39800 8852 39828
rect 7791 39797 7803 39800
rect 7745 39791 7803 39797
rect 8846 39788 8852 39800
rect 8904 39788 8910 39840
rect 1104 39738 9936 39760
rect 1104 39686 3610 39738
rect 3662 39686 3674 39738
rect 3726 39686 3738 39738
rect 3790 39686 3802 39738
rect 3854 39686 3866 39738
rect 3918 39686 5210 39738
rect 5262 39686 5274 39738
rect 5326 39686 5338 39738
rect 5390 39686 5402 39738
rect 5454 39686 5466 39738
rect 5518 39686 6810 39738
rect 6862 39686 6874 39738
rect 6926 39686 6938 39738
rect 6990 39686 7002 39738
rect 7054 39686 7066 39738
rect 7118 39686 8410 39738
rect 8462 39686 8474 39738
rect 8526 39686 8538 39738
rect 8590 39686 8602 39738
rect 8654 39686 8666 39738
rect 8718 39686 9936 39738
rect 1104 39664 9936 39686
rect 4338 39584 4344 39636
rect 4396 39624 4402 39636
rect 4433 39627 4491 39633
rect 4433 39624 4445 39627
rect 4396 39596 4445 39624
rect 4396 39584 4402 39596
rect 4433 39593 4445 39596
rect 4479 39593 4491 39627
rect 4433 39587 4491 39593
rect 5534 39584 5540 39636
rect 5592 39624 5598 39636
rect 6914 39624 6920 39636
rect 5592 39596 6920 39624
rect 5592 39584 5598 39596
rect 6914 39584 6920 39596
rect 6972 39584 6978 39636
rect 5442 39516 5448 39568
rect 5500 39556 5506 39568
rect 7377 39559 7435 39565
rect 7377 39556 7389 39559
rect 5500 39528 7389 39556
rect 5500 39516 5506 39528
rect 7377 39525 7389 39528
rect 7423 39525 7435 39559
rect 7377 39519 7435 39525
rect 7466 39516 7472 39568
rect 7524 39516 7530 39568
rect 7193 39491 7251 39497
rect 7193 39457 7205 39491
rect 7239 39488 7251 39491
rect 7484 39488 7512 39516
rect 7239 39460 7512 39488
rect 7239 39457 7251 39460
rect 7193 39451 7251 39457
rect 7558 39448 7564 39500
rect 7616 39448 7622 39500
rect 7650 39448 7656 39500
rect 7708 39448 7714 39500
rect 7834 39448 7840 39500
rect 7892 39448 7898 39500
rect 7929 39491 7987 39497
rect 7929 39457 7941 39491
rect 7975 39457 7987 39491
rect 7929 39451 7987 39457
rect 658 39380 664 39432
rect 716 39420 722 39432
rect 4341 39423 4399 39429
rect 4341 39420 4353 39423
rect 716 39392 4353 39420
rect 716 39380 722 39392
rect 4341 39389 4353 39392
rect 4387 39420 4399 39423
rect 5534 39420 5540 39432
rect 4387 39392 5540 39420
rect 4387 39389 4399 39392
rect 4341 39383 4399 39389
rect 5534 39380 5540 39392
rect 5592 39380 5598 39432
rect 6917 39423 6975 39429
rect 6917 39389 6929 39423
rect 6963 39420 6975 39423
rect 7282 39420 7288 39432
rect 6963 39392 7288 39420
rect 6963 39389 6975 39392
rect 6917 39383 6975 39389
rect 7282 39380 7288 39392
rect 7340 39380 7346 39432
rect 7009 39355 7067 39361
rect 7009 39321 7021 39355
rect 7055 39352 7067 39355
rect 7576 39352 7604 39448
rect 7668 39420 7696 39448
rect 7944 39420 7972 39451
rect 7668 39392 7972 39420
rect 7055 39324 7604 39352
rect 7055 39321 7067 39324
rect 7009 39315 7067 39321
rect 4154 39244 4160 39296
rect 4212 39284 4218 39296
rect 4801 39287 4859 39293
rect 4801 39284 4813 39287
rect 4212 39256 4813 39284
rect 4212 39244 4218 39256
rect 4801 39253 4813 39256
rect 4847 39253 4859 39287
rect 4801 39247 4859 39253
rect 5994 39244 6000 39296
rect 6052 39284 6058 39296
rect 6549 39287 6607 39293
rect 6549 39284 6561 39287
rect 6052 39256 6561 39284
rect 6052 39244 6058 39256
rect 6549 39253 6561 39256
rect 6595 39253 6607 39287
rect 6549 39247 6607 39253
rect 6914 39244 6920 39296
rect 6972 39284 6978 39296
rect 7558 39284 7564 39296
rect 6972 39256 7564 39284
rect 6972 39244 6978 39256
rect 7558 39244 7564 39256
rect 7616 39284 7622 39296
rect 7745 39287 7803 39293
rect 7745 39284 7757 39287
rect 7616 39256 7757 39284
rect 7616 39244 7622 39256
rect 7745 39253 7757 39256
rect 7791 39253 7803 39287
rect 7745 39247 7803 39253
rect 1104 39194 9936 39216
rect 1104 39142 2950 39194
rect 3002 39142 3014 39194
rect 3066 39142 3078 39194
rect 3130 39142 3142 39194
rect 3194 39142 3206 39194
rect 3258 39142 4550 39194
rect 4602 39142 4614 39194
rect 4666 39142 4678 39194
rect 4730 39142 4742 39194
rect 4794 39142 4806 39194
rect 4858 39142 6150 39194
rect 6202 39142 6214 39194
rect 6266 39142 6278 39194
rect 6330 39142 6342 39194
rect 6394 39142 6406 39194
rect 6458 39142 7750 39194
rect 7802 39142 7814 39194
rect 7866 39142 7878 39194
rect 7930 39142 7942 39194
rect 7994 39142 8006 39194
rect 8058 39142 9350 39194
rect 9402 39142 9414 39194
rect 9466 39142 9478 39194
rect 9530 39142 9542 39194
rect 9594 39142 9606 39194
rect 9658 39142 9936 39194
rect 1104 39120 9936 39142
rect 1302 39040 1308 39092
rect 1360 39080 1366 39092
rect 6641 39083 6699 39089
rect 6641 39080 6653 39083
rect 1360 39052 6653 39080
rect 1360 39040 1366 39052
rect 6641 39049 6653 39052
rect 6687 39080 6699 39083
rect 7469 39083 7527 39089
rect 7469 39080 7481 39083
rect 6687 39052 7481 39080
rect 6687 39049 6699 39052
rect 6641 39043 6699 39049
rect 7469 39049 7481 39052
rect 7515 39049 7527 39083
rect 7469 39043 7527 39049
rect 4062 38972 4068 39024
rect 4120 39012 4126 39024
rect 4120 38984 5672 39012
rect 4120 38972 4126 38984
rect 1026 38904 1032 38956
rect 1084 38944 1090 38956
rect 1489 38947 1547 38953
rect 1489 38944 1501 38947
rect 1084 38916 1501 38944
rect 1084 38904 1090 38916
rect 1489 38913 1501 38916
rect 1535 38913 1547 38947
rect 1489 38907 1547 38913
rect 5534 38904 5540 38956
rect 5592 38904 5598 38956
rect 5644 38944 5672 38984
rect 6730 38972 6736 39024
rect 6788 39012 6794 39024
rect 7837 39015 7895 39021
rect 7837 39012 7849 39015
rect 6788 38984 7849 39012
rect 6788 38972 6794 38984
rect 7837 38981 7849 38984
rect 7883 38981 7895 39015
rect 7837 38975 7895 38981
rect 7282 38944 7288 38956
rect 5644 38916 7288 38944
rect 7282 38904 7288 38916
rect 7340 38944 7346 38956
rect 7377 38947 7435 38953
rect 7377 38944 7389 38947
rect 7340 38916 7389 38944
rect 7340 38904 7346 38916
rect 7377 38913 7389 38916
rect 7423 38913 7435 38947
rect 7377 38907 7435 38913
rect 1765 38743 1823 38749
rect 1765 38709 1777 38743
rect 1811 38740 1823 38743
rect 2774 38740 2780 38752
rect 1811 38712 2780 38740
rect 1811 38709 1823 38712
rect 1765 38703 1823 38709
rect 2774 38700 2780 38712
rect 2832 38700 2838 38752
rect 5552 38740 5580 38904
rect 7650 38836 7656 38888
rect 7708 38836 7714 38888
rect 6822 38768 6828 38820
rect 6880 38808 6886 38820
rect 6880 38780 9352 38808
rect 6880 38768 6886 38780
rect 6638 38740 6644 38752
rect 5552 38712 6644 38740
rect 6638 38700 6644 38712
rect 6696 38700 6702 38752
rect 7009 38743 7067 38749
rect 7009 38709 7021 38743
rect 7055 38740 7067 38743
rect 9122 38740 9128 38752
rect 7055 38712 9128 38740
rect 7055 38709 7067 38712
rect 7009 38703 7067 38709
rect 9122 38700 9128 38712
rect 9180 38700 9186 38752
rect 9324 38749 9352 38780
rect 9309 38743 9367 38749
rect 9309 38709 9321 38743
rect 9355 38740 9367 38743
rect 11698 38740 11704 38752
rect 9355 38712 11704 38740
rect 9355 38709 9367 38712
rect 9309 38703 9367 38709
rect 11698 38700 11704 38712
rect 11756 38700 11762 38752
rect 1104 38650 9936 38672
rect 1104 38598 3610 38650
rect 3662 38598 3674 38650
rect 3726 38598 3738 38650
rect 3790 38598 3802 38650
rect 3854 38598 3866 38650
rect 3918 38598 5210 38650
rect 5262 38598 5274 38650
rect 5326 38598 5338 38650
rect 5390 38598 5402 38650
rect 5454 38598 5466 38650
rect 5518 38598 6810 38650
rect 6862 38598 6874 38650
rect 6926 38598 6938 38650
rect 6990 38598 7002 38650
rect 7054 38598 7066 38650
rect 7118 38598 8410 38650
rect 8462 38598 8474 38650
rect 8526 38598 8538 38650
rect 8590 38598 8602 38650
rect 8654 38598 8666 38650
rect 8718 38598 9936 38650
rect 1104 38576 9936 38598
rect 1854 38496 1860 38548
rect 1912 38536 1918 38548
rect 2866 38536 2872 38548
rect 1912 38508 2872 38536
rect 1912 38496 1918 38508
rect 2866 38496 2872 38508
rect 2924 38496 2930 38548
rect 7561 38471 7619 38477
rect 7561 38437 7573 38471
rect 7607 38468 7619 38471
rect 11514 38468 11520 38480
rect 7607 38440 11520 38468
rect 7607 38437 7619 38440
rect 7561 38431 7619 38437
rect 11514 38428 11520 38440
rect 11572 38428 11578 38480
rect 8113 38335 8171 38341
rect 8113 38332 8125 38335
rect 7668 38304 8125 38332
rect 7668 38276 7696 38304
rect 8113 38301 8125 38304
rect 8159 38301 8171 38335
rect 8113 38295 8171 38301
rect 7098 38224 7104 38276
rect 7156 38224 7162 38276
rect 7650 38224 7656 38276
rect 7708 38224 7714 38276
rect 7837 38267 7895 38273
rect 7837 38233 7849 38267
rect 7883 38233 7895 38267
rect 7837 38227 7895 38233
rect 7116 38196 7144 38224
rect 7852 38196 7880 38227
rect 7116 38168 7880 38196
rect 8021 38199 8079 38205
rect 8021 38165 8033 38199
rect 8067 38196 8079 38199
rect 8110 38196 8116 38208
rect 8067 38168 8116 38196
rect 8067 38165 8079 38168
rect 8021 38159 8079 38165
rect 8110 38156 8116 38168
rect 8168 38156 8174 38208
rect 1104 38106 9936 38128
rect 1104 38054 2950 38106
rect 3002 38054 3014 38106
rect 3066 38054 3078 38106
rect 3130 38054 3142 38106
rect 3194 38054 3206 38106
rect 3258 38054 4550 38106
rect 4602 38054 4614 38106
rect 4666 38054 4678 38106
rect 4730 38054 4742 38106
rect 4794 38054 4806 38106
rect 4858 38054 6150 38106
rect 6202 38054 6214 38106
rect 6266 38054 6278 38106
rect 6330 38054 6342 38106
rect 6394 38054 6406 38106
rect 6458 38054 7750 38106
rect 7802 38054 7814 38106
rect 7866 38054 7878 38106
rect 7930 38054 7942 38106
rect 7994 38054 8006 38106
rect 8058 38054 9350 38106
rect 9402 38054 9414 38106
rect 9466 38054 9478 38106
rect 9530 38054 9542 38106
rect 9594 38054 9606 38106
rect 9658 38054 9936 38106
rect 1104 38032 9936 38054
rect 7009 37995 7067 38001
rect 7009 37961 7021 37995
rect 7055 37992 7067 37995
rect 7190 37992 7196 38004
rect 7055 37964 7196 37992
rect 7055 37961 7067 37964
rect 7009 37955 7067 37961
rect 7190 37952 7196 37964
rect 7248 37952 7254 38004
rect 7374 37952 7380 38004
rect 7432 37952 7438 38004
rect 8021 37995 8079 38001
rect 8021 37961 8033 37995
rect 8067 37992 8079 37995
rect 8202 37992 8208 38004
rect 8067 37964 8208 37992
rect 8067 37961 8079 37964
rect 8021 37955 8079 37961
rect 8202 37952 8208 37964
rect 8260 37952 8266 38004
rect 7101 37927 7159 37933
rect 7101 37893 7113 37927
rect 7147 37924 7159 37927
rect 7392 37924 7420 37952
rect 7147 37896 7420 37924
rect 7147 37893 7159 37896
rect 7101 37887 7159 37893
rect 1026 37816 1032 37868
rect 1084 37856 1090 37868
rect 1489 37859 1547 37865
rect 1489 37856 1501 37859
rect 1084 37828 1501 37856
rect 1084 37816 1090 37828
rect 1489 37825 1501 37828
rect 1535 37825 1547 37859
rect 1489 37819 1547 37825
rect 7285 37791 7343 37797
rect 7285 37757 7297 37791
rect 7331 37788 7343 37791
rect 7466 37788 7472 37800
rect 7331 37760 7472 37788
rect 7331 37757 7343 37760
rect 7285 37751 7343 37757
rect 7466 37748 7472 37760
rect 7524 37748 7530 37800
rect 7929 37791 7987 37797
rect 7929 37757 7941 37791
rect 7975 37757 7987 37791
rect 7929 37751 7987 37757
rect 7944 37720 7972 37751
rect 8110 37748 8116 37800
rect 8168 37748 8174 37800
rect 7484 37692 7972 37720
rect 7484 37664 7512 37692
rect 1765 37655 1823 37661
rect 1765 37621 1777 37655
rect 1811 37652 1823 37655
rect 2314 37652 2320 37664
rect 1811 37624 2320 37652
rect 1811 37621 1823 37624
rect 1765 37615 1823 37621
rect 2314 37612 2320 37624
rect 2372 37612 2378 37664
rect 4338 37612 4344 37664
rect 4396 37652 4402 37664
rect 6641 37655 6699 37661
rect 6641 37652 6653 37655
rect 4396 37624 6653 37652
rect 4396 37612 4402 37624
rect 6641 37621 6653 37624
rect 6687 37621 6699 37655
rect 6641 37615 6699 37621
rect 7466 37612 7472 37664
rect 7524 37612 7530 37664
rect 7561 37655 7619 37661
rect 7561 37621 7573 37655
rect 7607 37652 7619 37655
rect 11974 37652 11980 37664
rect 7607 37624 11980 37652
rect 7607 37621 7619 37624
rect 7561 37615 7619 37621
rect 11974 37612 11980 37624
rect 12032 37612 12038 37664
rect 1104 37562 9936 37584
rect 1104 37510 3610 37562
rect 3662 37510 3674 37562
rect 3726 37510 3738 37562
rect 3790 37510 3802 37562
rect 3854 37510 3866 37562
rect 3918 37510 5210 37562
rect 5262 37510 5274 37562
rect 5326 37510 5338 37562
rect 5390 37510 5402 37562
rect 5454 37510 5466 37562
rect 5518 37510 6810 37562
rect 6862 37510 6874 37562
rect 6926 37510 6938 37562
rect 6990 37510 7002 37562
rect 7054 37510 7066 37562
rect 7118 37510 8410 37562
rect 8462 37510 8474 37562
rect 8526 37510 8538 37562
rect 8590 37510 8602 37562
rect 8654 37510 8666 37562
rect 8718 37510 9936 37562
rect 1104 37488 9936 37510
rect 2682 37408 2688 37460
rect 2740 37448 2746 37460
rect 7374 37448 7380 37460
rect 2740 37420 7380 37448
rect 2740 37408 2746 37420
rect 7374 37408 7380 37420
rect 7432 37408 7438 37460
rect 8846 37380 8852 37392
rect 5552 37352 8852 37380
rect 5552 37256 5580 37352
rect 8846 37340 8852 37352
rect 8904 37340 8910 37392
rect 6914 37272 6920 37324
rect 6972 37312 6978 37324
rect 7653 37315 7711 37321
rect 7653 37312 7665 37315
rect 6972 37284 7665 37312
rect 6972 37272 6978 37284
rect 7653 37281 7665 37284
rect 7699 37281 7711 37315
rect 7653 37275 7711 37281
rect 7742 37272 7748 37324
rect 7800 37272 7806 37324
rect 1026 37204 1032 37256
rect 1084 37244 1090 37256
rect 1397 37247 1455 37253
rect 1397 37244 1409 37247
rect 1084 37216 1409 37244
rect 1084 37204 1090 37216
rect 1397 37213 1409 37216
rect 1443 37213 1455 37247
rect 1397 37207 1455 37213
rect 1854 37204 1860 37256
rect 1912 37244 1918 37256
rect 4982 37244 4988 37256
rect 1912 37216 4988 37244
rect 1912 37204 1918 37216
rect 4982 37204 4988 37216
rect 5040 37204 5046 37256
rect 5534 37204 5540 37256
rect 5592 37204 5598 37256
rect 9766 37244 9772 37256
rect 7208 37216 9772 37244
rect 1673 37179 1731 37185
rect 1673 37145 1685 37179
rect 1719 37176 1731 37179
rect 2406 37176 2412 37188
rect 1719 37148 2412 37176
rect 1719 37145 1731 37148
rect 1673 37139 1731 37145
rect 2406 37136 2412 37148
rect 2464 37136 2470 37188
rect 474 37068 480 37120
rect 532 37108 538 37120
rect 7098 37108 7104 37120
rect 532 37080 7104 37108
rect 532 37068 538 37080
rect 7098 37068 7104 37080
rect 7156 37068 7162 37120
rect 7208 37117 7236 37216
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 7193 37111 7251 37117
rect 7193 37077 7205 37111
rect 7239 37077 7251 37111
rect 7193 37071 7251 37077
rect 7374 37068 7380 37120
rect 7432 37108 7438 37120
rect 7561 37111 7619 37117
rect 7561 37108 7573 37111
rect 7432 37080 7573 37108
rect 7432 37068 7438 37080
rect 7561 37077 7573 37080
rect 7607 37077 7619 37111
rect 7561 37071 7619 37077
rect 1104 37018 9936 37040
rect 1104 36966 2950 37018
rect 3002 36966 3014 37018
rect 3066 36966 3078 37018
rect 3130 36966 3142 37018
rect 3194 36966 3206 37018
rect 3258 36966 4550 37018
rect 4602 36966 4614 37018
rect 4666 36966 4678 37018
rect 4730 36966 4742 37018
rect 4794 36966 4806 37018
rect 4858 36966 6150 37018
rect 6202 36966 6214 37018
rect 6266 36966 6278 37018
rect 6330 36966 6342 37018
rect 6394 36966 6406 37018
rect 6458 36966 7750 37018
rect 7802 36966 7814 37018
rect 7866 36966 7878 37018
rect 7930 36966 7942 37018
rect 7994 36966 8006 37018
rect 8058 36966 9350 37018
rect 9402 36966 9414 37018
rect 9466 36966 9478 37018
rect 9530 36966 9542 37018
rect 9594 36966 9606 37018
rect 9658 36966 9936 37018
rect 1104 36944 9936 36966
rect 8294 36904 8300 36916
rect 7484 36876 8300 36904
rect 7098 36796 7104 36848
rect 7156 36836 7162 36848
rect 7484 36836 7512 36876
rect 8294 36864 8300 36876
rect 8352 36864 8358 36916
rect 8573 36907 8631 36913
rect 8573 36873 8585 36907
rect 8619 36904 8631 36907
rect 11606 36904 11612 36916
rect 8619 36876 11612 36904
rect 8619 36873 8631 36876
rect 8573 36867 8631 36873
rect 11606 36864 11612 36876
rect 11664 36864 11670 36916
rect 7156 36808 7512 36836
rect 7156 36796 7162 36808
rect 8573 36703 8631 36709
rect 8573 36669 8585 36703
rect 8619 36669 8631 36703
rect 8573 36663 8631 36669
rect 8665 36703 8723 36709
rect 8665 36669 8677 36703
rect 8711 36700 8723 36703
rect 8846 36700 8852 36712
rect 8711 36672 8852 36700
rect 8711 36669 8723 36672
rect 8665 36663 8723 36669
rect 4982 36592 4988 36644
rect 5040 36632 5046 36644
rect 5442 36632 5448 36644
rect 5040 36604 5448 36632
rect 5040 36592 5046 36604
rect 5442 36592 5448 36604
rect 5500 36592 5506 36644
rect 6454 36592 6460 36644
rect 6512 36632 6518 36644
rect 6638 36632 6644 36644
rect 6512 36604 6644 36632
rect 6512 36592 6518 36604
rect 6638 36592 6644 36604
rect 6696 36592 6702 36644
rect 8588 36632 8616 36663
rect 8846 36660 8852 36672
rect 8904 36660 8910 36712
rect 9214 36632 9220 36644
rect 8588 36604 9220 36632
rect 9214 36592 9220 36604
rect 9272 36592 9278 36644
rect 842 36524 848 36576
rect 900 36564 906 36576
rect 8113 36567 8171 36573
rect 8113 36564 8125 36567
rect 900 36536 8125 36564
rect 900 36524 906 36536
rect 8113 36533 8125 36536
rect 8159 36533 8171 36567
rect 8113 36527 8171 36533
rect 1104 36474 9936 36496
rect 1104 36422 3610 36474
rect 3662 36422 3674 36474
rect 3726 36422 3738 36474
rect 3790 36422 3802 36474
rect 3854 36422 3866 36474
rect 3918 36422 5210 36474
rect 5262 36422 5274 36474
rect 5326 36422 5338 36474
rect 5390 36422 5402 36474
rect 5454 36422 5466 36474
rect 5518 36422 6810 36474
rect 6862 36422 6874 36474
rect 6926 36422 6938 36474
rect 6990 36422 7002 36474
rect 7054 36422 7066 36474
rect 7118 36422 8410 36474
rect 8462 36422 8474 36474
rect 8526 36422 8538 36474
rect 8590 36422 8602 36474
rect 8654 36422 8666 36474
rect 8718 36422 9936 36474
rect 1104 36400 9936 36422
rect 1670 36184 1676 36236
rect 1728 36184 1734 36236
rect 8757 36227 8815 36233
rect 2746 36196 8156 36224
rect 1394 36116 1400 36168
rect 1452 36116 1458 36168
rect 1688 36156 1716 36184
rect 2746 36156 2774 36196
rect 8128 36165 8156 36196
rect 8220 36196 8708 36224
rect 1688 36128 2774 36156
rect 8021 36159 8079 36165
rect 8021 36125 8033 36159
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 8113 36159 8171 36165
rect 8113 36125 8125 36159
rect 8159 36125 8171 36159
rect 8113 36119 8171 36125
rect 1210 36048 1216 36100
rect 1268 36088 1274 36100
rect 1673 36091 1731 36097
rect 1673 36088 1685 36091
rect 1268 36060 1685 36088
rect 1268 36048 1274 36060
rect 1673 36057 1685 36060
rect 1719 36057 1731 36091
rect 1673 36051 1731 36057
rect 7377 36091 7435 36097
rect 7377 36057 7389 36091
rect 7423 36088 7435 36091
rect 8036 36088 8064 36119
rect 8220 36088 8248 36196
rect 8297 36159 8355 36165
rect 8297 36125 8309 36159
rect 8343 36125 8355 36159
rect 8680 36156 8708 36196
rect 8757 36193 8769 36227
rect 8803 36224 8815 36227
rect 8846 36224 8852 36236
rect 8803 36196 8852 36224
rect 8803 36193 8815 36196
rect 8757 36187 8815 36193
rect 8846 36184 8852 36196
rect 8904 36184 8910 36236
rect 9122 36156 9128 36168
rect 8680 36128 9128 36156
rect 8297 36119 8355 36125
rect 7423 36060 7972 36088
rect 8036 36060 8248 36088
rect 8312 36088 8340 36119
rect 9122 36116 9128 36128
rect 9180 36116 9186 36168
rect 8846 36088 8852 36100
rect 8312 36060 8852 36088
rect 7423 36057 7435 36060
rect 7377 36051 7435 36057
rect 6546 35980 6552 36032
rect 6604 36020 6610 36032
rect 7190 36020 7196 36032
rect 6604 35992 7196 36020
rect 6604 35980 6610 35992
rect 7190 35980 7196 35992
rect 7248 35980 7254 36032
rect 7469 36023 7527 36029
rect 7469 35989 7481 36023
rect 7515 36020 7527 36023
rect 7650 36020 7656 36032
rect 7515 35992 7656 36020
rect 7515 35989 7527 35992
rect 7469 35983 7527 35989
rect 7650 35980 7656 35992
rect 7708 35980 7714 36032
rect 7944 36020 7972 36060
rect 8312 36020 8340 36060
rect 8846 36048 8852 36060
rect 8904 36048 8910 36100
rect 7944 35992 8340 36020
rect 1104 35930 9936 35952
rect 1104 35878 2950 35930
rect 3002 35878 3014 35930
rect 3066 35878 3078 35930
rect 3130 35878 3142 35930
rect 3194 35878 3206 35930
rect 3258 35878 4550 35930
rect 4602 35878 4614 35930
rect 4666 35878 4678 35930
rect 4730 35878 4742 35930
rect 4794 35878 4806 35930
rect 4858 35878 6150 35930
rect 6202 35878 6214 35930
rect 6266 35878 6278 35930
rect 6330 35878 6342 35930
rect 6394 35878 6406 35930
rect 6458 35878 7750 35930
rect 7802 35878 7814 35930
rect 7866 35878 7878 35930
rect 7930 35878 7942 35930
rect 7994 35878 8006 35930
rect 8058 35878 9350 35930
rect 9402 35878 9414 35930
rect 9466 35878 9478 35930
rect 9530 35878 9542 35930
rect 9594 35878 9606 35930
rect 9658 35878 9936 35930
rect 1104 35856 9936 35878
rect 2222 35776 2228 35828
rect 2280 35816 2286 35828
rect 7190 35816 7196 35828
rect 2280 35788 7196 35816
rect 2280 35776 2286 35788
rect 7190 35776 7196 35788
rect 7248 35776 7254 35828
rect 1118 35708 1124 35760
rect 1176 35748 1182 35760
rect 8294 35748 8300 35760
rect 1176 35720 8300 35748
rect 1176 35708 1182 35720
rect 8294 35708 8300 35720
rect 8352 35708 8358 35760
rect 4062 35640 4068 35692
rect 4120 35680 4126 35692
rect 4890 35680 4896 35692
rect 4120 35652 4896 35680
rect 4120 35640 4126 35652
rect 4890 35640 4896 35652
rect 4948 35640 4954 35692
rect 1104 35386 9936 35408
rect 1104 35334 3610 35386
rect 3662 35334 3674 35386
rect 3726 35334 3738 35386
rect 3790 35334 3802 35386
rect 3854 35334 3866 35386
rect 3918 35334 5210 35386
rect 5262 35334 5274 35386
rect 5326 35334 5338 35386
rect 5390 35334 5402 35386
rect 5454 35334 5466 35386
rect 5518 35334 6810 35386
rect 6862 35334 6874 35386
rect 6926 35334 6938 35386
rect 6990 35334 7002 35386
rect 7054 35334 7066 35386
rect 7118 35334 8410 35386
rect 8462 35334 8474 35386
rect 8526 35334 8538 35386
rect 8590 35334 8602 35386
rect 8654 35334 8666 35386
rect 8718 35334 9936 35386
rect 1104 35312 9936 35334
rect 842 35232 848 35284
rect 900 35272 906 35284
rect 1302 35272 1308 35284
rect 900 35244 1308 35272
rect 900 35232 906 35244
rect 1302 35232 1308 35244
rect 1360 35232 1366 35284
rect 2682 35096 2688 35148
rect 2740 35136 2746 35148
rect 3326 35136 3332 35148
rect 2740 35108 3332 35136
rect 2740 35096 2746 35108
rect 3326 35096 3332 35108
rect 3384 35096 3390 35148
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 992 35040 1409 35068
rect 992 35028 998 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 2866 34932 2872 34944
rect 1627 34904 2872 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 2866 34892 2872 34904
rect 2924 34892 2930 34944
rect 1104 34842 9936 34864
rect 1104 34790 2950 34842
rect 3002 34790 3014 34842
rect 3066 34790 3078 34842
rect 3130 34790 3142 34842
rect 3194 34790 3206 34842
rect 3258 34790 4550 34842
rect 4602 34790 4614 34842
rect 4666 34790 4678 34842
rect 4730 34790 4742 34842
rect 4794 34790 4806 34842
rect 4858 34790 6150 34842
rect 6202 34790 6214 34842
rect 6266 34790 6278 34842
rect 6330 34790 6342 34842
rect 6394 34790 6406 34842
rect 6458 34790 7750 34842
rect 7802 34790 7814 34842
rect 7866 34790 7878 34842
rect 7930 34790 7942 34842
rect 7994 34790 8006 34842
rect 8058 34790 9350 34842
rect 9402 34790 9414 34842
rect 9466 34790 9478 34842
rect 9530 34790 9542 34842
rect 9594 34790 9606 34842
rect 9658 34790 9936 34842
rect 1104 34768 9936 34790
rect 8103 34731 8161 34737
rect 8103 34697 8115 34731
rect 8149 34728 8161 34731
rect 10686 34728 10692 34740
rect 8149 34700 10692 34728
rect 8149 34697 8161 34700
rect 8103 34691 8161 34697
rect 10686 34688 10692 34700
rect 10744 34688 10750 34740
rect 1762 34620 1768 34672
rect 1820 34660 1826 34672
rect 8573 34663 8631 34669
rect 8573 34660 8585 34663
rect 1820 34632 8585 34660
rect 1820 34620 1826 34632
rect 8573 34629 8585 34632
rect 8619 34629 8631 34663
rect 8573 34623 8631 34629
rect 9030 34592 9036 34604
rect 8588 34564 9036 34592
rect 8588 34533 8616 34564
rect 9030 34552 9036 34564
rect 9088 34552 9094 34604
rect 8573 34527 8631 34533
rect 8573 34493 8585 34527
rect 8619 34493 8631 34527
rect 8573 34487 8631 34493
rect 8665 34527 8723 34533
rect 8665 34493 8677 34527
rect 8711 34524 8723 34527
rect 8846 34524 8852 34536
rect 8711 34496 8852 34524
rect 8711 34493 8723 34496
rect 8665 34487 8723 34493
rect 8846 34484 8852 34496
rect 8904 34484 8910 34536
rect 1104 34298 9936 34320
rect 1104 34246 3610 34298
rect 3662 34246 3674 34298
rect 3726 34246 3738 34298
rect 3790 34246 3802 34298
rect 3854 34246 3866 34298
rect 3918 34246 5210 34298
rect 5262 34246 5274 34298
rect 5326 34246 5338 34298
rect 5390 34246 5402 34298
rect 5454 34246 5466 34298
rect 5518 34246 6810 34298
rect 6862 34246 6874 34298
rect 6926 34246 6938 34298
rect 6990 34246 7002 34298
rect 7054 34246 7066 34298
rect 7118 34246 8410 34298
rect 8462 34246 8474 34298
rect 8526 34246 8538 34298
rect 8590 34246 8602 34298
rect 8654 34246 8666 34298
rect 8718 34246 9936 34298
rect 1104 34224 9936 34246
rect 3326 34144 3332 34196
rect 3384 34184 3390 34196
rect 3878 34184 3884 34196
rect 3384 34156 3884 34184
rect 3384 34144 3390 34156
rect 3878 34144 3884 34156
rect 3936 34144 3942 34196
rect 8113 34119 8171 34125
rect 8113 34085 8125 34119
rect 8159 34116 8171 34119
rect 11882 34116 11888 34128
rect 8159 34088 11888 34116
rect 8159 34085 8171 34088
rect 8113 34079 8171 34085
rect 11882 34076 11888 34088
rect 11940 34076 11946 34128
rect 8570 34008 8576 34060
rect 8628 34008 8634 34060
rect 934 33940 940 33992
rect 992 33980 998 33992
rect 1397 33983 1455 33989
rect 1397 33980 1409 33983
rect 992 33952 1409 33980
rect 992 33940 998 33952
rect 1397 33949 1409 33952
rect 1443 33949 1455 33983
rect 1397 33943 1455 33949
rect 7190 33872 7196 33924
rect 7248 33912 7254 33924
rect 8573 33915 8631 33921
rect 8573 33912 8585 33915
rect 7248 33884 8585 33912
rect 7248 33872 7254 33884
rect 8573 33881 8585 33884
rect 8619 33881 8631 33915
rect 8573 33875 8631 33881
rect 8662 33872 8668 33924
rect 8720 33912 8726 33924
rect 8846 33912 8852 33924
rect 8720 33884 8852 33912
rect 8720 33872 8726 33884
rect 8846 33872 8852 33884
rect 8904 33872 8910 33924
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 3326 33844 3332 33856
rect 1627 33816 3332 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 3326 33804 3332 33816
rect 3384 33804 3390 33856
rect 8478 33804 8484 33856
rect 8536 33844 8542 33856
rect 8938 33844 8944 33856
rect 8536 33816 8944 33844
rect 8536 33804 8542 33816
rect 8938 33804 8944 33816
rect 8996 33804 9002 33856
rect 1104 33754 9936 33776
rect 1104 33702 2950 33754
rect 3002 33702 3014 33754
rect 3066 33702 3078 33754
rect 3130 33702 3142 33754
rect 3194 33702 3206 33754
rect 3258 33702 4550 33754
rect 4602 33702 4614 33754
rect 4666 33702 4678 33754
rect 4730 33702 4742 33754
rect 4794 33702 4806 33754
rect 4858 33702 6150 33754
rect 6202 33702 6214 33754
rect 6266 33702 6278 33754
rect 6330 33702 6342 33754
rect 6394 33702 6406 33754
rect 6458 33702 7750 33754
rect 7802 33702 7814 33754
rect 7866 33702 7878 33754
rect 7930 33702 7942 33754
rect 7994 33702 8006 33754
rect 8058 33702 9350 33754
rect 9402 33702 9414 33754
rect 9466 33702 9478 33754
rect 9530 33702 9542 33754
rect 9594 33702 9606 33754
rect 9658 33702 9936 33754
rect 1104 33680 9936 33702
rect 3878 33600 3884 33652
rect 3936 33640 3942 33652
rect 8573 33643 8631 33649
rect 8573 33640 8585 33643
rect 3936 33612 8585 33640
rect 3936 33600 3942 33612
rect 8573 33609 8585 33612
rect 8619 33609 8631 33643
rect 8573 33603 8631 33609
rect 8662 33600 8668 33652
rect 8720 33640 8726 33652
rect 9306 33640 9312 33652
rect 8720 33612 9312 33640
rect 8720 33600 8726 33612
rect 9306 33600 9312 33612
rect 9364 33600 9370 33652
rect 8110 33532 8116 33584
rect 8168 33572 8174 33584
rect 8168 33544 8708 33572
rect 8168 33532 8174 33544
rect 1486 33464 1492 33516
rect 1544 33464 1550 33516
rect 8386 33464 8392 33516
rect 8444 33464 8450 33516
rect 8680 33513 8708 33544
rect 8665 33507 8723 33513
rect 8665 33473 8677 33507
rect 8711 33504 8723 33507
rect 8938 33504 8944 33516
rect 8711 33476 8944 33504
rect 8711 33473 8723 33476
rect 8665 33467 8723 33473
rect 8938 33464 8944 33476
rect 8996 33464 9002 33516
rect 7282 33396 7288 33448
rect 7340 33436 7346 33448
rect 8478 33436 8484 33448
rect 7340 33408 8484 33436
rect 7340 33396 7346 33408
rect 8478 33396 8484 33408
rect 8536 33396 8542 33448
rect 1118 33328 1124 33380
rect 1176 33368 1182 33380
rect 8113 33371 8171 33377
rect 8113 33368 8125 33371
rect 1176 33340 8125 33368
rect 1176 33328 1182 33340
rect 8113 33337 8125 33340
rect 8159 33337 8171 33371
rect 8113 33331 8171 33337
rect 1765 33303 1823 33309
rect 1765 33269 1777 33303
rect 1811 33300 1823 33303
rect 7466 33300 7472 33312
rect 1811 33272 7472 33300
rect 1811 33269 1823 33272
rect 1765 33263 1823 33269
rect 7466 33260 7472 33272
rect 7524 33260 7530 33312
rect 1104 33210 9936 33232
rect 1104 33158 3610 33210
rect 3662 33158 3674 33210
rect 3726 33158 3738 33210
rect 3790 33158 3802 33210
rect 3854 33158 3866 33210
rect 3918 33158 5210 33210
rect 5262 33158 5274 33210
rect 5326 33158 5338 33210
rect 5390 33158 5402 33210
rect 5454 33158 5466 33210
rect 5518 33158 6810 33210
rect 6862 33158 6874 33210
rect 6926 33158 6938 33210
rect 6990 33158 7002 33210
rect 7054 33158 7066 33210
rect 7118 33158 8410 33210
rect 8462 33158 8474 33210
rect 8526 33158 8538 33210
rect 8590 33158 8602 33210
rect 8654 33158 8666 33210
rect 8718 33158 9936 33210
rect 1104 33136 9936 33158
rect 6546 33056 6552 33108
rect 6604 33096 6610 33108
rect 7098 33096 7104 33108
rect 6604 33068 7104 33096
rect 6604 33056 6610 33068
rect 7098 33056 7104 33068
rect 7156 33056 7162 33108
rect 8662 33056 8668 33108
rect 8720 33096 8726 33108
rect 9306 33096 9312 33108
rect 8720 33068 9312 33096
rect 8720 33056 8726 33068
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 8021 33031 8079 33037
rect 8021 32997 8033 33031
rect 8067 33028 8079 33031
rect 10502 33028 10508 33040
rect 8067 33000 10508 33028
rect 8067 32997 8079 33000
rect 8021 32991 8079 32997
rect 10502 32988 10508 33000
rect 10560 32988 10566 33040
rect 8573 32963 8631 32969
rect 8573 32929 8585 32963
rect 8619 32960 8631 32963
rect 8938 32960 8944 32972
rect 8619 32932 8944 32960
rect 8619 32929 8631 32932
rect 8573 32923 8631 32929
rect 8938 32920 8944 32932
rect 8996 32920 9002 32972
rect 2130 32852 2136 32904
rect 2188 32892 2194 32904
rect 8110 32892 8116 32904
rect 2188 32864 8116 32892
rect 2188 32852 2194 32864
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 6638 32784 6644 32836
rect 6696 32824 6702 32836
rect 8297 32827 8355 32833
rect 8297 32824 8309 32827
rect 6696 32796 8309 32824
rect 6696 32784 6702 32796
rect 8297 32793 8309 32796
rect 8343 32793 8355 32827
rect 8297 32787 8355 32793
rect 9858 32784 9864 32836
rect 9916 32784 9922 32836
rect 8481 32759 8539 32765
rect 8481 32725 8493 32759
rect 8527 32756 8539 32759
rect 9876 32756 9904 32784
rect 8527 32728 9904 32756
rect 8527 32725 8539 32728
rect 8481 32719 8539 32725
rect 1104 32666 9936 32688
rect 1104 32614 2950 32666
rect 3002 32614 3014 32666
rect 3066 32614 3078 32666
rect 3130 32614 3142 32666
rect 3194 32614 3206 32666
rect 3258 32614 4550 32666
rect 4602 32614 4614 32666
rect 4666 32614 4678 32666
rect 4730 32614 4742 32666
rect 4794 32614 4806 32666
rect 4858 32614 6150 32666
rect 6202 32614 6214 32666
rect 6266 32614 6278 32666
rect 6330 32614 6342 32666
rect 6394 32614 6406 32666
rect 6458 32614 7750 32666
rect 7802 32614 7814 32666
rect 7866 32614 7878 32666
rect 7930 32614 7942 32666
rect 7994 32614 8006 32666
rect 8058 32614 9350 32666
rect 9402 32614 9414 32666
rect 9466 32614 9478 32666
rect 9530 32614 9542 32666
rect 9594 32614 9606 32666
rect 9658 32614 9936 32666
rect 1104 32592 9936 32614
rect 7193 32555 7251 32561
rect 7193 32521 7205 32555
rect 7239 32552 7251 32555
rect 8202 32552 8208 32564
rect 7239 32524 8208 32552
rect 7239 32521 7251 32524
rect 7193 32515 7251 32521
rect 8202 32512 8208 32524
rect 8260 32512 8266 32564
rect 8662 32512 8668 32564
rect 8720 32552 8726 32564
rect 9306 32552 9312 32564
rect 8720 32524 9312 32552
rect 8720 32512 8726 32524
rect 9306 32512 9312 32524
rect 9364 32512 9370 32564
rect 6457 32487 6515 32493
rect 6457 32453 6469 32487
rect 6503 32484 6515 32487
rect 6546 32484 6552 32496
rect 6503 32456 6552 32484
rect 6503 32453 6515 32456
rect 6457 32447 6515 32453
rect 6546 32444 6552 32456
rect 6604 32444 6610 32496
rect 8018 32484 8024 32496
rect 7208 32456 8024 32484
rect 7208 32428 7236 32456
rect 8018 32444 8024 32456
rect 8076 32444 8082 32496
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1489 32419 1547 32425
rect 1489 32416 1501 32419
rect 992 32388 1501 32416
rect 992 32376 998 32388
rect 1489 32385 1501 32388
rect 1535 32385 1547 32419
rect 1489 32379 1547 32385
rect 7190 32376 7196 32428
rect 7248 32376 7254 32428
rect 7285 32419 7343 32425
rect 7285 32385 7297 32419
rect 7331 32416 7343 32419
rect 7466 32416 7472 32428
rect 7331 32388 7472 32416
rect 7331 32385 7343 32388
rect 7285 32379 7343 32385
rect 7466 32376 7472 32388
rect 7524 32416 7530 32428
rect 7524 32388 10640 32416
rect 7524 32376 7530 32388
rect 10612 32360 10640 32388
rect 7377 32351 7435 32357
rect 7377 32317 7389 32351
rect 7423 32348 7435 32351
rect 7742 32348 7748 32360
rect 7423 32320 7748 32348
rect 7423 32317 7435 32320
rect 7377 32311 7435 32317
rect 7742 32308 7748 32320
rect 7800 32308 7806 32360
rect 8202 32308 8208 32360
rect 8260 32348 8266 32360
rect 8846 32348 8852 32360
rect 8260 32320 8852 32348
rect 8260 32308 8266 32320
rect 8846 32308 8852 32320
rect 8904 32308 8910 32360
rect 10594 32308 10600 32360
rect 10652 32308 10658 32360
rect 1762 32172 1768 32224
rect 1820 32172 1826 32224
rect 4890 32172 4896 32224
rect 4948 32212 4954 32224
rect 6549 32215 6607 32221
rect 6549 32212 6561 32215
rect 4948 32184 6561 32212
rect 4948 32172 4954 32184
rect 6549 32181 6561 32184
rect 6595 32181 6607 32215
rect 6549 32175 6607 32181
rect 6825 32215 6883 32221
rect 6825 32181 6837 32215
rect 6871 32212 6883 32215
rect 7282 32212 7288 32224
rect 6871 32184 7288 32212
rect 6871 32181 6883 32184
rect 6825 32175 6883 32181
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 7834 32172 7840 32224
rect 7892 32212 7898 32224
rect 10778 32212 10784 32224
rect 7892 32184 10784 32212
rect 7892 32172 7898 32184
rect 10778 32172 10784 32184
rect 10836 32172 10842 32224
rect 1104 32122 9936 32144
rect 1104 32070 3610 32122
rect 3662 32070 3674 32122
rect 3726 32070 3738 32122
rect 3790 32070 3802 32122
rect 3854 32070 3866 32122
rect 3918 32070 5210 32122
rect 5262 32070 5274 32122
rect 5326 32070 5338 32122
rect 5390 32070 5402 32122
rect 5454 32070 5466 32122
rect 5518 32070 6810 32122
rect 6862 32070 6874 32122
rect 6926 32070 6938 32122
rect 6990 32070 7002 32122
rect 7054 32070 7066 32122
rect 7118 32070 8410 32122
rect 8462 32070 8474 32122
rect 8526 32070 8538 32122
rect 8590 32070 8602 32122
rect 8654 32070 8666 32122
rect 8718 32070 9936 32122
rect 1104 32048 9936 32070
rect 1026 31968 1032 32020
rect 1084 32008 1090 32020
rect 8021 32011 8079 32017
rect 8021 32008 8033 32011
rect 1084 31980 8033 32008
rect 1084 31968 1090 31980
rect 8021 31977 8033 31980
rect 8067 31977 8079 32011
rect 8021 31971 8079 31977
rect 8110 31968 8116 32020
rect 8168 32008 8174 32020
rect 8168 31980 9168 32008
rect 8168 31968 8174 31980
rect 5442 31900 5448 31952
rect 5500 31940 5506 31952
rect 5902 31940 5908 31952
rect 5500 31912 5908 31940
rect 5500 31900 5506 31912
rect 5902 31900 5908 31912
rect 5960 31900 5966 31952
rect 7009 31943 7067 31949
rect 7009 31909 7021 31943
rect 7055 31940 7067 31943
rect 7466 31940 7472 31952
rect 7055 31912 7472 31940
rect 7055 31909 7067 31912
rect 7009 31903 7067 31909
rect 7466 31900 7472 31912
rect 7524 31900 7530 31952
rect 7650 31900 7656 31952
rect 7708 31940 7714 31952
rect 9140 31940 9168 31980
rect 9214 31968 9220 32020
rect 9272 32008 9278 32020
rect 10134 32008 10140 32020
rect 9272 31980 10140 32008
rect 9272 31968 9278 31980
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 9582 31940 9588 31952
rect 7708 31912 8984 31940
rect 9140 31912 9588 31940
rect 7708 31900 7714 31912
rect 1762 31832 1768 31884
rect 1820 31832 1826 31884
rect 7561 31875 7619 31881
rect 7561 31841 7573 31875
rect 7607 31872 7619 31875
rect 7742 31872 7748 31884
rect 7607 31844 7748 31872
rect 7607 31841 7619 31844
rect 7561 31835 7619 31841
rect 7742 31832 7748 31844
rect 7800 31832 7806 31884
rect 8110 31832 8116 31884
rect 8168 31832 8174 31884
rect 1780 31804 1808 31832
rect 7190 31804 7196 31816
rect 1780 31776 7196 31804
rect 7190 31764 7196 31776
rect 7248 31804 7254 31816
rect 7469 31807 7527 31813
rect 7469 31804 7481 31807
rect 7248 31776 7481 31804
rect 7248 31764 7254 31776
rect 7469 31773 7481 31776
rect 7515 31804 7527 31807
rect 7834 31804 7840 31816
rect 7515 31776 7840 31804
rect 7515 31773 7527 31776
rect 7469 31767 7527 31773
rect 7834 31764 7840 31776
rect 7892 31764 7898 31816
rect 8128 31804 8156 31832
rect 8297 31807 8355 31813
rect 8297 31804 8309 31807
rect 8128 31776 8309 31804
rect 8297 31773 8309 31776
rect 8343 31773 8355 31807
rect 8297 31767 8355 31773
rect 8573 31807 8631 31813
rect 8573 31773 8585 31807
rect 8619 31804 8631 31807
rect 8956 31804 8984 31912
rect 9582 31900 9588 31912
rect 9640 31900 9646 31952
rect 8619 31776 8984 31804
rect 8619 31773 8631 31776
rect 8573 31767 8631 31773
rect 7377 31739 7435 31745
rect 7377 31705 7389 31739
rect 7423 31736 7435 31739
rect 8202 31736 8208 31748
rect 7423 31708 8208 31736
rect 7423 31705 7435 31708
rect 7377 31699 7435 31705
rect 8202 31696 8208 31708
rect 8260 31696 8266 31748
rect 8481 31739 8539 31745
rect 8481 31705 8493 31739
rect 8527 31736 8539 31739
rect 10042 31736 10048 31748
rect 8527 31708 10048 31736
rect 8527 31705 8539 31708
rect 8481 31699 8539 31705
rect 10042 31696 10048 31708
rect 10100 31696 10106 31748
rect 7558 31628 7564 31680
rect 7616 31668 7622 31680
rect 7742 31668 7748 31680
rect 7616 31640 7748 31668
rect 7616 31628 7622 31640
rect 7742 31628 7748 31640
rect 7800 31628 7806 31680
rect 1104 31578 9936 31600
rect 1104 31526 2950 31578
rect 3002 31526 3014 31578
rect 3066 31526 3078 31578
rect 3130 31526 3142 31578
rect 3194 31526 3206 31578
rect 3258 31526 4550 31578
rect 4602 31526 4614 31578
rect 4666 31526 4678 31578
rect 4730 31526 4742 31578
rect 4794 31526 4806 31578
rect 4858 31526 6150 31578
rect 6202 31526 6214 31578
rect 6266 31526 6278 31578
rect 6330 31526 6342 31578
rect 6394 31526 6406 31578
rect 6458 31526 7750 31578
rect 7802 31526 7814 31578
rect 7866 31526 7878 31578
rect 7930 31526 7942 31578
rect 7994 31526 8006 31578
rect 8058 31526 9350 31578
rect 9402 31526 9414 31578
rect 9466 31526 9478 31578
rect 9530 31526 9542 31578
rect 9594 31526 9606 31578
rect 9658 31526 9936 31578
rect 1104 31504 9936 31526
rect 7374 31424 7380 31476
rect 7432 31464 7438 31476
rect 8110 31464 8116 31476
rect 7432 31436 8116 31464
rect 7432 31424 7438 31436
rect 8110 31424 8116 31436
rect 8168 31424 8174 31476
rect 5902 31356 5908 31408
rect 5960 31396 5966 31408
rect 7006 31396 7012 31408
rect 5960 31368 7012 31396
rect 5960 31356 5966 31368
rect 7006 31356 7012 31368
rect 7064 31356 7070 31408
rect 934 31288 940 31340
rect 992 31328 998 31340
rect 1581 31331 1639 31337
rect 1581 31328 1593 31331
rect 992 31300 1593 31328
rect 992 31288 998 31300
rect 1581 31297 1593 31300
rect 1627 31297 1639 31331
rect 1581 31291 1639 31297
rect 5442 31288 5448 31340
rect 5500 31328 5506 31340
rect 6086 31328 6092 31340
rect 5500 31300 6092 31328
rect 5500 31288 5506 31300
rect 6086 31288 6092 31300
rect 6144 31288 6150 31340
rect 7558 31288 7564 31340
rect 7616 31288 7622 31340
rect 7576 31260 7604 31288
rect 7392 31232 7604 31260
rect 7392 31204 7420 31232
rect 1578 31152 1584 31204
rect 1636 31192 1642 31204
rect 2682 31192 2688 31204
rect 1636 31164 2688 31192
rect 1636 31152 1642 31164
rect 2682 31152 2688 31164
rect 2740 31152 2746 31204
rect 7374 31152 7380 31204
rect 7432 31152 7438 31204
rect 1397 31127 1455 31133
rect 1397 31093 1409 31127
rect 1443 31124 1455 31127
rect 7466 31124 7472 31136
rect 1443 31096 7472 31124
rect 1443 31093 1455 31096
rect 1397 31087 1455 31093
rect 7466 31084 7472 31096
rect 7524 31084 7530 31136
rect 1104 31034 9936 31056
rect 1104 30982 3610 31034
rect 3662 30982 3674 31034
rect 3726 30982 3738 31034
rect 3790 30982 3802 31034
rect 3854 30982 3866 31034
rect 3918 30982 5210 31034
rect 5262 30982 5274 31034
rect 5326 30982 5338 31034
rect 5390 30982 5402 31034
rect 5454 30982 5466 31034
rect 5518 30982 6810 31034
rect 6862 30982 6874 31034
rect 6926 30982 6938 31034
rect 6990 30982 7002 31034
rect 7054 30982 7066 31034
rect 7118 30982 8410 31034
rect 8462 30982 8474 31034
rect 8526 30982 8538 31034
rect 8590 30982 8602 31034
rect 8654 30982 8666 31034
rect 8718 30982 9936 31034
rect 1104 30960 9936 30982
rect 1104 30490 9936 30512
rect 1104 30438 2950 30490
rect 3002 30438 3014 30490
rect 3066 30438 3078 30490
rect 3130 30438 3142 30490
rect 3194 30438 3206 30490
rect 3258 30438 4550 30490
rect 4602 30438 4614 30490
rect 4666 30438 4678 30490
rect 4730 30438 4742 30490
rect 4794 30438 4806 30490
rect 4858 30438 6150 30490
rect 6202 30438 6214 30490
rect 6266 30438 6278 30490
rect 6330 30438 6342 30490
rect 6394 30438 6406 30490
rect 6458 30438 7750 30490
rect 7802 30438 7814 30490
rect 7866 30438 7878 30490
rect 7930 30438 7942 30490
rect 7994 30438 8006 30490
rect 8058 30438 9350 30490
rect 9402 30438 9414 30490
rect 9466 30438 9478 30490
rect 9530 30438 9542 30490
rect 9594 30438 9606 30490
rect 9658 30438 9936 30490
rect 1104 30416 9936 30438
rect 4154 30268 4160 30320
rect 4212 30308 4218 30320
rect 4798 30308 4804 30320
rect 4212 30280 4804 30308
rect 4212 30268 4218 30280
rect 4798 30268 4804 30280
rect 4856 30268 4862 30320
rect 7653 30311 7711 30317
rect 7653 30277 7665 30311
rect 7699 30308 7711 30311
rect 9214 30308 9220 30320
rect 7699 30280 9220 30308
rect 7699 30277 7711 30280
rect 7653 30271 7711 30277
rect 9214 30268 9220 30280
rect 9272 30268 9278 30320
rect 934 30200 940 30252
rect 992 30240 998 30252
rect 1581 30243 1639 30249
rect 1581 30240 1593 30243
rect 992 30212 1593 30240
rect 992 30200 998 30212
rect 1581 30209 1593 30212
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 7282 30200 7288 30252
rect 7340 30240 7346 30252
rect 7469 30243 7527 30249
rect 7469 30240 7481 30243
rect 7340 30212 7481 30240
rect 7340 30200 7346 30212
rect 7469 30209 7481 30212
rect 7515 30209 7527 30243
rect 7469 30203 7527 30209
rect 4154 30132 4160 30184
rect 4212 30172 4218 30184
rect 4982 30172 4988 30184
rect 4212 30144 4988 30172
rect 4212 30132 4218 30144
rect 4982 30132 4988 30144
rect 5040 30132 5046 30184
rect 1397 30039 1455 30045
rect 1397 30005 1409 30039
rect 1443 30036 1455 30039
rect 4982 30036 4988 30048
rect 1443 30008 4988 30036
rect 1443 30005 1455 30008
rect 1397 29999 1455 30005
rect 4982 29996 4988 30008
rect 5040 29996 5046 30048
rect 1104 29946 9936 29968
rect 1104 29894 3610 29946
rect 3662 29894 3674 29946
rect 3726 29894 3738 29946
rect 3790 29894 3802 29946
rect 3854 29894 3866 29946
rect 3918 29894 5210 29946
rect 5262 29894 5274 29946
rect 5326 29894 5338 29946
rect 5390 29894 5402 29946
rect 5454 29894 5466 29946
rect 5518 29894 6810 29946
rect 6862 29894 6874 29946
rect 6926 29894 6938 29946
rect 6990 29894 7002 29946
rect 7054 29894 7066 29946
rect 7118 29894 8410 29946
rect 8462 29894 8474 29946
rect 8526 29894 8538 29946
rect 8590 29894 8602 29946
rect 8654 29894 8666 29946
rect 8718 29894 9936 29946
rect 1104 29872 9936 29894
rect 5626 29656 5632 29708
rect 5684 29656 5690 29708
rect 5718 29656 5724 29708
rect 5776 29696 5782 29708
rect 6822 29696 6828 29708
rect 5776 29668 6828 29696
rect 5776 29656 5782 29668
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 934 29588 940 29640
rect 992 29628 998 29640
rect 1581 29631 1639 29637
rect 1581 29628 1593 29631
rect 992 29600 1593 29628
rect 992 29588 998 29600
rect 1581 29597 1593 29600
rect 1627 29597 1639 29631
rect 1581 29591 1639 29597
rect 4798 29520 4804 29572
rect 4856 29560 4862 29572
rect 5166 29560 5172 29572
rect 4856 29532 5172 29560
rect 4856 29520 4862 29532
rect 5166 29520 5172 29532
rect 5224 29520 5230 29572
rect 5644 29504 5672 29656
rect 1397 29495 1455 29501
rect 1397 29461 1409 29495
rect 1443 29492 1455 29495
rect 5534 29492 5540 29504
rect 1443 29464 5540 29492
rect 1443 29461 1455 29464
rect 1397 29455 1455 29461
rect 5534 29452 5540 29464
rect 5592 29452 5598 29504
rect 5626 29452 5632 29504
rect 5684 29452 5690 29504
rect 1104 29402 9936 29424
rect 1104 29350 2950 29402
rect 3002 29350 3014 29402
rect 3066 29350 3078 29402
rect 3130 29350 3142 29402
rect 3194 29350 3206 29402
rect 3258 29350 4550 29402
rect 4602 29350 4614 29402
rect 4666 29350 4678 29402
rect 4730 29350 4742 29402
rect 4794 29350 4806 29402
rect 4858 29350 6150 29402
rect 6202 29350 6214 29402
rect 6266 29350 6278 29402
rect 6330 29350 6342 29402
rect 6394 29350 6406 29402
rect 6458 29350 7750 29402
rect 7802 29350 7814 29402
rect 7866 29350 7878 29402
rect 7930 29350 7942 29402
rect 7994 29350 8006 29402
rect 8058 29350 9350 29402
rect 9402 29350 9414 29402
rect 9466 29350 9478 29402
rect 9530 29350 9542 29402
rect 9594 29350 9606 29402
rect 9658 29350 9936 29402
rect 1104 29328 9936 29350
rect 6730 29248 6736 29300
rect 6788 29288 6794 29300
rect 8757 29291 8815 29297
rect 8757 29288 8769 29291
rect 6788 29260 8769 29288
rect 6788 29248 6794 29260
rect 8757 29257 8769 29260
rect 8803 29257 8815 29291
rect 8757 29251 8815 29257
rect 7469 29223 7527 29229
rect 7469 29189 7481 29223
rect 7515 29220 7527 29223
rect 8846 29220 8852 29232
rect 7515 29192 8852 29220
rect 7515 29189 7527 29192
rect 7469 29183 7527 29189
rect 8846 29180 8852 29192
rect 8904 29180 8910 29232
rect 8938 29180 8944 29232
rect 8996 29220 9002 29232
rect 9858 29220 9864 29232
rect 8996 29192 9864 29220
rect 8996 29180 9002 29192
rect 9858 29180 9864 29192
rect 9916 29180 9922 29232
rect 7282 29112 7288 29164
rect 7340 29112 7346 29164
rect 11882 29152 11888 29164
rect 8312 29124 11888 29152
rect 8312 29025 8340 29124
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 8757 29087 8815 29093
rect 8757 29053 8769 29087
rect 8803 29053 8815 29087
rect 8757 29047 8815 29053
rect 8297 29019 8355 29025
rect 8297 28985 8309 29019
rect 8343 28985 8355 29019
rect 8772 29016 8800 29047
rect 8772 28988 9076 29016
rect 8297 28979 8355 28985
rect 9048 28960 9076 28988
rect 4798 28908 4804 28960
rect 4856 28948 4862 28960
rect 5166 28948 5172 28960
rect 4856 28920 5172 28948
rect 4856 28908 4862 28920
rect 5166 28908 5172 28920
rect 5224 28908 5230 28960
rect 6822 28908 6828 28960
rect 6880 28948 6886 28960
rect 7834 28948 7840 28960
rect 6880 28920 7840 28948
rect 6880 28908 6886 28920
rect 7834 28908 7840 28920
rect 7892 28908 7898 28960
rect 9030 28908 9036 28960
rect 9088 28908 9094 28960
rect 1104 28858 9936 28880
rect 1104 28806 3610 28858
rect 3662 28806 3674 28858
rect 3726 28806 3738 28858
rect 3790 28806 3802 28858
rect 3854 28806 3866 28858
rect 3918 28806 5210 28858
rect 5262 28806 5274 28858
rect 5326 28806 5338 28858
rect 5390 28806 5402 28858
rect 5454 28806 5466 28858
rect 5518 28806 6810 28858
rect 6862 28806 6874 28858
rect 6926 28806 6938 28858
rect 6990 28806 7002 28858
rect 7054 28806 7066 28858
rect 7118 28806 8410 28858
rect 8462 28806 8474 28858
rect 8526 28806 8538 28858
rect 8590 28806 8602 28858
rect 8654 28806 8666 28858
rect 8718 28806 9936 28858
rect 1104 28784 9936 28806
rect 6086 28704 6092 28756
rect 6144 28744 6150 28756
rect 7006 28744 7012 28756
rect 6144 28716 7012 28744
rect 6144 28704 6150 28716
rect 7006 28704 7012 28716
rect 7064 28704 7070 28756
rect 7101 28747 7159 28753
rect 7101 28713 7113 28747
rect 7147 28744 7159 28747
rect 9214 28744 9220 28756
rect 7147 28716 9220 28744
rect 7147 28713 7159 28716
rect 7101 28707 7159 28713
rect 9214 28704 9220 28716
rect 9272 28704 9278 28756
rect 7190 28636 7196 28688
rect 7248 28676 7254 28688
rect 7248 28648 7788 28676
rect 7248 28636 7254 28648
rect 7650 28568 7656 28620
rect 7708 28568 7714 28620
rect 934 28500 940 28552
rect 992 28540 998 28552
rect 1581 28543 1639 28549
rect 1581 28540 1593 28543
rect 992 28512 1593 28540
rect 992 28500 998 28512
rect 1581 28509 1593 28512
rect 1627 28509 1639 28543
rect 1581 28503 1639 28509
rect 6086 28500 6092 28552
rect 6144 28540 6150 28552
rect 6822 28540 6828 28552
rect 6144 28512 6828 28540
rect 6144 28500 6150 28512
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 7466 28500 7472 28552
rect 7524 28500 7530 28552
rect 7760 28540 7788 28648
rect 7834 28636 7840 28688
rect 7892 28636 7898 28688
rect 8113 28679 8171 28685
rect 8113 28645 8125 28679
rect 8159 28676 8171 28679
rect 10318 28676 10324 28688
rect 8159 28648 10324 28676
rect 8159 28645 8171 28648
rect 8113 28639 8171 28645
rect 10318 28636 10324 28648
rect 10376 28636 10382 28688
rect 7852 28608 7880 28636
rect 7852 28580 8064 28608
rect 7760 28512 7972 28540
rect 1394 28364 1400 28416
rect 1452 28364 1458 28416
rect 4798 28364 4804 28416
rect 4856 28404 4862 28416
rect 5442 28404 5448 28416
rect 4856 28376 5448 28404
rect 4856 28364 4862 28376
rect 5442 28364 5448 28376
rect 5500 28364 5506 28416
rect 5810 28364 5816 28416
rect 5868 28404 5874 28416
rect 5994 28404 6000 28416
rect 5868 28376 6000 28404
rect 5868 28364 5874 28376
rect 5994 28364 6000 28376
rect 6052 28364 6058 28416
rect 7190 28364 7196 28416
rect 7248 28404 7254 28416
rect 7561 28407 7619 28413
rect 7561 28404 7573 28407
rect 7248 28376 7573 28404
rect 7248 28364 7254 28376
rect 7561 28373 7573 28376
rect 7607 28404 7619 28407
rect 7742 28404 7748 28416
rect 7607 28376 7748 28404
rect 7607 28373 7619 28376
rect 7561 28367 7619 28373
rect 7742 28364 7748 28376
rect 7800 28364 7806 28416
rect 7944 28404 7972 28512
rect 8036 28472 8064 28580
rect 8202 28568 8208 28620
rect 8260 28608 8266 28620
rect 8478 28608 8484 28620
rect 8260 28580 8484 28608
rect 8260 28568 8266 28580
rect 8478 28568 8484 28580
rect 8536 28568 8542 28620
rect 8573 28611 8631 28617
rect 8573 28577 8585 28611
rect 8619 28608 8631 28611
rect 8846 28608 8852 28620
rect 8619 28580 8852 28608
rect 8619 28577 8631 28580
rect 8573 28571 8631 28577
rect 8846 28568 8852 28580
rect 8904 28568 8910 28620
rect 8665 28543 8723 28549
rect 8665 28509 8677 28543
rect 8711 28540 8723 28543
rect 8754 28540 8760 28552
rect 8711 28512 8760 28540
rect 8711 28509 8723 28512
rect 8665 28503 8723 28509
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 8573 28475 8631 28481
rect 8573 28472 8585 28475
rect 8036 28444 8585 28472
rect 8573 28441 8585 28444
rect 8619 28441 8631 28475
rect 8573 28435 8631 28441
rect 8110 28404 8116 28416
rect 7944 28376 8116 28404
rect 8110 28364 8116 28376
rect 8168 28364 8174 28416
rect 1104 28314 9936 28336
rect 1104 28262 2950 28314
rect 3002 28262 3014 28314
rect 3066 28262 3078 28314
rect 3130 28262 3142 28314
rect 3194 28262 3206 28314
rect 3258 28262 4550 28314
rect 4602 28262 4614 28314
rect 4666 28262 4678 28314
rect 4730 28262 4742 28314
rect 4794 28262 4806 28314
rect 4858 28262 6150 28314
rect 6202 28262 6214 28314
rect 6266 28262 6278 28314
rect 6330 28262 6342 28314
rect 6394 28262 6406 28314
rect 6458 28262 7750 28314
rect 7802 28262 7814 28314
rect 7866 28262 7878 28314
rect 7930 28262 7942 28314
rect 7994 28262 8006 28314
rect 8058 28262 9350 28314
rect 9402 28262 9414 28314
rect 9466 28262 9478 28314
rect 9530 28262 9542 28314
rect 9594 28262 9606 28314
rect 9658 28262 9936 28314
rect 1104 28240 9936 28262
rect 1394 28160 1400 28212
rect 1452 28200 1458 28212
rect 5810 28200 5816 28212
rect 1452 28172 5816 28200
rect 1452 28160 1458 28172
rect 5810 28160 5816 28172
rect 5868 28160 5874 28212
rect 2590 27820 2596 27872
rect 2648 27860 2654 27872
rect 3326 27860 3332 27872
rect 2648 27832 3332 27860
rect 2648 27820 2654 27832
rect 3326 27820 3332 27832
rect 3384 27820 3390 27872
rect 1104 27770 9936 27792
rect 1104 27718 3610 27770
rect 3662 27718 3674 27770
rect 3726 27718 3738 27770
rect 3790 27718 3802 27770
rect 3854 27718 3866 27770
rect 3918 27718 5210 27770
rect 5262 27718 5274 27770
rect 5326 27718 5338 27770
rect 5390 27718 5402 27770
rect 5454 27718 5466 27770
rect 5518 27718 6810 27770
rect 6862 27718 6874 27770
rect 6926 27718 6938 27770
rect 6990 27718 7002 27770
rect 7054 27718 7066 27770
rect 7118 27718 8410 27770
rect 8462 27718 8474 27770
rect 8526 27718 8538 27770
rect 8590 27718 8602 27770
rect 8654 27718 8666 27770
rect 8718 27718 9936 27770
rect 1104 27696 9936 27718
rect 3326 27616 3332 27668
rect 3384 27656 3390 27668
rect 4154 27656 4160 27668
rect 3384 27628 4160 27656
rect 3384 27616 3390 27628
rect 4154 27616 4160 27628
rect 4212 27616 4218 27668
rect 7377 27659 7435 27665
rect 7377 27625 7389 27659
rect 7423 27656 7435 27659
rect 7650 27656 7656 27668
rect 7423 27628 7656 27656
rect 7423 27625 7435 27628
rect 7377 27619 7435 27625
rect 7650 27616 7656 27628
rect 7708 27616 7714 27668
rect 934 27412 940 27464
rect 992 27452 998 27464
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 992 27424 1409 27452
rect 992 27412 998 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 1670 27344 1676 27396
rect 1728 27344 1734 27396
rect 6914 27344 6920 27396
rect 6972 27384 6978 27396
rect 7285 27387 7343 27393
rect 7285 27384 7297 27387
rect 6972 27356 7297 27384
rect 6972 27344 6978 27356
rect 7285 27353 7297 27356
rect 7331 27384 7343 27387
rect 7374 27384 7380 27396
rect 7331 27356 7380 27384
rect 7331 27353 7343 27356
rect 7285 27347 7343 27353
rect 7374 27344 7380 27356
rect 7432 27344 7438 27396
rect 1104 27226 9936 27248
rect 1104 27174 2950 27226
rect 3002 27174 3014 27226
rect 3066 27174 3078 27226
rect 3130 27174 3142 27226
rect 3194 27174 3206 27226
rect 3258 27174 4550 27226
rect 4602 27174 4614 27226
rect 4666 27174 4678 27226
rect 4730 27174 4742 27226
rect 4794 27174 4806 27226
rect 4858 27174 6150 27226
rect 6202 27174 6214 27226
rect 6266 27174 6278 27226
rect 6330 27174 6342 27226
rect 6394 27174 6406 27226
rect 6458 27174 7750 27226
rect 7802 27174 7814 27226
rect 7866 27174 7878 27226
rect 7930 27174 7942 27226
rect 7994 27174 8006 27226
rect 8058 27174 9350 27226
rect 9402 27174 9414 27226
rect 9466 27174 9478 27226
rect 9530 27174 9542 27226
rect 9594 27174 9606 27226
rect 9658 27174 9936 27226
rect 1104 27152 9936 27174
rect 5534 27072 5540 27124
rect 5592 27112 5598 27124
rect 7653 27115 7711 27121
rect 7653 27112 7665 27115
rect 5592 27084 7665 27112
rect 5592 27072 5598 27084
rect 7653 27081 7665 27084
rect 7699 27081 7711 27115
rect 7653 27075 7711 27081
rect 7745 27115 7803 27121
rect 7745 27081 7757 27115
rect 7791 27112 7803 27115
rect 8202 27112 8208 27124
rect 7791 27084 8208 27112
rect 7791 27081 7803 27084
rect 7745 27075 7803 27081
rect 7009 27047 7067 27053
rect 7009 27013 7021 27047
rect 7055 27044 7067 27047
rect 7760 27044 7788 27075
rect 8202 27072 8208 27084
rect 8260 27112 8266 27124
rect 11606 27112 11612 27124
rect 8260 27084 11612 27112
rect 8260 27072 8266 27084
rect 11606 27072 11612 27084
rect 11664 27072 11670 27124
rect 7055 27016 7788 27044
rect 7055 27013 7067 27016
rect 7009 27007 7067 27013
rect 6454 26936 6460 26988
rect 6512 26976 6518 26988
rect 7098 26976 7104 26988
rect 6512 26948 7104 26976
rect 6512 26936 6518 26948
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 7668 26948 7880 26976
rect 7668 26920 7696 26948
rect 6086 26868 6092 26920
rect 6144 26908 6150 26920
rect 6914 26908 6920 26920
rect 6144 26880 6920 26908
rect 6144 26868 6150 26880
rect 6914 26868 6920 26880
rect 6972 26868 6978 26920
rect 7650 26868 7656 26920
rect 7708 26868 7714 26920
rect 7852 26917 7880 26948
rect 7837 26911 7895 26917
rect 7837 26877 7849 26911
rect 7883 26877 7895 26911
rect 7837 26871 7895 26877
rect 750 26800 756 26852
rect 808 26840 814 26852
rect 9490 26840 9496 26852
rect 808 26812 9496 26840
rect 808 26800 814 26812
rect 9490 26800 9496 26812
rect 9548 26800 9554 26852
rect 6638 26732 6644 26784
rect 6696 26772 6702 26784
rect 6822 26772 6828 26784
rect 6696 26744 6828 26772
rect 6696 26732 6702 26744
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7285 26775 7343 26781
rect 7285 26741 7297 26775
rect 7331 26772 7343 26775
rect 8202 26772 8208 26784
rect 7331 26744 8208 26772
rect 7331 26741 7343 26744
rect 7285 26735 7343 26741
rect 8202 26732 8208 26744
rect 8260 26732 8266 26784
rect 8938 26732 8944 26784
rect 8996 26772 9002 26784
rect 10042 26772 10048 26784
rect 8996 26744 10048 26772
rect 8996 26732 9002 26744
rect 10042 26732 10048 26744
rect 10100 26732 10106 26784
rect 1104 26682 9936 26704
rect 1104 26630 3610 26682
rect 3662 26630 3674 26682
rect 3726 26630 3738 26682
rect 3790 26630 3802 26682
rect 3854 26630 3866 26682
rect 3918 26630 5210 26682
rect 5262 26630 5274 26682
rect 5326 26630 5338 26682
rect 5390 26630 5402 26682
rect 5454 26630 5466 26682
rect 5518 26630 6810 26682
rect 6862 26630 6874 26682
rect 6926 26630 6938 26682
rect 6990 26630 7002 26682
rect 7054 26630 7066 26682
rect 7118 26630 8410 26682
rect 8462 26630 8474 26682
rect 8526 26630 8538 26682
rect 8590 26630 8602 26682
rect 8654 26630 8666 26682
rect 8718 26630 9936 26682
rect 1104 26608 9936 26630
rect 6549 26571 6607 26577
rect 6549 26537 6561 26571
rect 6595 26568 6607 26571
rect 7374 26568 7380 26580
rect 6595 26540 7380 26568
rect 6595 26537 6607 26540
rect 6549 26531 6607 26537
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 7558 26528 7564 26580
rect 7616 26568 7622 26580
rect 7616 26540 9260 26568
rect 7616 26528 7622 26540
rect 5350 26460 5356 26512
rect 5408 26500 5414 26512
rect 6454 26500 6460 26512
rect 5408 26472 6460 26500
rect 5408 26460 5414 26472
rect 6454 26460 6460 26472
rect 6512 26460 6518 26512
rect 7285 26503 7343 26509
rect 7285 26469 7297 26503
rect 7331 26500 7343 26503
rect 8938 26500 8944 26512
rect 7331 26472 8944 26500
rect 7331 26469 7343 26472
rect 7285 26463 7343 26469
rect 8938 26460 8944 26472
rect 8996 26460 9002 26512
rect 2746 26404 5580 26432
rect 934 26324 940 26376
rect 992 26364 998 26376
rect 1397 26367 1455 26373
rect 1397 26364 1409 26367
rect 992 26336 1409 26364
rect 992 26324 998 26336
rect 1397 26333 1409 26336
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 1673 26299 1731 26305
rect 1673 26265 1685 26299
rect 1719 26296 1731 26299
rect 2746 26296 2774 26404
rect 5552 26376 5580 26404
rect 7098 26392 7104 26444
rect 7156 26432 7162 26444
rect 7466 26432 7472 26444
rect 7156 26404 7472 26432
rect 7156 26392 7162 26404
rect 7466 26392 7472 26404
rect 7524 26392 7530 26444
rect 7650 26392 7656 26444
rect 7708 26432 7714 26444
rect 7837 26435 7895 26441
rect 7837 26432 7849 26435
rect 7708 26404 7849 26432
rect 7708 26392 7714 26404
rect 7837 26401 7849 26404
rect 7883 26401 7895 26435
rect 7837 26395 7895 26401
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 6546 26324 6552 26376
rect 6604 26364 6610 26376
rect 6825 26367 6883 26373
rect 6825 26364 6837 26367
rect 6604 26336 6837 26364
rect 6604 26324 6610 26336
rect 6825 26333 6837 26336
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 6914 26324 6920 26376
rect 6972 26324 6978 26376
rect 7006 26324 7012 26376
rect 7064 26324 7070 26376
rect 7190 26324 7196 26376
rect 7248 26324 7254 26376
rect 9232 26373 9260 26540
rect 9490 26528 9496 26580
rect 9548 26568 9554 26580
rect 10134 26568 10140 26580
rect 9548 26540 10140 26568
rect 9548 26528 9554 26540
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9217 26327 9275 26333
rect 5000 26296 5028 26324
rect 7653 26299 7711 26305
rect 7653 26296 7665 26299
rect 1719 26268 2774 26296
rect 4080 26268 4292 26296
rect 5000 26268 7665 26296
rect 1719 26265 1731 26268
rect 1673 26259 1731 26265
rect 2866 26188 2872 26240
rect 2924 26228 2930 26240
rect 4080 26228 4108 26268
rect 2924 26200 4108 26228
rect 2924 26188 2930 26200
rect 4154 26188 4160 26240
rect 4212 26188 4218 26240
rect 4264 26228 4292 26268
rect 7653 26265 7665 26268
rect 7699 26265 7711 26299
rect 7653 26259 7711 26265
rect 7745 26299 7803 26305
rect 7745 26265 7757 26299
rect 7791 26296 7803 26299
rect 9582 26296 9588 26308
rect 7791 26268 9588 26296
rect 7791 26265 7803 26268
rect 7745 26259 7803 26265
rect 9582 26256 9588 26268
rect 9640 26296 9646 26308
rect 10410 26296 10416 26308
rect 9640 26268 10416 26296
rect 9640 26256 9646 26268
rect 10410 26256 10416 26268
rect 10468 26256 10474 26308
rect 8386 26228 8392 26240
rect 4264 26200 8392 26228
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 1104 26138 9936 26160
rect 1104 26086 2950 26138
rect 3002 26086 3014 26138
rect 3066 26086 3078 26138
rect 3130 26086 3142 26138
rect 3194 26086 3206 26138
rect 3258 26086 4550 26138
rect 4602 26086 4614 26138
rect 4666 26086 4678 26138
rect 4730 26086 4742 26138
rect 4794 26086 4806 26138
rect 4858 26086 6150 26138
rect 6202 26086 6214 26138
rect 6266 26086 6278 26138
rect 6330 26086 6342 26138
rect 6394 26086 6406 26138
rect 6458 26086 7750 26138
rect 7802 26086 7814 26138
rect 7866 26086 7878 26138
rect 7930 26086 7942 26138
rect 7994 26086 8006 26138
rect 8058 26086 9350 26138
rect 9402 26086 9414 26138
rect 9466 26086 9478 26138
rect 9530 26086 9542 26138
rect 9594 26086 9606 26138
rect 9658 26086 9936 26138
rect 1104 26064 9936 26086
rect 1578 25984 1584 26036
rect 1636 25984 1642 26036
rect 4982 25984 4988 26036
rect 5040 26024 5046 26036
rect 5350 26024 5356 26036
rect 5040 25996 5356 26024
rect 5040 25984 5046 25996
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 5810 25984 5816 26036
rect 5868 26024 5874 26036
rect 7561 26027 7619 26033
rect 7561 26024 7573 26027
rect 5868 25996 7573 26024
rect 5868 25984 5874 25996
rect 7561 25993 7573 25996
rect 7607 25993 7619 26027
rect 7561 25987 7619 25993
rect 7650 25984 7656 26036
rect 7708 25984 7714 26036
rect 8386 25984 8392 26036
rect 8444 25984 8450 26036
rect 9122 25984 9128 26036
rect 9180 25984 9186 26036
rect 5902 25956 5908 25968
rect 4172 25928 5908 25956
rect 934 25848 940 25900
rect 992 25888 998 25900
rect 4172 25897 4200 25928
rect 5902 25916 5908 25928
rect 5960 25916 5966 25968
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 6972 25928 7604 25956
rect 6972 25916 6978 25928
rect 7576 25900 7604 25928
rect 1489 25891 1547 25897
rect 1489 25888 1501 25891
rect 992 25860 1501 25888
rect 992 25848 998 25860
rect 1489 25857 1501 25860
rect 1535 25857 1547 25891
rect 1489 25851 1547 25857
rect 4157 25891 4215 25897
rect 4157 25857 4169 25891
rect 4203 25857 4215 25891
rect 4157 25851 4215 25857
rect 5534 25848 5540 25900
rect 5592 25848 5598 25900
rect 5810 25848 5816 25900
rect 5868 25848 5874 25900
rect 5991 25892 6049 25897
rect 5991 25891 6132 25892
rect 5991 25857 6003 25891
rect 6037 25888 6132 25891
rect 6178 25888 6184 25900
rect 6037 25864 6184 25888
rect 6037 25857 6049 25864
rect 6104 25860 6184 25864
rect 5991 25851 6049 25857
rect 6178 25848 6184 25860
rect 6236 25888 6242 25900
rect 7006 25888 7012 25900
rect 6236 25860 7012 25888
rect 6236 25848 6242 25860
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7558 25848 7564 25900
rect 7616 25848 7622 25900
rect 7668 25888 7696 25984
rect 8110 25916 8116 25968
rect 8168 25956 8174 25968
rect 9033 25959 9091 25965
rect 9033 25956 9045 25959
rect 8168 25928 9045 25956
rect 8168 25916 8174 25928
rect 9033 25925 9045 25928
rect 9079 25925 9091 25959
rect 9033 25919 9091 25925
rect 7668 25860 7788 25888
rect 5552 25820 5580 25848
rect 5902 25820 5908 25832
rect 5552 25792 5908 25820
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25820 6975 25823
rect 7098 25820 7104 25832
rect 6963 25792 7104 25820
rect 6963 25789 6975 25792
rect 6917 25783 6975 25789
rect 7098 25780 7104 25792
rect 7156 25820 7162 25832
rect 7650 25820 7656 25832
rect 7156 25792 7656 25820
rect 7156 25780 7162 25792
rect 7650 25780 7656 25792
rect 7708 25780 7714 25832
rect 7760 25829 7788 25860
rect 8018 25848 8024 25900
rect 8076 25888 8082 25900
rect 8076 25860 8708 25888
rect 8076 25848 8082 25860
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25789 7803 25823
rect 7745 25783 7803 25789
rect 5813 25755 5871 25761
rect 5813 25721 5825 25755
rect 5859 25752 5871 25755
rect 7282 25752 7288 25764
rect 5859 25724 7288 25752
rect 5859 25721 5871 25724
rect 5813 25715 5871 25721
rect 7282 25712 7288 25724
rect 7340 25712 7346 25764
rect 7760 25752 7788 25783
rect 7834 25780 7840 25832
rect 7892 25820 7898 25832
rect 8481 25823 8539 25829
rect 8481 25820 8493 25823
rect 7892 25792 8493 25820
rect 7892 25780 7898 25792
rect 8481 25789 8493 25792
rect 8527 25789 8539 25823
rect 8481 25783 8539 25789
rect 8573 25823 8631 25829
rect 8573 25789 8585 25823
rect 8619 25789 8631 25823
rect 8680 25820 8708 25860
rect 8754 25820 8760 25832
rect 8680 25792 8760 25820
rect 8573 25783 8631 25789
rect 8588 25752 8616 25783
rect 8754 25780 8760 25792
rect 8812 25780 8818 25832
rect 7760 25724 8616 25752
rect 1762 25644 1768 25696
rect 1820 25684 1826 25696
rect 4341 25687 4399 25693
rect 4341 25684 4353 25687
rect 1820 25656 4353 25684
rect 1820 25644 1826 25656
rect 4341 25653 4353 25656
rect 4387 25653 4399 25687
rect 4341 25647 4399 25653
rect 7193 25687 7251 25693
rect 7193 25653 7205 25687
rect 7239 25684 7251 25687
rect 7650 25684 7656 25696
rect 7239 25656 7656 25684
rect 7239 25653 7251 25656
rect 7193 25647 7251 25653
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 8021 25687 8079 25693
rect 8021 25653 8033 25687
rect 8067 25684 8079 25687
rect 8754 25684 8760 25696
rect 8067 25656 8760 25684
rect 8067 25653 8079 25656
rect 8021 25647 8079 25653
rect 8754 25644 8760 25656
rect 8812 25644 8818 25696
rect 1104 25594 9936 25616
rect 1104 25542 3610 25594
rect 3662 25542 3674 25594
rect 3726 25542 3738 25594
rect 3790 25542 3802 25594
rect 3854 25542 3866 25594
rect 3918 25542 5210 25594
rect 5262 25542 5274 25594
rect 5326 25542 5338 25594
rect 5390 25542 5402 25594
rect 5454 25542 5466 25594
rect 5518 25542 6810 25594
rect 6862 25542 6874 25594
rect 6926 25542 6938 25594
rect 6990 25542 7002 25594
rect 7054 25542 7066 25594
rect 7118 25542 8410 25594
rect 8462 25542 8474 25594
rect 8526 25542 8538 25594
rect 8590 25542 8602 25594
rect 8654 25542 8666 25594
rect 8718 25542 9936 25594
rect 1104 25520 9936 25542
rect 2774 25440 2780 25492
rect 2832 25440 2838 25492
rect 7190 25440 7196 25492
rect 7248 25480 7254 25492
rect 7561 25483 7619 25489
rect 7561 25480 7573 25483
rect 7248 25452 7573 25480
rect 7248 25440 7254 25452
rect 7561 25449 7573 25452
rect 7607 25449 7619 25483
rect 7561 25443 7619 25449
rect 2792 25412 2820 25440
rect 7834 25412 7840 25424
rect 2792 25384 7840 25412
rect 7834 25372 7840 25384
rect 7892 25412 7898 25424
rect 9582 25412 9588 25424
rect 7892 25384 9588 25412
rect 7892 25372 7898 25384
rect 9582 25372 9588 25384
rect 9640 25372 9646 25424
rect 1578 25304 1584 25356
rect 1636 25344 1642 25356
rect 6178 25344 6184 25356
rect 1636 25316 6184 25344
rect 1636 25304 1642 25316
rect 5000 25152 5028 25316
rect 6178 25304 6184 25316
rect 6236 25304 6242 25356
rect 7469 25279 7527 25285
rect 7469 25276 7481 25279
rect 7300 25248 7481 25276
rect 7300 25152 7328 25248
rect 7469 25245 7481 25248
rect 7515 25245 7527 25279
rect 7469 25239 7527 25245
rect 4982 25100 4988 25152
rect 5040 25100 5046 25152
rect 7282 25100 7288 25152
rect 7340 25100 7346 25152
rect 1104 25050 9936 25072
rect 1104 24998 2950 25050
rect 3002 24998 3014 25050
rect 3066 24998 3078 25050
rect 3130 24998 3142 25050
rect 3194 24998 3206 25050
rect 3258 24998 4550 25050
rect 4602 24998 4614 25050
rect 4666 24998 4678 25050
rect 4730 24998 4742 25050
rect 4794 24998 4806 25050
rect 4858 24998 6150 25050
rect 6202 24998 6214 25050
rect 6266 24998 6278 25050
rect 6330 24998 6342 25050
rect 6394 24998 6406 25050
rect 6458 24998 7750 25050
rect 7802 24998 7814 25050
rect 7866 24998 7878 25050
rect 7930 24998 7942 25050
rect 7994 24998 8006 25050
rect 8058 24998 9350 25050
rect 9402 24998 9414 25050
rect 9466 24998 9478 25050
rect 9530 24998 9542 25050
rect 9594 24998 9606 25050
rect 9658 24998 9936 25050
rect 1104 24976 9936 24998
rect 5534 24896 5540 24948
rect 5592 24936 5598 24948
rect 7926 24936 7932 24948
rect 5592 24908 7932 24936
rect 5592 24896 5598 24908
rect 7926 24896 7932 24908
rect 7984 24896 7990 24948
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 992 24772 1409 24800
rect 992 24760 998 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 6638 24760 6644 24812
rect 6696 24800 6702 24812
rect 11054 24800 11060 24812
rect 6696 24772 11060 24800
rect 6696 24760 6702 24772
rect 11054 24760 11060 24772
rect 11112 24760 11118 24812
rect 2314 24692 2320 24744
rect 2372 24732 2378 24744
rect 7742 24732 7748 24744
rect 2372 24704 7748 24732
rect 2372 24692 2378 24704
rect 7742 24692 7748 24704
rect 7800 24692 7806 24744
rect 8110 24692 8116 24744
rect 8168 24732 8174 24744
rect 9306 24732 9312 24744
rect 8168 24704 9312 24732
rect 8168 24692 8174 24704
rect 9306 24692 9312 24704
rect 9364 24692 9370 24744
rect 842 24556 848 24608
rect 900 24596 906 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 900 24568 1593 24596
rect 900 24556 906 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 1104 24506 9936 24528
rect 1104 24454 3610 24506
rect 3662 24454 3674 24506
rect 3726 24454 3738 24506
rect 3790 24454 3802 24506
rect 3854 24454 3866 24506
rect 3918 24454 5210 24506
rect 5262 24454 5274 24506
rect 5326 24454 5338 24506
rect 5390 24454 5402 24506
rect 5454 24454 5466 24506
rect 5518 24454 6810 24506
rect 6862 24454 6874 24506
rect 6926 24454 6938 24506
rect 6990 24454 7002 24506
rect 7054 24454 7066 24506
rect 7118 24454 8410 24506
rect 8462 24454 8474 24506
rect 8526 24454 8538 24506
rect 8590 24454 8602 24506
rect 8654 24454 8666 24506
rect 8718 24454 9936 24506
rect 1104 24432 9936 24454
rect 7374 24352 7380 24404
rect 7432 24392 7438 24404
rect 7834 24392 7840 24404
rect 7432 24364 7840 24392
rect 7432 24352 7438 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 9309 24395 9367 24401
rect 9309 24392 9321 24395
rect 8352 24364 9321 24392
rect 8352 24352 8358 24364
rect 9309 24361 9321 24364
rect 9355 24392 9367 24395
rect 10870 24392 10876 24404
rect 9355 24364 10876 24392
rect 9355 24361 9367 24364
rect 9309 24355 9367 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 7285 24327 7343 24333
rect 7285 24293 7297 24327
rect 7331 24324 7343 24327
rect 7466 24324 7472 24336
rect 7331 24296 7472 24324
rect 7331 24293 7343 24296
rect 7285 24287 7343 24293
rect 7466 24284 7472 24296
rect 7524 24284 7530 24336
rect 8110 24284 8116 24336
rect 8168 24284 8174 24336
rect 9214 24284 9220 24336
rect 9272 24284 9278 24336
rect 7837 24259 7895 24265
rect 7837 24256 7849 24259
rect 2608 24228 5856 24256
rect 2608 24200 2636 24228
rect 2590 24148 2596 24200
rect 2648 24148 2654 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 5718 24188 5724 24200
rect 4203 24160 5724 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 5718 24148 5724 24160
rect 5776 24148 5782 24200
rect 5828 24188 5856 24228
rect 7576 24228 7849 24256
rect 7101 24191 7159 24197
rect 5828 24160 7052 24188
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 5810 24120 5816 24132
rect 2924 24092 5816 24120
rect 2924 24080 2930 24092
rect 5810 24080 5816 24092
rect 5868 24120 5874 24132
rect 6917 24123 6975 24129
rect 6917 24120 6929 24123
rect 5868 24092 6929 24120
rect 5868 24080 5874 24092
rect 6917 24089 6929 24092
rect 6963 24089 6975 24123
rect 6917 24083 6975 24089
rect 2222 24012 2228 24064
rect 2280 24052 2286 24064
rect 4341 24055 4399 24061
rect 4341 24052 4353 24055
rect 2280 24024 4353 24052
rect 2280 24012 2286 24024
rect 4341 24021 4353 24024
rect 4387 24021 4399 24055
rect 4341 24015 4399 24021
rect 4982 24012 4988 24064
rect 5040 24052 5046 24064
rect 5718 24052 5724 24064
rect 5040 24024 5724 24052
rect 5040 24012 5046 24024
rect 5718 24012 5724 24024
rect 5776 24012 5782 24064
rect 7024 24052 7052 24160
rect 7101 24157 7113 24191
rect 7147 24188 7159 24191
rect 7147 24184 7236 24188
rect 7282 24184 7288 24200
rect 7147 24160 7288 24184
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 7208 24156 7288 24160
rect 7282 24148 7288 24156
rect 7340 24182 7346 24200
rect 7576 24182 7604 24228
rect 7837 24225 7849 24228
rect 7883 24225 7895 24259
rect 7837 24219 7895 24225
rect 7340 24154 7604 24182
rect 7340 24148 7346 24154
rect 7742 24148 7748 24200
rect 7800 24148 7806 24200
rect 7852 24188 7880 24219
rect 7926 24216 7932 24268
rect 7984 24256 7990 24268
rect 7984 24228 8432 24256
rect 7984 24216 7990 24228
rect 8404 24197 8432 24228
rect 9232 24197 9260 24284
rect 8297 24191 8355 24197
rect 8297 24188 8309 24191
rect 7852 24160 8309 24188
rect 8297 24157 8309 24160
rect 8343 24157 8355 24191
rect 8297 24151 8355 24157
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 7834 24080 7840 24132
rect 7892 24120 7898 24132
rect 8113 24123 8171 24129
rect 8113 24120 8125 24123
rect 7892 24092 8125 24120
rect 7892 24080 7898 24092
rect 8113 24089 8125 24092
rect 8159 24089 8171 24123
rect 8113 24083 8171 24089
rect 7653 24055 7711 24061
rect 7653 24052 7665 24055
rect 7024 24024 7665 24052
rect 7653 24021 7665 24024
rect 7699 24021 7711 24055
rect 7653 24015 7711 24021
rect 7742 24012 7748 24064
rect 7800 24052 7806 24064
rect 8386 24052 8392 24064
rect 7800 24024 8392 24052
rect 7800 24012 7806 24024
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 1104 23962 9936 23984
rect 1104 23910 2950 23962
rect 3002 23910 3014 23962
rect 3066 23910 3078 23962
rect 3130 23910 3142 23962
rect 3194 23910 3206 23962
rect 3258 23910 4550 23962
rect 4602 23910 4614 23962
rect 4666 23910 4678 23962
rect 4730 23910 4742 23962
rect 4794 23910 4806 23962
rect 4858 23910 6150 23962
rect 6202 23910 6214 23962
rect 6266 23910 6278 23962
rect 6330 23910 6342 23962
rect 6394 23910 6406 23962
rect 6458 23910 7750 23962
rect 7802 23910 7814 23962
rect 7866 23910 7878 23962
rect 7930 23910 7942 23962
rect 7994 23910 8006 23962
rect 8058 23910 9350 23962
rect 9402 23910 9414 23962
rect 9466 23910 9478 23962
rect 9530 23910 9542 23962
rect 9594 23910 9606 23962
rect 9658 23910 9936 23962
rect 1104 23888 9936 23910
rect 1578 23808 1584 23860
rect 1636 23808 1642 23860
rect 7466 23808 7472 23860
rect 7524 23848 7530 23860
rect 8294 23848 8300 23860
rect 7524 23820 8300 23848
rect 7524 23808 7530 23820
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 934 23672 940 23724
rect 992 23712 998 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 992 23684 1409 23712
rect 992 23672 998 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 4341 23715 4399 23721
rect 4341 23681 4353 23715
rect 4387 23712 4399 23715
rect 5626 23712 5632 23724
rect 4387 23684 5632 23712
rect 4387 23681 4399 23684
rect 4341 23675 4399 23681
rect 5626 23672 5632 23684
rect 5684 23672 5690 23724
rect 8386 23604 8392 23656
rect 8444 23644 8450 23656
rect 9306 23644 9312 23656
rect 8444 23616 9312 23644
rect 8444 23604 8450 23616
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 2406 23536 2412 23588
rect 2464 23576 2470 23588
rect 4982 23576 4988 23588
rect 2464 23548 4988 23576
rect 2464 23536 2470 23548
rect 4982 23536 4988 23548
rect 5040 23536 5046 23588
rect 3326 23468 3332 23520
rect 3384 23508 3390 23520
rect 4525 23511 4583 23517
rect 4525 23508 4537 23511
rect 3384 23480 4537 23508
rect 3384 23468 3390 23480
rect 4525 23477 4537 23480
rect 4571 23477 4583 23511
rect 4525 23471 4583 23477
rect 1104 23418 9936 23440
rect 1104 23366 3610 23418
rect 3662 23366 3674 23418
rect 3726 23366 3738 23418
rect 3790 23366 3802 23418
rect 3854 23366 3866 23418
rect 3918 23366 5210 23418
rect 5262 23366 5274 23418
rect 5326 23366 5338 23418
rect 5390 23366 5402 23418
rect 5454 23366 5466 23418
rect 5518 23366 6810 23418
rect 6862 23366 6874 23418
rect 6926 23366 6938 23418
rect 6990 23366 7002 23418
rect 7054 23366 7066 23418
rect 7118 23366 8410 23418
rect 8462 23366 8474 23418
rect 8526 23366 8538 23418
rect 8590 23366 8602 23418
rect 8654 23366 8666 23418
rect 8718 23366 9936 23418
rect 1104 23344 9936 23366
rect 3234 23264 3240 23316
rect 3292 23304 3298 23316
rect 3602 23304 3608 23316
rect 3292 23276 3608 23304
rect 3292 23264 3298 23276
rect 3602 23264 3608 23276
rect 3660 23264 3666 23316
rect 8665 23307 8723 23313
rect 8665 23273 8677 23307
rect 8711 23304 8723 23307
rect 9214 23304 9220 23316
rect 8711 23276 9220 23304
rect 8711 23273 8723 23276
rect 8665 23267 8723 23273
rect 9214 23264 9220 23276
rect 9272 23304 9278 23316
rect 11422 23304 11428 23316
rect 9272 23276 11428 23304
rect 9272 23264 9278 23276
rect 11422 23264 11428 23276
rect 11480 23264 11486 23316
rect 5810 23196 5816 23248
rect 5868 23236 5874 23248
rect 9493 23239 9551 23245
rect 9493 23236 9505 23239
rect 5868 23208 9505 23236
rect 5868 23196 5874 23208
rect 9493 23205 9505 23208
rect 9539 23236 9551 23239
rect 10042 23236 10048 23248
rect 9539 23208 10048 23236
rect 9539 23205 9551 23208
rect 9493 23199 9551 23205
rect 10042 23196 10048 23208
rect 10100 23196 10106 23248
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 5994 23100 6000 23112
rect 4203 23072 6000 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 8202 23060 8208 23112
rect 8260 23100 8266 23112
rect 8481 23103 8539 23109
rect 8481 23100 8493 23103
rect 8260 23072 8493 23100
rect 8260 23060 8266 23072
rect 8481 23069 8493 23072
rect 8527 23069 8539 23103
rect 8481 23063 8539 23069
rect 8938 23060 8944 23112
rect 8996 23100 9002 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8996 23072 9229 23100
rect 8996 23060 9002 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9582 23032 9588 23044
rect 8956 23004 9588 23032
rect 8956 22976 8984 23004
rect 9582 22992 9588 23004
rect 9640 22992 9646 23044
rect 2314 22924 2320 22976
rect 2372 22964 2378 22976
rect 4341 22967 4399 22973
rect 4341 22964 4353 22967
rect 2372 22936 4353 22964
rect 2372 22924 2378 22936
rect 4341 22933 4353 22936
rect 4387 22933 4399 22967
rect 4341 22927 4399 22933
rect 7374 22924 7380 22976
rect 7432 22964 7438 22976
rect 8202 22964 8208 22976
rect 7432 22936 8208 22964
rect 7432 22924 7438 22936
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 8938 22924 8944 22976
rect 8996 22924 9002 22976
rect 1104 22874 9936 22896
rect 1104 22822 2950 22874
rect 3002 22822 3014 22874
rect 3066 22822 3078 22874
rect 3130 22822 3142 22874
rect 3194 22822 3206 22874
rect 3258 22822 4550 22874
rect 4602 22822 4614 22874
rect 4666 22822 4678 22874
rect 4730 22822 4742 22874
rect 4794 22822 4806 22874
rect 4858 22822 6150 22874
rect 6202 22822 6214 22874
rect 6266 22822 6278 22874
rect 6330 22822 6342 22874
rect 6394 22822 6406 22874
rect 6458 22822 7750 22874
rect 7802 22822 7814 22874
rect 7866 22822 7878 22874
rect 7930 22822 7942 22874
rect 7994 22822 8006 22874
rect 8058 22822 9350 22874
rect 9402 22822 9414 22874
rect 9466 22822 9478 22874
rect 9530 22822 9542 22874
rect 9594 22822 9606 22874
rect 9658 22822 9936 22874
rect 1104 22800 9936 22822
rect 3050 22720 3056 22772
rect 3108 22760 3114 22772
rect 3510 22760 3516 22772
rect 3108 22732 3516 22760
rect 3108 22720 3114 22732
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4246 22720 4252 22772
rect 4304 22760 4310 22772
rect 4522 22760 4528 22772
rect 4304 22732 4528 22760
rect 4304 22720 4310 22732
rect 4522 22720 4528 22732
rect 4580 22720 4586 22772
rect 1673 22695 1731 22701
rect 1673 22661 1685 22695
rect 1719 22692 1731 22695
rect 2866 22692 2872 22704
rect 1719 22664 2872 22692
rect 1719 22661 1731 22664
rect 1673 22655 1731 22661
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 6546 22692 6552 22704
rect 4080 22664 6552 22692
rect 934 22584 940 22636
rect 992 22624 998 22636
rect 4080 22633 4108 22664
rect 6546 22652 6552 22664
rect 6604 22652 6610 22704
rect 7190 22652 7196 22704
rect 7248 22692 7254 22704
rect 7745 22695 7803 22701
rect 7745 22692 7757 22695
rect 7248 22664 7757 22692
rect 7248 22652 7254 22664
rect 7745 22661 7757 22664
rect 7791 22661 7803 22695
rect 7745 22655 7803 22661
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 992 22596 1501 22624
rect 992 22584 998 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 1489 22587 1547 22593
rect 4065 22627 4123 22633
rect 4065 22593 4077 22627
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22624 4399 22627
rect 9950 22624 9956 22636
rect 4387 22596 9956 22624
rect 4387 22593 4399 22596
rect 4341 22587 4399 22593
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 3970 22380 3976 22432
rect 4028 22420 4034 22432
rect 4249 22423 4307 22429
rect 4249 22420 4261 22423
rect 4028 22392 4261 22420
rect 4028 22380 4034 22392
rect 4249 22389 4261 22392
rect 4295 22389 4307 22423
rect 4249 22383 4307 22389
rect 4525 22423 4583 22429
rect 4525 22389 4537 22423
rect 4571 22420 4583 22423
rect 4614 22420 4620 22432
rect 4571 22392 4620 22420
rect 4571 22389 4583 22392
rect 4525 22383 4583 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 7834 22380 7840 22432
rect 7892 22380 7898 22432
rect 1104 22330 9936 22352
rect 1104 22278 3610 22330
rect 3662 22278 3674 22330
rect 3726 22278 3738 22330
rect 3790 22278 3802 22330
rect 3854 22278 3866 22330
rect 3918 22278 5210 22330
rect 5262 22278 5274 22330
rect 5326 22278 5338 22330
rect 5390 22278 5402 22330
rect 5454 22278 5466 22330
rect 5518 22278 6810 22330
rect 6862 22278 6874 22330
rect 6926 22278 6938 22330
rect 6990 22278 7002 22330
rect 7054 22278 7066 22330
rect 7118 22278 8410 22330
rect 8462 22278 8474 22330
rect 8526 22278 8538 22330
rect 8590 22278 8602 22330
rect 8654 22278 8666 22330
rect 8718 22278 9936 22330
rect 1104 22256 9936 22278
rect 4246 22108 4252 22160
rect 4304 22148 4310 22160
rect 4614 22148 4620 22160
rect 4304 22120 4620 22148
rect 4304 22108 4310 22120
rect 4614 22108 4620 22120
rect 4672 22108 4678 22160
rect 7650 22040 7656 22092
rect 7708 22080 7714 22092
rect 7708 22052 9352 22080
rect 7708 22040 7714 22052
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4522 22012 4528 22024
rect 4111 21984 4528 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 9324 22021 9352 22052
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 1673 21947 1731 21953
rect 1673 21913 1685 21947
rect 1719 21944 1731 21947
rect 5902 21944 5908 21956
rect 1719 21916 5908 21944
rect 1719 21913 1731 21916
rect 1673 21907 1731 21913
rect 5902 21904 5908 21916
rect 5960 21904 5966 21956
rect 6748 21916 9536 21944
rect 6748 21888 6776 21916
rect 2130 21836 2136 21888
rect 2188 21876 2194 21888
rect 4249 21879 4307 21885
rect 4249 21876 4261 21879
rect 2188 21848 4261 21876
rect 2188 21836 2194 21848
rect 4249 21845 4261 21848
rect 4295 21845 4307 21879
rect 4249 21839 4307 21845
rect 6730 21836 6736 21888
rect 6788 21836 6794 21888
rect 9508 21885 9536 21916
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21845 9551 21879
rect 9493 21839 9551 21845
rect 1104 21786 9936 21808
rect 1104 21734 2950 21786
rect 3002 21734 3014 21786
rect 3066 21734 3078 21786
rect 3130 21734 3142 21786
rect 3194 21734 3206 21786
rect 3258 21734 4550 21786
rect 4602 21734 4614 21786
rect 4666 21734 4678 21786
rect 4730 21734 4742 21786
rect 4794 21734 4806 21786
rect 4858 21734 6150 21786
rect 6202 21734 6214 21786
rect 6266 21734 6278 21786
rect 6330 21734 6342 21786
rect 6394 21734 6406 21786
rect 6458 21734 7750 21786
rect 7802 21734 7814 21786
rect 7866 21734 7878 21786
rect 7930 21734 7942 21786
rect 7994 21734 8006 21786
rect 8058 21734 9350 21786
rect 9402 21734 9414 21786
rect 9466 21734 9478 21786
rect 9530 21734 9542 21786
rect 9594 21734 9606 21786
rect 9658 21734 9936 21786
rect 1104 21712 9936 21734
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 5776 21508 7205 21536
rect 5776 21496 5782 21508
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 7340 21508 7389 21536
rect 7340 21496 7346 21508
rect 7377 21505 7389 21508
rect 7423 21536 7435 21539
rect 7423 21508 7512 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7484 21480 7512 21508
rect 7466 21428 7472 21480
rect 7524 21428 7530 21480
rect 7558 21292 7564 21344
rect 7616 21292 7622 21344
rect 1104 21242 9936 21264
rect 1104 21190 3610 21242
rect 3662 21190 3674 21242
rect 3726 21190 3738 21242
rect 3790 21190 3802 21242
rect 3854 21190 3866 21242
rect 3918 21190 5210 21242
rect 5262 21190 5274 21242
rect 5326 21190 5338 21242
rect 5390 21190 5402 21242
rect 5454 21190 5466 21242
rect 5518 21190 6810 21242
rect 6862 21190 6874 21242
rect 6926 21190 6938 21242
rect 6990 21190 7002 21242
rect 7054 21190 7066 21242
rect 7118 21190 8410 21242
rect 8462 21190 8474 21242
rect 8526 21190 8538 21242
rect 8590 21190 8602 21242
rect 8654 21190 8666 21242
rect 8718 21190 9936 21242
rect 1104 21168 9936 21190
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 1673 20859 1731 20865
rect 1673 20825 1685 20859
rect 1719 20856 1731 20859
rect 5994 20856 6000 20868
rect 1719 20828 6000 20856
rect 1719 20825 1731 20828
rect 1673 20819 1731 20825
rect 5994 20816 6000 20828
rect 6052 20816 6058 20868
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 7374 20788 7380 20800
rect 6788 20760 7380 20788
rect 6788 20748 6794 20760
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 1104 20698 9936 20720
rect 1104 20646 2950 20698
rect 3002 20646 3014 20698
rect 3066 20646 3078 20698
rect 3130 20646 3142 20698
rect 3194 20646 3206 20698
rect 3258 20646 4550 20698
rect 4602 20646 4614 20698
rect 4666 20646 4678 20698
rect 4730 20646 4742 20698
rect 4794 20646 4806 20698
rect 4858 20646 6150 20698
rect 6202 20646 6214 20698
rect 6266 20646 6278 20698
rect 6330 20646 6342 20698
rect 6394 20646 6406 20698
rect 6458 20646 7750 20698
rect 7802 20646 7814 20698
rect 7866 20646 7878 20698
rect 7930 20646 7942 20698
rect 7994 20646 8006 20698
rect 8058 20646 9350 20698
rect 9402 20646 9414 20698
rect 9466 20646 9478 20698
rect 9530 20646 9542 20698
rect 9594 20646 9606 20698
rect 9658 20646 9936 20698
rect 1104 20624 9936 20646
rect 8754 20408 8760 20460
rect 8812 20448 8818 20460
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 8812 20420 9321 20448
rect 8812 20408 8818 20420
rect 9309 20417 9321 20420
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 9493 20247 9551 20253
rect 9493 20244 9505 20247
rect 8904 20216 9505 20244
rect 8904 20204 8910 20216
rect 9493 20213 9505 20216
rect 9539 20244 9551 20247
rect 9582 20244 9588 20256
rect 9539 20216 9588 20244
rect 9539 20213 9551 20216
rect 9493 20207 9551 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 1104 20154 9936 20176
rect 1104 20102 3610 20154
rect 3662 20102 3674 20154
rect 3726 20102 3738 20154
rect 3790 20102 3802 20154
rect 3854 20102 3866 20154
rect 3918 20102 5210 20154
rect 5262 20102 5274 20154
rect 5326 20102 5338 20154
rect 5390 20102 5402 20154
rect 5454 20102 5466 20154
rect 5518 20102 6810 20154
rect 6862 20102 6874 20154
rect 6926 20102 6938 20154
rect 6990 20102 7002 20154
rect 7054 20102 7066 20154
rect 7118 20102 8410 20154
rect 8462 20102 8474 20154
rect 8526 20102 8538 20154
rect 8590 20102 8602 20154
rect 8654 20102 8666 20154
rect 8718 20102 9936 20154
rect 1104 20080 9936 20102
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 8352 19808 9321 19836
rect 8352 19796 8358 19808
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 1673 19771 1731 19777
rect 1673 19737 1685 19771
rect 1719 19768 1731 19771
rect 5718 19768 5724 19780
rect 1719 19740 5724 19768
rect 1719 19737 1731 19740
rect 1673 19731 1731 19737
rect 5718 19728 5724 19740
rect 5776 19728 5782 19780
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 9088 19672 9505 19700
rect 9088 19660 9094 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 9493 19663 9551 19669
rect 1104 19610 9936 19632
rect 1104 19558 2950 19610
rect 3002 19558 3014 19610
rect 3066 19558 3078 19610
rect 3130 19558 3142 19610
rect 3194 19558 3206 19610
rect 3258 19558 4550 19610
rect 4602 19558 4614 19610
rect 4666 19558 4678 19610
rect 4730 19558 4742 19610
rect 4794 19558 4806 19610
rect 4858 19558 6150 19610
rect 6202 19558 6214 19610
rect 6266 19558 6278 19610
rect 6330 19558 6342 19610
rect 6394 19558 6406 19610
rect 6458 19558 7750 19610
rect 7802 19558 7814 19610
rect 7866 19558 7878 19610
rect 7930 19558 7942 19610
rect 7994 19558 8006 19610
rect 8058 19558 9350 19610
rect 9402 19558 9414 19610
rect 9466 19558 9478 19610
rect 9530 19558 9542 19610
rect 9594 19558 9606 19610
rect 9658 19558 9936 19610
rect 1104 19536 9936 19558
rect 1104 19066 9936 19088
rect 1104 19014 3610 19066
rect 3662 19014 3674 19066
rect 3726 19014 3738 19066
rect 3790 19014 3802 19066
rect 3854 19014 3866 19066
rect 3918 19014 5210 19066
rect 5262 19014 5274 19066
rect 5326 19014 5338 19066
rect 5390 19014 5402 19066
rect 5454 19014 5466 19066
rect 5518 19014 6810 19066
rect 6862 19014 6874 19066
rect 6926 19014 6938 19066
rect 6990 19014 7002 19066
rect 7054 19014 7066 19066
rect 7118 19014 8410 19066
rect 8462 19014 8474 19066
rect 8526 19014 8538 19066
rect 8590 19014 8602 19066
rect 8654 19014 8666 19066
rect 8718 19014 9936 19066
rect 1104 18992 9936 19014
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7650 18952 7656 18964
rect 7340 18924 7656 18952
rect 7340 18912 7346 18924
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 7190 18844 7196 18896
rect 7248 18884 7254 18896
rect 7742 18884 7748 18896
rect 7248 18856 7748 18884
rect 7248 18844 7254 18856
rect 7742 18844 7748 18856
rect 7800 18844 7806 18896
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 3418 18816 3424 18828
rect 2271 18788 3424 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 7282 18776 7288 18828
rect 7340 18776 7346 18828
rect 7760 18816 7788 18844
rect 7668 18788 7788 18816
rect 4890 18708 4896 18760
rect 4948 18708 4954 18760
rect 7300 18748 7328 18776
rect 7668 18757 7696 18788
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 7300 18720 7389 18748
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18717 7711 18751
rect 7653 18711 7711 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18748 7803 18751
rect 8202 18748 8208 18760
rect 7791 18720 8208 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1397 18683 1455 18689
rect 1397 18680 1409 18683
rect 992 18652 1409 18680
rect 992 18640 998 18652
rect 1397 18649 1409 18652
rect 1443 18649 1455 18683
rect 4908 18680 4936 18708
rect 7282 18680 7288 18692
rect 4908 18652 7288 18680
rect 1397 18643 1455 18649
rect 7282 18640 7288 18652
rect 7340 18680 7346 18692
rect 7484 18680 7512 18711
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 7340 18652 7512 18680
rect 7340 18640 7346 18652
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 6788 18584 7205 18612
rect 6788 18572 6794 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7193 18575 7251 18581
rect 1104 18522 9936 18544
rect 1104 18470 2950 18522
rect 3002 18470 3014 18522
rect 3066 18470 3078 18522
rect 3130 18470 3142 18522
rect 3194 18470 3206 18522
rect 3258 18470 4550 18522
rect 4602 18470 4614 18522
rect 4666 18470 4678 18522
rect 4730 18470 4742 18522
rect 4794 18470 4806 18522
rect 4858 18470 6150 18522
rect 6202 18470 6214 18522
rect 6266 18470 6278 18522
rect 6330 18470 6342 18522
rect 6394 18470 6406 18522
rect 6458 18470 7750 18522
rect 7802 18470 7814 18522
rect 7866 18470 7878 18522
rect 7930 18470 7942 18522
rect 7994 18470 8006 18522
rect 8058 18470 9350 18522
rect 9402 18470 9414 18522
rect 9466 18470 9478 18522
rect 9530 18470 9542 18522
rect 9594 18470 9606 18522
rect 9658 18470 9936 18522
rect 1104 18448 9936 18470
rect 1489 18343 1547 18349
rect 1489 18309 1501 18343
rect 1535 18340 1547 18343
rect 2590 18340 2596 18352
rect 1535 18312 2596 18340
rect 1535 18309 1547 18312
rect 1489 18303 1547 18309
rect 2590 18300 2596 18312
rect 2648 18300 2654 18352
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 1104 17978 9936 18000
rect 1104 17926 3610 17978
rect 3662 17926 3674 17978
rect 3726 17926 3738 17978
rect 3790 17926 3802 17978
rect 3854 17926 3866 17978
rect 3918 17926 5210 17978
rect 5262 17926 5274 17978
rect 5326 17926 5338 17978
rect 5390 17926 5402 17978
rect 5454 17926 5466 17978
rect 5518 17926 6810 17978
rect 6862 17926 6874 17978
rect 6926 17926 6938 17978
rect 6990 17926 7002 17978
rect 7054 17926 7066 17978
rect 7118 17926 8410 17978
rect 8462 17926 8474 17978
rect 8526 17926 8538 17978
rect 8590 17926 8602 17978
rect 8654 17926 8666 17978
rect 8718 17926 9936 17978
rect 1104 17904 9936 17926
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 7466 17688 7472 17740
rect 7524 17728 7530 17740
rect 7524 17700 7880 17728
rect 7524 17688 7530 17700
rect 7300 17660 7328 17688
rect 7852 17669 7880 17700
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 7300 17632 7665 17660
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8294 17524 8300 17536
rect 7883 17496 8300 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 1104 17434 9936 17456
rect 1104 17382 2950 17434
rect 3002 17382 3014 17434
rect 3066 17382 3078 17434
rect 3130 17382 3142 17434
rect 3194 17382 3206 17434
rect 3258 17382 4550 17434
rect 4602 17382 4614 17434
rect 4666 17382 4678 17434
rect 4730 17382 4742 17434
rect 4794 17382 4806 17434
rect 4858 17382 6150 17434
rect 6202 17382 6214 17434
rect 6266 17382 6278 17434
rect 6330 17382 6342 17434
rect 6394 17382 6406 17434
rect 6458 17382 7750 17434
rect 7802 17382 7814 17434
rect 7866 17382 7878 17434
rect 7930 17382 7942 17434
rect 7994 17382 8006 17434
rect 8058 17382 9350 17434
rect 9402 17382 9414 17434
rect 9466 17382 9478 17434
rect 9530 17382 9542 17434
rect 9594 17382 9606 17434
rect 9658 17382 9936 17434
rect 1104 17360 9936 17382
rect 7558 17280 7564 17332
rect 7616 17280 7622 17332
rect 1489 17255 1547 17261
rect 1489 17221 1501 17255
rect 1535 17252 1547 17255
rect 2038 17252 2044 17264
rect 1535 17224 2044 17252
rect 1535 17221 1547 17224
rect 1489 17215 1547 17221
rect 2038 17212 2044 17224
rect 2096 17212 2102 17264
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 7576 17184 7604 17280
rect 7515 17156 7604 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 934 16940 940 16992
rect 992 16980 998 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 992 16952 1593 16980
rect 992 16940 998 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 7616 16952 7665 16980
rect 7616 16940 7622 16952
rect 7653 16949 7665 16952
rect 7699 16949 7711 16983
rect 7653 16943 7711 16949
rect 1104 16890 9936 16912
rect 1104 16838 3610 16890
rect 3662 16838 3674 16890
rect 3726 16838 3738 16890
rect 3790 16838 3802 16890
rect 3854 16838 3866 16890
rect 3918 16838 5210 16890
rect 5262 16838 5274 16890
rect 5326 16838 5338 16890
rect 5390 16838 5402 16890
rect 5454 16838 5466 16890
rect 5518 16838 6810 16890
rect 6862 16838 6874 16890
rect 6926 16838 6938 16890
rect 6990 16838 7002 16890
rect 7054 16838 7066 16890
rect 7118 16838 8410 16890
rect 8462 16838 8474 16890
rect 8526 16838 8538 16890
rect 8590 16838 8602 16890
rect 8654 16838 8666 16890
rect 8718 16838 9936 16890
rect 1104 16816 9936 16838
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7285 16779 7343 16785
rect 7285 16776 7297 16779
rect 7248 16748 7297 16776
rect 7248 16736 7254 16748
rect 7285 16745 7297 16748
rect 7331 16776 7343 16779
rect 7331 16748 8248 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 8220 16720 8248 16748
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 7668 16680 8125 16708
rect 7668 16584 7696 16680
rect 8113 16677 8125 16680
rect 8159 16677 8171 16711
rect 8113 16671 8171 16677
rect 8202 16668 8208 16720
rect 8260 16668 8266 16720
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16572 7619 16575
rect 7650 16572 7656 16584
rect 7607 16544 7656 16572
rect 7607 16541 7619 16544
rect 7561 16535 7619 16541
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7745 16575 7803 16581
rect 7745 16541 7757 16575
rect 7791 16572 7803 16575
rect 8021 16575 8079 16581
rect 8021 16572 8033 16575
rect 7791 16544 8033 16572
rect 7791 16541 7803 16544
rect 7745 16535 7803 16541
rect 8021 16541 8033 16544
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 7760 16504 7788 16535
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 9858 16572 9864 16584
rect 9355 16544 9864 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 8846 16504 8852 16516
rect 7300 16476 7788 16504
rect 7852 16476 8852 16504
rect 7300 16448 7328 16476
rect 7282 16396 7288 16448
rect 7340 16396 7346 16448
rect 7466 16396 7472 16448
rect 7524 16396 7530 16448
rect 7852 16445 7880 16476
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 7837 16439 7895 16445
rect 7837 16405 7849 16439
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 9493 16439 9551 16445
rect 9493 16436 9505 16439
rect 8352 16408 9505 16436
rect 8352 16396 8358 16408
rect 9493 16405 9505 16408
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 1104 16346 9936 16368
rect 1104 16294 2950 16346
rect 3002 16294 3014 16346
rect 3066 16294 3078 16346
rect 3130 16294 3142 16346
rect 3194 16294 3206 16346
rect 3258 16294 4550 16346
rect 4602 16294 4614 16346
rect 4666 16294 4678 16346
rect 4730 16294 4742 16346
rect 4794 16294 4806 16346
rect 4858 16294 6150 16346
rect 6202 16294 6214 16346
rect 6266 16294 6278 16346
rect 6330 16294 6342 16346
rect 6394 16294 6406 16346
rect 6458 16294 7750 16346
rect 7802 16294 7814 16346
rect 7866 16294 7878 16346
rect 7930 16294 7942 16346
rect 7994 16294 8006 16346
rect 8058 16294 9350 16346
rect 9402 16294 9414 16346
rect 9466 16294 9478 16346
rect 9530 16294 9542 16346
rect 9594 16294 9606 16346
rect 9658 16294 9936 16346
rect 1104 16272 9936 16294
rect 7650 16192 7656 16244
rect 7708 16192 7714 16244
rect 9858 16232 9864 16244
rect 9232 16204 9864 16232
rect 1489 16167 1547 16173
rect 1489 16133 1501 16167
rect 1535 16164 1547 16167
rect 4338 16164 4344 16176
rect 1535 16136 4344 16164
rect 1535 16133 1547 16136
rect 1489 16127 1547 16133
rect 4338 16124 4344 16136
rect 4396 16124 4402 16176
rect 7668 16096 7696 16192
rect 8754 16124 8760 16176
rect 8812 16164 8818 16176
rect 9232 16173 9260 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 9217 16167 9275 16173
rect 9217 16164 9229 16167
rect 8812 16136 9229 16164
rect 8812 16124 8818 16136
rect 9217 16133 9229 16136
rect 9263 16133 9275 16167
rect 9401 16167 9459 16173
rect 9401 16164 9413 16167
rect 9217 16127 9275 16133
rect 9324 16136 9413 16164
rect 9324 16096 9352 16136
rect 9401 16133 9413 16136
rect 9447 16133 9459 16167
rect 9401 16127 9459 16133
rect 7668 16068 9352 16096
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 8260 16000 9505 16028
rect 8260 15988 8266 16000
rect 9493 15997 9505 16000
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 992 15864 1593 15892
rect 992 15852 998 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 8941 15895 8999 15901
rect 8941 15892 8953 15895
rect 5684 15864 8953 15892
rect 5684 15852 5690 15864
rect 8941 15861 8953 15864
rect 8987 15861 8999 15895
rect 8941 15855 8999 15861
rect 1104 15802 9936 15824
rect 1104 15750 3610 15802
rect 3662 15750 3674 15802
rect 3726 15750 3738 15802
rect 3790 15750 3802 15802
rect 3854 15750 3866 15802
rect 3918 15750 5210 15802
rect 5262 15750 5274 15802
rect 5326 15750 5338 15802
rect 5390 15750 5402 15802
rect 5454 15750 5466 15802
rect 5518 15750 6810 15802
rect 6862 15750 6874 15802
rect 6926 15750 6938 15802
rect 6990 15750 7002 15802
rect 7054 15750 7066 15802
rect 7118 15750 8410 15802
rect 8462 15750 8474 15802
rect 8526 15750 8538 15802
rect 8590 15750 8602 15802
rect 8654 15750 8666 15802
rect 8718 15750 9936 15802
rect 1104 15728 9936 15750
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9214 15552 9220 15564
rect 9088 15524 9220 15552
rect 9088 15512 9094 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 3568 15456 9321 15484
rect 3568 15444 3574 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9493 15351 9551 15357
rect 9493 15348 9505 15351
rect 9272 15320 9505 15348
rect 9272 15308 9278 15320
rect 9493 15317 9505 15320
rect 9539 15317 9551 15351
rect 9493 15311 9551 15317
rect 1104 15258 9936 15280
rect 1104 15206 2950 15258
rect 3002 15206 3014 15258
rect 3066 15206 3078 15258
rect 3130 15206 3142 15258
rect 3194 15206 3206 15258
rect 3258 15206 4550 15258
rect 4602 15206 4614 15258
rect 4666 15206 4678 15258
rect 4730 15206 4742 15258
rect 4794 15206 4806 15258
rect 4858 15206 6150 15258
rect 6202 15206 6214 15258
rect 6266 15206 6278 15258
rect 6330 15206 6342 15258
rect 6394 15206 6406 15258
rect 6458 15206 7750 15258
rect 7802 15206 7814 15258
rect 7866 15206 7878 15258
rect 7930 15206 7942 15258
rect 7994 15206 8006 15258
rect 8058 15206 9350 15258
rect 9402 15206 9414 15258
rect 9466 15206 9478 15258
rect 9530 15206 9542 15258
rect 9594 15206 9606 15258
rect 9658 15206 9936 15258
rect 1104 15184 9936 15206
rect 1489 15079 1547 15085
rect 1489 15045 1501 15079
rect 1535 15076 1547 15079
rect 4430 15076 4436 15088
rect 1535 15048 4436 15076
rect 1535 15045 1547 15048
rect 1489 15039 1547 15045
rect 4430 15036 4436 15048
rect 4488 15036 4494 15088
rect 934 14764 940 14816
rect 992 14804 998 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 992 14776 1593 14804
rect 992 14764 998 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 1104 14714 9936 14736
rect 1104 14662 3610 14714
rect 3662 14662 3674 14714
rect 3726 14662 3738 14714
rect 3790 14662 3802 14714
rect 3854 14662 3866 14714
rect 3918 14662 5210 14714
rect 5262 14662 5274 14714
rect 5326 14662 5338 14714
rect 5390 14662 5402 14714
rect 5454 14662 5466 14714
rect 5518 14662 6810 14714
rect 6862 14662 6874 14714
rect 6926 14662 6938 14714
rect 6990 14662 7002 14714
rect 7054 14662 7066 14714
rect 7118 14662 8410 14714
rect 8462 14662 8474 14714
rect 8526 14662 8538 14714
rect 8590 14662 8602 14714
rect 8654 14662 8666 14714
rect 8718 14662 9936 14714
rect 1104 14640 9936 14662
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 8113 14535 8171 14541
rect 8113 14532 8125 14535
rect 7708 14504 8125 14532
rect 7708 14492 7714 14504
rect 8113 14501 8125 14504
rect 8159 14501 8171 14535
rect 8113 14495 8171 14501
rect 8202 14424 8208 14476
rect 8260 14424 8266 14476
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 8754 14464 8760 14476
rect 8619 14436 8760 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 8754 14424 8760 14436
rect 8812 14464 8818 14476
rect 9030 14464 9036 14476
rect 8812 14436 9036 14464
rect 8812 14424 8818 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 1489 14399 1547 14405
rect 1489 14365 1501 14399
rect 1535 14396 1547 14399
rect 4062 14396 4068 14408
rect 1535 14368 4068 14396
rect 1535 14365 1547 14368
rect 1489 14359 1547 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 8220 14396 8248 14424
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8220 14368 8677 14396
rect 8665 14365 8677 14368
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14396 9367 14399
rect 9766 14396 9772 14408
rect 9355 14368 9772 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 7282 14288 7288 14340
rect 7340 14328 7346 14340
rect 8573 14331 8631 14337
rect 8573 14328 8585 14331
rect 7340 14300 8585 14328
rect 7340 14288 7346 14300
rect 8573 14297 8585 14300
rect 8619 14297 8631 14331
rect 8573 14291 8631 14297
rect 934 14220 940 14272
rect 992 14260 998 14272
rect 1581 14263 1639 14269
rect 1581 14260 1593 14263
rect 992 14232 1593 14260
rect 992 14220 998 14232
rect 1581 14229 1593 14232
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 9088 14232 9505 14260
rect 9088 14220 9094 14232
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9493 14223 9551 14229
rect 1104 14170 9936 14192
rect 1104 14118 2950 14170
rect 3002 14118 3014 14170
rect 3066 14118 3078 14170
rect 3130 14118 3142 14170
rect 3194 14118 3206 14170
rect 3258 14118 4550 14170
rect 4602 14118 4614 14170
rect 4666 14118 4678 14170
rect 4730 14118 4742 14170
rect 4794 14118 4806 14170
rect 4858 14118 6150 14170
rect 6202 14118 6214 14170
rect 6266 14118 6278 14170
rect 6330 14118 6342 14170
rect 6394 14118 6406 14170
rect 6458 14118 7750 14170
rect 7802 14118 7814 14170
rect 7866 14118 7878 14170
rect 7930 14118 7942 14170
rect 7994 14118 8006 14170
rect 8058 14118 9350 14170
rect 9402 14118 9414 14170
rect 9466 14118 9478 14170
rect 9530 14118 9542 14170
rect 9594 14118 9606 14170
rect 9658 14118 9936 14170
rect 1104 14096 9936 14118
rect 1104 13626 9936 13648
rect 1104 13574 3610 13626
rect 3662 13574 3674 13626
rect 3726 13574 3738 13626
rect 3790 13574 3802 13626
rect 3854 13574 3866 13626
rect 3918 13574 5210 13626
rect 5262 13574 5274 13626
rect 5326 13574 5338 13626
rect 5390 13574 5402 13626
rect 5454 13574 5466 13626
rect 5518 13574 6810 13626
rect 6862 13574 6874 13626
rect 6926 13574 6938 13626
rect 6990 13574 7002 13626
rect 7054 13574 7066 13626
rect 7118 13574 8410 13626
rect 8462 13574 8474 13626
rect 8526 13574 8538 13626
rect 8590 13574 8602 13626
rect 8654 13574 8666 13626
rect 8718 13574 9936 13626
rect 1104 13552 9936 13574
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 7558 13376 7564 13388
rect 7432 13348 7564 13376
rect 7432 13336 7438 13348
rect 7558 13336 7564 13348
rect 7616 13376 7622 13388
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 7616 13348 7757 13376
rect 7616 13336 7622 13348
rect 7745 13345 7757 13348
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13308 1547 13311
rect 1854 13308 1860 13320
rect 1535 13280 1860 13308
rect 1535 13277 1547 13280
rect 1489 13271 1547 13277
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 8018 13268 8024 13320
rect 8076 13268 8082 13320
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7558 13240 7564 13252
rect 7340 13212 7564 13240
rect 7340 13200 7346 13212
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 992 13144 1593 13172
rect 992 13132 998 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 10962 13172 10968 13184
rect 8803 13144 10968 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 1104 13082 9936 13104
rect 1104 13030 2950 13082
rect 3002 13030 3014 13082
rect 3066 13030 3078 13082
rect 3130 13030 3142 13082
rect 3194 13030 3206 13082
rect 3258 13030 4550 13082
rect 4602 13030 4614 13082
rect 4666 13030 4678 13082
rect 4730 13030 4742 13082
rect 4794 13030 4806 13082
rect 4858 13030 6150 13082
rect 6202 13030 6214 13082
rect 6266 13030 6278 13082
rect 6330 13030 6342 13082
rect 6394 13030 6406 13082
rect 6458 13030 7750 13082
rect 7802 13030 7814 13082
rect 7866 13030 7878 13082
rect 7930 13030 7942 13082
rect 7994 13030 8006 13082
rect 8058 13030 9350 13082
rect 9402 13030 9414 13082
rect 9466 13030 9478 13082
rect 9530 13030 9542 13082
rect 9594 13030 9606 13082
rect 9658 13030 9936 13082
rect 1104 13008 9936 13030
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9214 12764 9220 12776
rect 8996 12736 9220 12764
rect 8996 12724 9002 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9674 12628 9680 12640
rect 8996 12600 9680 12628
rect 8996 12588 9002 12600
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 1104 12538 9936 12560
rect 1104 12486 3610 12538
rect 3662 12486 3674 12538
rect 3726 12486 3738 12538
rect 3790 12486 3802 12538
rect 3854 12486 3866 12538
rect 3918 12486 5210 12538
rect 5262 12486 5274 12538
rect 5326 12486 5338 12538
rect 5390 12486 5402 12538
rect 5454 12486 5466 12538
rect 5518 12486 6810 12538
rect 6862 12486 6874 12538
rect 6926 12486 6938 12538
rect 6990 12486 7002 12538
rect 7054 12486 7066 12538
rect 7118 12486 8410 12538
rect 8462 12486 8474 12538
rect 8526 12486 8538 12538
rect 8590 12486 8602 12538
rect 8654 12486 8666 12538
rect 8718 12486 9936 12538
rect 1104 12464 9936 12486
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 1946 12220 1952 12232
rect 1535 12192 1952 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 934 12044 940 12096
rect 992 12084 998 12096
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 992 12056 1593 12084
rect 992 12044 998 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 1104 11994 9936 12016
rect 1104 11942 2950 11994
rect 3002 11942 3014 11994
rect 3066 11942 3078 11994
rect 3130 11942 3142 11994
rect 3194 11942 3206 11994
rect 3258 11942 4550 11994
rect 4602 11942 4614 11994
rect 4666 11942 4678 11994
rect 4730 11942 4742 11994
rect 4794 11942 4806 11994
rect 4858 11942 6150 11994
rect 6202 11942 6214 11994
rect 6266 11942 6278 11994
rect 6330 11942 6342 11994
rect 6394 11942 6406 11994
rect 6458 11942 7750 11994
rect 7802 11942 7814 11994
rect 7866 11942 7878 11994
rect 7930 11942 7942 11994
rect 7994 11942 8006 11994
rect 8058 11942 9350 11994
rect 9402 11942 9414 11994
rect 9466 11942 9478 11994
rect 9530 11942 9542 11994
rect 9594 11942 9606 11994
rect 9658 11942 9936 11994
rect 1104 11920 9936 11942
rect 6730 11840 6736 11892
rect 6788 11840 6794 11892
rect 6748 11812 6776 11840
rect 6748 11784 8892 11812
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 8864 11753 8892 11784
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 7392 11676 7420 11704
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 7392 11648 8585 11676
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 8168 11512 9597 11540
rect 8168 11500 8174 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 1104 11450 9936 11472
rect 1104 11398 3610 11450
rect 3662 11398 3674 11450
rect 3726 11398 3738 11450
rect 3790 11398 3802 11450
rect 3854 11398 3866 11450
rect 3918 11398 5210 11450
rect 5262 11398 5274 11450
rect 5326 11398 5338 11450
rect 5390 11398 5402 11450
rect 5454 11398 5466 11450
rect 5518 11398 6810 11450
rect 6862 11398 6874 11450
rect 6926 11398 6938 11450
rect 6990 11398 7002 11450
rect 7054 11398 7066 11450
rect 7118 11398 8410 11450
rect 8462 11398 8474 11450
rect 8526 11398 8538 11450
rect 8590 11398 8602 11450
rect 8654 11398 8666 11450
rect 8718 11398 9936 11450
rect 1104 11376 9936 11398
rect 934 11296 940 11348
rect 992 11336 998 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 992 11308 1593 11336
rect 992 11296 998 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 1581 11299 1639 11305
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 9582 11336 9588 11348
rect 5592 11308 9588 11336
rect 5592 11296 5598 11308
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 8757 11271 8815 11277
rect 8757 11237 8769 11271
rect 8803 11268 8815 11271
rect 10226 11268 10232 11280
rect 8803 11240 10232 11268
rect 8803 11237 8815 11240
rect 8757 11231 8815 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7432 11172 7757 11200
rect 7432 11160 7438 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 2498 11132 2504 11144
rect 1535 11104 2504 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 8036 11064 8064 11095
rect 7524 11036 8064 11064
rect 7524 11024 7530 11036
rect 1104 10906 9936 10928
rect 1104 10854 2950 10906
rect 3002 10854 3014 10906
rect 3066 10854 3078 10906
rect 3130 10854 3142 10906
rect 3194 10854 3206 10906
rect 3258 10854 4550 10906
rect 4602 10854 4614 10906
rect 4666 10854 4678 10906
rect 4730 10854 4742 10906
rect 4794 10854 4806 10906
rect 4858 10854 6150 10906
rect 6202 10854 6214 10906
rect 6266 10854 6278 10906
rect 6330 10854 6342 10906
rect 6394 10854 6406 10906
rect 6458 10854 7750 10906
rect 7802 10854 7814 10906
rect 7866 10854 7878 10906
rect 7930 10854 7942 10906
rect 7994 10854 8006 10906
rect 8058 10854 9350 10906
rect 9402 10854 9414 10906
rect 9466 10854 9478 10906
rect 9530 10854 9542 10906
rect 9594 10854 9606 10906
rect 9658 10854 9936 10906
rect 1104 10832 9936 10854
rect 1489 10727 1547 10733
rect 1489 10693 1501 10727
rect 1535 10724 1547 10727
rect 2222 10724 2228 10736
rect 1535 10696 2228 10724
rect 1535 10693 1547 10696
rect 1489 10687 1547 10693
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 992 10424 1593 10452
rect 992 10412 998 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 1104 10362 9936 10384
rect 1104 10310 3610 10362
rect 3662 10310 3674 10362
rect 3726 10310 3738 10362
rect 3790 10310 3802 10362
rect 3854 10310 3866 10362
rect 3918 10310 5210 10362
rect 5262 10310 5274 10362
rect 5326 10310 5338 10362
rect 5390 10310 5402 10362
rect 5454 10310 5466 10362
rect 5518 10310 6810 10362
rect 6862 10310 6874 10362
rect 6926 10310 6938 10362
rect 6990 10310 7002 10362
rect 7054 10310 7066 10362
rect 7118 10310 8410 10362
rect 8462 10310 8474 10362
rect 8526 10310 8538 10362
rect 8590 10310 8602 10362
rect 8654 10310 8666 10362
rect 8718 10310 9936 10362
rect 1104 10288 9936 10310
rect 1104 9818 9936 9840
rect 1104 9766 2950 9818
rect 3002 9766 3014 9818
rect 3066 9766 3078 9818
rect 3130 9766 3142 9818
rect 3194 9766 3206 9818
rect 3258 9766 4550 9818
rect 4602 9766 4614 9818
rect 4666 9766 4678 9818
rect 4730 9766 4742 9818
rect 4794 9766 4806 9818
rect 4858 9766 6150 9818
rect 6202 9766 6214 9818
rect 6266 9766 6278 9818
rect 6330 9766 6342 9818
rect 6394 9766 6406 9818
rect 6458 9766 7750 9818
rect 7802 9766 7814 9818
rect 7866 9766 7878 9818
rect 7930 9766 7942 9818
rect 7994 9766 8006 9818
rect 8058 9766 9350 9818
rect 9402 9766 9414 9818
rect 9466 9766 9478 9818
rect 9530 9766 9542 9818
rect 9594 9766 9606 9818
rect 9658 9766 9936 9818
rect 1104 9744 9936 9766
rect 1489 9639 1547 9645
rect 1489 9605 1501 9639
rect 1535 9636 1547 9639
rect 4154 9636 4160 9648
rect 1535 9608 4160 9636
rect 1535 9605 1547 9608
rect 1489 9599 1547 9605
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 7432 9472 8585 9500
rect 7432 9460 7438 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 992 9336 1593 9364
rect 992 9324 998 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 8260 9336 9597 9364
rect 8260 9324 8266 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 1104 9274 9936 9296
rect 1104 9222 3610 9274
rect 3662 9222 3674 9274
rect 3726 9222 3738 9274
rect 3790 9222 3802 9274
rect 3854 9222 3866 9274
rect 3918 9222 5210 9274
rect 5262 9222 5274 9274
rect 5326 9222 5338 9274
rect 5390 9222 5402 9274
rect 5454 9222 5466 9274
rect 5518 9222 6810 9274
rect 6862 9222 6874 9274
rect 6926 9222 6938 9274
rect 6990 9222 7002 9274
rect 7054 9222 7066 9274
rect 7118 9222 8410 9274
rect 8462 9222 8474 9274
rect 8526 9222 8538 9274
rect 8590 9222 8602 9274
rect 8654 9222 8666 9274
rect 8718 9222 9936 9274
rect 1104 9200 9936 9222
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 9582 8956 9588 8968
rect 8352 8928 9588 8956
rect 8352 8916 8358 8928
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 1104 8730 9936 8752
rect 1104 8678 2950 8730
rect 3002 8678 3014 8730
rect 3066 8678 3078 8730
rect 3130 8678 3142 8730
rect 3194 8678 3206 8730
rect 3258 8678 4550 8730
rect 4602 8678 4614 8730
rect 4666 8678 4678 8730
rect 4730 8678 4742 8730
rect 4794 8678 4806 8730
rect 4858 8678 6150 8730
rect 6202 8678 6214 8730
rect 6266 8678 6278 8730
rect 6330 8678 6342 8730
rect 6394 8678 6406 8730
rect 6458 8678 7750 8730
rect 7802 8678 7814 8730
rect 7866 8678 7878 8730
rect 7930 8678 7942 8730
rect 7994 8678 8006 8730
rect 8058 8678 9350 8730
rect 9402 8678 9414 8730
rect 9466 8678 9478 8730
rect 9530 8678 9542 8730
rect 9594 8678 9606 8730
rect 9658 8678 9936 8730
rect 1104 8656 9936 8678
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 1762 8548 1768 8560
rect 1535 8520 1768 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 1673 8347 1731 8353
rect 1673 8344 1685 8347
rect 1452 8316 1685 8344
rect 1452 8304 1458 8316
rect 1673 8313 1685 8316
rect 1719 8313 1731 8347
rect 1673 8307 1731 8313
rect 1104 8186 9936 8208
rect 1104 8134 3610 8186
rect 3662 8134 3674 8186
rect 3726 8134 3738 8186
rect 3790 8134 3802 8186
rect 3854 8134 3866 8186
rect 3918 8134 5210 8186
rect 5262 8134 5274 8186
rect 5326 8134 5338 8186
rect 5390 8134 5402 8186
rect 5454 8134 5466 8186
rect 5518 8134 6810 8186
rect 6862 8134 6874 8186
rect 6926 8134 6938 8186
rect 6990 8134 7002 8186
rect 7054 8134 7066 8186
rect 7118 8134 8410 8186
rect 8462 8134 8474 8186
rect 8526 8134 8538 8186
rect 8590 8134 8602 8186
rect 8654 8134 8666 8186
rect 8718 8134 9936 8186
rect 1104 8112 9936 8134
rect 1104 7642 9936 7664
rect 1104 7590 2950 7642
rect 3002 7590 3014 7642
rect 3066 7590 3078 7642
rect 3130 7590 3142 7642
rect 3194 7590 3206 7642
rect 3258 7590 4550 7642
rect 4602 7590 4614 7642
rect 4666 7590 4678 7642
rect 4730 7590 4742 7642
rect 4794 7590 4806 7642
rect 4858 7590 6150 7642
rect 6202 7590 6214 7642
rect 6266 7590 6278 7642
rect 6330 7590 6342 7642
rect 6394 7590 6406 7642
rect 6458 7590 7750 7642
rect 7802 7590 7814 7642
rect 7866 7590 7878 7642
rect 7930 7590 7942 7642
rect 7994 7590 8006 7642
rect 8058 7590 9350 7642
rect 9402 7590 9414 7642
rect 9466 7590 9478 7642
rect 9530 7590 9542 7642
rect 9594 7590 9606 7642
rect 9658 7590 9936 7642
rect 1104 7568 9936 7590
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7460 1547 7463
rect 3326 7460 3332 7472
rect 1535 7432 3332 7460
rect 1535 7429 1547 7432
rect 1489 7423 1547 7429
rect 3326 7420 3332 7432
rect 3384 7420 3390 7472
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 992 7160 1593 7188
rect 992 7148 998 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 1581 7151 1639 7157
rect 1104 7098 9936 7120
rect 1104 7046 3610 7098
rect 3662 7046 3674 7098
rect 3726 7046 3738 7098
rect 3790 7046 3802 7098
rect 3854 7046 3866 7098
rect 3918 7046 5210 7098
rect 5262 7046 5274 7098
rect 5326 7046 5338 7098
rect 5390 7046 5402 7098
rect 5454 7046 5466 7098
rect 5518 7046 6810 7098
rect 6862 7046 6874 7098
rect 6926 7046 6938 7098
rect 6990 7046 7002 7098
rect 7054 7046 7066 7098
rect 7118 7046 8410 7098
rect 8462 7046 8474 7098
rect 8526 7046 8538 7098
rect 8590 7046 8602 7098
rect 8654 7046 8666 7098
rect 8718 7046 9936 7098
rect 1104 7024 9936 7046
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 2130 6780 2136 6792
rect 1535 6752 2136 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 934 6604 940 6656
rect 992 6644 998 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 992 6616 1593 6644
rect 992 6604 998 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 1104 6554 9936 6576
rect 1104 6502 2950 6554
rect 3002 6502 3014 6554
rect 3066 6502 3078 6554
rect 3130 6502 3142 6554
rect 3194 6502 3206 6554
rect 3258 6502 4550 6554
rect 4602 6502 4614 6554
rect 4666 6502 4678 6554
rect 4730 6502 4742 6554
rect 4794 6502 4806 6554
rect 4858 6502 6150 6554
rect 6202 6502 6214 6554
rect 6266 6502 6278 6554
rect 6330 6502 6342 6554
rect 6394 6502 6406 6554
rect 6458 6502 7750 6554
rect 7802 6502 7814 6554
rect 7866 6502 7878 6554
rect 7930 6502 7942 6554
rect 7994 6502 8006 6554
rect 8058 6502 9350 6554
rect 9402 6502 9414 6554
rect 9466 6502 9478 6554
rect 9530 6502 9542 6554
rect 9594 6502 9606 6554
rect 9658 6502 9936 6554
rect 1104 6480 9936 6502
rect 1104 6010 9936 6032
rect 1104 5958 3610 6010
rect 3662 5958 3674 6010
rect 3726 5958 3738 6010
rect 3790 5958 3802 6010
rect 3854 5958 3866 6010
rect 3918 5958 5210 6010
rect 5262 5958 5274 6010
rect 5326 5958 5338 6010
rect 5390 5958 5402 6010
rect 5454 5958 5466 6010
rect 5518 5958 6810 6010
rect 6862 5958 6874 6010
rect 6926 5958 6938 6010
rect 6990 5958 7002 6010
rect 7054 5958 7066 6010
rect 7118 5958 8410 6010
rect 8462 5958 8474 6010
rect 8526 5958 8538 6010
rect 8590 5958 8602 6010
rect 8654 5958 8666 6010
rect 8718 5958 9936 6010
rect 1104 5936 9936 5958
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5692 1547 5695
rect 3970 5692 3976 5704
rect 1535 5664 3976 5692
rect 1535 5661 1547 5664
rect 1489 5655 1547 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 1104 5466 9936 5488
rect 1104 5414 2950 5466
rect 3002 5414 3014 5466
rect 3066 5414 3078 5466
rect 3130 5414 3142 5466
rect 3194 5414 3206 5466
rect 3258 5414 4550 5466
rect 4602 5414 4614 5466
rect 4666 5414 4678 5466
rect 4730 5414 4742 5466
rect 4794 5414 4806 5466
rect 4858 5414 6150 5466
rect 6202 5414 6214 5466
rect 6266 5414 6278 5466
rect 6330 5414 6342 5466
rect 6394 5414 6406 5466
rect 6458 5414 7750 5466
rect 7802 5414 7814 5466
rect 7866 5414 7878 5466
rect 7930 5414 7942 5466
rect 7994 5414 8006 5466
rect 8058 5414 9350 5466
rect 9402 5414 9414 5466
rect 9466 5414 9478 5466
rect 9530 5414 9542 5466
rect 9594 5414 9606 5466
rect 9658 5414 9936 5466
rect 1104 5392 9936 5414
rect 1104 4922 9936 4944
rect 1104 4870 3610 4922
rect 3662 4870 3674 4922
rect 3726 4870 3738 4922
rect 3790 4870 3802 4922
rect 3854 4870 3866 4922
rect 3918 4870 5210 4922
rect 5262 4870 5274 4922
rect 5326 4870 5338 4922
rect 5390 4870 5402 4922
rect 5454 4870 5466 4922
rect 5518 4870 6810 4922
rect 6862 4870 6874 4922
rect 6926 4870 6938 4922
rect 6990 4870 7002 4922
rect 7054 4870 7066 4922
rect 7118 4870 8410 4922
rect 8462 4870 8474 4922
rect 8526 4870 8538 4922
rect 8590 4870 8602 4922
rect 8654 4870 8666 4922
rect 8718 4870 9936 4922
rect 1104 4848 9936 4870
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 4246 4604 4252 4616
rect 1535 4576 4252 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 934 4428 940 4480
rect 992 4468 998 4480
rect 1581 4471 1639 4477
rect 1581 4468 1593 4471
rect 992 4440 1593 4468
rect 992 4428 998 4440
rect 1581 4437 1593 4440
rect 1627 4437 1639 4471
rect 1581 4431 1639 4437
rect 1104 4378 9936 4400
rect 1104 4326 2950 4378
rect 3002 4326 3014 4378
rect 3066 4326 3078 4378
rect 3130 4326 3142 4378
rect 3194 4326 3206 4378
rect 3258 4326 4550 4378
rect 4602 4326 4614 4378
rect 4666 4326 4678 4378
rect 4730 4326 4742 4378
rect 4794 4326 4806 4378
rect 4858 4326 6150 4378
rect 6202 4326 6214 4378
rect 6266 4326 6278 4378
rect 6330 4326 6342 4378
rect 6394 4326 6406 4378
rect 6458 4326 7750 4378
rect 7802 4326 7814 4378
rect 7866 4326 7878 4378
rect 7930 4326 7942 4378
rect 7994 4326 8006 4378
rect 8058 4326 9350 4378
rect 9402 4326 9414 4378
rect 9466 4326 9478 4378
rect 9530 4326 9542 4378
rect 9594 4326 9606 4378
rect 9658 4326 9936 4378
rect 1104 4304 9936 4326
rect 11698 3952 11704 4004
rect 11756 3992 11762 4004
rect 17862 3992 17868 4004
rect 11756 3964 17868 3992
rect 11756 3952 11762 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 54386 3924 54392 3936
rect 9088 3896 54392 3924
rect 9088 3884 9094 3896
rect 54386 3884 54392 3896
rect 54444 3884 54450 3936
rect 1104 3834 9936 3856
rect 1104 3782 3610 3834
rect 3662 3782 3674 3834
rect 3726 3782 3738 3834
rect 3790 3782 3802 3834
rect 3854 3782 3866 3834
rect 3918 3782 5210 3834
rect 5262 3782 5274 3834
rect 5326 3782 5338 3834
rect 5390 3782 5402 3834
rect 5454 3782 5466 3834
rect 5518 3782 6810 3834
rect 6862 3782 6874 3834
rect 6926 3782 6938 3834
rect 6990 3782 7002 3834
rect 7054 3782 7066 3834
rect 7118 3782 8410 3834
rect 8462 3782 8474 3834
rect 8526 3782 8538 3834
rect 8590 3782 8602 3834
rect 8654 3782 8666 3834
rect 8718 3782 9936 3834
rect 11422 3816 11428 3868
rect 11480 3856 11486 3868
rect 46106 3856 46112 3868
rect 11480 3828 46112 3856
rect 11480 3816 11486 3828
rect 46106 3816 46112 3828
rect 46164 3816 46170 3868
rect 1104 3760 9936 3782
rect 10778 3748 10784 3800
rect 10836 3788 10842 3800
rect 40310 3788 40316 3800
rect 10836 3760 40316 3788
rect 10836 3748 10842 3760
rect 40310 3748 40316 3760
rect 40368 3748 40374 3800
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 50890 3720 50896 3732
rect 9180 3692 50896 3720
rect 9180 3680 9186 3692
rect 50890 3680 50896 3692
rect 50948 3680 50954 3732
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 45002 3652 45008 3664
rect 7616 3624 45008 3652
rect 7616 3612 7622 3624
rect 45002 3612 45008 3624
rect 45060 3612 45066 3664
rect 5074 3544 5080 3596
rect 5132 3584 5138 3596
rect 39206 3584 39212 3596
rect 5132 3556 39212 3584
rect 5132 3544 5138 3556
rect 39206 3544 39212 3556
rect 39264 3544 39270 3596
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2314 3516 2320 3528
rect 1535 3488 2320 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 29822 3516 29828 3528
rect 11020 3488 29828 3516
rect 11020 3476 11026 3488
rect 29822 3476 29828 3488
rect 29880 3476 29886 3528
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 54570 3448 54576 3460
rect 6696 3420 54576 3448
rect 6696 3408 6702 3420
rect 54570 3408 54576 3420
rect 54628 3408 54634 3460
rect 934 3340 940 3392
rect 992 3380 998 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 992 3352 1593 3380
rect 992 3340 998 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 28718 3380 28724 3392
rect 10284 3352 28724 3380
rect 10284 3340 10290 3352
rect 28718 3340 28724 3352
rect 28776 3340 28782 3392
rect 1104 3290 9936 3312
rect 1104 3238 2950 3290
rect 3002 3238 3014 3290
rect 3066 3238 3078 3290
rect 3130 3238 3142 3290
rect 3194 3238 3206 3290
rect 3258 3238 4550 3290
rect 4602 3238 4614 3290
rect 4666 3238 4678 3290
rect 4730 3238 4742 3290
rect 4794 3238 4806 3290
rect 4858 3238 6150 3290
rect 6202 3238 6214 3290
rect 6266 3238 6278 3290
rect 6330 3238 6342 3290
rect 6394 3238 6406 3290
rect 6458 3238 7750 3290
rect 7802 3238 7814 3290
rect 7866 3238 7878 3290
rect 7930 3238 7942 3290
rect 7994 3238 8006 3290
rect 8058 3238 9350 3290
rect 9402 3238 9414 3290
rect 9466 3238 9478 3290
rect 9530 3238 9542 3290
rect 9594 3238 9606 3290
rect 9658 3238 9936 3290
rect 10318 3272 10324 3324
rect 10376 3312 10382 3324
rect 32122 3312 32128 3324
rect 10376 3284 32128 3312
rect 10376 3272 10382 3284
rect 32122 3272 32128 3284
rect 32180 3272 32186 3324
rect 1104 3216 9936 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 47486 3176 47492 3188
rect 5868 3148 47492 3176
rect 5868 3136 5874 3148
rect 47486 3136 47492 3148
rect 47544 3136 47550 3188
rect 1104 2746 9936 2768
rect 1104 2694 3610 2746
rect 3662 2694 3674 2746
rect 3726 2694 3738 2746
rect 3790 2694 3802 2746
rect 3854 2694 3866 2746
rect 3918 2694 5210 2746
rect 5262 2694 5274 2746
rect 5326 2694 5338 2746
rect 5390 2694 5402 2746
rect 5454 2694 5466 2746
rect 5518 2694 6810 2746
rect 6862 2694 6874 2746
rect 6926 2694 6938 2746
rect 6990 2694 7002 2746
rect 7054 2694 7066 2746
rect 7118 2694 8410 2746
rect 8462 2694 8474 2746
rect 8526 2694 8538 2746
rect 8590 2694 8602 2746
rect 8654 2694 8666 2746
rect 8718 2694 9936 2746
rect 11882 2728 11888 2780
rect 11940 2768 11946 2780
rect 27522 2768 27528 2780
rect 11940 2740 27528 2768
rect 11940 2728 11946 2740
rect 27522 2728 27528 2740
rect 27580 2728 27586 2780
rect 1104 2672 9936 2694
rect 11790 2660 11796 2712
rect 11848 2700 11854 2712
rect 34698 2700 34704 2712
rect 11848 2672 34704 2700
rect 11848 2660 11854 2672
rect 34698 2660 34704 2672
rect 34756 2660 34762 2712
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 107930 2632 107936 2644
rect 6052 2604 107936 2632
rect 6052 2592 6058 2604
rect 107930 2592 107936 2604
rect 107988 2592 107994 2644
rect 8110 2524 8116 2576
rect 8168 2564 8174 2576
rect 32030 2564 32036 2576
rect 8168 2536 32036 2564
rect 8168 2524 8174 2536
rect 32030 2524 32036 2536
rect 32088 2524 32094 2576
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 43806 2496 43812 2508
rect 8996 2468 43812 2496
rect 8996 2456 9002 2468
rect 43806 2456 43812 2468
rect 43864 2456 43870 2508
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 55398 2428 55404 2440
rect 8812 2400 55404 2428
rect 8812 2388 8818 2400
rect 55398 2388 55404 2400
rect 55456 2388 55462 2440
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 57974 2360 57980 2372
rect 8352 2332 57980 2360
rect 8352 2320 8358 2332
rect 57974 2320 57980 2332
rect 58032 2320 58038 2372
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 49694 2292 49700 2304
rect 900 2264 49700 2292
rect 900 2252 906 2264
rect 49694 2252 49700 2264
rect 49752 2252 49758 2304
rect 1104 2202 9936 2224
rect 1104 2150 2950 2202
rect 3002 2150 3014 2202
rect 3066 2150 3078 2202
rect 3130 2150 3142 2202
rect 3194 2150 3206 2202
rect 3258 2150 4550 2202
rect 4602 2150 4614 2202
rect 4666 2150 4678 2202
rect 4730 2150 4742 2202
rect 4794 2150 4806 2202
rect 4858 2150 6150 2202
rect 6202 2150 6214 2202
rect 6266 2150 6278 2202
rect 6330 2150 6342 2202
rect 6394 2150 6406 2202
rect 6458 2150 7750 2202
rect 7802 2150 7814 2202
rect 7866 2150 7878 2202
rect 7930 2150 7942 2202
rect 7994 2150 8006 2202
rect 8058 2150 9350 2202
rect 9402 2150 9414 2202
rect 9466 2150 9478 2202
rect 9530 2150 9542 2202
rect 9594 2150 9606 2202
rect 9658 2150 9936 2202
rect 11606 2184 11612 2236
rect 11664 2224 11670 2236
rect 36998 2224 37004 2236
rect 11664 2196 37004 2224
rect 11664 2184 11670 2196
rect 36998 2184 37004 2196
rect 37056 2184 37062 2236
rect 1104 2128 9936 2150
rect 10870 2116 10876 2168
rect 10928 2156 10934 2168
rect 48590 2156 48596 2168
rect 10928 2128 48596 2156
rect 10928 2116 10934 2128
rect 48590 2116 48596 2128
rect 48648 2116 48654 2168
rect 6546 2048 6552 2100
rect 6604 2088 6610 2100
rect 94958 2088 94964 2100
rect 6604 2060 94964 2088
rect 6604 2048 6610 2060
rect 94958 2048 94964 2060
rect 95016 2048 95022 2100
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 42794 2020 42800 2032
rect 9272 1992 42800 2020
rect 9272 1980 9278 1992
rect 42794 1980 42800 1992
rect 42852 1980 42858 2032
rect 1104 1658 108836 1680
rect 1104 1606 3610 1658
rect 3662 1606 3674 1658
rect 3726 1606 3738 1658
rect 3790 1606 3802 1658
rect 3854 1606 3866 1658
rect 3918 1606 5210 1658
rect 5262 1606 5274 1658
rect 5326 1606 5338 1658
rect 5390 1606 5402 1658
rect 5454 1606 5466 1658
rect 5518 1606 6810 1658
rect 6862 1606 6874 1658
rect 6926 1606 6938 1658
rect 6990 1606 7002 1658
rect 7054 1606 7066 1658
rect 7118 1606 8410 1658
rect 8462 1606 8474 1658
rect 8526 1606 8538 1658
rect 8590 1606 8602 1658
rect 8654 1606 8666 1658
rect 8718 1606 10010 1658
rect 10062 1606 10074 1658
rect 10126 1606 10138 1658
rect 10190 1606 10202 1658
rect 10254 1606 10266 1658
rect 10318 1606 11610 1658
rect 11662 1606 11674 1658
rect 11726 1606 11738 1658
rect 11790 1606 11802 1658
rect 11854 1606 11866 1658
rect 11918 1606 13210 1658
rect 13262 1606 13274 1658
rect 13326 1606 13338 1658
rect 13390 1606 13402 1658
rect 13454 1606 13466 1658
rect 13518 1606 14810 1658
rect 14862 1606 14874 1658
rect 14926 1606 14938 1658
rect 14990 1606 15002 1658
rect 15054 1606 15066 1658
rect 15118 1606 16410 1658
rect 16462 1606 16474 1658
rect 16526 1606 16538 1658
rect 16590 1606 16602 1658
rect 16654 1606 16666 1658
rect 16718 1606 18010 1658
rect 18062 1606 18074 1658
rect 18126 1606 18138 1658
rect 18190 1606 18202 1658
rect 18254 1606 18266 1658
rect 18318 1606 19610 1658
rect 19662 1606 19674 1658
rect 19726 1606 19738 1658
rect 19790 1606 19802 1658
rect 19854 1606 19866 1658
rect 19918 1606 21210 1658
rect 21262 1606 21274 1658
rect 21326 1606 21338 1658
rect 21390 1606 21402 1658
rect 21454 1606 21466 1658
rect 21518 1606 22810 1658
rect 22862 1606 22874 1658
rect 22926 1606 22938 1658
rect 22990 1606 23002 1658
rect 23054 1606 23066 1658
rect 23118 1606 24410 1658
rect 24462 1606 24474 1658
rect 24526 1606 24538 1658
rect 24590 1606 24602 1658
rect 24654 1606 24666 1658
rect 24718 1606 26010 1658
rect 26062 1606 26074 1658
rect 26126 1606 26138 1658
rect 26190 1606 26202 1658
rect 26254 1606 26266 1658
rect 26318 1606 27610 1658
rect 27662 1606 27674 1658
rect 27726 1606 27738 1658
rect 27790 1606 27802 1658
rect 27854 1606 27866 1658
rect 27918 1606 29210 1658
rect 29262 1606 29274 1658
rect 29326 1606 29338 1658
rect 29390 1606 29402 1658
rect 29454 1606 29466 1658
rect 29518 1606 30810 1658
rect 30862 1606 30874 1658
rect 30926 1606 30938 1658
rect 30990 1606 31002 1658
rect 31054 1606 31066 1658
rect 31118 1606 32410 1658
rect 32462 1606 32474 1658
rect 32526 1606 32538 1658
rect 32590 1606 32602 1658
rect 32654 1606 32666 1658
rect 32718 1606 34010 1658
rect 34062 1606 34074 1658
rect 34126 1606 34138 1658
rect 34190 1606 34202 1658
rect 34254 1606 34266 1658
rect 34318 1606 35610 1658
rect 35662 1606 35674 1658
rect 35726 1606 35738 1658
rect 35790 1606 35802 1658
rect 35854 1606 35866 1658
rect 35918 1606 37210 1658
rect 37262 1606 37274 1658
rect 37326 1606 37338 1658
rect 37390 1606 37402 1658
rect 37454 1606 37466 1658
rect 37518 1606 38810 1658
rect 38862 1606 38874 1658
rect 38926 1606 38938 1658
rect 38990 1606 39002 1658
rect 39054 1606 39066 1658
rect 39118 1606 40410 1658
rect 40462 1606 40474 1658
rect 40526 1606 40538 1658
rect 40590 1606 40602 1658
rect 40654 1606 40666 1658
rect 40718 1606 42010 1658
rect 42062 1606 42074 1658
rect 42126 1606 42138 1658
rect 42190 1606 42202 1658
rect 42254 1606 42266 1658
rect 42318 1606 43610 1658
rect 43662 1606 43674 1658
rect 43726 1606 43738 1658
rect 43790 1606 43802 1658
rect 43854 1606 43866 1658
rect 43918 1606 45210 1658
rect 45262 1606 45274 1658
rect 45326 1606 45338 1658
rect 45390 1606 45402 1658
rect 45454 1606 45466 1658
rect 45518 1606 46810 1658
rect 46862 1606 46874 1658
rect 46926 1606 46938 1658
rect 46990 1606 47002 1658
rect 47054 1606 47066 1658
rect 47118 1606 48410 1658
rect 48462 1606 48474 1658
rect 48526 1606 48538 1658
rect 48590 1606 48602 1658
rect 48654 1606 48666 1658
rect 48718 1606 50010 1658
rect 50062 1606 50074 1658
rect 50126 1606 50138 1658
rect 50190 1606 50202 1658
rect 50254 1606 50266 1658
rect 50318 1606 51610 1658
rect 51662 1606 51674 1658
rect 51726 1606 51738 1658
rect 51790 1606 51802 1658
rect 51854 1606 51866 1658
rect 51918 1606 53210 1658
rect 53262 1606 53274 1658
rect 53326 1606 53338 1658
rect 53390 1606 53402 1658
rect 53454 1606 53466 1658
rect 53518 1606 54810 1658
rect 54862 1606 54874 1658
rect 54926 1606 54938 1658
rect 54990 1606 55002 1658
rect 55054 1606 55066 1658
rect 55118 1606 56410 1658
rect 56462 1606 56474 1658
rect 56526 1606 56538 1658
rect 56590 1606 56602 1658
rect 56654 1606 56666 1658
rect 56718 1606 58010 1658
rect 58062 1606 58074 1658
rect 58126 1606 58138 1658
rect 58190 1606 58202 1658
rect 58254 1606 58266 1658
rect 58318 1606 59610 1658
rect 59662 1606 59674 1658
rect 59726 1606 59738 1658
rect 59790 1606 59802 1658
rect 59854 1606 59866 1658
rect 59918 1606 61210 1658
rect 61262 1606 61274 1658
rect 61326 1606 61338 1658
rect 61390 1606 61402 1658
rect 61454 1606 61466 1658
rect 61518 1606 62810 1658
rect 62862 1606 62874 1658
rect 62926 1606 62938 1658
rect 62990 1606 63002 1658
rect 63054 1606 63066 1658
rect 63118 1606 64410 1658
rect 64462 1606 64474 1658
rect 64526 1606 64538 1658
rect 64590 1606 64602 1658
rect 64654 1606 64666 1658
rect 64718 1606 66010 1658
rect 66062 1606 66074 1658
rect 66126 1606 66138 1658
rect 66190 1606 66202 1658
rect 66254 1606 66266 1658
rect 66318 1606 67610 1658
rect 67662 1606 67674 1658
rect 67726 1606 67738 1658
rect 67790 1606 67802 1658
rect 67854 1606 67866 1658
rect 67918 1606 69210 1658
rect 69262 1606 69274 1658
rect 69326 1606 69338 1658
rect 69390 1606 69402 1658
rect 69454 1606 69466 1658
rect 69518 1606 70810 1658
rect 70862 1606 70874 1658
rect 70926 1606 70938 1658
rect 70990 1606 71002 1658
rect 71054 1606 71066 1658
rect 71118 1606 72410 1658
rect 72462 1606 72474 1658
rect 72526 1606 72538 1658
rect 72590 1606 72602 1658
rect 72654 1606 72666 1658
rect 72718 1606 74010 1658
rect 74062 1606 74074 1658
rect 74126 1606 74138 1658
rect 74190 1606 74202 1658
rect 74254 1606 74266 1658
rect 74318 1606 75610 1658
rect 75662 1606 75674 1658
rect 75726 1606 75738 1658
rect 75790 1606 75802 1658
rect 75854 1606 75866 1658
rect 75918 1606 77210 1658
rect 77262 1606 77274 1658
rect 77326 1606 77338 1658
rect 77390 1606 77402 1658
rect 77454 1606 77466 1658
rect 77518 1606 78810 1658
rect 78862 1606 78874 1658
rect 78926 1606 78938 1658
rect 78990 1606 79002 1658
rect 79054 1606 79066 1658
rect 79118 1606 80410 1658
rect 80462 1606 80474 1658
rect 80526 1606 80538 1658
rect 80590 1606 80602 1658
rect 80654 1606 80666 1658
rect 80718 1606 82010 1658
rect 82062 1606 82074 1658
rect 82126 1606 82138 1658
rect 82190 1606 82202 1658
rect 82254 1606 82266 1658
rect 82318 1606 83610 1658
rect 83662 1606 83674 1658
rect 83726 1606 83738 1658
rect 83790 1606 83802 1658
rect 83854 1606 83866 1658
rect 83918 1606 85210 1658
rect 85262 1606 85274 1658
rect 85326 1606 85338 1658
rect 85390 1606 85402 1658
rect 85454 1606 85466 1658
rect 85518 1606 86810 1658
rect 86862 1606 86874 1658
rect 86926 1606 86938 1658
rect 86990 1606 87002 1658
rect 87054 1606 87066 1658
rect 87118 1606 88410 1658
rect 88462 1606 88474 1658
rect 88526 1606 88538 1658
rect 88590 1606 88602 1658
rect 88654 1606 88666 1658
rect 88718 1606 90010 1658
rect 90062 1606 90074 1658
rect 90126 1606 90138 1658
rect 90190 1606 90202 1658
rect 90254 1606 90266 1658
rect 90318 1606 91610 1658
rect 91662 1606 91674 1658
rect 91726 1606 91738 1658
rect 91790 1606 91802 1658
rect 91854 1606 91866 1658
rect 91918 1606 93210 1658
rect 93262 1606 93274 1658
rect 93326 1606 93338 1658
rect 93390 1606 93402 1658
rect 93454 1606 93466 1658
rect 93518 1606 94810 1658
rect 94862 1606 94874 1658
rect 94926 1606 94938 1658
rect 94990 1606 95002 1658
rect 95054 1606 95066 1658
rect 95118 1606 96410 1658
rect 96462 1606 96474 1658
rect 96526 1606 96538 1658
rect 96590 1606 96602 1658
rect 96654 1606 96666 1658
rect 96718 1606 98010 1658
rect 98062 1606 98074 1658
rect 98126 1606 98138 1658
rect 98190 1606 98202 1658
rect 98254 1606 98266 1658
rect 98318 1606 99610 1658
rect 99662 1606 99674 1658
rect 99726 1606 99738 1658
rect 99790 1606 99802 1658
rect 99854 1606 99866 1658
rect 99918 1606 101210 1658
rect 101262 1606 101274 1658
rect 101326 1606 101338 1658
rect 101390 1606 101402 1658
rect 101454 1606 101466 1658
rect 101518 1606 102810 1658
rect 102862 1606 102874 1658
rect 102926 1606 102938 1658
rect 102990 1606 103002 1658
rect 103054 1606 103066 1658
rect 103118 1606 104410 1658
rect 104462 1606 104474 1658
rect 104526 1606 104538 1658
rect 104590 1606 104602 1658
rect 104654 1606 104666 1658
rect 104718 1606 106010 1658
rect 106062 1606 106074 1658
rect 106126 1606 106138 1658
rect 106190 1606 106202 1658
rect 106254 1606 106266 1658
rect 106318 1606 107610 1658
rect 107662 1606 107674 1658
rect 107726 1606 107738 1658
rect 107790 1606 107802 1658
rect 107854 1606 107866 1658
rect 107918 1606 108836 1658
rect 1104 1584 108836 1606
rect 23658 1436 23664 1488
rect 23716 1476 23722 1488
rect 23716 1448 28488 1476
rect 23716 1436 23722 1448
rect 17236 1380 17632 1408
rect 11514 1300 11520 1352
rect 11572 1340 11578 1352
rect 17236 1340 17264 1380
rect 11572 1312 17264 1340
rect 11572 1300 11578 1312
rect 1026 1232 1032 1284
rect 1084 1272 1090 1284
rect 17604 1272 17632 1380
rect 23198 1368 23204 1420
rect 23256 1408 23262 1420
rect 23256 1380 27108 1408
rect 23256 1368 23262 1380
rect 22833 1343 22891 1349
rect 22833 1340 22845 1343
rect 22066 1312 22845 1340
rect 22066 1272 22094 1312
rect 22833 1309 22845 1312
rect 22879 1309 22891 1343
rect 22833 1303 22891 1309
rect 24118 1300 24124 1352
rect 24176 1340 24182 1352
rect 26145 1343 26203 1349
rect 26145 1340 26157 1343
rect 24176 1312 26157 1340
rect 24176 1300 24182 1312
rect 26145 1309 26157 1312
rect 26191 1309 26203 1343
rect 26145 1303 26203 1309
rect 23201 1275 23259 1281
rect 23201 1272 23213 1275
rect 1084 1244 17356 1272
rect 17604 1244 22094 1272
rect 22848 1244 23213 1272
rect 1084 1232 1090 1244
rect 1118 1164 1124 1216
rect 1176 1204 1182 1216
rect 17218 1204 17224 1216
rect 1176 1176 17224 1204
rect 1176 1164 1182 1176
rect 17218 1164 17224 1176
rect 17276 1164 17282 1216
rect 17328 1204 17356 1244
rect 22848 1204 22876 1244
rect 23201 1241 23213 1244
rect 23247 1241 23259 1275
rect 23201 1235 23259 1241
rect 23385 1275 23443 1281
rect 23385 1241 23397 1275
rect 23431 1241 23443 1275
rect 23385 1235 23443 1241
rect 17328 1176 22876 1204
rect 22922 1164 22928 1216
rect 22980 1164 22986 1216
rect 23400 1204 23428 1235
rect 23474 1232 23480 1284
rect 23532 1272 23538 1284
rect 27080 1281 27108 1380
rect 27522 1368 27528 1420
rect 27580 1368 27586 1420
rect 27798 1300 27804 1352
rect 27856 1300 27862 1352
rect 28460 1349 28488 1448
rect 34698 1368 34704 1420
rect 34756 1408 34762 1420
rect 35805 1411 35863 1417
rect 35805 1408 35817 1411
rect 34756 1380 35817 1408
rect 34756 1368 34762 1380
rect 35805 1377 35817 1380
rect 35851 1377 35863 1411
rect 35805 1371 35863 1377
rect 28445 1343 28503 1349
rect 28445 1309 28457 1343
rect 28491 1309 28503 1343
rect 28445 1303 28503 1309
rect 29638 1300 29644 1352
rect 29696 1300 29702 1352
rect 30484 1312 31754 1340
rect 24489 1275 24547 1281
rect 24489 1272 24501 1275
rect 23532 1244 24501 1272
rect 23532 1232 23538 1244
rect 24489 1241 24501 1244
rect 24535 1241 24547 1275
rect 24489 1235 24547 1241
rect 24673 1275 24731 1281
rect 24673 1241 24685 1275
rect 24719 1272 24731 1275
rect 27065 1275 27123 1281
rect 24719 1244 27016 1272
rect 24719 1241 24731 1244
rect 24673 1235 24731 1241
rect 26234 1204 26240 1216
rect 23400 1176 26240 1204
rect 26234 1164 26240 1176
rect 26292 1164 26298 1216
rect 26326 1164 26332 1216
rect 26384 1164 26390 1216
rect 26988 1204 27016 1244
rect 27065 1241 27077 1275
rect 27111 1241 27123 1275
rect 27065 1235 27123 1241
rect 27249 1275 27307 1281
rect 27249 1241 27261 1275
rect 27295 1272 27307 1275
rect 27338 1272 27344 1284
rect 27295 1244 27344 1272
rect 27295 1241 27307 1244
rect 27249 1235 27307 1241
rect 27338 1232 27344 1244
rect 27396 1232 27402 1284
rect 30484 1272 30512 1312
rect 27448 1244 30512 1272
rect 30561 1275 30619 1281
rect 27448 1204 27476 1244
rect 30561 1241 30573 1275
rect 30607 1241 30619 1275
rect 31726 1272 31754 1312
rect 32122 1300 32128 1352
rect 32180 1300 32186 1352
rect 32398 1300 32404 1352
rect 32456 1300 32462 1352
rect 33134 1300 33140 1352
rect 33192 1340 33198 1352
rect 33597 1343 33655 1349
rect 33597 1340 33609 1343
rect 33192 1312 33609 1340
rect 33192 1300 33198 1312
rect 33597 1309 33609 1312
rect 33643 1309 33655 1343
rect 33597 1303 33655 1309
rect 33870 1300 33876 1352
rect 33928 1300 33934 1352
rect 34977 1343 35035 1349
rect 34977 1309 34989 1343
rect 35023 1340 35035 1343
rect 37366 1340 37372 1352
rect 35023 1312 37372 1340
rect 35023 1309 35035 1312
rect 34977 1303 35035 1309
rect 37366 1300 37372 1312
rect 37424 1300 37430 1352
rect 37461 1343 37519 1349
rect 37461 1309 37473 1343
rect 37507 1340 37519 1343
rect 37550 1340 37556 1352
rect 37507 1312 37556 1340
rect 37507 1309 37519 1312
rect 37461 1303 37519 1309
rect 37550 1300 37556 1312
rect 37608 1300 37614 1352
rect 37734 1300 37740 1352
rect 37792 1300 37798 1352
rect 59354 1272 59360 1284
rect 31726 1244 59360 1272
rect 30561 1235 30619 1241
rect 26988 1176 27476 1204
rect 28629 1207 28687 1213
rect 28629 1173 28641 1207
rect 28675 1204 28687 1207
rect 29454 1204 29460 1216
rect 28675 1176 29460 1204
rect 28675 1173 28687 1176
rect 28629 1167 28687 1173
rect 29454 1164 29460 1176
rect 29512 1164 29518 1216
rect 29730 1164 29736 1216
rect 29788 1164 29794 1216
rect 29822 1164 29828 1216
rect 29880 1204 29886 1216
rect 30101 1207 30159 1213
rect 30101 1204 30113 1207
rect 29880 1176 30113 1204
rect 29880 1164 29886 1176
rect 30101 1173 30113 1176
rect 30147 1204 30159 1207
rect 30576 1204 30604 1235
rect 59354 1232 59360 1244
rect 59412 1232 59418 1284
rect 30147 1176 30604 1204
rect 30147 1173 30159 1176
rect 30101 1167 30159 1173
rect 30650 1164 30656 1216
rect 30708 1164 30714 1216
rect 32306 1164 32312 1216
rect 32364 1204 32370 1216
rect 37274 1204 37280 1216
rect 32364 1176 37280 1204
rect 32364 1164 32370 1176
rect 37274 1164 37280 1176
rect 37332 1164 37338 1216
rect 37550 1164 37556 1216
rect 37608 1204 37614 1216
rect 38565 1207 38623 1213
rect 38565 1204 38577 1207
rect 37608 1176 38577 1204
rect 37608 1164 37614 1176
rect 38565 1173 38577 1176
rect 38611 1173 38623 1207
rect 38565 1167 38623 1173
rect 1104 1114 108864 1136
rect 1104 1062 2950 1114
rect 3002 1062 3014 1114
rect 3066 1062 3078 1114
rect 3130 1062 3142 1114
rect 3194 1062 3206 1114
rect 3258 1062 4550 1114
rect 4602 1062 4614 1114
rect 4666 1062 4678 1114
rect 4730 1062 4742 1114
rect 4794 1062 4806 1114
rect 4858 1062 6150 1114
rect 6202 1062 6214 1114
rect 6266 1062 6278 1114
rect 6330 1062 6342 1114
rect 6394 1062 6406 1114
rect 6458 1062 7750 1114
rect 7802 1062 7814 1114
rect 7866 1062 7878 1114
rect 7930 1062 7942 1114
rect 7994 1062 8006 1114
rect 8058 1062 9350 1114
rect 9402 1062 9414 1114
rect 9466 1062 9478 1114
rect 9530 1062 9542 1114
rect 9594 1062 9606 1114
rect 9658 1062 10950 1114
rect 11002 1062 11014 1114
rect 11066 1062 11078 1114
rect 11130 1062 11142 1114
rect 11194 1062 11206 1114
rect 11258 1062 12550 1114
rect 12602 1062 12614 1114
rect 12666 1062 12678 1114
rect 12730 1062 12742 1114
rect 12794 1062 12806 1114
rect 12858 1062 14150 1114
rect 14202 1062 14214 1114
rect 14266 1062 14278 1114
rect 14330 1062 14342 1114
rect 14394 1062 14406 1114
rect 14458 1062 15750 1114
rect 15802 1062 15814 1114
rect 15866 1062 15878 1114
rect 15930 1062 15942 1114
rect 15994 1062 16006 1114
rect 16058 1062 17350 1114
rect 17402 1062 17414 1114
rect 17466 1062 17478 1114
rect 17530 1062 17542 1114
rect 17594 1062 17606 1114
rect 17658 1062 18950 1114
rect 19002 1062 19014 1114
rect 19066 1062 19078 1114
rect 19130 1062 19142 1114
rect 19194 1062 19206 1114
rect 19258 1062 20550 1114
rect 20602 1062 20614 1114
rect 20666 1062 20678 1114
rect 20730 1062 20742 1114
rect 20794 1062 20806 1114
rect 20858 1062 22150 1114
rect 22202 1062 22214 1114
rect 22266 1062 22278 1114
rect 22330 1062 22342 1114
rect 22394 1062 22406 1114
rect 22458 1062 23750 1114
rect 23802 1062 23814 1114
rect 23866 1062 23878 1114
rect 23930 1062 23942 1114
rect 23994 1062 24006 1114
rect 24058 1062 25350 1114
rect 25402 1062 25414 1114
rect 25466 1062 25478 1114
rect 25530 1062 25542 1114
rect 25594 1062 25606 1114
rect 25658 1062 26950 1114
rect 27002 1062 27014 1114
rect 27066 1062 27078 1114
rect 27130 1062 27142 1114
rect 27194 1062 27206 1114
rect 27258 1062 28550 1114
rect 28602 1062 28614 1114
rect 28666 1062 28678 1114
rect 28730 1062 28742 1114
rect 28794 1062 28806 1114
rect 28858 1062 30150 1114
rect 30202 1062 30214 1114
rect 30266 1062 30278 1114
rect 30330 1062 30342 1114
rect 30394 1062 30406 1114
rect 30458 1062 31750 1114
rect 31802 1062 31814 1114
rect 31866 1062 31878 1114
rect 31930 1062 31942 1114
rect 31994 1062 32006 1114
rect 32058 1062 33350 1114
rect 33402 1062 33414 1114
rect 33466 1062 33478 1114
rect 33530 1062 33542 1114
rect 33594 1062 33606 1114
rect 33658 1062 34950 1114
rect 35002 1062 35014 1114
rect 35066 1062 35078 1114
rect 35130 1062 35142 1114
rect 35194 1062 35206 1114
rect 35258 1062 36550 1114
rect 36602 1062 36614 1114
rect 36666 1062 36678 1114
rect 36730 1062 36742 1114
rect 36794 1062 36806 1114
rect 36858 1062 38150 1114
rect 38202 1062 38214 1114
rect 38266 1062 38278 1114
rect 38330 1062 38342 1114
rect 38394 1062 38406 1114
rect 38458 1062 39750 1114
rect 39802 1062 39814 1114
rect 39866 1062 39878 1114
rect 39930 1062 39942 1114
rect 39994 1062 40006 1114
rect 40058 1062 41350 1114
rect 41402 1062 41414 1114
rect 41466 1062 41478 1114
rect 41530 1062 41542 1114
rect 41594 1062 41606 1114
rect 41658 1062 42950 1114
rect 43002 1062 43014 1114
rect 43066 1062 43078 1114
rect 43130 1062 43142 1114
rect 43194 1062 43206 1114
rect 43258 1062 44550 1114
rect 44602 1062 44614 1114
rect 44666 1062 44678 1114
rect 44730 1062 44742 1114
rect 44794 1062 44806 1114
rect 44858 1062 46150 1114
rect 46202 1062 46214 1114
rect 46266 1062 46278 1114
rect 46330 1062 46342 1114
rect 46394 1062 46406 1114
rect 46458 1062 47750 1114
rect 47802 1062 47814 1114
rect 47866 1062 47878 1114
rect 47930 1062 47942 1114
rect 47994 1062 48006 1114
rect 48058 1062 49350 1114
rect 49402 1062 49414 1114
rect 49466 1062 49478 1114
rect 49530 1062 49542 1114
rect 49594 1062 49606 1114
rect 49658 1062 50950 1114
rect 51002 1062 51014 1114
rect 51066 1062 51078 1114
rect 51130 1062 51142 1114
rect 51194 1062 51206 1114
rect 51258 1062 52550 1114
rect 52602 1062 52614 1114
rect 52666 1062 52678 1114
rect 52730 1062 52742 1114
rect 52794 1062 52806 1114
rect 52858 1062 54150 1114
rect 54202 1062 54214 1114
rect 54266 1062 54278 1114
rect 54330 1062 54342 1114
rect 54394 1062 54406 1114
rect 54458 1062 55750 1114
rect 55802 1062 55814 1114
rect 55866 1062 55878 1114
rect 55930 1062 55942 1114
rect 55994 1062 56006 1114
rect 56058 1062 57350 1114
rect 57402 1062 57414 1114
rect 57466 1062 57478 1114
rect 57530 1062 57542 1114
rect 57594 1062 57606 1114
rect 57658 1062 58950 1114
rect 59002 1062 59014 1114
rect 59066 1062 59078 1114
rect 59130 1062 59142 1114
rect 59194 1062 59206 1114
rect 59258 1062 60550 1114
rect 60602 1062 60614 1114
rect 60666 1062 60678 1114
rect 60730 1062 60742 1114
rect 60794 1062 60806 1114
rect 60858 1062 62150 1114
rect 62202 1062 62214 1114
rect 62266 1062 62278 1114
rect 62330 1062 62342 1114
rect 62394 1062 62406 1114
rect 62458 1062 63750 1114
rect 63802 1062 63814 1114
rect 63866 1062 63878 1114
rect 63930 1062 63942 1114
rect 63994 1062 64006 1114
rect 64058 1062 65350 1114
rect 65402 1062 65414 1114
rect 65466 1062 65478 1114
rect 65530 1062 65542 1114
rect 65594 1062 65606 1114
rect 65658 1062 66950 1114
rect 67002 1062 67014 1114
rect 67066 1062 67078 1114
rect 67130 1062 67142 1114
rect 67194 1062 67206 1114
rect 67258 1062 68550 1114
rect 68602 1062 68614 1114
rect 68666 1062 68678 1114
rect 68730 1062 68742 1114
rect 68794 1062 68806 1114
rect 68858 1062 70150 1114
rect 70202 1062 70214 1114
rect 70266 1062 70278 1114
rect 70330 1062 70342 1114
rect 70394 1062 70406 1114
rect 70458 1062 71750 1114
rect 71802 1062 71814 1114
rect 71866 1062 71878 1114
rect 71930 1062 71942 1114
rect 71994 1062 72006 1114
rect 72058 1062 73350 1114
rect 73402 1062 73414 1114
rect 73466 1062 73478 1114
rect 73530 1062 73542 1114
rect 73594 1062 73606 1114
rect 73658 1062 74950 1114
rect 75002 1062 75014 1114
rect 75066 1062 75078 1114
rect 75130 1062 75142 1114
rect 75194 1062 75206 1114
rect 75258 1062 76550 1114
rect 76602 1062 76614 1114
rect 76666 1062 76678 1114
rect 76730 1062 76742 1114
rect 76794 1062 76806 1114
rect 76858 1062 78150 1114
rect 78202 1062 78214 1114
rect 78266 1062 78278 1114
rect 78330 1062 78342 1114
rect 78394 1062 78406 1114
rect 78458 1062 79750 1114
rect 79802 1062 79814 1114
rect 79866 1062 79878 1114
rect 79930 1062 79942 1114
rect 79994 1062 80006 1114
rect 80058 1062 81350 1114
rect 81402 1062 81414 1114
rect 81466 1062 81478 1114
rect 81530 1062 81542 1114
rect 81594 1062 81606 1114
rect 81658 1062 82950 1114
rect 83002 1062 83014 1114
rect 83066 1062 83078 1114
rect 83130 1062 83142 1114
rect 83194 1062 83206 1114
rect 83258 1062 84550 1114
rect 84602 1062 84614 1114
rect 84666 1062 84678 1114
rect 84730 1062 84742 1114
rect 84794 1062 84806 1114
rect 84858 1062 86150 1114
rect 86202 1062 86214 1114
rect 86266 1062 86278 1114
rect 86330 1062 86342 1114
rect 86394 1062 86406 1114
rect 86458 1062 87750 1114
rect 87802 1062 87814 1114
rect 87866 1062 87878 1114
rect 87930 1062 87942 1114
rect 87994 1062 88006 1114
rect 88058 1062 89350 1114
rect 89402 1062 89414 1114
rect 89466 1062 89478 1114
rect 89530 1062 89542 1114
rect 89594 1062 89606 1114
rect 89658 1062 90950 1114
rect 91002 1062 91014 1114
rect 91066 1062 91078 1114
rect 91130 1062 91142 1114
rect 91194 1062 91206 1114
rect 91258 1062 92550 1114
rect 92602 1062 92614 1114
rect 92666 1062 92678 1114
rect 92730 1062 92742 1114
rect 92794 1062 92806 1114
rect 92858 1062 94150 1114
rect 94202 1062 94214 1114
rect 94266 1062 94278 1114
rect 94330 1062 94342 1114
rect 94394 1062 94406 1114
rect 94458 1062 95750 1114
rect 95802 1062 95814 1114
rect 95866 1062 95878 1114
rect 95930 1062 95942 1114
rect 95994 1062 96006 1114
rect 96058 1062 97350 1114
rect 97402 1062 97414 1114
rect 97466 1062 97478 1114
rect 97530 1062 97542 1114
rect 97594 1062 97606 1114
rect 97658 1062 98950 1114
rect 99002 1062 99014 1114
rect 99066 1062 99078 1114
rect 99130 1062 99142 1114
rect 99194 1062 99206 1114
rect 99258 1062 100550 1114
rect 100602 1062 100614 1114
rect 100666 1062 100678 1114
rect 100730 1062 100742 1114
rect 100794 1062 100806 1114
rect 100858 1062 102150 1114
rect 102202 1062 102214 1114
rect 102266 1062 102278 1114
rect 102330 1062 102342 1114
rect 102394 1062 102406 1114
rect 102458 1062 103750 1114
rect 103802 1062 103814 1114
rect 103866 1062 103878 1114
rect 103930 1062 103942 1114
rect 103994 1062 104006 1114
rect 104058 1062 105350 1114
rect 105402 1062 105414 1114
rect 105466 1062 105478 1114
rect 105530 1062 105542 1114
rect 105594 1062 105606 1114
rect 105658 1062 106950 1114
rect 107002 1062 107014 1114
rect 107066 1062 107078 1114
rect 107130 1062 107142 1114
rect 107194 1062 107206 1114
rect 107258 1062 108550 1114
rect 108602 1062 108614 1114
rect 108666 1062 108678 1114
rect 108730 1062 108742 1114
rect 108794 1062 108806 1114
rect 108858 1062 108864 1114
rect 1104 1040 108864 1062
rect 5626 960 5632 1012
rect 5684 1000 5690 1012
rect 5684 972 12434 1000
rect 5684 960 5690 972
rect 12406 864 12434 972
rect 17218 960 17224 1012
rect 17276 1000 17282 1012
rect 17276 972 26096 1000
rect 17276 960 17282 972
rect 24118 932 24124 944
rect 22066 904 24124 932
rect 22066 864 22094 904
rect 24118 892 24124 904
rect 24176 892 24182 944
rect 12406 836 22094 864
rect 8202 756 8208 808
rect 8260 796 8266 808
rect 24394 796 24400 808
rect 8260 768 24400 796
rect 8260 756 8266 768
rect 24394 756 24400 768
rect 24452 756 24458 808
rect 26068 796 26096 972
rect 26234 960 26240 1012
rect 26292 1000 26298 1012
rect 26292 972 29592 1000
rect 26292 960 26298 972
rect 29564 864 29592 972
rect 29730 960 29736 1012
rect 29788 1000 29794 1012
rect 65150 1000 65156 1012
rect 29788 972 65156 1000
rect 29788 960 29794 972
rect 65150 960 65156 972
rect 65208 960 65214 1012
rect 33870 892 33876 944
rect 33928 932 33934 944
rect 67634 932 67640 944
rect 33928 904 67640 932
rect 33928 892 33934 904
rect 67634 892 67640 904
rect 67692 892 67698 944
rect 56594 864 56600 876
rect 29564 836 56600 864
rect 56594 824 56600 836
rect 56652 824 56658 876
rect 29546 796 29552 808
rect 26068 768 29552 796
rect 29546 756 29552 768
rect 29604 756 29610 808
rect 30650 756 30656 808
rect 30708 796 30714 808
rect 64874 796 64880 808
rect 30708 768 64880 796
rect 30708 756 30714 768
rect 64874 756 64880 768
rect 64932 756 64938 808
rect 11974 688 11980 740
rect 12032 728 12038 740
rect 23474 728 23480 740
rect 12032 700 23480 728
rect 12032 688 12038 700
rect 23474 688 23480 700
rect 23532 688 23538 740
rect 24504 700 28994 728
rect 10410 620 10416 672
rect 10468 660 10474 672
rect 24504 660 24532 700
rect 10468 632 24532 660
rect 28966 660 28994 700
rect 29454 688 29460 740
rect 29512 728 29518 740
rect 32214 728 32220 740
rect 29512 700 32220 728
rect 29512 688 29518 700
rect 32214 688 32220 700
rect 32272 688 32278 740
rect 32306 688 32312 740
rect 32364 688 32370 740
rect 60918 728 60924 740
rect 35866 700 60924 728
rect 32324 660 32352 688
rect 28966 632 32352 660
rect 10468 620 10474 632
rect 8846 552 8852 604
rect 8904 592 8910 604
rect 8904 564 24348 592
rect 8904 552 8910 564
rect 7650 484 7656 536
rect 7708 524 7714 536
rect 23658 524 23664 536
rect 7708 496 23664 524
rect 7708 484 7714 496
rect 23658 484 23664 496
rect 23716 484 23722 536
rect 10502 416 10508 468
rect 10560 456 10566 468
rect 23198 456 23204 468
rect 10560 428 23204 456
rect 10560 416 10566 428
rect 23198 416 23204 428
rect 23256 416 23262 468
rect 9858 280 9864 332
rect 9916 320 9922 332
rect 24320 320 24348 564
rect 27338 552 27344 604
rect 27396 552 27402 604
rect 27798 552 27804 604
rect 27856 592 27862 604
rect 35866 592 35894 700
rect 60918 688 60924 700
rect 60976 688 60982 740
rect 37734 620 37740 672
rect 37792 660 37798 672
rect 69014 660 69020 672
rect 37792 632 69020 660
rect 37792 620 37798 632
rect 69014 620 69020 632
rect 69072 620 69078 672
rect 27856 564 35894 592
rect 27856 552 27862 564
rect 37366 552 37372 604
rect 37424 592 37430 604
rect 66254 592 66260 604
rect 37424 564 66260 592
rect 37424 552 37430 564
rect 66254 552 66260 564
rect 66312 552 66318 604
rect 27356 388 27384 552
rect 32398 484 32404 536
rect 32456 524 32462 536
rect 62482 524 62488 536
rect 32456 496 62488 524
rect 32456 484 32462 496
rect 62482 484 62488 496
rect 62540 484 62546 536
rect 63494 388 63500 400
rect 27356 360 63500 388
rect 63494 348 63500 360
rect 63552 348 63558 400
rect 33226 320 33232 332
rect 9916 292 22094 320
rect 24320 292 33232 320
rect 9916 280 9922 292
rect 22066 184 22094 292
rect 33226 280 33232 292
rect 33284 280 33290 332
rect 34514 280 34520 332
rect 34572 280 34578 332
rect 24394 212 24400 264
rect 24452 252 24458 264
rect 30558 252 30564 264
rect 24452 224 30564 252
rect 24452 212 24458 224
rect 30558 212 30564 224
rect 30616 212 30622 264
rect 34532 184 34560 280
rect 57974 252 57980 264
rect 22066 156 34560 184
rect 35866 224 57980 252
rect 22922 76 22928 128
rect 22980 116 22986 128
rect 35866 116 35894 224
rect 57974 212 57980 224
rect 58032 212 58038 264
rect 22980 88 35894 116
rect 22980 76 22986 88
<< via1 >>
rect 36544 87592 36596 87644
rect 47308 87592 47360 87644
rect 27528 87524 27580 87576
rect 41696 87524 41748 87576
rect 33876 87456 33928 87508
rect 47860 87456 47912 87508
rect 37648 87388 37700 87440
rect 53564 87388 53616 87440
rect 3424 87320 3476 87372
rect 91284 87320 91336 87372
rect 11336 87252 11388 87304
rect 30196 87252 30248 87304
rect 30380 87252 30432 87304
rect 44824 87252 44876 87304
rect 1308 87184 1360 87236
rect 17316 87184 17368 87236
rect 44916 87184 44968 87236
rect 45100 87184 45152 87236
rect 63500 87184 63552 87236
rect 9036 87116 9088 87168
rect 24768 87116 24820 87168
rect 35348 87116 35400 87168
rect 10784 87048 10836 87100
rect 41788 87048 41840 87100
rect 72148 87116 72200 87168
rect 10416 86980 10468 87032
rect 36544 86980 36596 87032
rect 44916 86980 44968 87032
rect 77668 87048 77720 87100
rect 11428 86912 11480 86964
rect 50804 86912 50856 86964
rect 10508 86844 10560 86896
rect 62488 86844 62540 86896
rect 4896 86776 4948 86828
rect 58348 86776 58400 86828
rect 5540 86708 5592 86760
rect 61016 86708 61068 86760
rect 11520 86640 11572 86692
rect 68100 86640 68152 86692
rect 10600 86572 10652 86624
rect 68008 86572 68060 86624
rect 3610 86470 3662 86522
rect 3674 86470 3726 86522
rect 3738 86470 3790 86522
rect 3802 86470 3854 86522
rect 3866 86470 3918 86522
rect 5210 86470 5262 86522
rect 5274 86470 5326 86522
rect 5338 86470 5390 86522
rect 5402 86470 5454 86522
rect 5466 86470 5518 86522
rect 6810 86470 6862 86522
rect 6874 86470 6926 86522
rect 6938 86470 6990 86522
rect 7002 86470 7054 86522
rect 7066 86470 7118 86522
rect 8410 86470 8462 86522
rect 8474 86470 8526 86522
rect 8538 86470 8590 86522
rect 8602 86470 8654 86522
rect 8666 86470 8718 86522
rect 10010 86470 10062 86522
rect 10074 86470 10126 86522
rect 10138 86470 10190 86522
rect 10202 86470 10254 86522
rect 10266 86470 10318 86522
rect 11610 86470 11662 86522
rect 11674 86470 11726 86522
rect 11738 86470 11790 86522
rect 11802 86470 11854 86522
rect 11866 86470 11918 86522
rect 13210 86470 13262 86522
rect 13274 86470 13326 86522
rect 13338 86470 13390 86522
rect 13402 86470 13454 86522
rect 13466 86470 13518 86522
rect 14810 86470 14862 86522
rect 14874 86470 14926 86522
rect 14938 86470 14990 86522
rect 15002 86470 15054 86522
rect 15066 86470 15118 86522
rect 16410 86470 16462 86522
rect 16474 86470 16526 86522
rect 16538 86470 16590 86522
rect 16602 86470 16654 86522
rect 16666 86470 16718 86522
rect 18010 86470 18062 86522
rect 18074 86470 18126 86522
rect 18138 86470 18190 86522
rect 18202 86470 18254 86522
rect 18266 86470 18318 86522
rect 19610 86470 19662 86522
rect 19674 86470 19726 86522
rect 19738 86470 19790 86522
rect 19802 86470 19854 86522
rect 19866 86470 19918 86522
rect 21210 86470 21262 86522
rect 21274 86470 21326 86522
rect 21338 86470 21390 86522
rect 21402 86470 21454 86522
rect 21466 86470 21518 86522
rect 22810 86470 22862 86522
rect 22874 86470 22926 86522
rect 22938 86470 22990 86522
rect 23002 86470 23054 86522
rect 23066 86470 23118 86522
rect 24410 86470 24462 86522
rect 24474 86470 24526 86522
rect 24538 86470 24590 86522
rect 24602 86470 24654 86522
rect 24666 86470 24718 86522
rect 26010 86470 26062 86522
rect 26074 86470 26126 86522
rect 26138 86470 26190 86522
rect 26202 86470 26254 86522
rect 26266 86470 26318 86522
rect 27610 86470 27662 86522
rect 27674 86470 27726 86522
rect 27738 86470 27790 86522
rect 27802 86470 27854 86522
rect 27866 86470 27918 86522
rect 29210 86470 29262 86522
rect 29274 86470 29326 86522
rect 29338 86470 29390 86522
rect 29402 86470 29454 86522
rect 29466 86470 29518 86522
rect 30810 86470 30862 86522
rect 30874 86470 30926 86522
rect 30938 86470 30990 86522
rect 31002 86470 31054 86522
rect 31066 86470 31118 86522
rect 32410 86470 32462 86522
rect 32474 86470 32526 86522
rect 32538 86470 32590 86522
rect 32602 86470 32654 86522
rect 32666 86470 32718 86522
rect 34010 86470 34062 86522
rect 34074 86470 34126 86522
rect 34138 86470 34190 86522
rect 34202 86470 34254 86522
rect 34266 86470 34318 86522
rect 35610 86470 35662 86522
rect 35674 86470 35726 86522
rect 35738 86470 35790 86522
rect 35802 86470 35854 86522
rect 35866 86470 35918 86522
rect 37210 86470 37262 86522
rect 37274 86470 37326 86522
rect 37338 86470 37390 86522
rect 37402 86470 37454 86522
rect 37466 86470 37518 86522
rect 38810 86470 38862 86522
rect 38874 86470 38926 86522
rect 38938 86470 38990 86522
rect 39002 86470 39054 86522
rect 39066 86470 39118 86522
rect 40410 86470 40462 86522
rect 40474 86470 40526 86522
rect 40538 86470 40590 86522
rect 40602 86470 40654 86522
rect 40666 86470 40718 86522
rect 42010 86470 42062 86522
rect 42074 86470 42126 86522
rect 42138 86470 42190 86522
rect 42202 86470 42254 86522
rect 42266 86470 42318 86522
rect 43610 86470 43662 86522
rect 43674 86470 43726 86522
rect 43738 86470 43790 86522
rect 43802 86470 43854 86522
rect 43866 86470 43918 86522
rect 45210 86470 45262 86522
rect 45274 86470 45326 86522
rect 45338 86470 45390 86522
rect 45402 86470 45454 86522
rect 45466 86470 45518 86522
rect 46810 86470 46862 86522
rect 46874 86470 46926 86522
rect 46938 86470 46990 86522
rect 47002 86470 47054 86522
rect 47066 86470 47118 86522
rect 48410 86470 48462 86522
rect 48474 86470 48526 86522
rect 48538 86470 48590 86522
rect 48602 86470 48654 86522
rect 48666 86470 48718 86522
rect 50010 86470 50062 86522
rect 50074 86470 50126 86522
rect 50138 86470 50190 86522
rect 50202 86470 50254 86522
rect 50266 86470 50318 86522
rect 51610 86470 51662 86522
rect 51674 86470 51726 86522
rect 51738 86470 51790 86522
rect 51802 86470 51854 86522
rect 51866 86470 51918 86522
rect 53210 86470 53262 86522
rect 53274 86470 53326 86522
rect 53338 86470 53390 86522
rect 53402 86470 53454 86522
rect 53466 86470 53518 86522
rect 54810 86470 54862 86522
rect 54874 86470 54926 86522
rect 54938 86470 54990 86522
rect 55002 86470 55054 86522
rect 55066 86470 55118 86522
rect 56410 86470 56462 86522
rect 56474 86470 56526 86522
rect 56538 86470 56590 86522
rect 56602 86470 56654 86522
rect 56666 86470 56718 86522
rect 58010 86470 58062 86522
rect 58074 86470 58126 86522
rect 58138 86470 58190 86522
rect 58202 86470 58254 86522
rect 58266 86470 58318 86522
rect 59610 86470 59662 86522
rect 59674 86470 59726 86522
rect 59738 86470 59790 86522
rect 59802 86470 59854 86522
rect 59866 86470 59918 86522
rect 61210 86470 61262 86522
rect 61274 86470 61326 86522
rect 61338 86470 61390 86522
rect 61402 86470 61454 86522
rect 61466 86470 61518 86522
rect 62810 86470 62862 86522
rect 62874 86470 62926 86522
rect 62938 86470 62990 86522
rect 63002 86470 63054 86522
rect 63066 86470 63118 86522
rect 64410 86470 64462 86522
rect 64474 86470 64526 86522
rect 64538 86470 64590 86522
rect 64602 86470 64654 86522
rect 64666 86470 64718 86522
rect 66010 86470 66062 86522
rect 66074 86470 66126 86522
rect 66138 86470 66190 86522
rect 66202 86470 66254 86522
rect 66266 86470 66318 86522
rect 67610 86470 67662 86522
rect 67674 86470 67726 86522
rect 67738 86470 67790 86522
rect 67802 86470 67854 86522
rect 67866 86470 67918 86522
rect 69210 86470 69262 86522
rect 69274 86470 69326 86522
rect 69338 86470 69390 86522
rect 69402 86470 69454 86522
rect 69466 86470 69518 86522
rect 70810 86470 70862 86522
rect 70874 86470 70926 86522
rect 70938 86470 70990 86522
rect 71002 86470 71054 86522
rect 71066 86470 71118 86522
rect 72410 86470 72462 86522
rect 72474 86470 72526 86522
rect 72538 86470 72590 86522
rect 72602 86470 72654 86522
rect 72666 86470 72718 86522
rect 74010 86470 74062 86522
rect 74074 86470 74126 86522
rect 74138 86470 74190 86522
rect 74202 86470 74254 86522
rect 74266 86470 74318 86522
rect 75610 86470 75662 86522
rect 75674 86470 75726 86522
rect 75738 86470 75790 86522
rect 75802 86470 75854 86522
rect 75866 86470 75918 86522
rect 77210 86470 77262 86522
rect 77274 86470 77326 86522
rect 77338 86470 77390 86522
rect 77402 86470 77454 86522
rect 77466 86470 77518 86522
rect 78810 86470 78862 86522
rect 78874 86470 78926 86522
rect 78938 86470 78990 86522
rect 79002 86470 79054 86522
rect 79066 86470 79118 86522
rect 80410 86470 80462 86522
rect 80474 86470 80526 86522
rect 80538 86470 80590 86522
rect 80602 86470 80654 86522
rect 80666 86470 80718 86522
rect 82010 86470 82062 86522
rect 82074 86470 82126 86522
rect 82138 86470 82190 86522
rect 82202 86470 82254 86522
rect 82266 86470 82318 86522
rect 83610 86470 83662 86522
rect 83674 86470 83726 86522
rect 83738 86470 83790 86522
rect 83802 86470 83854 86522
rect 83866 86470 83918 86522
rect 85210 86470 85262 86522
rect 85274 86470 85326 86522
rect 85338 86470 85390 86522
rect 85402 86470 85454 86522
rect 85466 86470 85518 86522
rect 86810 86470 86862 86522
rect 86874 86470 86926 86522
rect 86938 86470 86990 86522
rect 87002 86470 87054 86522
rect 87066 86470 87118 86522
rect 88410 86470 88462 86522
rect 88474 86470 88526 86522
rect 88538 86470 88590 86522
rect 88602 86470 88654 86522
rect 88666 86470 88718 86522
rect 90010 86470 90062 86522
rect 90074 86470 90126 86522
rect 90138 86470 90190 86522
rect 90202 86470 90254 86522
rect 90266 86470 90318 86522
rect 91610 86470 91662 86522
rect 91674 86470 91726 86522
rect 91738 86470 91790 86522
rect 91802 86470 91854 86522
rect 91866 86470 91918 86522
rect 93210 86470 93262 86522
rect 93274 86470 93326 86522
rect 93338 86470 93390 86522
rect 93402 86470 93454 86522
rect 93466 86470 93518 86522
rect 94810 86470 94862 86522
rect 94874 86470 94926 86522
rect 94938 86470 94990 86522
rect 95002 86470 95054 86522
rect 95066 86470 95118 86522
rect 96410 86470 96462 86522
rect 96474 86470 96526 86522
rect 96538 86470 96590 86522
rect 96602 86470 96654 86522
rect 96666 86470 96718 86522
rect 98010 86470 98062 86522
rect 98074 86470 98126 86522
rect 98138 86470 98190 86522
rect 98202 86470 98254 86522
rect 98266 86470 98318 86522
rect 99610 86470 99662 86522
rect 99674 86470 99726 86522
rect 99738 86470 99790 86522
rect 99802 86470 99854 86522
rect 99866 86470 99918 86522
rect 101210 86470 101262 86522
rect 101274 86470 101326 86522
rect 101338 86470 101390 86522
rect 101402 86470 101454 86522
rect 101466 86470 101518 86522
rect 102810 86470 102862 86522
rect 102874 86470 102926 86522
rect 102938 86470 102990 86522
rect 103002 86470 103054 86522
rect 103066 86470 103118 86522
rect 104410 86470 104462 86522
rect 104474 86470 104526 86522
rect 104538 86470 104590 86522
rect 104602 86470 104654 86522
rect 104666 86470 104718 86522
rect 106010 86470 106062 86522
rect 106074 86470 106126 86522
rect 106138 86470 106190 86522
rect 106202 86470 106254 86522
rect 106266 86470 106318 86522
rect 107610 86470 107662 86522
rect 107674 86470 107726 86522
rect 107738 86470 107790 86522
rect 107802 86470 107854 86522
rect 107866 86470 107918 86522
rect 6000 86368 6052 86420
rect 13728 86368 13780 86420
rect 5908 86300 5960 86352
rect 4344 86232 4396 86284
rect 16948 86232 17000 86284
rect 4988 86164 5040 86216
rect 17224 86232 17276 86284
rect 34796 86300 34848 86352
rect 37372 86343 37424 86352
rect 37372 86309 37381 86343
rect 37381 86309 37415 86343
rect 37415 86309 37424 86343
rect 37372 86300 37424 86309
rect 25044 86275 25096 86284
rect 25044 86241 25053 86275
rect 25053 86241 25087 86275
rect 25087 86241 25096 86275
rect 25044 86232 25096 86241
rect 27160 86232 27212 86284
rect 11980 86096 12032 86148
rect 26792 86164 26844 86216
rect 17316 86096 17368 86148
rect 19708 86139 19760 86148
rect 19708 86105 19717 86139
rect 19717 86105 19751 86139
rect 19751 86105 19760 86139
rect 19708 86096 19760 86105
rect 19800 86096 19852 86148
rect 19984 86139 20036 86148
rect 19984 86105 19993 86139
rect 19993 86105 20027 86139
rect 20027 86105 20036 86139
rect 19984 86096 20036 86105
rect 24768 86139 24820 86148
rect 24768 86105 24777 86139
rect 24777 86105 24811 86139
rect 24811 86105 24820 86139
rect 24768 86096 24820 86105
rect 8760 86028 8812 86080
rect 24952 86071 25004 86080
rect 24952 86037 24961 86071
rect 24961 86037 24995 86071
rect 24995 86037 25004 86071
rect 24952 86028 25004 86037
rect 26792 86028 26844 86080
rect 27620 86207 27672 86216
rect 27620 86173 27629 86207
rect 27629 86173 27663 86207
rect 27663 86173 27672 86207
rect 27620 86164 27672 86173
rect 30012 86164 30064 86216
rect 30196 86139 30248 86148
rect 30196 86105 30205 86139
rect 30205 86105 30239 86139
rect 30239 86105 30248 86139
rect 30196 86096 30248 86105
rect 27252 86028 27304 86080
rect 27528 86071 27580 86080
rect 27528 86037 27537 86071
rect 27537 86037 27571 86071
rect 27571 86037 27580 86071
rect 27528 86028 27580 86037
rect 27620 86028 27672 86080
rect 33876 86139 33928 86148
rect 33876 86105 33885 86139
rect 33885 86105 33919 86139
rect 33919 86105 33928 86139
rect 33876 86096 33928 86105
rect 33968 86096 34020 86148
rect 34796 86164 34848 86216
rect 36084 86232 36136 86284
rect 40408 86275 40460 86284
rect 40408 86241 40417 86275
rect 40417 86241 40451 86275
rect 40451 86241 40460 86275
rect 40408 86232 40460 86241
rect 40776 86368 40828 86420
rect 41696 86368 41748 86420
rect 48964 86368 49016 86420
rect 50712 86411 50764 86420
rect 50712 86377 50721 86411
rect 50721 86377 50755 86411
rect 50755 86377 50764 86411
rect 50712 86368 50764 86377
rect 50804 86368 50856 86420
rect 58348 86368 58400 86420
rect 44824 86343 44876 86352
rect 44824 86309 44833 86343
rect 44833 86309 44867 86343
rect 44867 86309 44876 86343
rect 44824 86300 44876 86309
rect 47860 86343 47912 86352
rect 47860 86309 47869 86343
rect 47869 86309 47903 86343
rect 47903 86309 47912 86343
rect 47860 86300 47912 86309
rect 42708 86232 42760 86284
rect 42800 86232 42852 86284
rect 35348 86139 35400 86148
rect 35348 86105 35382 86139
rect 35382 86105 35400 86139
rect 30380 86071 30432 86080
rect 30380 86037 30389 86071
rect 30389 86037 30423 86071
rect 30423 86037 30432 86071
rect 30380 86028 30432 86037
rect 35348 86096 35400 86105
rect 36452 86071 36504 86080
rect 36452 86037 36461 86071
rect 36461 86037 36495 86071
rect 36495 86037 36504 86071
rect 36452 86028 36504 86037
rect 37648 86139 37700 86148
rect 37648 86105 37657 86139
rect 37657 86105 37691 86139
rect 37691 86105 37700 86139
rect 37648 86096 37700 86105
rect 38844 86139 38896 86148
rect 38844 86105 38853 86139
rect 38853 86105 38887 86139
rect 38887 86105 38896 86139
rect 38844 86096 38896 86105
rect 37832 86071 37884 86080
rect 37832 86037 37841 86071
rect 37841 86037 37875 86071
rect 37875 86037 37884 86071
rect 37832 86028 37884 86037
rect 40868 86139 40920 86148
rect 40868 86105 40902 86139
rect 40902 86105 40920 86139
rect 40868 86096 40920 86105
rect 42800 86028 42852 86080
rect 44916 86096 44968 86148
rect 48872 86096 48924 86148
rect 48964 86139 49016 86148
rect 48964 86105 48982 86139
rect 48982 86105 49016 86139
rect 48964 86096 49016 86105
rect 49240 86028 49292 86080
rect 49884 86071 49936 86080
rect 49884 86037 49893 86071
rect 49893 86037 49927 86071
rect 49927 86037 49936 86071
rect 49884 86028 49936 86037
rect 50712 86096 50764 86148
rect 52000 86071 52052 86080
rect 52000 86037 52009 86071
rect 52009 86037 52043 86071
rect 52043 86037 52052 86071
rect 52000 86028 52052 86037
rect 53012 86071 53064 86080
rect 53012 86037 53021 86071
rect 53021 86037 53055 86071
rect 53055 86037 53064 86071
rect 53012 86028 53064 86037
rect 55312 86207 55364 86216
rect 55312 86173 55321 86207
rect 55321 86173 55355 86207
rect 55355 86173 55364 86207
rect 55312 86164 55364 86173
rect 100944 86164 100996 86216
rect 108028 86207 108080 86216
rect 108028 86173 108037 86207
rect 108037 86173 108071 86207
rect 108071 86173 108080 86207
rect 108028 86164 108080 86173
rect 53564 86096 53616 86148
rect 74632 86096 74684 86148
rect 56692 86071 56744 86080
rect 56692 86037 56701 86071
rect 56701 86037 56735 86071
rect 56735 86037 56744 86071
rect 56692 86028 56744 86037
rect 2950 85926 3002 85978
rect 3014 85926 3066 85978
rect 3078 85926 3130 85978
rect 3142 85926 3194 85978
rect 3206 85926 3258 85978
rect 4550 85926 4602 85978
rect 4614 85926 4666 85978
rect 4678 85926 4730 85978
rect 4742 85926 4794 85978
rect 4806 85926 4858 85978
rect 6150 85926 6202 85978
rect 6214 85926 6266 85978
rect 6278 85926 6330 85978
rect 6342 85926 6394 85978
rect 6406 85926 6458 85978
rect 7750 85926 7802 85978
rect 7814 85926 7866 85978
rect 7878 85926 7930 85978
rect 7942 85926 7994 85978
rect 8006 85926 8058 85978
rect 9350 85926 9402 85978
rect 9414 85926 9466 85978
rect 9478 85926 9530 85978
rect 9542 85926 9594 85978
rect 9606 85926 9658 85978
rect 10950 85926 11002 85978
rect 11014 85926 11066 85978
rect 11078 85926 11130 85978
rect 11142 85926 11194 85978
rect 11206 85926 11258 85978
rect 12550 85926 12602 85978
rect 12614 85926 12666 85978
rect 12678 85926 12730 85978
rect 12742 85926 12794 85978
rect 12806 85926 12858 85978
rect 14150 85926 14202 85978
rect 14214 85926 14266 85978
rect 14278 85926 14330 85978
rect 14342 85926 14394 85978
rect 14406 85926 14458 85978
rect 15750 85926 15802 85978
rect 15814 85926 15866 85978
rect 15878 85926 15930 85978
rect 15942 85926 15994 85978
rect 16006 85926 16058 85978
rect 17350 85926 17402 85978
rect 17414 85926 17466 85978
rect 17478 85926 17530 85978
rect 17542 85926 17594 85978
rect 17606 85926 17658 85978
rect 18950 85926 19002 85978
rect 19014 85926 19066 85978
rect 19078 85926 19130 85978
rect 19142 85926 19194 85978
rect 19206 85926 19258 85978
rect 20550 85926 20602 85978
rect 20614 85926 20666 85978
rect 20678 85926 20730 85978
rect 20742 85926 20794 85978
rect 20806 85926 20858 85978
rect 22150 85926 22202 85978
rect 22214 85926 22266 85978
rect 22278 85926 22330 85978
rect 22342 85926 22394 85978
rect 22406 85926 22458 85978
rect 23750 85926 23802 85978
rect 23814 85926 23866 85978
rect 23878 85926 23930 85978
rect 23942 85926 23994 85978
rect 24006 85926 24058 85978
rect 25350 85926 25402 85978
rect 25414 85926 25466 85978
rect 25478 85926 25530 85978
rect 25542 85926 25594 85978
rect 25606 85926 25658 85978
rect 26950 85926 27002 85978
rect 27014 85926 27066 85978
rect 27078 85926 27130 85978
rect 27142 85926 27194 85978
rect 27206 85926 27258 85978
rect 28550 85926 28602 85978
rect 28614 85926 28666 85978
rect 28678 85926 28730 85978
rect 28742 85926 28794 85978
rect 28806 85926 28858 85978
rect 30150 85926 30202 85978
rect 30214 85926 30266 85978
rect 30278 85926 30330 85978
rect 30342 85926 30394 85978
rect 30406 85926 30458 85978
rect 31750 85926 31802 85978
rect 31814 85926 31866 85978
rect 31878 85926 31930 85978
rect 31942 85926 31994 85978
rect 32006 85926 32058 85978
rect 33350 85926 33402 85978
rect 33414 85926 33466 85978
rect 33478 85926 33530 85978
rect 33542 85926 33594 85978
rect 33606 85926 33658 85978
rect 34950 85926 35002 85978
rect 35014 85926 35066 85978
rect 35078 85926 35130 85978
rect 35142 85926 35194 85978
rect 35206 85926 35258 85978
rect 36550 85926 36602 85978
rect 36614 85926 36666 85978
rect 36678 85926 36730 85978
rect 36742 85926 36794 85978
rect 36806 85926 36858 85978
rect 38150 85926 38202 85978
rect 38214 85926 38266 85978
rect 38278 85926 38330 85978
rect 38342 85926 38394 85978
rect 38406 85926 38458 85978
rect 39750 85926 39802 85978
rect 39814 85926 39866 85978
rect 39878 85926 39930 85978
rect 39942 85926 39994 85978
rect 40006 85926 40058 85978
rect 41350 85926 41402 85978
rect 41414 85926 41466 85978
rect 41478 85926 41530 85978
rect 41542 85926 41594 85978
rect 41606 85926 41658 85978
rect 42950 85926 43002 85978
rect 43014 85926 43066 85978
rect 43078 85926 43130 85978
rect 43142 85926 43194 85978
rect 43206 85926 43258 85978
rect 44550 85926 44602 85978
rect 44614 85926 44666 85978
rect 44678 85926 44730 85978
rect 44742 85926 44794 85978
rect 44806 85926 44858 85978
rect 46150 85926 46202 85978
rect 46214 85926 46266 85978
rect 46278 85926 46330 85978
rect 46342 85926 46394 85978
rect 46406 85926 46458 85978
rect 47750 85926 47802 85978
rect 47814 85926 47866 85978
rect 47878 85926 47930 85978
rect 47942 85926 47994 85978
rect 48006 85926 48058 85978
rect 49350 85926 49402 85978
rect 49414 85926 49466 85978
rect 49478 85926 49530 85978
rect 49542 85926 49594 85978
rect 49606 85926 49658 85978
rect 50950 85926 51002 85978
rect 51014 85926 51066 85978
rect 51078 85926 51130 85978
rect 51142 85926 51194 85978
rect 51206 85926 51258 85978
rect 52550 85926 52602 85978
rect 52614 85926 52666 85978
rect 52678 85926 52730 85978
rect 52742 85926 52794 85978
rect 52806 85926 52858 85978
rect 54150 85926 54202 85978
rect 54214 85926 54266 85978
rect 54278 85926 54330 85978
rect 54342 85926 54394 85978
rect 54406 85926 54458 85978
rect 55750 85926 55802 85978
rect 55814 85926 55866 85978
rect 55878 85926 55930 85978
rect 55942 85926 55994 85978
rect 56006 85926 56058 85978
rect 57350 85926 57402 85978
rect 57414 85926 57466 85978
rect 57478 85926 57530 85978
rect 57542 85926 57594 85978
rect 57606 85926 57658 85978
rect 58950 85926 59002 85978
rect 59014 85926 59066 85978
rect 59078 85926 59130 85978
rect 59142 85926 59194 85978
rect 59206 85926 59258 85978
rect 60550 85926 60602 85978
rect 60614 85926 60666 85978
rect 60678 85926 60730 85978
rect 60742 85926 60794 85978
rect 60806 85926 60858 85978
rect 62150 85926 62202 85978
rect 62214 85926 62266 85978
rect 62278 85926 62330 85978
rect 62342 85926 62394 85978
rect 62406 85926 62458 85978
rect 63750 85926 63802 85978
rect 63814 85926 63866 85978
rect 63878 85926 63930 85978
rect 63942 85926 63994 85978
rect 64006 85926 64058 85978
rect 65350 85926 65402 85978
rect 65414 85926 65466 85978
rect 65478 85926 65530 85978
rect 65542 85926 65594 85978
rect 65606 85926 65658 85978
rect 66950 85926 67002 85978
rect 67014 85926 67066 85978
rect 67078 85926 67130 85978
rect 67142 85926 67194 85978
rect 67206 85926 67258 85978
rect 68550 85926 68602 85978
rect 68614 85926 68666 85978
rect 68678 85926 68730 85978
rect 68742 85926 68794 85978
rect 68806 85926 68858 85978
rect 70150 85926 70202 85978
rect 70214 85926 70266 85978
rect 70278 85926 70330 85978
rect 70342 85926 70394 85978
rect 70406 85926 70458 85978
rect 71750 85926 71802 85978
rect 71814 85926 71866 85978
rect 71878 85926 71930 85978
rect 71942 85926 71994 85978
rect 72006 85926 72058 85978
rect 73350 85926 73402 85978
rect 73414 85926 73466 85978
rect 73478 85926 73530 85978
rect 73542 85926 73594 85978
rect 73606 85926 73658 85978
rect 74950 85926 75002 85978
rect 75014 85926 75066 85978
rect 75078 85926 75130 85978
rect 75142 85926 75194 85978
rect 75206 85926 75258 85978
rect 76550 85926 76602 85978
rect 76614 85926 76666 85978
rect 76678 85926 76730 85978
rect 76742 85926 76794 85978
rect 76806 85926 76858 85978
rect 78150 85926 78202 85978
rect 78214 85926 78266 85978
rect 78278 85926 78330 85978
rect 78342 85926 78394 85978
rect 78406 85926 78458 85978
rect 79750 85926 79802 85978
rect 79814 85926 79866 85978
rect 79878 85926 79930 85978
rect 79942 85926 79994 85978
rect 80006 85926 80058 85978
rect 81350 85926 81402 85978
rect 81414 85926 81466 85978
rect 81478 85926 81530 85978
rect 81542 85926 81594 85978
rect 81606 85926 81658 85978
rect 82950 85926 83002 85978
rect 83014 85926 83066 85978
rect 83078 85926 83130 85978
rect 83142 85926 83194 85978
rect 83206 85926 83258 85978
rect 84550 85926 84602 85978
rect 84614 85926 84666 85978
rect 84678 85926 84730 85978
rect 84742 85926 84794 85978
rect 84806 85926 84858 85978
rect 86150 85926 86202 85978
rect 86214 85926 86266 85978
rect 86278 85926 86330 85978
rect 86342 85926 86394 85978
rect 86406 85926 86458 85978
rect 87750 85926 87802 85978
rect 87814 85926 87866 85978
rect 87878 85926 87930 85978
rect 87942 85926 87994 85978
rect 88006 85926 88058 85978
rect 89350 85926 89402 85978
rect 89414 85926 89466 85978
rect 89478 85926 89530 85978
rect 89542 85926 89594 85978
rect 89606 85926 89658 85978
rect 90950 85926 91002 85978
rect 91014 85926 91066 85978
rect 91078 85926 91130 85978
rect 91142 85926 91194 85978
rect 91206 85926 91258 85978
rect 92550 85926 92602 85978
rect 92614 85926 92666 85978
rect 92678 85926 92730 85978
rect 92742 85926 92794 85978
rect 92806 85926 92858 85978
rect 94150 85926 94202 85978
rect 94214 85926 94266 85978
rect 94278 85926 94330 85978
rect 94342 85926 94394 85978
rect 94406 85926 94458 85978
rect 95750 85926 95802 85978
rect 95814 85926 95866 85978
rect 95878 85926 95930 85978
rect 95942 85926 95994 85978
rect 96006 85926 96058 85978
rect 97350 85926 97402 85978
rect 97414 85926 97466 85978
rect 97478 85926 97530 85978
rect 97542 85926 97594 85978
rect 97606 85926 97658 85978
rect 98950 85926 99002 85978
rect 99014 85926 99066 85978
rect 99078 85926 99130 85978
rect 99142 85926 99194 85978
rect 99206 85926 99258 85978
rect 100550 85926 100602 85978
rect 100614 85926 100666 85978
rect 100678 85926 100730 85978
rect 100742 85926 100794 85978
rect 100806 85926 100858 85978
rect 102150 85926 102202 85978
rect 102214 85926 102266 85978
rect 102278 85926 102330 85978
rect 102342 85926 102394 85978
rect 102406 85926 102458 85978
rect 103750 85926 103802 85978
rect 103814 85926 103866 85978
rect 103878 85926 103930 85978
rect 103942 85926 103994 85978
rect 104006 85926 104058 85978
rect 105350 85926 105402 85978
rect 105414 85926 105466 85978
rect 105478 85926 105530 85978
rect 105542 85926 105594 85978
rect 105606 85926 105658 85978
rect 106950 85926 107002 85978
rect 107014 85926 107066 85978
rect 107078 85926 107130 85978
rect 107142 85926 107194 85978
rect 107206 85926 107258 85978
rect 108550 85926 108602 85978
rect 108614 85926 108666 85978
rect 108678 85926 108730 85978
rect 108742 85926 108794 85978
rect 108806 85926 108858 85978
rect 4436 85824 4488 85876
rect 25044 85824 25096 85876
rect 27620 85824 27672 85876
rect 30012 85824 30064 85876
rect 33876 85824 33928 85876
rect 36084 85824 36136 85876
rect 40408 85824 40460 85876
rect 42800 85824 42852 85876
rect 9220 85756 9272 85808
rect 19800 85756 19852 85808
rect 37648 85756 37700 85808
rect 8944 85688 8996 85740
rect 19984 85688 20036 85740
rect 24952 85688 25004 85740
rect 36452 85688 36504 85740
rect 13728 85620 13780 85672
rect 19708 85620 19760 85672
rect 9128 85552 9180 85604
rect 26792 85552 26844 85604
rect 26976 85620 27028 85672
rect 40868 85756 40920 85808
rect 75920 85824 75972 85876
rect 46572 85756 46624 85808
rect 49884 85756 49936 85808
rect 37832 85688 37884 85740
rect 56692 85756 56744 85808
rect 52000 85688 52052 85740
rect 73160 85688 73212 85740
rect 40776 85620 40828 85672
rect 42708 85620 42760 85672
rect 55220 85620 55272 85672
rect 38844 85552 38896 85604
rect 42800 85552 42852 85604
rect 46940 85552 46992 85604
rect 55680 85552 55732 85604
rect 1032 85484 1084 85536
rect 40040 85484 40092 85536
rect 3610 85382 3662 85434
rect 3674 85382 3726 85434
rect 3738 85382 3790 85434
rect 3802 85382 3854 85434
rect 3866 85382 3918 85434
rect 5210 85382 5262 85434
rect 5274 85382 5326 85434
rect 5338 85382 5390 85434
rect 5402 85382 5454 85434
rect 5466 85382 5518 85434
rect 6810 85382 6862 85434
rect 6874 85382 6926 85434
rect 6938 85382 6990 85434
rect 7002 85382 7054 85434
rect 7066 85382 7118 85434
rect 8410 85382 8462 85434
rect 8474 85382 8526 85434
rect 8538 85382 8590 85434
rect 8602 85382 8654 85434
rect 8666 85382 8718 85434
rect 10324 85416 10376 85468
rect 46572 85416 46624 85468
rect 11704 85348 11756 85400
rect 49240 85348 49292 85400
rect 10140 85280 10192 85332
rect 52460 85280 52512 85332
rect 8208 85212 8260 85264
rect 53840 85212 53892 85264
rect 8116 85144 8168 85196
rect 51172 85144 51224 85196
rect 7472 85076 7524 85128
rect 66260 85076 66312 85128
rect 7196 85008 7248 85060
rect 71228 85008 71280 85060
rect 6552 84940 6604 84992
rect 34796 84940 34848 84992
rect 2950 84838 3002 84890
rect 3014 84838 3066 84890
rect 3078 84838 3130 84890
rect 3142 84838 3194 84890
rect 3206 84838 3258 84890
rect 4550 84838 4602 84890
rect 4614 84838 4666 84890
rect 4678 84838 4730 84890
rect 4742 84838 4794 84890
rect 4806 84838 4858 84890
rect 6150 84838 6202 84890
rect 6214 84838 6266 84890
rect 6278 84838 6330 84890
rect 6342 84838 6394 84890
rect 6406 84838 6458 84890
rect 7750 84838 7802 84890
rect 7814 84838 7866 84890
rect 7878 84838 7930 84890
rect 7942 84838 7994 84890
rect 8006 84838 8058 84890
rect 9350 84838 9402 84890
rect 9414 84838 9466 84890
rect 9478 84838 9530 84890
rect 9542 84838 9594 84890
rect 9606 84838 9658 84890
rect 10876 84872 10928 84924
rect 57612 84872 57664 84924
rect 10692 84804 10744 84856
rect 78680 84804 78732 84856
rect 11796 84736 11848 84788
rect 44732 84736 44784 84788
rect 11888 84668 11940 84720
rect 42524 84668 42576 84720
rect 940 84600 992 84652
rect 4160 84600 4212 84652
rect 27344 84600 27396 84652
rect 1676 84507 1728 84516
rect 1676 84473 1685 84507
rect 1685 84473 1719 84507
rect 1719 84473 1728 84507
rect 1676 84464 1728 84473
rect 3610 84294 3662 84346
rect 3674 84294 3726 84346
rect 3738 84294 3790 84346
rect 3802 84294 3854 84346
rect 3866 84294 3918 84346
rect 5210 84294 5262 84346
rect 5274 84294 5326 84346
rect 5338 84294 5390 84346
rect 5402 84294 5454 84346
rect 5466 84294 5518 84346
rect 6810 84294 6862 84346
rect 6874 84294 6926 84346
rect 6938 84294 6990 84346
rect 7002 84294 7054 84346
rect 7066 84294 7118 84346
rect 8410 84294 8462 84346
rect 8474 84294 8526 84346
rect 8538 84294 8590 84346
rect 8602 84294 8654 84346
rect 8666 84294 8718 84346
rect 6644 83852 6696 83904
rect 37372 83852 37424 83904
rect 2950 83750 3002 83802
rect 3014 83750 3066 83802
rect 3078 83750 3130 83802
rect 3142 83750 3194 83802
rect 3206 83750 3258 83802
rect 4550 83750 4602 83802
rect 4614 83750 4666 83802
rect 4678 83750 4730 83802
rect 4742 83750 4794 83802
rect 4806 83750 4858 83802
rect 6150 83750 6202 83802
rect 6214 83750 6266 83802
rect 6278 83750 6330 83802
rect 6342 83750 6394 83802
rect 6406 83750 6458 83802
rect 7750 83750 7802 83802
rect 7814 83750 7866 83802
rect 7878 83750 7930 83802
rect 7942 83750 7994 83802
rect 8006 83750 8058 83802
rect 9350 83750 9402 83802
rect 9414 83750 9466 83802
rect 9478 83750 9530 83802
rect 9542 83750 9594 83802
rect 9606 83750 9658 83802
rect 7380 83648 7432 83700
rect 45100 83648 45152 83700
rect 8300 83580 8352 83632
rect 46940 83580 46992 83632
rect 940 83512 992 83564
rect 10968 83512 11020 83564
rect 59912 83512 59964 83564
rect 10232 83444 10284 83496
rect 70216 83444 70268 83496
rect 3976 83376 4028 83428
rect 3610 83206 3662 83258
rect 3674 83206 3726 83258
rect 3738 83206 3790 83258
rect 3802 83206 3854 83258
rect 3866 83206 3918 83258
rect 5210 83206 5262 83258
rect 5274 83206 5326 83258
rect 5338 83206 5390 83258
rect 5402 83206 5454 83258
rect 5466 83206 5518 83258
rect 6810 83206 6862 83258
rect 6874 83206 6926 83258
rect 6938 83206 6990 83258
rect 7002 83206 7054 83258
rect 7066 83206 7118 83258
rect 8410 83206 8462 83258
rect 8474 83206 8526 83258
rect 8538 83206 8590 83258
rect 8602 83206 8654 83258
rect 8666 83206 8718 83258
rect 1492 82875 1544 82884
rect 1492 82841 1501 82875
rect 1501 82841 1535 82875
rect 1535 82841 1544 82875
rect 1492 82832 1544 82841
rect 2228 82832 2280 82884
rect 2950 82662 3002 82714
rect 3014 82662 3066 82714
rect 3078 82662 3130 82714
rect 3142 82662 3194 82714
rect 3206 82662 3258 82714
rect 4550 82662 4602 82714
rect 4614 82662 4666 82714
rect 4678 82662 4730 82714
rect 4742 82662 4794 82714
rect 4806 82662 4858 82714
rect 6150 82662 6202 82714
rect 6214 82662 6266 82714
rect 6278 82662 6330 82714
rect 6342 82662 6394 82714
rect 6406 82662 6458 82714
rect 7750 82662 7802 82714
rect 7814 82662 7866 82714
rect 7878 82662 7930 82714
rect 7942 82662 7994 82714
rect 8006 82662 8058 82714
rect 9350 82662 9402 82714
rect 9414 82662 9466 82714
rect 9478 82662 9530 82714
rect 9542 82662 9594 82714
rect 9606 82662 9658 82714
rect 3610 82118 3662 82170
rect 3674 82118 3726 82170
rect 3738 82118 3790 82170
rect 3802 82118 3854 82170
rect 3866 82118 3918 82170
rect 5210 82118 5262 82170
rect 5274 82118 5326 82170
rect 5338 82118 5390 82170
rect 5402 82118 5454 82170
rect 5466 82118 5518 82170
rect 6810 82118 6862 82170
rect 6874 82118 6926 82170
rect 6938 82118 6990 82170
rect 7002 82118 7054 82170
rect 7066 82118 7118 82170
rect 8410 82118 8462 82170
rect 8474 82118 8526 82170
rect 8538 82118 8590 82170
rect 8602 82118 8654 82170
rect 8666 82118 8718 82170
rect 940 81744 992 81796
rect 1768 81744 1820 81796
rect 2950 81574 3002 81626
rect 3014 81574 3066 81626
rect 3078 81574 3130 81626
rect 3142 81574 3194 81626
rect 3206 81574 3258 81626
rect 4550 81574 4602 81626
rect 4614 81574 4666 81626
rect 4678 81574 4730 81626
rect 4742 81574 4794 81626
rect 4806 81574 4858 81626
rect 6150 81574 6202 81626
rect 6214 81574 6266 81626
rect 6278 81574 6330 81626
rect 6342 81574 6394 81626
rect 6406 81574 6458 81626
rect 7750 81574 7802 81626
rect 7814 81574 7866 81626
rect 7878 81574 7930 81626
rect 7942 81574 7994 81626
rect 8006 81574 8058 81626
rect 9350 81574 9402 81626
rect 9414 81574 9466 81626
rect 9478 81574 9530 81626
rect 9542 81574 9594 81626
rect 9606 81574 9658 81626
rect 3610 81030 3662 81082
rect 3674 81030 3726 81082
rect 3738 81030 3790 81082
rect 3802 81030 3854 81082
rect 3866 81030 3918 81082
rect 5210 81030 5262 81082
rect 5274 81030 5326 81082
rect 5338 81030 5390 81082
rect 5402 81030 5454 81082
rect 5466 81030 5518 81082
rect 6810 81030 6862 81082
rect 6874 81030 6926 81082
rect 6938 81030 6990 81082
rect 7002 81030 7054 81082
rect 7066 81030 7118 81082
rect 8410 81030 8462 81082
rect 8474 81030 8526 81082
rect 8538 81030 8590 81082
rect 8602 81030 8654 81082
rect 8666 81030 8718 81082
rect 940 80656 992 80708
rect 1860 80656 1912 80708
rect 2950 80486 3002 80538
rect 3014 80486 3066 80538
rect 3078 80486 3130 80538
rect 3142 80486 3194 80538
rect 3206 80486 3258 80538
rect 4550 80486 4602 80538
rect 4614 80486 4666 80538
rect 4678 80486 4730 80538
rect 4742 80486 4794 80538
rect 4806 80486 4858 80538
rect 6150 80486 6202 80538
rect 6214 80486 6266 80538
rect 6278 80486 6330 80538
rect 6342 80486 6394 80538
rect 6406 80486 6458 80538
rect 7750 80486 7802 80538
rect 7814 80486 7866 80538
rect 7878 80486 7930 80538
rect 7942 80486 7994 80538
rect 8006 80486 8058 80538
rect 9350 80486 9402 80538
rect 9414 80486 9466 80538
rect 9478 80486 9530 80538
rect 9542 80486 9594 80538
rect 9606 80486 9658 80538
rect 3610 79942 3662 79994
rect 3674 79942 3726 79994
rect 3738 79942 3790 79994
rect 3802 79942 3854 79994
rect 3866 79942 3918 79994
rect 5210 79942 5262 79994
rect 5274 79942 5326 79994
rect 5338 79942 5390 79994
rect 5402 79942 5454 79994
rect 5466 79942 5518 79994
rect 6810 79942 6862 79994
rect 6874 79942 6926 79994
rect 6938 79942 6990 79994
rect 7002 79942 7054 79994
rect 7066 79942 7118 79994
rect 8410 79942 8462 79994
rect 8474 79942 8526 79994
rect 8538 79942 8590 79994
rect 8602 79942 8654 79994
rect 8666 79942 8718 79994
rect 940 79568 992 79620
rect 2044 79568 2096 79620
rect 4160 79500 4212 79552
rect 4988 79500 5040 79552
rect 2950 79398 3002 79450
rect 3014 79398 3066 79450
rect 3078 79398 3130 79450
rect 3142 79398 3194 79450
rect 3206 79398 3258 79450
rect 4550 79398 4602 79450
rect 4614 79398 4666 79450
rect 4678 79398 4730 79450
rect 4742 79398 4794 79450
rect 4806 79398 4858 79450
rect 6150 79398 6202 79450
rect 6214 79398 6266 79450
rect 6278 79398 6330 79450
rect 6342 79398 6394 79450
rect 6406 79398 6458 79450
rect 7750 79398 7802 79450
rect 7814 79398 7866 79450
rect 7878 79398 7930 79450
rect 7942 79398 7994 79450
rect 8006 79398 8058 79450
rect 9350 79398 9402 79450
rect 9414 79398 9466 79450
rect 9478 79398 9530 79450
rect 9542 79398 9594 79450
rect 9606 79398 9658 79450
rect 940 79160 992 79212
rect 1216 78956 1268 79008
rect 3610 78854 3662 78906
rect 3674 78854 3726 78906
rect 3738 78854 3790 78906
rect 3802 78854 3854 78906
rect 3866 78854 3918 78906
rect 5210 78854 5262 78906
rect 5274 78854 5326 78906
rect 5338 78854 5390 78906
rect 5402 78854 5454 78906
rect 5466 78854 5518 78906
rect 6810 78854 6862 78906
rect 6874 78854 6926 78906
rect 6938 78854 6990 78906
rect 7002 78854 7054 78906
rect 7066 78854 7118 78906
rect 8410 78854 8462 78906
rect 8474 78854 8526 78906
rect 8538 78854 8590 78906
rect 8602 78854 8654 78906
rect 8666 78854 8718 78906
rect 2950 78310 3002 78362
rect 3014 78310 3066 78362
rect 3078 78310 3130 78362
rect 3142 78310 3194 78362
rect 3206 78310 3258 78362
rect 4550 78310 4602 78362
rect 4614 78310 4666 78362
rect 4678 78310 4730 78362
rect 4742 78310 4794 78362
rect 4806 78310 4858 78362
rect 6150 78310 6202 78362
rect 6214 78310 6266 78362
rect 6278 78310 6330 78362
rect 6342 78310 6394 78362
rect 6406 78310 6458 78362
rect 7750 78310 7802 78362
rect 7814 78310 7866 78362
rect 7878 78310 7930 78362
rect 7942 78310 7994 78362
rect 8006 78310 8058 78362
rect 9350 78310 9402 78362
rect 9414 78310 9466 78362
rect 9478 78310 9530 78362
rect 9542 78310 9594 78362
rect 9606 78310 9658 78362
rect 940 78072 992 78124
rect 3332 77868 3384 77920
rect 3610 77766 3662 77818
rect 3674 77766 3726 77818
rect 3738 77766 3790 77818
rect 3802 77766 3854 77818
rect 3866 77766 3918 77818
rect 5210 77766 5262 77818
rect 5274 77766 5326 77818
rect 5338 77766 5390 77818
rect 5402 77766 5454 77818
rect 5466 77766 5518 77818
rect 6810 77766 6862 77818
rect 6874 77766 6926 77818
rect 6938 77766 6990 77818
rect 7002 77766 7054 77818
rect 7066 77766 7118 77818
rect 8410 77766 8462 77818
rect 8474 77766 8526 77818
rect 8538 77766 8590 77818
rect 8602 77766 8654 77818
rect 8666 77766 8718 77818
rect 2950 77222 3002 77274
rect 3014 77222 3066 77274
rect 3078 77222 3130 77274
rect 3142 77222 3194 77274
rect 3206 77222 3258 77274
rect 4550 77222 4602 77274
rect 4614 77222 4666 77274
rect 4678 77222 4730 77274
rect 4742 77222 4794 77274
rect 4806 77222 4858 77274
rect 6150 77222 6202 77274
rect 6214 77222 6266 77274
rect 6278 77222 6330 77274
rect 6342 77222 6394 77274
rect 6406 77222 6458 77274
rect 7750 77222 7802 77274
rect 7814 77222 7866 77274
rect 7878 77222 7930 77274
rect 7942 77222 7994 77274
rect 8006 77222 8058 77274
rect 9350 77222 9402 77274
rect 9414 77222 9466 77274
rect 9478 77222 9530 77274
rect 9542 77222 9594 77274
rect 9606 77222 9658 77274
rect 9036 77120 9088 77172
rect 940 76984 992 77036
rect 7656 76984 7708 77036
rect 10140 76984 10192 77036
rect 8944 76916 8996 76968
rect 2596 76848 2648 76900
rect 2504 76780 2556 76832
rect 3610 76678 3662 76730
rect 3674 76678 3726 76730
rect 3738 76678 3790 76730
rect 3802 76678 3854 76730
rect 3866 76678 3918 76730
rect 5210 76678 5262 76730
rect 5274 76678 5326 76730
rect 5338 76678 5390 76730
rect 5402 76678 5454 76730
rect 5466 76678 5518 76730
rect 6810 76678 6862 76730
rect 6874 76678 6926 76730
rect 6938 76678 6990 76730
rect 7002 76678 7054 76730
rect 7066 76678 7118 76730
rect 8410 76678 8462 76730
rect 8474 76678 8526 76730
rect 8538 76678 8590 76730
rect 8602 76678 8654 76730
rect 8666 76678 8718 76730
rect 8760 76440 8812 76492
rect 8944 76440 8996 76492
rect 8208 76372 8260 76424
rect 8852 76304 8904 76356
rect 1124 76236 1176 76288
rect 2950 76134 3002 76186
rect 3014 76134 3066 76186
rect 3078 76134 3130 76186
rect 3142 76134 3194 76186
rect 3206 76134 3258 76186
rect 4550 76134 4602 76186
rect 4614 76134 4666 76186
rect 4678 76134 4730 76186
rect 4742 76134 4794 76186
rect 4806 76134 4858 76186
rect 6150 76134 6202 76186
rect 6214 76134 6266 76186
rect 6278 76134 6330 76186
rect 6342 76134 6394 76186
rect 6406 76134 6458 76186
rect 7750 76134 7802 76186
rect 7814 76134 7866 76186
rect 7878 76134 7930 76186
rect 7942 76134 7994 76186
rect 8006 76134 8058 76186
rect 9350 76134 9402 76186
rect 9414 76134 9466 76186
rect 9478 76134 9530 76186
rect 9542 76134 9594 76186
rect 9606 76134 9658 76186
rect 1492 75939 1544 75948
rect 1492 75905 1501 75939
rect 1501 75905 1535 75939
rect 1535 75905 1544 75939
rect 1492 75896 1544 75905
rect 4068 75760 4120 75812
rect 3610 75590 3662 75642
rect 3674 75590 3726 75642
rect 3738 75590 3790 75642
rect 3802 75590 3854 75642
rect 3866 75590 3918 75642
rect 5210 75590 5262 75642
rect 5274 75590 5326 75642
rect 5338 75590 5390 75642
rect 5402 75590 5454 75642
rect 5466 75590 5518 75642
rect 6810 75590 6862 75642
rect 6874 75590 6926 75642
rect 6938 75590 6990 75642
rect 7002 75590 7054 75642
rect 7066 75590 7118 75642
rect 8410 75590 8462 75642
rect 8474 75590 8526 75642
rect 8538 75590 8590 75642
rect 8602 75590 8654 75642
rect 8666 75590 8718 75642
rect 4436 75352 4488 75404
rect 5724 75352 5776 75404
rect 8484 75352 8536 75404
rect 9220 75327 9272 75336
rect 9220 75293 9229 75327
rect 9229 75293 9263 75327
rect 9263 75293 9272 75327
rect 9220 75284 9272 75293
rect 940 75216 992 75268
rect 2688 75216 2740 75268
rect 7196 75216 7248 75268
rect 9496 75284 9548 75336
rect 4436 75148 4488 75200
rect 4896 75148 4948 75200
rect 5632 75148 5684 75200
rect 2950 75046 3002 75098
rect 3014 75046 3066 75098
rect 3078 75046 3130 75098
rect 3142 75046 3194 75098
rect 3206 75046 3258 75098
rect 4550 75046 4602 75098
rect 4614 75046 4666 75098
rect 4678 75046 4730 75098
rect 4742 75046 4794 75098
rect 4806 75046 4858 75098
rect 6150 75046 6202 75098
rect 6214 75046 6266 75098
rect 6278 75046 6330 75098
rect 6342 75046 6394 75098
rect 6406 75046 6458 75098
rect 7750 75046 7802 75098
rect 7814 75046 7866 75098
rect 7878 75046 7930 75098
rect 7942 75046 7994 75098
rect 8006 75046 8058 75098
rect 9350 75046 9402 75098
rect 9414 75046 9466 75098
rect 9478 75046 9530 75098
rect 9542 75046 9594 75098
rect 9606 75046 9658 75098
rect 4252 74944 4304 74996
rect 4896 74944 4948 74996
rect 8760 74944 8812 74996
rect 8484 74851 8536 74860
rect 8484 74817 8493 74851
rect 8493 74817 8527 74851
rect 8527 74817 8536 74851
rect 8484 74808 8536 74817
rect 9588 74876 9640 74928
rect 7564 74740 7616 74792
rect 8300 74672 8352 74724
rect 8760 74672 8812 74724
rect 9312 74783 9364 74792
rect 9312 74749 9321 74783
rect 9321 74749 9355 74783
rect 9355 74749 9364 74783
rect 9312 74740 9364 74749
rect 9404 74783 9456 74792
rect 9404 74749 9413 74783
rect 9413 74749 9447 74783
rect 9447 74749 9456 74783
rect 9404 74740 9456 74749
rect 5908 74604 5960 74656
rect 8208 74604 8260 74656
rect 8484 74604 8536 74656
rect 9680 74604 9732 74656
rect 3610 74502 3662 74554
rect 3674 74502 3726 74554
rect 3738 74502 3790 74554
rect 3802 74502 3854 74554
rect 3866 74502 3918 74554
rect 5210 74502 5262 74554
rect 5274 74502 5326 74554
rect 5338 74502 5390 74554
rect 5402 74502 5454 74554
rect 5466 74502 5518 74554
rect 6810 74502 6862 74554
rect 6874 74502 6926 74554
rect 6938 74502 6990 74554
rect 7002 74502 7054 74554
rect 7066 74502 7118 74554
rect 8410 74502 8462 74554
rect 8474 74502 8526 74554
rect 8538 74502 8590 74554
rect 8602 74502 8654 74554
rect 8666 74502 8718 74554
rect 7288 74400 7340 74452
rect 9312 74400 9364 74452
rect 8944 74332 8996 74384
rect 9220 74332 9272 74384
rect 940 74196 992 74248
rect 6920 74196 6972 74248
rect 7196 74196 7248 74248
rect 8208 74196 8260 74248
rect 9036 74196 9088 74248
rect 9588 74239 9640 74248
rect 9128 74128 9180 74180
rect 9588 74205 9597 74239
rect 9597 74205 9631 74239
rect 9631 74205 9640 74239
rect 9588 74196 9640 74205
rect 1952 74060 2004 74112
rect 8944 74103 8996 74112
rect 8944 74069 8953 74103
rect 8953 74069 8987 74103
rect 8987 74069 8996 74103
rect 8944 74060 8996 74069
rect 9036 74060 9088 74112
rect 9404 74060 9456 74112
rect 9772 74060 9824 74112
rect 2950 73958 3002 74010
rect 3014 73958 3066 74010
rect 3078 73958 3130 74010
rect 3142 73958 3194 74010
rect 3206 73958 3258 74010
rect 4550 73958 4602 74010
rect 4614 73958 4666 74010
rect 4678 73958 4730 74010
rect 4742 73958 4794 74010
rect 4806 73958 4858 74010
rect 6150 73958 6202 74010
rect 6214 73958 6266 74010
rect 6278 73958 6330 74010
rect 6342 73958 6394 74010
rect 6406 73958 6458 74010
rect 7750 73958 7802 74010
rect 7814 73958 7866 74010
rect 7878 73958 7930 74010
rect 7942 73958 7994 74010
rect 8006 73958 8058 74010
rect 9350 73958 9402 74010
rect 9414 73958 9466 74010
rect 9478 73958 9530 74010
rect 9542 73958 9594 74010
rect 9606 73958 9658 74010
rect 3516 73856 3568 73908
rect 6828 73788 6880 73840
rect 6736 73720 6788 73772
rect 7840 73763 7892 73772
rect 7840 73729 7849 73763
rect 7849 73729 7883 73763
rect 7883 73729 7892 73763
rect 7840 73720 7892 73729
rect 8024 73720 8076 73772
rect 8116 73763 8168 73772
rect 8116 73729 8125 73763
rect 8125 73729 8159 73763
rect 8159 73729 8168 73763
rect 8116 73720 8168 73729
rect 8392 73720 8444 73772
rect 6460 73652 6512 73704
rect 7196 73652 7248 73704
rect 7472 73652 7524 73704
rect 9956 73584 10008 73636
rect 6920 73516 6972 73568
rect 8300 73516 8352 73568
rect 8392 73516 8444 73568
rect 9312 73516 9364 73568
rect 3610 73414 3662 73466
rect 3674 73414 3726 73466
rect 3738 73414 3790 73466
rect 3802 73414 3854 73466
rect 3866 73414 3918 73466
rect 5210 73414 5262 73466
rect 5274 73414 5326 73466
rect 5338 73414 5390 73466
rect 5402 73414 5454 73466
rect 5466 73414 5518 73466
rect 6810 73414 6862 73466
rect 6874 73414 6926 73466
rect 6938 73414 6990 73466
rect 7002 73414 7054 73466
rect 7066 73414 7118 73466
rect 8410 73414 8462 73466
rect 8474 73414 8526 73466
rect 8538 73414 8590 73466
rect 8602 73414 8654 73466
rect 8666 73414 8718 73466
rect 4988 73312 5040 73364
rect 7380 73312 7432 73364
rect 8116 73312 8168 73364
rect 8484 73312 8536 73364
rect 7840 73244 7892 73296
rect 6644 73176 6696 73228
rect 6460 73108 6512 73160
rect 6920 73176 6972 73228
rect 6828 73108 6880 73160
rect 7748 73176 7800 73228
rect 7932 73219 7984 73228
rect 7932 73185 7941 73219
rect 7941 73185 7975 73219
rect 7975 73185 7984 73219
rect 7932 73176 7984 73185
rect 8208 73244 8260 73296
rect 8392 73244 8444 73296
rect 7564 73108 7616 73160
rect 940 73040 992 73092
rect 4344 73040 4396 73092
rect 7104 73040 7156 73092
rect 7472 73040 7524 73092
rect 1584 73015 1636 73024
rect 1584 72981 1593 73015
rect 1593 72981 1627 73015
rect 1627 72981 1636 73015
rect 1584 72972 1636 72981
rect 7656 73040 7708 73092
rect 8392 73151 8444 73160
rect 8392 73117 8401 73151
rect 8401 73117 8435 73151
rect 8435 73117 8444 73151
rect 8392 73108 8444 73117
rect 8852 73108 8904 73160
rect 10140 73108 10192 73160
rect 10508 73108 10560 73160
rect 8484 72972 8536 73024
rect 9312 72972 9364 73024
rect 2950 72870 3002 72922
rect 3014 72870 3066 72922
rect 3078 72870 3130 72922
rect 3142 72870 3194 72922
rect 3206 72870 3258 72922
rect 4550 72870 4602 72922
rect 4614 72870 4666 72922
rect 4678 72870 4730 72922
rect 4742 72870 4794 72922
rect 4806 72870 4858 72922
rect 6150 72870 6202 72922
rect 6214 72870 6266 72922
rect 6278 72870 6330 72922
rect 6342 72870 6394 72922
rect 6406 72870 6458 72922
rect 7750 72870 7802 72922
rect 7814 72870 7866 72922
rect 7878 72870 7930 72922
rect 7942 72870 7994 72922
rect 8006 72870 8058 72922
rect 9350 72870 9402 72922
rect 9414 72870 9466 72922
rect 9478 72870 9530 72922
rect 9542 72870 9594 72922
rect 9606 72870 9658 72922
rect 8484 72768 8536 72820
rect 6000 72700 6052 72752
rect 2044 72632 2096 72684
rect 4252 72632 4304 72684
rect 6460 72675 6512 72684
rect 6460 72641 6469 72675
rect 6469 72641 6503 72675
rect 6503 72641 6512 72675
rect 6460 72632 6512 72641
rect 6828 72632 6880 72684
rect 7196 72632 7248 72684
rect 7380 72675 7432 72684
rect 7380 72641 7389 72675
rect 7389 72641 7423 72675
rect 7423 72641 7432 72675
rect 7380 72632 7432 72641
rect 7472 72675 7524 72684
rect 7472 72641 7481 72675
rect 7481 72641 7515 72675
rect 7515 72641 7524 72675
rect 7472 72632 7524 72641
rect 7656 72632 7708 72684
rect 7932 72632 7984 72684
rect 6000 72564 6052 72616
rect 6920 72564 6972 72616
rect 7104 72564 7156 72616
rect 8024 72564 8076 72616
rect 8392 72675 8444 72684
rect 8392 72641 8401 72675
rect 8401 72641 8435 72675
rect 8435 72641 8444 72675
rect 8392 72632 8444 72641
rect 8484 72675 8536 72684
rect 8484 72641 8493 72675
rect 8493 72641 8527 72675
rect 8527 72641 8536 72675
rect 8484 72632 8536 72641
rect 8852 72675 8904 72684
rect 8852 72641 8861 72675
rect 8861 72641 8895 72675
rect 8895 72641 8904 72675
rect 8852 72632 8904 72641
rect 4896 72496 4948 72548
rect 6828 72471 6880 72480
rect 6828 72437 6837 72471
rect 6837 72437 6871 72471
rect 6871 72437 6880 72471
rect 6828 72428 6880 72437
rect 7012 72471 7064 72480
rect 7012 72437 7021 72471
rect 7021 72437 7055 72471
rect 7055 72437 7064 72471
rect 7012 72428 7064 72437
rect 7472 72428 7524 72480
rect 7748 72428 7800 72480
rect 8208 72496 8260 72548
rect 9404 72564 9456 72616
rect 10140 72564 10192 72616
rect 8576 72471 8628 72480
rect 8576 72437 8585 72471
rect 8585 72437 8619 72471
rect 8619 72437 8628 72471
rect 8576 72428 8628 72437
rect 9404 72471 9456 72480
rect 9404 72437 9413 72471
rect 9413 72437 9447 72471
rect 9447 72437 9456 72471
rect 9404 72428 9456 72437
rect 3610 72326 3662 72378
rect 3674 72326 3726 72378
rect 3738 72326 3790 72378
rect 3802 72326 3854 72378
rect 3866 72326 3918 72378
rect 5210 72326 5262 72378
rect 5274 72326 5326 72378
rect 5338 72326 5390 72378
rect 5402 72326 5454 72378
rect 5466 72326 5518 72378
rect 6810 72326 6862 72378
rect 6874 72326 6926 72378
rect 6938 72326 6990 72378
rect 7002 72326 7054 72378
rect 7066 72326 7118 72378
rect 8410 72326 8462 72378
rect 8474 72326 8526 72378
rect 8538 72326 8590 72378
rect 8602 72326 8654 72378
rect 8666 72326 8718 72378
rect 5540 72224 5592 72276
rect 6460 72088 6512 72140
rect 5540 72020 5592 72072
rect 940 71952 992 72004
rect 5724 72020 5776 72072
rect 6276 71952 6328 72004
rect 7196 72088 7248 72140
rect 7656 72224 7708 72276
rect 7932 72156 7984 72208
rect 9772 72156 9824 72208
rect 8576 72088 8628 72140
rect 1584 71927 1636 71936
rect 1584 71893 1593 71927
rect 1593 71893 1627 71927
rect 1627 71893 1636 71927
rect 1584 71884 1636 71893
rect 6000 71884 6052 71936
rect 8024 72020 8076 72072
rect 8392 71884 8444 71936
rect 2950 71782 3002 71834
rect 3014 71782 3066 71834
rect 3078 71782 3130 71834
rect 3142 71782 3194 71834
rect 3206 71782 3258 71834
rect 4550 71782 4602 71834
rect 4614 71782 4666 71834
rect 4678 71782 4730 71834
rect 4742 71782 4794 71834
rect 4806 71782 4858 71834
rect 6150 71782 6202 71834
rect 6214 71782 6266 71834
rect 6278 71782 6330 71834
rect 6342 71782 6394 71834
rect 6406 71782 6458 71834
rect 7750 71782 7802 71834
rect 7814 71782 7866 71834
rect 7878 71782 7930 71834
rect 7942 71782 7994 71834
rect 8006 71782 8058 71834
rect 9350 71782 9402 71834
rect 9414 71782 9466 71834
rect 9478 71782 9530 71834
rect 9542 71782 9594 71834
rect 9606 71782 9658 71834
rect 4344 71680 4396 71732
rect 6828 71680 6880 71732
rect 7288 71680 7340 71732
rect 664 71612 716 71664
rect 1124 71612 1176 71664
rect 4896 71612 4948 71664
rect 940 71544 992 71596
rect 6368 71587 6420 71596
rect 6368 71553 6377 71587
rect 6377 71553 6411 71587
rect 6411 71553 6420 71587
rect 6368 71544 6420 71553
rect 6460 71544 6512 71596
rect 7104 71544 7156 71596
rect 7196 71544 7248 71596
rect 7748 71544 7800 71596
rect 9128 71612 9180 71664
rect 10876 71680 10928 71732
rect 11336 71680 11388 71732
rect 8208 71587 8260 71596
rect 8208 71553 8217 71587
rect 8217 71553 8251 71587
rect 8251 71553 8260 71587
rect 8208 71544 8260 71553
rect 1124 71476 1176 71528
rect 1308 71476 1360 71528
rect 7380 71476 7432 71528
rect 9036 71544 9088 71596
rect 8576 71476 8628 71528
rect 11152 71476 11204 71528
rect 9036 71408 9088 71460
rect 572 71340 624 71392
rect 5540 71340 5592 71392
rect 6736 71340 6788 71392
rect 7104 71340 7156 71392
rect 7932 71340 7984 71392
rect 11244 71340 11296 71392
rect 3610 71238 3662 71290
rect 3674 71238 3726 71290
rect 3738 71238 3790 71290
rect 3802 71238 3854 71290
rect 3866 71238 3918 71290
rect 5210 71238 5262 71290
rect 5274 71238 5326 71290
rect 5338 71238 5390 71290
rect 5402 71238 5454 71290
rect 5466 71238 5518 71290
rect 6810 71238 6862 71290
rect 6874 71238 6926 71290
rect 6938 71238 6990 71290
rect 7002 71238 7054 71290
rect 7066 71238 7118 71290
rect 8410 71238 8462 71290
rect 8474 71238 8526 71290
rect 8538 71238 8590 71290
rect 8602 71238 8654 71290
rect 8666 71238 8718 71290
rect 6460 71136 6512 71188
rect 6920 71136 6972 71188
rect 7012 71136 7064 71188
rect 7288 71136 7340 71188
rect 7840 71136 7892 71188
rect 6828 71068 6880 71120
rect 7564 71068 7616 71120
rect 9772 71068 9824 71120
rect 5724 71000 5776 71052
rect 7932 71000 7984 71052
rect 8392 71000 8444 71052
rect 8484 71043 8536 71052
rect 8484 71009 8493 71043
rect 8493 71009 8527 71043
rect 8527 71009 8536 71043
rect 8484 71000 8536 71009
rect 9220 71000 9272 71052
rect 5540 70932 5592 70984
rect 6552 70975 6604 70984
rect 6552 70941 6561 70975
rect 6561 70941 6595 70975
rect 6595 70941 6604 70975
rect 6552 70932 6604 70941
rect 7012 70932 7064 70984
rect 7104 70932 7156 70984
rect 10232 70932 10284 70984
rect 2780 70864 2832 70916
rect 8576 70864 8628 70916
rect 2412 70796 2464 70848
rect 3516 70796 3568 70848
rect 7196 70796 7248 70848
rect 7380 70796 7432 70848
rect 8484 70796 8536 70848
rect 8852 70796 8904 70848
rect 9128 70796 9180 70848
rect 2950 70694 3002 70746
rect 3014 70694 3066 70746
rect 3078 70694 3130 70746
rect 3142 70694 3194 70746
rect 3206 70694 3258 70746
rect 4550 70694 4602 70746
rect 4614 70694 4666 70746
rect 4678 70694 4730 70746
rect 4742 70694 4794 70746
rect 4806 70694 4858 70746
rect 6150 70694 6202 70746
rect 6214 70694 6266 70746
rect 6278 70694 6330 70746
rect 6342 70694 6394 70746
rect 6406 70694 6458 70746
rect 7750 70694 7802 70746
rect 7814 70694 7866 70746
rect 7878 70694 7930 70746
rect 7942 70694 7994 70746
rect 8006 70694 8058 70746
rect 9350 70694 9402 70746
rect 9414 70694 9466 70746
rect 9478 70694 9530 70746
rect 9542 70694 9594 70746
rect 9606 70694 9658 70746
rect 664 70592 716 70644
rect 6368 70592 6420 70644
rect 6828 70592 6880 70644
rect 6552 70524 6604 70576
rect 7012 70524 7064 70576
rect 1400 70499 1452 70508
rect 1400 70465 1409 70499
rect 1409 70465 1443 70499
rect 1443 70465 1452 70499
rect 1400 70456 1452 70465
rect 2044 70456 2096 70508
rect 3516 70456 3568 70508
rect 4344 70456 4396 70508
rect 6460 70456 6512 70508
rect 6920 70456 6972 70508
rect 7104 70499 7156 70508
rect 7104 70465 7113 70499
rect 7113 70465 7147 70499
rect 7147 70465 7156 70499
rect 7104 70456 7156 70465
rect 7748 70592 7800 70644
rect 8576 70592 8628 70644
rect 9128 70592 9180 70644
rect 10048 70592 10100 70644
rect 6000 70388 6052 70440
rect 5724 70320 5776 70372
rect 5816 70320 5868 70372
rect 1308 70252 1360 70304
rect 4436 70252 4488 70304
rect 4712 70252 4764 70304
rect 6092 70252 6144 70304
rect 6184 70252 6236 70304
rect 7380 70456 7432 70508
rect 7656 70456 7708 70508
rect 7656 70295 7708 70304
rect 7656 70261 7665 70295
rect 7665 70261 7699 70295
rect 7699 70261 7708 70295
rect 7656 70252 7708 70261
rect 8024 70320 8076 70372
rect 8208 70456 8260 70508
rect 8392 70456 8444 70508
rect 8576 70499 8628 70508
rect 8576 70465 8585 70499
rect 8585 70465 8619 70499
rect 8619 70465 8628 70499
rect 8576 70456 8628 70465
rect 9404 70524 9456 70576
rect 11428 70524 11480 70576
rect 9220 70456 9272 70508
rect 11336 70456 11388 70508
rect 9588 70320 9640 70372
rect 11520 70320 11572 70372
rect 3610 70150 3662 70202
rect 3674 70150 3726 70202
rect 3738 70150 3790 70202
rect 3802 70150 3854 70202
rect 3866 70150 3918 70202
rect 5210 70150 5262 70202
rect 5274 70150 5326 70202
rect 5338 70150 5390 70202
rect 5402 70150 5454 70202
rect 5466 70150 5518 70202
rect 6810 70150 6862 70202
rect 6874 70150 6926 70202
rect 6938 70150 6990 70202
rect 7002 70150 7054 70202
rect 7066 70150 7118 70202
rect 8410 70150 8462 70202
rect 8474 70150 8526 70202
rect 8538 70150 8590 70202
rect 8602 70150 8654 70202
rect 8666 70150 8718 70202
rect 4988 70048 5040 70100
rect 5172 70048 5224 70100
rect 5724 70091 5776 70100
rect 5724 70057 5733 70091
rect 5733 70057 5767 70091
rect 5767 70057 5776 70091
rect 5724 70048 5776 70057
rect 6184 70048 6236 70100
rect 6368 70091 6420 70100
rect 6368 70057 6377 70091
rect 6377 70057 6411 70091
rect 6411 70057 6420 70091
rect 6368 70048 6420 70057
rect 6920 70048 6972 70100
rect 9036 70048 9088 70100
rect 4620 69912 4672 69964
rect 7196 69980 7248 70032
rect 7288 69980 7340 70032
rect 6184 69912 6236 69964
rect 6828 69912 6880 69964
rect 5448 69844 5500 69896
rect 4252 69776 4304 69828
rect 4712 69776 4764 69828
rect 4988 69776 5040 69828
rect 7196 69844 7248 69896
rect 7288 69887 7340 69896
rect 7288 69853 7297 69887
rect 7297 69853 7331 69887
rect 7331 69853 7340 69887
rect 7288 69844 7340 69853
rect 7380 69844 7432 69896
rect 7932 69912 7984 69964
rect 8208 69980 8260 70032
rect 8392 69980 8444 70032
rect 9312 70048 9364 70100
rect 9588 70048 9640 70100
rect 8668 69912 8720 69964
rect 9220 69912 9272 69964
rect 9680 69912 9732 69964
rect 10876 69912 10928 69964
rect 6736 69776 6788 69828
rect 5448 69708 5500 69760
rect 6092 69708 6144 69760
rect 6276 69708 6328 69760
rect 7104 69708 7156 69760
rect 7748 69708 7800 69760
rect 8484 69887 8536 69896
rect 8484 69853 8503 69887
rect 8503 69853 8536 69887
rect 8484 69844 8536 69853
rect 9680 69776 9732 69828
rect 8484 69708 8536 69760
rect 9220 69708 9272 69760
rect 9588 69708 9640 69760
rect 10968 69708 11020 69760
rect 2950 69606 3002 69658
rect 3014 69606 3066 69658
rect 3078 69606 3130 69658
rect 3142 69606 3194 69658
rect 3206 69606 3258 69658
rect 4550 69606 4602 69658
rect 4614 69606 4666 69658
rect 4678 69606 4730 69658
rect 4742 69606 4794 69658
rect 4806 69606 4858 69658
rect 6150 69606 6202 69658
rect 6214 69606 6266 69658
rect 6278 69606 6330 69658
rect 6342 69606 6394 69658
rect 6406 69606 6458 69658
rect 7750 69606 7802 69658
rect 7814 69606 7866 69658
rect 7878 69606 7930 69658
rect 7942 69606 7994 69658
rect 8006 69606 8058 69658
rect 9350 69606 9402 69658
rect 9414 69606 9466 69658
rect 9478 69606 9530 69658
rect 9542 69606 9594 69658
rect 9606 69606 9658 69658
rect 4344 69504 4396 69556
rect 4804 69504 4856 69556
rect 5172 69504 5224 69556
rect 6552 69504 6604 69556
rect 6828 69547 6880 69556
rect 6828 69513 6837 69547
rect 6837 69513 6871 69547
rect 6871 69513 6880 69547
rect 6828 69504 6880 69513
rect 6920 69504 6972 69556
rect 7748 69504 7800 69556
rect 8760 69504 8812 69556
rect 10784 69504 10836 69556
rect 8024 69436 8076 69488
rect 8208 69436 8260 69488
rect 8576 69436 8628 69488
rect 940 69368 992 69420
rect 1584 69368 1636 69420
rect 6368 69368 6420 69420
rect 2136 69232 2188 69284
rect 7104 69368 7156 69420
rect 6920 69343 6972 69352
rect 6920 69309 6929 69343
rect 6929 69309 6963 69343
rect 6963 69309 6972 69343
rect 6920 69300 6972 69309
rect 7380 69368 7432 69420
rect 9128 69411 9180 69420
rect 9128 69377 9137 69411
rect 9137 69377 9171 69411
rect 9171 69377 9180 69411
rect 9128 69368 9180 69377
rect 9312 69411 9364 69420
rect 9312 69377 9321 69411
rect 9321 69377 9355 69411
rect 9355 69377 9364 69411
rect 9312 69368 9364 69377
rect 9404 69411 9456 69420
rect 9404 69377 9413 69411
rect 9413 69377 9447 69411
rect 9447 69377 9456 69411
rect 9404 69368 9456 69377
rect 9956 69368 10008 69420
rect 7932 69300 7984 69352
rect 8392 69300 8444 69352
rect 6552 69232 6604 69284
rect 4620 69164 4672 69216
rect 4712 69164 4764 69216
rect 5448 69164 5500 69216
rect 6092 69164 6144 69216
rect 6460 69164 6512 69216
rect 6920 69164 6972 69216
rect 8208 69164 8260 69216
rect 9036 69164 9088 69216
rect 3610 69062 3662 69114
rect 3674 69062 3726 69114
rect 3738 69062 3790 69114
rect 3802 69062 3854 69114
rect 3866 69062 3918 69114
rect 5210 69062 5262 69114
rect 5274 69062 5326 69114
rect 5338 69062 5390 69114
rect 5402 69062 5454 69114
rect 5466 69062 5518 69114
rect 6810 69062 6862 69114
rect 6874 69062 6926 69114
rect 6938 69062 6990 69114
rect 7002 69062 7054 69114
rect 7066 69062 7118 69114
rect 8410 69062 8462 69114
rect 8474 69062 8526 69114
rect 8538 69062 8590 69114
rect 8602 69062 8654 69114
rect 8666 69062 8718 69114
rect 4252 69003 4304 69012
rect 4252 68969 4261 69003
rect 4261 68969 4295 69003
rect 4295 68969 4304 69003
rect 4252 68960 4304 68969
rect 4344 68960 4396 69012
rect 5356 68892 5408 68944
rect 5908 68892 5960 68944
rect 7012 68892 7064 68944
rect 7104 68892 7156 68944
rect 7564 68960 7616 69012
rect 8484 68960 8536 69012
rect 9404 68960 9456 69012
rect 3884 68824 3936 68876
rect 4344 68799 4396 68808
rect 4344 68765 4353 68799
rect 4353 68765 4387 68799
rect 4387 68765 4396 68799
rect 4344 68756 4396 68765
rect 5816 68756 5868 68808
rect 4712 68688 4764 68740
rect 4804 68688 4856 68740
rect 5264 68688 5316 68740
rect 4252 68620 4304 68672
rect 4620 68620 4672 68672
rect 5172 68620 5224 68672
rect 5540 68620 5592 68672
rect 6092 68620 6144 68672
rect 6460 68756 6512 68808
rect 6736 68756 6788 68808
rect 7012 68756 7064 68808
rect 8576 68892 8628 68944
rect 9036 68824 9088 68876
rect 8392 68756 8444 68808
rect 7932 68688 7984 68740
rect 9312 68688 9364 68740
rect 6736 68620 6788 68672
rect 8024 68620 8076 68672
rect 8392 68620 8444 68672
rect 9128 68663 9180 68672
rect 9128 68629 9137 68663
rect 9137 68629 9171 68663
rect 9171 68629 9180 68663
rect 9128 68620 9180 68629
rect 2950 68518 3002 68570
rect 3014 68518 3066 68570
rect 3078 68518 3130 68570
rect 3142 68518 3194 68570
rect 3206 68518 3258 68570
rect 4550 68518 4602 68570
rect 4614 68518 4666 68570
rect 4678 68518 4730 68570
rect 4742 68518 4794 68570
rect 4806 68518 4858 68570
rect 6150 68518 6202 68570
rect 6214 68518 6266 68570
rect 6278 68518 6330 68570
rect 6342 68518 6394 68570
rect 6406 68518 6458 68570
rect 7750 68518 7802 68570
rect 7814 68518 7866 68570
rect 7878 68518 7930 68570
rect 7942 68518 7994 68570
rect 8006 68518 8058 68570
rect 9350 68518 9402 68570
rect 9414 68518 9466 68570
rect 9478 68518 9530 68570
rect 9542 68518 9594 68570
rect 9606 68518 9658 68570
rect 4988 68459 5040 68468
rect 4988 68425 4997 68459
rect 4997 68425 5031 68459
rect 5031 68425 5040 68459
rect 4988 68416 5040 68425
rect 5264 68416 5316 68468
rect 6276 68416 6328 68468
rect 6736 68416 6788 68468
rect 7932 68416 7984 68468
rect 8944 68416 8996 68468
rect 5080 68348 5132 68400
rect 940 68280 992 68332
rect 4528 68280 4580 68332
rect 4804 68323 4856 68332
rect 4804 68289 4813 68323
rect 4813 68289 4847 68323
rect 4847 68289 4856 68323
rect 4804 68280 4856 68289
rect 5632 68348 5684 68400
rect 6460 68280 6512 68332
rect 4436 68212 4488 68264
rect 6184 68212 6236 68264
rect 7012 68348 7064 68400
rect 848 68144 900 68196
rect 296 68076 348 68128
rect 2504 68076 2556 68128
rect 2872 68076 2924 68128
rect 3884 68076 3936 68128
rect 4436 68119 4488 68128
rect 4436 68085 4445 68119
rect 4445 68085 4479 68119
rect 4479 68085 4488 68119
rect 4436 68076 4488 68085
rect 5356 68144 5408 68196
rect 5724 68144 5776 68196
rect 6552 68144 6604 68196
rect 6828 68144 6880 68196
rect 7380 68280 7432 68332
rect 7932 68326 7984 68332
rect 7932 68292 7940 68326
rect 7940 68292 7974 68326
rect 7974 68292 7984 68326
rect 7932 68280 7984 68292
rect 8024 68323 8076 68332
rect 8024 68289 8033 68323
rect 8033 68289 8067 68323
rect 8067 68289 8076 68323
rect 8024 68280 8076 68289
rect 8944 68280 8996 68332
rect 11888 68280 11940 68332
rect 9128 68212 9180 68264
rect 11796 68212 11848 68264
rect 11520 68144 11572 68196
rect 8024 68076 8076 68128
rect 8392 68076 8444 68128
rect 3610 67974 3662 68026
rect 3674 67974 3726 68026
rect 3738 67974 3790 68026
rect 3802 67974 3854 68026
rect 3866 67974 3918 68026
rect 5210 67974 5262 68026
rect 5274 67974 5326 68026
rect 5338 67974 5390 68026
rect 5402 67974 5454 68026
rect 5466 67974 5518 68026
rect 6810 67974 6862 68026
rect 6874 67974 6926 68026
rect 6938 67974 6990 68026
rect 7002 67974 7054 68026
rect 7066 67974 7118 68026
rect 8410 67974 8462 68026
rect 8474 67974 8526 68026
rect 8538 67974 8590 68026
rect 8602 67974 8654 68026
rect 8666 67974 8718 68026
rect 4896 67872 4948 67924
rect 5080 67872 5132 67924
rect 5264 67872 5316 67924
rect 5356 67872 5408 67924
rect 7932 67872 7984 67924
rect 9036 67872 9088 67924
rect 4252 67804 4304 67856
rect 5908 67804 5960 67856
rect 756 67736 808 67788
rect 4620 67736 4672 67788
rect 6552 67736 6604 67788
rect 5540 67668 5592 67720
rect 6092 67668 6144 67720
rect 7472 67736 7524 67788
rect 1492 67643 1544 67652
rect 1492 67609 1501 67643
rect 1501 67609 1535 67643
rect 1535 67609 1544 67643
rect 1492 67600 1544 67609
rect 2320 67600 2372 67652
rect 4804 67600 4856 67652
rect 5080 67600 5132 67652
rect 5448 67600 5500 67652
rect 7380 67668 7432 67720
rect 8300 67736 8352 67788
rect 8392 67736 8444 67788
rect 9220 67736 9272 67788
rect 6920 67600 6972 67652
rect 7012 67600 7064 67652
rect 7104 67600 7156 67652
rect 8760 67668 8812 67720
rect 10784 67600 10836 67652
rect 8576 67532 8628 67584
rect 2950 67430 3002 67482
rect 3014 67430 3066 67482
rect 3078 67430 3130 67482
rect 3142 67430 3194 67482
rect 3206 67430 3258 67482
rect 4550 67430 4602 67482
rect 4614 67430 4666 67482
rect 4678 67430 4730 67482
rect 4742 67430 4794 67482
rect 4806 67430 4858 67482
rect 6150 67430 6202 67482
rect 6214 67430 6266 67482
rect 6278 67430 6330 67482
rect 6342 67430 6394 67482
rect 6406 67430 6458 67482
rect 7750 67430 7802 67482
rect 7814 67430 7866 67482
rect 7878 67430 7930 67482
rect 7942 67430 7994 67482
rect 8006 67430 8058 67482
rect 9350 67430 9402 67482
rect 9414 67430 9466 67482
rect 9478 67430 9530 67482
rect 9542 67430 9594 67482
rect 9606 67430 9658 67482
rect 5264 67328 5316 67380
rect 5908 67328 5960 67380
rect 6460 67328 6512 67380
rect 6552 67328 6604 67380
rect 7012 67328 7064 67380
rect 4344 67260 4396 67312
rect 3884 67192 3936 67244
rect 4620 67192 4672 67244
rect 4252 67167 4304 67176
rect 4252 67133 4261 67167
rect 4261 67133 4295 67167
rect 4295 67133 4304 67167
rect 4252 67124 4304 67133
rect 4712 67124 4764 67176
rect 5356 67192 5408 67244
rect 7196 67192 7248 67244
rect 6092 67124 6144 67176
rect 6736 67124 6788 67176
rect 9128 67328 9180 67380
rect 10324 67328 10376 67380
rect 7380 67260 7432 67312
rect 7656 67192 7708 67244
rect 7748 67192 7800 67244
rect 8760 67192 8812 67244
rect 10140 67192 10192 67244
rect 7932 67124 7984 67176
rect 8484 67124 8536 67176
rect 9036 67124 9088 67176
rect 9128 67167 9180 67176
rect 9128 67133 9137 67167
rect 9137 67133 9171 67167
rect 9171 67133 9180 67167
rect 9128 67124 9180 67133
rect 6000 67056 6052 67108
rect 5080 66988 5132 67040
rect 5448 66988 5500 67040
rect 5908 66988 5960 67040
rect 6736 66988 6788 67040
rect 7656 67056 7708 67108
rect 7840 67099 7892 67108
rect 7840 67065 7849 67099
rect 7849 67065 7883 67099
rect 7883 67065 7892 67099
rect 7840 67056 7892 67065
rect 9404 67124 9456 67176
rect 9864 67124 9916 67176
rect 9864 66988 9916 67040
rect 10600 66988 10652 67040
rect 3610 66886 3662 66938
rect 3674 66886 3726 66938
rect 3738 66886 3790 66938
rect 3802 66886 3854 66938
rect 3866 66886 3918 66938
rect 5210 66886 5262 66938
rect 5274 66886 5326 66938
rect 5338 66886 5390 66938
rect 5402 66886 5454 66938
rect 5466 66886 5518 66938
rect 6810 66886 6862 66938
rect 6874 66886 6926 66938
rect 6938 66886 6990 66938
rect 7002 66886 7054 66938
rect 7066 66886 7118 66938
rect 8410 66886 8462 66938
rect 8474 66886 8526 66938
rect 8538 66886 8590 66938
rect 8602 66886 8654 66938
rect 8666 66886 8718 66938
rect 1032 66784 1084 66836
rect 4896 66716 4948 66768
rect 5172 66716 5224 66768
rect 5356 66716 5408 66768
rect 5908 66716 5960 66768
rect 4528 66648 4580 66700
rect 7196 66716 7248 66768
rect 6460 66648 6512 66700
rect 3976 66580 4028 66632
rect 5908 66580 5960 66632
rect 7012 66580 7064 66632
rect 7380 66623 7432 66632
rect 940 66512 992 66564
rect 4252 66512 4304 66564
rect 5264 66512 5316 66564
rect 6184 66512 6236 66564
rect 6552 66512 6604 66564
rect 7380 66589 7388 66623
rect 7388 66589 7422 66623
rect 7422 66589 7432 66623
rect 7380 66580 7432 66589
rect 8484 66784 8536 66836
rect 9220 66784 9272 66836
rect 7932 66716 7984 66768
rect 8116 66648 8168 66700
rect 8576 66648 8628 66700
rect 9036 66648 9088 66700
rect 4436 66444 4488 66496
rect 6092 66444 6144 66496
rect 7196 66444 7248 66496
rect 7748 66444 7800 66496
rect 8944 66580 8996 66632
rect 9220 66623 9272 66632
rect 9220 66589 9243 66623
rect 9243 66589 9272 66623
rect 9220 66580 9272 66589
rect 9312 66623 9364 66632
rect 9312 66589 9321 66623
rect 9321 66589 9355 66623
rect 9355 66589 9364 66623
rect 9312 66580 9364 66589
rect 9588 66623 9640 66632
rect 9588 66589 9597 66623
rect 9597 66589 9631 66623
rect 9631 66589 9640 66623
rect 9588 66580 9640 66589
rect 10692 66580 10744 66632
rect 8392 66444 8444 66496
rect 8760 66444 8812 66496
rect 8944 66487 8996 66496
rect 8944 66453 8953 66487
rect 8953 66453 8987 66487
rect 8987 66453 8996 66487
rect 8944 66444 8996 66453
rect 11428 66444 11480 66496
rect 2950 66342 3002 66394
rect 3014 66342 3066 66394
rect 3078 66342 3130 66394
rect 3142 66342 3194 66394
rect 3206 66342 3258 66394
rect 4550 66342 4602 66394
rect 4614 66342 4666 66394
rect 4678 66342 4730 66394
rect 4742 66342 4794 66394
rect 4806 66342 4858 66394
rect 6150 66342 6202 66394
rect 6214 66342 6266 66394
rect 6278 66342 6330 66394
rect 6342 66342 6394 66394
rect 6406 66342 6458 66394
rect 7750 66342 7802 66394
rect 7814 66342 7866 66394
rect 7878 66342 7930 66394
rect 7942 66342 7994 66394
rect 8006 66342 8058 66394
rect 9350 66342 9402 66394
rect 9414 66342 9466 66394
rect 9478 66342 9530 66394
rect 9542 66342 9594 66394
rect 9606 66342 9658 66394
rect 4344 66240 4396 66292
rect 5540 66240 5592 66292
rect 4988 66172 5040 66224
rect 5724 66172 5776 66224
rect 7656 66240 7708 66292
rect 7840 66240 7892 66292
rect 8024 66240 8076 66292
rect 8392 66240 8444 66292
rect 8668 66240 8720 66292
rect 9128 66240 9180 66292
rect 9312 66240 9364 66292
rect 9864 66240 9916 66292
rect 5172 66147 5224 66156
rect 5172 66113 5181 66147
rect 5181 66113 5215 66147
rect 5215 66113 5224 66147
rect 5172 66104 5224 66113
rect 5356 66147 5408 66156
rect 5356 66113 5365 66147
rect 5365 66113 5399 66147
rect 5399 66113 5408 66147
rect 5356 66104 5408 66113
rect 5816 66147 5868 66156
rect 5816 66113 5825 66147
rect 5825 66113 5859 66147
rect 5859 66113 5868 66147
rect 5816 66104 5868 66113
rect 6000 66104 6052 66156
rect 4988 66036 5040 66088
rect 5264 66036 5316 66088
rect 6276 66036 6328 66088
rect 7932 66172 7984 66224
rect 7288 66147 7340 66156
rect 7288 66113 7294 66147
rect 7294 66113 7328 66147
rect 7328 66113 7340 66147
rect 7288 66104 7340 66113
rect 7840 66147 7892 66156
rect 7840 66113 7849 66147
rect 7849 66113 7883 66147
rect 7883 66113 7892 66147
rect 7840 66104 7892 66113
rect 7564 66079 7616 66088
rect 7564 66045 7573 66079
rect 7573 66045 7607 66079
rect 7607 66045 7616 66079
rect 7564 66036 7616 66045
rect 3976 65968 4028 66020
rect 5816 65968 5868 66020
rect 8300 66036 8352 66088
rect 8852 66104 8904 66156
rect 9036 66104 9088 66156
rect 7012 65900 7064 65952
rect 8392 65968 8444 66020
rect 8852 65968 8904 66020
rect 9036 65968 9088 66020
rect 10968 66172 11020 66224
rect 9864 65900 9916 65952
rect 3610 65798 3662 65850
rect 3674 65798 3726 65850
rect 3738 65798 3790 65850
rect 3802 65798 3854 65850
rect 3866 65798 3918 65850
rect 5210 65798 5262 65850
rect 5274 65798 5326 65850
rect 5338 65798 5390 65850
rect 5402 65798 5454 65850
rect 5466 65798 5518 65850
rect 6810 65798 6862 65850
rect 6874 65798 6926 65850
rect 6938 65798 6990 65850
rect 7002 65798 7054 65850
rect 7066 65798 7118 65850
rect 8410 65798 8462 65850
rect 8474 65798 8526 65850
rect 8538 65798 8590 65850
rect 8602 65798 8654 65850
rect 8666 65798 8718 65850
rect 3332 65696 3384 65748
rect 5632 65696 5684 65748
rect 7104 65696 7156 65748
rect 7472 65696 7524 65748
rect 7564 65696 7616 65748
rect 7932 65696 7984 65748
rect 2412 65628 2464 65680
rect 3608 65628 3660 65680
rect 4896 65560 4948 65612
rect 5724 65560 5776 65612
rect 2412 65492 2464 65544
rect 2688 65492 2740 65544
rect 3516 65492 3568 65544
rect 6000 65492 6052 65544
rect 7288 65560 7340 65612
rect 7472 65560 7524 65612
rect 940 65424 992 65476
rect 2136 65424 2188 65476
rect 2780 65424 2832 65476
rect 3332 65424 3384 65476
rect 5080 65467 5132 65476
rect 5080 65433 5089 65467
rect 5089 65433 5123 65467
rect 5123 65433 5132 65467
rect 5080 65424 5132 65433
rect 5632 65424 5684 65476
rect 7012 65424 7064 65476
rect 9956 65424 10008 65476
rect 296 65356 348 65408
rect 1216 65356 1268 65408
rect 4620 65356 4672 65408
rect 5172 65399 5224 65408
rect 5172 65365 5181 65399
rect 5181 65365 5215 65399
rect 5215 65365 5224 65399
rect 5172 65356 5224 65365
rect 6276 65356 6328 65408
rect 6828 65356 6880 65408
rect 7288 65399 7340 65408
rect 7288 65365 7297 65399
rect 7297 65365 7331 65399
rect 7331 65365 7340 65399
rect 7288 65356 7340 65365
rect 7564 65356 7616 65408
rect 8024 65356 8076 65408
rect 8484 65356 8536 65408
rect 9312 65356 9364 65408
rect 2950 65254 3002 65306
rect 3014 65254 3066 65306
rect 3078 65254 3130 65306
rect 3142 65254 3194 65306
rect 3206 65254 3258 65306
rect 4550 65254 4602 65306
rect 4614 65254 4666 65306
rect 4678 65254 4730 65306
rect 4742 65254 4794 65306
rect 4806 65254 4858 65306
rect 6150 65254 6202 65306
rect 6214 65254 6266 65306
rect 6278 65254 6330 65306
rect 6342 65254 6394 65306
rect 6406 65254 6458 65306
rect 7750 65254 7802 65306
rect 7814 65254 7866 65306
rect 7878 65254 7930 65306
rect 7942 65254 7994 65306
rect 8006 65254 8058 65306
rect 9350 65254 9402 65306
rect 9414 65254 9466 65306
rect 9478 65254 9530 65306
rect 9542 65254 9594 65306
rect 9606 65254 9658 65306
rect 10048 65288 10100 65340
rect 10324 65288 10376 65340
rect 5080 65152 5132 65204
rect 9128 65152 9180 65204
rect 2504 65084 2556 65136
rect 2596 65016 2648 65068
rect 2136 64948 2188 65000
rect 4712 65016 4764 65068
rect 6552 65016 6604 65068
rect 7472 65059 7524 65068
rect 7472 65025 7481 65059
rect 7481 65025 7515 65059
rect 7515 65025 7524 65059
rect 7472 65016 7524 65025
rect 3240 64948 3292 65000
rect 5172 64948 5224 65000
rect 7656 65059 7708 65068
rect 7656 65025 7665 65059
rect 7665 65025 7699 65059
rect 7699 65025 7708 65059
rect 7656 65016 7708 65025
rect 8024 65059 8076 65068
rect 8024 65025 8033 65059
rect 8033 65025 8067 65059
rect 8067 65025 8076 65059
rect 8024 65016 8076 65025
rect 8208 65016 8260 65068
rect 8484 65016 8536 65068
rect 9864 65016 9916 65068
rect 10232 65016 10284 65068
rect 5356 64880 5408 64932
rect 6092 64880 6144 64932
rect 7104 64880 7156 64932
rect 7656 64880 7708 64932
rect 2872 64812 2924 64864
rect 4160 64812 4212 64864
rect 4896 64812 4948 64864
rect 5080 64812 5132 64864
rect 6552 64812 6604 64864
rect 6828 64812 6880 64864
rect 7472 64812 7524 64864
rect 8300 64948 8352 65000
rect 8760 64948 8812 65000
rect 9036 64948 9088 65000
rect 9312 64991 9364 65000
rect 9312 64957 9321 64991
rect 9321 64957 9355 64991
rect 9355 64957 9364 64991
rect 9312 64948 9364 64957
rect 9496 64991 9548 65000
rect 9496 64957 9505 64991
rect 9505 64957 9539 64991
rect 9539 64957 9548 64991
rect 9496 64948 9548 64957
rect 11152 64948 11204 65000
rect 10140 64880 10192 64932
rect 9496 64812 9548 64864
rect 3610 64710 3662 64762
rect 3674 64710 3726 64762
rect 3738 64710 3790 64762
rect 3802 64710 3854 64762
rect 3866 64710 3918 64762
rect 5210 64710 5262 64762
rect 5274 64710 5326 64762
rect 5338 64710 5390 64762
rect 5402 64710 5454 64762
rect 5466 64710 5518 64762
rect 6810 64710 6862 64762
rect 6874 64710 6926 64762
rect 6938 64710 6990 64762
rect 7002 64710 7054 64762
rect 7066 64710 7118 64762
rect 8410 64710 8462 64762
rect 8474 64710 8526 64762
rect 8538 64710 8590 64762
rect 8602 64710 8654 64762
rect 8666 64710 8718 64762
rect 2412 64608 2464 64660
rect 2780 64608 2832 64660
rect 4804 64608 4856 64660
rect 5172 64608 5224 64660
rect 4160 64472 4212 64524
rect 5080 64472 5132 64524
rect 5724 64515 5776 64524
rect 5724 64481 5733 64515
rect 5733 64481 5767 64515
rect 5767 64481 5776 64515
rect 5724 64472 5776 64481
rect 7472 64472 7524 64524
rect 8576 64515 8628 64524
rect 8576 64481 8585 64515
rect 8585 64481 8619 64515
rect 8619 64481 8628 64515
rect 8576 64472 8628 64481
rect 8668 64472 8720 64524
rect 9036 64472 9088 64524
rect 2688 64404 2740 64456
rect 3240 64404 3292 64456
rect 5816 64404 5868 64456
rect 7104 64404 7156 64456
rect 8024 64404 8076 64456
rect 10416 64404 10468 64456
rect 940 64336 992 64388
rect 8852 64336 8904 64388
rect 9036 64336 9088 64388
rect 1584 64311 1636 64320
rect 1584 64277 1593 64311
rect 1593 64277 1627 64311
rect 1627 64277 1636 64311
rect 1584 64268 1636 64277
rect 4712 64268 4764 64320
rect 5080 64268 5132 64320
rect 5816 64268 5868 64320
rect 6092 64268 6144 64320
rect 7564 64268 7616 64320
rect 8024 64311 8076 64320
rect 8024 64277 8033 64311
rect 8033 64277 8067 64311
rect 8067 64277 8076 64311
rect 8024 64268 8076 64277
rect 9128 64268 9180 64320
rect 9864 64268 9916 64320
rect 2950 64166 3002 64218
rect 3014 64166 3066 64218
rect 3078 64166 3130 64218
rect 3142 64166 3194 64218
rect 3206 64166 3258 64218
rect 4550 64166 4602 64218
rect 4614 64166 4666 64218
rect 4678 64166 4730 64218
rect 4742 64166 4794 64218
rect 4806 64166 4858 64218
rect 6150 64166 6202 64218
rect 6214 64166 6266 64218
rect 6278 64166 6330 64218
rect 6342 64166 6394 64218
rect 6406 64166 6458 64218
rect 7750 64166 7802 64218
rect 7814 64166 7866 64218
rect 7878 64166 7930 64218
rect 7942 64166 7994 64218
rect 8006 64166 8058 64218
rect 9350 64166 9402 64218
rect 9414 64166 9466 64218
rect 9478 64166 9530 64218
rect 9542 64166 9594 64218
rect 9606 64166 9658 64218
rect 1584 64064 1636 64116
rect 4804 64064 4856 64116
rect 5172 64064 5224 64116
rect 5816 64064 5868 64116
rect 6276 64064 6328 64116
rect 8852 64107 8904 64116
rect 8852 64073 8861 64107
rect 8861 64073 8895 64107
rect 8895 64073 8904 64107
rect 8852 64064 8904 64073
rect 11704 64064 11756 64116
rect 1492 63971 1544 63980
rect 1492 63937 1501 63971
rect 1501 63937 1535 63971
rect 1535 63937 1544 63971
rect 1492 63928 1544 63937
rect 5724 63928 5776 63980
rect 6092 63928 6144 63980
rect 7196 63928 7248 63980
rect 7748 63928 7800 63980
rect 7932 63928 7984 63980
rect 8300 63928 8352 63980
rect 8576 63860 8628 63912
rect 8668 63860 8720 63912
rect 10600 63928 10652 63980
rect 8300 63792 8352 63844
rect 1584 63767 1636 63776
rect 1584 63733 1593 63767
rect 1593 63733 1627 63767
rect 1627 63733 1636 63767
rect 1584 63724 1636 63733
rect 5540 63724 5592 63776
rect 5816 63724 5868 63776
rect 6368 63724 6420 63776
rect 6828 63724 6880 63776
rect 8116 63724 8168 63776
rect 9220 63724 9272 63776
rect 3610 63622 3662 63674
rect 3674 63622 3726 63674
rect 3738 63622 3790 63674
rect 3802 63622 3854 63674
rect 3866 63622 3918 63674
rect 5210 63622 5262 63674
rect 5274 63622 5326 63674
rect 5338 63622 5390 63674
rect 5402 63622 5454 63674
rect 5466 63622 5518 63674
rect 6810 63622 6862 63674
rect 6874 63622 6926 63674
rect 6938 63622 6990 63674
rect 7002 63622 7054 63674
rect 7066 63622 7118 63674
rect 8410 63622 8462 63674
rect 8474 63622 8526 63674
rect 8538 63622 8590 63674
rect 8602 63622 8654 63674
rect 8666 63622 8718 63674
rect 1584 63520 1636 63572
rect 10416 63520 10468 63572
rect 2136 63452 2188 63504
rect 2504 63452 2556 63504
rect 4804 63452 4856 63504
rect 5172 63452 5224 63504
rect 6000 63452 6052 63504
rect 6552 63452 6604 63504
rect 7656 63452 7708 63504
rect 1216 63384 1268 63436
rect 3608 63384 3660 63436
rect 5448 63384 5500 63436
rect 6092 63384 6144 63436
rect 6736 63384 6788 63436
rect 9680 63452 9732 63504
rect 6276 63316 6328 63368
rect 7196 63316 7248 63368
rect 7932 63316 7984 63368
rect 8392 63427 8444 63436
rect 8392 63393 8401 63427
rect 8401 63393 8435 63427
rect 8435 63393 8444 63427
rect 8392 63384 8444 63393
rect 8944 63384 8996 63436
rect 9036 63384 9088 63436
rect 5540 63180 5592 63232
rect 6828 63180 6880 63232
rect 8852 63316 8904 63368
rect 8760 63223 8812 63232
rect 8760 63189 8769 63223
rect 8769 63189 8803 63223
rect 8803 63189 8812 63223
rect 8760 63180 8812 63189
rect 8944 63180 8996 63232
rect 2950 63078 3002 63130
rect 3014 63078 3066 63130
rect 3078 63078 3130 63130
rect 3142 63078 3194 63130
rect 3206 63078 3258 63130
rect 4550 63078 4602 63130
rect 4614 63078 4666 63130
rect 4678 63078 4730 63130
rect 4742 63078 4794 63130
rect 4806 63078 4858 63130
rect 6150 63078 6202 63130
rect 6214 63078 6266 63130
rect 6278 63078 6330 63130
rect 6342 63078 6394 63130
rect 6406 63078 6458 63130
rect 7750 63078 7802 63130
rect 7814 63078 7866 63130
rect 7878 63078 7930 63130
rect 7942 63078 7994 63130
rect 8006 63078 8058 63130
rect 9350 63078 9402 63130
rect 9414 63078 9466 63130
rect 9478 63078 9530 63130
rect 9542 63078 9594 63130
rect 9606 63078 9658 63130
rect 6000 62976 6052 63028
rect 6736 62976 6788 63028
rect 8300 62976 8352 63028
rect 8760 62976 8812 63028
rect 1032 62908 1084 62960
rect 2320 62908 2372 62960
rect 940 62840 992 62892
rect 2320 62772 2372 62824
rect 4804 62840 4856 62892
rect 6092 62840 6144 62892
rect 6552 62883 6604 62892
rect 5172 62772 5224 62824
rect 5448 62772 5500 62824
rect 6552 62849 6561 62883
rect 6561 62849 6595 62883
rect 6595 62849 6604 62883
rect 6552 62840 6604 62849
rect 6828 62883 6880 62892
rect 6828 62849 6862 62883
rect 6862 62849 6880 62883
rect 6828 62840 6880 62849
rect 7104 62840 7156 62892
rect 7656 62840 7708 62892
rect 8668 62840 8720 62892
rect 7840 62772 7892 62824
rect 8484 62772 8536 62824
rect 8760 62772 8812 62824
rect 10048 62772 10100 62824
rect 7656 62636 7708 62688
rect 9956 62636 10008 62688
rect 10048 62636 10100 62688
rect 3610 62534 3662 62586
rect 3674 62534 3726 62586
rect 3738 62534 3790 62586
rect 3802 62534 3854 62586
rect 3866 62534 3918 62586
rect 5210 62534 5262 62586
rect 5274 62534 5326 62586
rect 5338 62534 5390 62586
rect 5402 62534 5454 62586
rect 5466 62534 5518 62586
rect 6810 62534 6862 62586
rect 6874 62534 6926 62586
rect 6938 62534 6990 62586
rect 7002 62534 7054 62586
rect 7066 62534 7118 62586
rect 8410 62534 8462 62586
rect 8474 62534 8526 62586
rect 8538 62534 8590 62586
rect 8602 62534 8654 62586
rect 8666 62534 8718 62586
rect 6460 62432 6512 62484
rect 4344 62364 4396 62416
rect 2504 62160 2556 62212
rect 4344 62160 4396 62212
rect 4712 62160 4764 62212
rect 5448 62160 5500 62212
rect 6092 62160 6144 62212
rect 8852 62432 8904 62484
rect 7196 62339 7248 62348
rect 7196 62305 7205 62339
rect 7205 62305 7239 62339
rect 7239 62305 7248 62339
rect 7196 62296 7248 62305
rect 7288 62296 7340 62348
rect 7564 62296 7616 62348
rect 7840 62271 7892 62280
rect 7840 62237 7849 62271
rect 7849 62237 7883 62271
rect 7883 62237 7892 62271
rect 7840 62228 7892 62237
rect 1584 62092 1636 62144
rect 6000 62092 6052 62144
rect 8760 62228 8812 62280
rect 11336 62092 11388 62144
rect 2950 61990 3002 62042
rect 3014 61990 3066 62042
rect 3078 61990 3130 62042
rect 3142 61990 3194 62042
rect 3206 61990 3258 62042
rect 4550 61990 4602 62042
rect 4614 61990 4666 62042
rect 4678 61990 4730 62042
rect 4742 61990 4794 62042
rect 4806 61990 4858 62042
rect 6150 61990 6202 62042
rect 6214 61990 6266 62042
rect 6278 61990 6330 62042
rect 6342 61990 6394 62042
rect 6406 61990 6458 62042
rect 7750 61990 7802 62042
rect 7814 61990 7866 62042
rect 7878 61990 7930 62042
rect 7942 61990 7994 62042
rect 8006 61990 8058 62042
rect 9350 61990 9402 62042
rect 9414 61990 9466 62042
rect 9478 61990 9530 62042
rect 9542 61990 9594 62042
rect 9606 61990 9658 62042
rect 5448 61888 5500 61940
rect 8300 61888 8352 61940
rect 940 61752 992 61804
rect 6552 61752 6604 61804
rect 7748 61752 7800 61804
rect 8208 61752 8260 61804
rect 8392 61820 8444 61872
rect 8760 61820 8812 61872
rect 8300 61684 8352 61736
rect 9312 61752 9364 61804
rect 8760 61684 8812 61736
rect 8944 61616 8996 61668
rect 8024 61591 8076 61600
rect 8024 61557 8033 61591
rect 8033 61557 8067 61591
rect 8067 61557 8076 61591
rect 8024 61548 8076 61557
rect 8116 61591 8168 61600
rect 8116 61557 8125 61591
rect 8125 61557 8159 61591
rect 8159 61557 8168 61591
rect 8116 61548 8168 61557
rect 3610 61446 3662 61498
rect 3674 61446 3726 61498
rect 3738 61446 3790 61498
rect 3802 61446 3854 61498
rect 3866 61446 3918 61498
rect 5210 61446 5262 61498
rect 5274 61446 5326 61498
rect 5338 61446 5390 61498
rect 5402 61446 5454 61498
rect 5466 61446 5518 61498
rect 6810 61446 6862 61498
rect 6874 61446 6926 61498
rect 6938 61446 6990 61498
rect 7002 61446 7054 61498
rect 7066 61446 7118 61498
rect 8410 61446 8462 61498
rect 8474 61446 8526 61498
rect 8538 61446 8590 61498
rect 8602 61446 8654 61498
rect 8666 61446 8718 61498
rect 7196 61344 7248 61396
rect 7472 61344 7524 61396
rect 7656 61251 7708 61260
rect 7656 61217 7665 61251
rect 7665 61217 7699 61251
rect 7699 61217 7708 61251
rect 7656 61208 7708 61217
rect 8024 61344 8076 61396
rect 8944 61344 8996 61396
rect 5264 61140 5316 61192
rect 5816 61140 5868 61192
rect 7288 61140 7340 61192
rect 8760 61208 8812 61260
rect 9128 61208 9180 61260
rect 9772 61208 9824 61260
rect 8944 61183 8996 61192
rect 8944 61149 8953 61183
rect 8953 61149 8987 61183
rect 8987 61149 8996 61183
rect 8944 61140 8996 61149
rect 5172 61072 5224 61124
rect 5816 61004 5868 61056
rect 8760 61072 8812 61124
rect 9312 61072 9364 61124
rect 9128 61047 9180 61056
rect 9128 61013 9137 61047
rect 9137 61013 9171 61047
rect 9171 61013 9180 61047
rect 9128 61004 9180 61013
rect 2950 60902 3002 60954
rect 3014 60902 3066 60954
rect 3078 60902 3130 60954
rect 3142 60902 3194 60954
rect 3206 60902 3258 60954
rect 4550 60902 4602 60954
rect 4614 60902 4666 60954
rect 4678 60902 4730 60954
rect 4742 60902 4794 60954
rect 4806 60902 4858 60954
rect 6150 60902 6202 60954
rect 6214 60902 6266 60954
rect 6278 60902 6330 60954
rect 6342 60902 6394 60954
rect 6406 60902 6458 60954
rect 7750 60902 7802 60954
rect 7814 60902 7866 60954
rect 7878 60902 7930 60954
rect 7942 60902 7994 60954
rect 8006 60902 8058 60954
rect 9350 60902 9402 60954
rect 9414 60902 9466 60954
rect 9478 60902 9530 60954
rect 9542 60902 9594 60954
rect 9606 60902 9658 60954
rect 480 60800 532 60852
rect 8944 60800 8996 60852
rect 9404 60800 9456 60852
rect 9864 60800 9916 60852
rect 4804 60732 4856 60784
rect 7656 60732 7708 60784
rect 940 60664 992 60716
rect 2688 60664 2740 60716
rect 4436 60707 4488 60716
rect 4436 60673 4445 60707
rect 4445 60673 4479 60707
rect 4479 60673 4488 60707
rect 4436 60664 4488 60673
rect 6552 60664 6604 60716
rect 7288 60664 7340 60716
rect 8300 60528 8352 60580
rect 2780 60460 2832 60512
rect 4436 60460 4488 60512
rect 4896 60460 4948 60512
rect 5264 60460 5316 60512
rect 5356 60460 5408 60512
rect 6552 60460 6604 60512
rect 3610 60358 3662 60410
rect 3674 60358 3726 60410
rect 3738 60358 3790 60410
rect 3802 60358 3854 60410
rect 3866 60358 3918 60410
rect 5210 60358 5262 60410
rect 5274 60358 5326 60410
rect 5338 60358 5390 60410
rect 5402 60358 5454 60410
rect 5466 60358 5518 60410
rect 6810 60358 6862 60410
rect 6874 60358 6926 60410
rect 6938 60358 6990 60410
rect 7002 60358 7054 60410
rect 7066 60358 7118 60410
rect 8410 60358 8462 60410
rect 8474 60358 8526 60410
rect 8538 60358 8590 60410
rect 8602 60358 8654 60410
rect 8666 60358 8718 60410
rect 4804 60256 4856 60308
rect 5080 60256 5132 60308
rect 7656 60256 7708 60308
rect 8208 60256 8260 60308
rect 8852 60188 8904 60240
rect 9220 60188 9272 60240
rect 2780 60120 2832 60172
rect 3884 60120 3936 60172
rect 7288 60163 7340 60172
rect 7288 60129 7297 60163
rect 7297 60129 7331 60163
rect 7331 60129 7340 60163
rect 7288 60120 7340 60129
rect 9404 60120 9456 60172
rect 1492 60027 1544 60036
rect 1492 59993 1501 60027
rect 1501 59993 1535 60027
rect 1535 59993 1544 60027
rect 1492 59984 1544 59993
rect 8208 59984 8260 60036
rect 940 59916 992 59968
rect 8300 59916 8352 59968
rect 2950 59814 3002 59866
rect 3014 59814 3066 59866
rect 3078 59814 3130 59866
rect 3142 59814 3194 59866
rect 3206 59814 3258 59866
rect 4550 59814 4602 59866
rect 4614 59814 4666 59866
rect 4678 59814 4730 59866
rect 4742 59814 4794 59866
rect 4806 59814 4858 59866
rect 6150 59814 6202 59866
rect 6214 59814 6266 59866
rect 6278 59814 6330 59866
rect 6342 59814 6394 59866
rect 6406 59814 6458 59866
rect 7750 59814 7802 59866
rect 7814 59814 7866 59866
rect 7878 59814 7930 59866
rect 7942 59814 7994 59866
rect 8006 59814 8058 59866
rect 9350 59814 9402 59866
rect 9414 59814 9466 59866
rect 9478 59814 9530 59866
rect 9542 59814 9594 59866
rect 9606 59814 9658 59866
rect 1492 59712 1544 59764
rect 7380 59712 7432 59764
rect 1216 59644 1268 59696
rect 3976 59619 4028 59628
rect 3976 59585 3985 59619
rect 3985 59585 4019 59619
rect 4019 59585 4028 59619
rect 3976 59576 4028 59585
rect 5724 59644 5776 59696
rect 11612 59644 11664 59696
rect 4896 59551 4948 59560
rect 4896 59517 4905 59551
rect 4905 59517 4939 59551
rect 4939 59517 4948 59551
rect 4896 59508 4948 59517
rect 7288 59508 7340 59560
rect 2780 59372 2832 59424
rect 4528 59372 4580 59424
rect 11152 59372 11204 59424
rect 11980 59372 12032 59424
rect 3610 59270 3662 59322
rect 3674 59270 3726 59322
rect 3738 59270 3790 59322
rect 3802 59270 3854 59322
rect 3866 59270 3918 59322
rect 5210 59270 5262 59322
rect 5274 59270 5326 59322
rect 5338 59270 5390 59322
rect 5402 59270 5454 59322
rect 5466 59270 5518 59322
rect 6810 59270 6862 59322
rect 6874 59270 6926 59322
rect 6938 59270 6990 59322
rect 7002 59270 7054 59322
rect 7066 59270 7118 59322
rect 8410 59270 8462 59322
rect 8474 59270 8526 59322
rect 8538 59270 8590 59322
rect 8602 59270 8654 59322
rect 8666 59270 8718 59322
rect 4252 59168 4304 59220
rect 6552 59100 6604 59152
rect 4344 59032 4396 59084
rect 296 58964 348 59016
rect 2872 58964 2924 59016
rect 4252 58964 4304 59016
rect 4528 58964 4580 59016
rect 4896 58964 4948 59016
rect 6828 59032 6880 59084
rect 6552 58964 6604 59016
rect 7380 59168 7432 59220
rect 7656 58964 7708 59016
rect 9588 58964 9640 59016
rect 5724 58939 5776 58948
rect 5724 58905 5736 58939
rect 5736 58905 5776 58939
rect 5724 58896 5776 58905
rect 5908 58896 5960 58948
rect 6828 58896 6880 58948
rect 940 58828 992 58880
rect 5080 58828 5132 58880
rect 7380 58828 7432 58880
rect 7748 58828 7800 58880
rect 8392 58828 8444 58880
rect 2950 58726 3002 58778
rect 3014 58726 3066 58778
rect 3078 58726 3130 58778
rect 3142 58726 3194 58778
rect 3206 58726 3258 58778
rect 4550 58726 4602 58778
rect 4614 58726 4666 58778
rect 4678 58726 4730 58778
rect 4742 58726 4794 58778
rect 4806 58726 4858 58778
rect 6150 58726 6202 58778
rect 6214 58726 6266 58778
rect 6278 58726 6330 58778
rect 6342 58726 6394 58778
rect 6406 58726 6458 58778
rect 7750 58726 7802 58778
rect 7814 58726 7866 58778
rect 7878 58726 7930 58778
rect 7942 58726 7994 58778
rect 8006 58726 8058 58778
rect 9350 58726 9402 58778
rect 9414 58726 9466 58778
rect 9478 58726 9530 58778
rect 9542 58726 9594 58778
rect 9606 58726 9658 58778
rect 5724 58624 5776 58676
rect 6092 58624 6144 58676
rect 6368 58624 6420 58676
rect 6920 58624 6972 58676
rect 8300 58624 8352 58676
rect 9036 58624 9088 58676
rect 9312 58624 9364 58676
rect 4896 58488 4948 58540
rect 10324 58556 10376 58608
rect 6828 58488 6880 58540
rect 7196 58531 7248 58540
rect 7196 58497 7205 58531
rect 7205 58497 7239 58531
rect 7239 58497 7248 58531
rect 7196 58488 7248 58497
rect 8208 58488 8260 58540
rect 10876 58488 10928 58540
rect 4896 58352 4948 58404
rect 5172 58352 5224 58404
rect 5724 58352 5776 58404
rect 7472 58420 7524 58472
rect 7656 58420 7708 58472
rect 8760 58420 8812 58472
rect 7196 58352 7248 58404
rect 5908 58284 5960 58336
rect 6460 58284 6512 58336
rect 7472 58284 7524 58336
rect 8208 58352 8260 58404
rect 8760 58327 8812 58336
rect 8760 58293 8769 58327
rect 8769 58293 8803 58327
rect 8803 58293 8812 58327
rect 8760 58284 8812 58293
rect 3610 58182 3662 58234
rect 3674 58182 3726 58234
rect 3738 58182 3790 58234
rect 3802 58182 3854 58234
rect 3866 58182 3918 58234
rect 5210 58182 5262 58234
rect 5274 58182 5326 58234
rect 5338 58182 5390 58234
rect 5402 58182 5454 58234
rect 5466 58182 5518 58234
rect 6810 58182 6862 58234
rect 6874 58182 6926 58234
rect 6938 58182 6990 58234
rect 7002 58182 7054 58234
rect 7066 58182 7118 58234
rect 8410 58182 8462 58234
rect 8474 58182 8526 58234
rect 8538 58182 8590 58234
rect 8602 58182 8654 58234
rect 8666 58182 8718 58234
rect 4896 58080 4948 58132
rect 5172 58080 5224 58132
rect 7196 58080 7248 58132
rect 7288 58080 7340 58132
rect 8300 57944 8352 57996
rect 2688 57876 2740 57928
rect 6368 57876 6420 57928
rect 7564 57876 7616 57928
rect 7748 57876 7800 57928
rect 8208 57808 8260 57860
rect 1584 57783 1636 57792
rect 1584 57749 1593 57783
rect 1593 57749 1627 57783
rect 1627 57749 1636 57783
rect 1584 57740 1636 57749
rect 5448 57740 5500 57792
rect 6092 57740 6144 57792
rect 7196 57740 7248 57792
rect 7288 57740 7340 57792
rect 8576 57740 8628 57792
rect 11244 57876 11296 57928
rect 8852 57740 8904 57792
rect 9128 57783 9180 57792
rect 9128 57749 9137 57783
rect 9137 57749 9171 57783
rect 9171 57749 9180 57783
rect 9128 57740 9180 57749
rect 2950 57638 3002 57690
rect 3014 57638 3066 57690
rect 3078 57638 3130 57690
rect 3142 57638 3194 57690
rect 3206 57638 3258 57690
rect 4550 57638 4602 57690
rect 4614 57638 4666 57690
rect 4678 57638 4730 57690
rect 4742 57638 4794 57690
rect 4806 57638 4858 57690
rect 6150 57638 6202 57690
rect 6214 57638 6266 57690
rect 6278 57638 6330 57690
rect 6342 57638 6394 57690
rect 6406 57638 6458 57690
rect 7750 57638 7802 57690
rect 7814 57638 7866 57690
rect 7878 57638 7930 57690
rect 7942 57638 7994 57690
rect 8006 57638 8058 57690
rect 9350 57638 9402 57690
rect 9414 57638 9466 57690
rect 9478 57638 9530 57690
rect 9542 57638 9594 57690
rect 9606 57638 9658 57690
rect 2596 57536 2648 57588
rect 4160 57536 4212 57588
rect 5172 57536 5224 57588
rect 6276 57536 6328 57588
rect 6368 57536 6420 57588
rect 6552 57536 6604 57588
rect 4436 57468 4488 57520
rect 4896 57468 4948 57520
rect 7104 57468 7156 57520
rect 6368 57443 6420 57452
rect 6368 57409 6377 57443
rect 6377 57409 6411 57443
rect 6411 57409 6420 57443
rect 6368 57400 6420 57409
rect 7196 57400 7248 57452
rect 8944 57400 8996 57452
rect 7564 57332 7616 57384
rect 4344 57264 4396 57316
rect 4436 57264 4488 57316
rect 5356 57264 5408 57316
rect 5632 57264 5684 57316
rect 6368 57264 6420 57316
rect 7380 57264 7432 57316
rect 8576 57264 8628 57316
rect 8944 57264 8996 57316
rect 4252 57196 4304 57248
rect 3610 57094 3662 57146
rect 3674 57094 3726 57146
rect 3738 57094 3790 57146
rect 3802 57094 3854 57146
rect 3866 57094 3918 57146
rect 5210 57094 5262 57146
rect 5274 57094 5326 57146
rect 5338 57094 5390 57146
rect 5402 57094 5454 57146
rect 5466 57094 5518 57146
rect 6810 57094 6862 57146
rect 6874 57094 6926 57146
rect 6938 57094 6990 57146
rect 7002 57094 7054 57146
rect 7066 57094 7118 57146
rect 8410 57094 8462 57146
rect 8474 57094 8526 57146
rect 8538 57094 8590 57146
rect 8602 57094 8654 57146
rect 8666 57094 8718 57146
rect 6276 56856 6328 56908
rect 6828 56856 6880 56908
rect 3516 56788 3568 56840
rect 6736 56788 6788 56840
rect 9220 56788 9272 56840
rect 6644 56720 6696 56772
rect 11060 56720 11112 56772
rect 940 56652 992 56704
rect 3516 56652 3568 56704
rect 6368 56652 6420 56704
rect 6736 56652 6788 56704
rect 7196 56652 7248 56704
rect 2950 56550 3002 56602
rect 3014 56550 3066 56602
rect 3078 56550 3130 56602
rect 3142 56550 3194 56602
rect 3206 56550 3258 56602
rect 4550 56550 4602 56602
rect 4614 56550 4666 56602
rect 4678 56550 4730 56602
rect 4742 56550 4794 56602
rect 4806 56550 4858 56602
rect 6150 56550 6202 56602
rect 6214 56550 6266 56602
rect 6278 56550 6330 56602
rect 6342 56550 6394 56602
rect 6406 56550 6458 56602
rect 7750 56550 7802 56602
rect 7814 56550 7866 56602
rect 7878 56550 7930 56602
rect 7942 56550 7994 56602
rect 8006 56550 8058 56602
rect 9350 56550 9402 56602
rect 9414 56550 9466 56602
rect 9478 56550 9530 56602
rect 9542 56550 9594 56602
rect 9606 56550 9658 56602
rect 7656 56448 7708 56500
rect 3332 56380 3384 56432
rect 4436 56312 4488 56364
rect 4988 56312 5040 56364
rect 5080 56312 5132 56364
rect 8852 56312 8904 56364
rect 3332 56244 3384 56296
rect 3516 56244 3568 56296
rect 1492 56176 1544 56228
rect 6644 56244 6696 56296
rect 8208 56244 8260 56296
rect 940 56108 992 56160
rect 2688 56108 2740 56160
rect 5080 56108 5132 56160
rect 6828 56108 6880 56160
rect 7656 56108 7708 56160
rect 3610 56006 3662 56058
rect 3674 56006 3726 56058
rect 3738 56006 3790 56058
rect 3802 56006 3854 56058
rect 3866 56006 3918 56058
rect 5210 56006 5262 56058
rect 5274 56006 5326 56058
rect 5338 56006 5390 56058
rect 5402 56006 5454 56058
rect 5466 56006 5518 56058
rect 6810 56006 6862 56058
rect 6874 56006 6926 56058
rect 6938 56006 6990 56058
rect 7002 56006 7054 56058
rect 7066 56006 7118 56058
rect 8410 56006 8462 56058
rect 8474 56006 8526 56058
rect 8538 56006 8590 56058
rect 8602 56006 8654 56058
rect 8666 56006 8718 56058
rect 1216 55904 1268 55956
rect 2136 55836 2188 55888
rect 9680 55836 9732 55888
rect 8208 55768 8260 55820
rect 4436 55632 4488 55684
rect 7564 55743 7616 55752
rect 7564 55709 7573 55743
rect 7573 55709 7607 55743
rect 7607 55709 7616 55743
rect 7564 55700 7616 55709
rect 8116 55700 8168 55752
rect 5540 55564 5592 55616
rect 8208 55564 8260 55616
rect 2950 55462 3002 55514
rect 3014 55462 3066 55514
rect 3078 55462 3130 55514
rect 3142 55462 3194 55514
rect 3206 55462 3258 55514
rect 4550 55462 4602 55514
rect 4614 55462 4666 55514
rect 4678 55462 4730 55514
rect 4742 55462 4794 55514
rect 4806 55462 4858 55514
rect 6150 55462 6202 55514
rect 6214 55462 6266 55514
rect 6278 55462 6330 55514
rect 6342 55462 6394 55514
rect 6406 55462 6458 55514
rect 7750 55462 7802 55514
rect 7814 55462 7866 55514
rect 7878 55462 7930 55514
rect 7942 55462 7994 55514
rect 8006 55462 8058 55514
rect 9350 55462 9402 55514
rect 9414 55462 9466 55514
rect 9478 55462 9530 55514
rect 9542 55462 9594 55514
rect 9606 55462 9658 55514
rect 7564 55360 7616 55412
rect 8116 55360 8168 55412
rect 2412 55292 2464 55344
rect 9680 55224 9732 55276
rect 9864 55224 9916 55276
rect 940 55020 992 55072
rect 3610 54918 3662 54970
rect 3674 54918 3726 54970
rect 3738 54918 3790 54970
rect 3802 54918 3854 54970
rect 3866 54918 3918 54970
rect 5210 54918 5262 54970
rect 5274 54918 5326 54970
rect 5338 54918 5390 54970
rect 5402 54918 5454 54970
rect 5466 54918 5518 54970
rect 6810 54918 6862 54970
rect 6874 54918 6926 54970
rect 6938 54918 6990 54970
rect 7002 54918 7054 54970
rect 7066 54918 7118 54970
rect 8410 54918 8462 54970
rect 8474 54918 8526 54970
rect 8538 54918 8590 54970
rect 8602 54918 8654 54970
rect 8666 54918 8718 54970
rect 6644 54612 6696 54664
rect 8944 54612 8996 54664
rect 9220 54544 9272 54596
rect 2872 54476 2924 54528
rect 2950 54374 3002 54426
rect 3014 54374 3066 54426
rect 3078 54374 3130 54426
rect 3142 54374 3194 54426
rect 3206 54374 3258 54426
rect 4550 54374 4602 54426
rect 4614 54374 4666 54426
rect 4678 54374 4730 54426
rect 4742 54374 4794 54426
rect 4806 54374 4858 54426
rect 6150 54374 6202 54426
rect 6214 54374 6266 54426
rect 6278 54374 6330 54426
rect 6342 54374 6394 54426
rect 6406 54374 6458 54426
rect 7750 54374 7802 54426
rect 7814 54374 7866 54426
rect 7878 54374 7930 54426
rect 7942 54374 7994 54426
rect 8006 54374 8058 54426
rect 9350 54374 9402 54426
rect 9414 54374 9466 54426
rect 9478 54374 9530 54426
rect 9542 54374 9594 54426
rect 9606 54374 9658 54426
rect 1400 54204 1452 54256
rect 5816 54204 5868 54256
rect 6000 54136 6052 54188
rect 6644 54136 6696 54188
rect 2596 54000 2648 54052
rect 9680 54272 9732 54324
rect 7472 54204 7524 54256
rect 10784 54204 10836 54256
rect 7840 54179 7892 54188
rect 7840 54145 7847 54179
rect 7847 54145 7881 54179
rect 7881 54145 7892 54179
rect 7840 54136 7892 54145
rect 8944 54136 8996 54188
rect 11520 54000 11572 54052
rect 940 53932 992 53984
rect 2688 53932 2740 53984
rect 7564 53975 7616 53984
rect 7564 53941 7573 53975
rect 7573 53941 7607 53975
rect 7607 53941 7616 53975
rect 7564 53932 7616 53941
rect 7656 53932 7708 53984
rect 3610 53830 3662 53882
rect 3674 53830 3726 53882
rect 3738 53830 3790 53882
rect 3802 53830 3854 53882
rect 3866 53830 3918 53882
rect 5210 53830 5262 53882
rect 5274 53830 5326 53882
rect 5338 53830 5390 53882
rect 5402 53830 5454 53882
rect 5466 53830 5518 53882
rect 6810 53830 6862 53882
rect 6874 53830 6926 53882
rect 6938 53830 6990 53882
rect 7002 53830 7054 53882
rect 7066 53830 7118 53882
rect 8410 53830 8462 53882
rect 8474 53830 8526 53882
rect 8538 53830 8590 53882
rect 8602 53830 8654 53882
rect 8666 53830 8718 53882
rect 4896 53728 4948 53780
rect 7012 53728 7064 53780
rect 10232 53728 10284 53780
rect 11428 53728 11480 53780
rect 4804 53660 4856 53712
rect 2136 53524 2188 53576
rect 4160 53524 4212 53576
rect 4436 53524 4488 53576
rect 3976 53456 4028 53508
rect 7104 53524 7156 53576
rect 7288 53524 7340 53576
rect 7380 53524 7432 53576
rect 7748 53567 7800 53576
rect 7748 53533 7757 53567
rect 7757 53533 7791 53567
rect 7791 53533 7800 53567
rect 7748 53524 7800 53533
rect 3516 53388 3568 53440
rect 7104 53388 7156 53440
rect 7380 53431 7432 53440
rect 7380 53397 7389 53431
rect 7389 53397 7423 53431
rect 7423 53397 7432 53431
rect 7380 53388 7432 53397
rect 7472 53388 7524 53440
rect 2950 53286 3002 53338
rect 3014 53286 3066 53338
rect 3078 53286 3130 53338
rect 3142 53286 3194 53338
rect 3206 53286 3258 53338
rect 4550 53286 4602 53338
rect 4614 53286 4666 53338
rect 4678 53286 4730 53338
rect 4742 53286 4794 53338
rect 4806 53286 4858 53338
rect 6150 53286 6202 53338
rect 6214 53286 6266 53338
rect 6278 53286 6330 53338
rect 6342 53286 6394 53338
rect 6406 53286 6458 53338
rect 7750 53286 7802 53338
rect 7814 53286 7866 53338
rect 7878 53286 7930 53338
rect 7942 53286 7994 53338
rect 8006 53286 8058 53338
rect 9350 53286 9402 53338
rect 9414 53286 9466 53338
rect 9478 53286 9530 53338
rect 9542 53286 9594 53338
rect 9606 53286 9658 53338
rect 5724 53184 5776 53236
rect 7012 53184 7064 53236
rect 7196 53184 7248 53236
rect 2780 53116 2832 53168
rect 5080 53116 5132 53168
rect 756 53048 808 53100
rect 4160 53048 4212 53100
rect 4804 53091 4856 53100
rect 1124 52980 1176 53032
rect 4804 53057 4813 53091
rect 4813 53057 4847 53091
rect 4847 53057 4856 53091
rect 4804 53048 4856 53057
rect 5632 52980 5684 53032
rect 2780 52912 2832 52964
rect 3792 52912 3844 52964
rect 6460 53048 6512 53100
rect 6644 53048 6696 53100
rect 7104 53116 7156 53168
rect 7380 53184 7432 53236
rect 7564 53184 7616 53236
rect 7656 53091 7708 53100
rect 7656 53057 7665 53091
rect 7665 53057 7699 53091
rect 7699 53057 7708 53091
rect 7656 53048 7708 53057
rect 9772 53116 9824 53168
rect 10048 53116 10100 53168
rect 8300 52980 8352 53032
rect 940 52844 992 52896
rect 2412 52844 2464 52896
rect 7288 52912 7340 52964
rect 7564 52912 7616 52964
rect 4804 52844 4856 52896
rect 5080 52844 5132 52896
rect 6184 52844 6236 52896
rect 7472 52887 7524 52896
rect 7472 52853 7481 52887
rect 7481 52853 7515 52887
rect 7515 52853 7524 52887
rect 7472 52844 7524 52853
rect 7748 52887 7800 52896
rect 7748 52853 7757 52887
rect 7757 52853 7791 52887
rect 7791 52853 7800 52887
rect 7748 52844 7800 52853
rect 3610 52742 3662 52794
rect 3674 52742 3726 52794
rect 3738 52742 3790 52794
rect 3802 52742 3854 52794
rect 3866 52742 3918 52794
rect 5210 52742 5262 52794
rect 5274 52742 5326 52794
rect 5338 52742 5390 52794
rect 5402 52742 5454 52794
rect 5466 52742 5518 52794
rect 6810 52742 6862 52794
rect 6874 52742 6926 52794
rect 6938 52742 6990 52794
rect 7002 52742 7054 52794
rect 7066 52742 7118 52794
rect 8410 52742 8462 52794
rect 8474 52742 8526 52794
rect 8538 52742 8590 52794
rect 8602 52742 8654 52794
rect 8666 52742 8718 52794
rect 5724 52640 5776 52692
rect 5908 52640 5960 52692
rect 6644 52640 6696 52692
rect 6184 52479 6236 52488
rect 6184 52445 6193 52479
rect 6193 52445 6227 52479
rect 6227 52445 6236 52479
rect 6184 52436 6236 52445
rect 6736 52479 6788 52488
rect 6736 52445 6745 52479
rect 6745 52445 6779 52479
rect 6779 52445 6788 52479
rect 6736 52436 6788 52445
rect 4252 52368 4304 52420
rect 1584 52343 1636 52352
rect 1584 52309 1593 52343
rect 1593 52309 1627 52343
rect 1627 52309 1636 52343
rect 1584 52300 1636 52309
rect 5908 52300 5960 52352
rect 6460 52300 6512 52352
rect 7288 52300 7340 52352
rect 7748 52300 7800 52352
rect 2950 52198 3002 52250
rect 3014 52198 3066 52250
rect 3078 52198 3130 52250
rect 3142 52198 3194 52250
rect 3206 52198 3258 52250
rect 4550 52198 4602 52250
rect 4614 52198 4666 52250
rect 4678 52198 4730 52250
rect 4742 52198 4794 52250
rect 4806 52198 4858 52250
rect 6150 52198 6202 52250
rect 6214 52198 6266 52250
rect 6278 52198 6330 52250
rect 6342 52198 6394 52250
rect 6406 52198 6458 52250
rect 7750 52198 7802 52250
rect 7814 52198 7866 52250
rect 7878 52198 7930 52250
rect 7942 52198 7994 52250
rect 8006 52198 8058 52250
rect 9350 52198 9402 52250
rect 9414 52198 9466 52250
rect 9478 52198 9530 52250
rect 9542 52198 9594 52250
rect 9606 52198 9658 52250
rect 4804 52096 4856 52148
rect 5908 52096 5960 52148
rect 7564 52028 7616 52080
rect 6460 51960 6512 52012
rect 6552 51892 6604 51944
rect 6828 51960 6880 52012
rect 7472 51960 7524 52012
rect 7748 51960 7800 52012
rect 10140 51960 10192 52012
rect 6736 51935 6788 51944
rect 6736 51901 6745 51935
rect 6745 51901 6779 51935
rect 6779 51901 6788 51935
rect 6736 51892 6788 51901
rect 1584 51756 1636 51808
rect 6368 51756 6420 51808
rect 8116 51799 8168 51808
rect 8116 51765 8125 51799
rect 8125 51765 8159 51799
rect 8159 51765 8168 51799
rect 8116 51756 8168 51765
rect 3610 51654 3662 51706
rect 3674 51654 3726 51706
rect 3738 51654 3790 51706
rect 3802 51654 3854 51706
rect 3866 51654 3918 51706
rect 5210 51654 5262 51706
rect 5274 51654 5326 51706
rect 5338 51654 5390 51706
rect 5402 51654 5454 51706
rect 5466 51654 5518 51706
rect 6810 51654 6862 51706
rect 6874 51654 6926 51706
rect 6938 51654 6990 51706
rect 7002 51654 7054 51706
rect 7066 51654 7118 51706
rect 8410 51654 8462 51706
rect 8474 51654 8526 51706
rect 8538 51654 8590 51706
rect 8602 51654 8654 51706
rect 8666 51654 8718 51706
rect 7012 51552 7064 51604
rect 8668 51552 8720 51604
rect 9588 51552 9640 51604
rect 4896 51416 4948 51468
rect 1492 51391 1544 51400
rect 1492 51357 1501 51391
rect 1501 51357 1535 51391
rect 1535 51357 1544 51391
rect 1492 51348 1544 51357
rect 5080 51348 5132 51400
rect 5908 51348 5960 51400
rect 6368 51348 6420 51400
rect 6736 51391 6788 51400
rect 6736 51357 6745 51391
rect 6745 51357 6779 51391
rect 6779 51357 6788 51391
rect 6736 51348 6788 51357
rect 8208 51348 8260 51400
rect 8300 51348 8352 51400
rect 8852 51348 8904 51400
rect 940 51212 992 51264
rect 4252 51212 4304 51264
rect 7288 51280 7340 51332
rect 7472 51280 7524 51332
rect 7748 51280 7800 51332
rect 8576 51280 8628 51332
rect 8208 51255 8260 51264
rect 8208 51221 8217 51255
rect 8217 51221 8251 51255
rect 8251 51221 8260 51255
rect 8208 51212 8260 51221
rect 8300 51212 8352 51264
rect 9220 51212 9272 51264
rect 2950 51110 3002 51162
rect 3014 51110 3066 51162
rect 3078 51110 3130 51162
rect 3142 51110 3194 51162
rect 3206 51110 3258 51162
rect 4550 51110 4602 51162
rect 4614 51110 4666 51162
rect 4678 51110 4730 51162
rect 4742 51110 4794 51162
rect 4806 51110 4858 51162
rect 6150 51110 6202 51162
rect 6214 51110 6266 51162
rect 6278 51110 6330 51162
rect 6342 51110 6394 51162
rect 6406 51110 6458 51162
rect 7750 51110 7802 51162
rect 7814 51110 7866 51162
rect 7878 51110 7930 51162
rect 7942 51110 7994 51162
rect 8006 51110 8058 51162
rect 9350 51110 9402 51162
rect 9414 51110 9466 51162
rect 9478 51110 9530 51162
rect 9542 51110 9594 51162
rect 9606 51110 9658 51162
rect 2228 51008 2280 51060
rect 2504 51008 2556 51060
rect 2596 51008 2648 51060
rect 2412 50940 2464 50992
rect 2412 50736 2464 50788
rect 6000 50940 6052 50992
rect 7012 51008 7064 51060
rect 7472 50940 7524 50992
rect 5632 50872 5684 50924
rect 6736 50872 6788 50924
rect 8668 50804 8720 50856
rect 9588 50804 9640 50856
rect 2504 50668 2556 50720
rect 7012 50668 7064 50720
rect 7288 50668 7340 50720
rect 3610 50566 3662 50618
rect 3674 50566 3726 50618
rect 3738 50566 3790 50618
rect 3802 50566 3854 50618
rect 3866 50566 3918 50618
rect 5210 50566 5262 50618
rect 5274 50566 5326 50618
rect 5338 50566 5390 50618
rect 5402 50566 5454 50618
rect 5466 50566 5518 50618
rect 6810 50566 6862 50618
rect 6874 50566 6926 50618
rect 6938 50566 6990 50618
rect 7002 50566 7054 50618
rect 7066 50566 7118 50618
rect 8410 50566 8462 50618
rect 8474 50566 8526 50618
rect 8538 50566 8590 50618
rect 8602 50566 8654 50618
rect 8666 50566 8718 50618
rect 3332 50260 3384 50312
rect 3792 50192 3844 50244
rect 4344 50192 4396 50244
rect 940 50124 992 50176
rect 5632 50124 5684 50176
rect 6092 50124 6144 50176
rect 2950 50022 3002 50074
rect 3014 50022 3066 50074
rect 3078 50022 3130 50074
rect 3142 50022 3194 50074
rect 3206 50022 3258 50074
rect 4550 50022 4602 50074
rect 4614 50022 4666 50074
rect 4678 50022 4730 50074
rect 4742 50022 4794 50074
rect 4806 50022 4858 50074
rect 6150 50022 6202 50074
rect 6214 50022 6266 50074
rect 6278 50022 6330 50074
rect 6342 50022 6394 50074
rect 6406 50022 6458 50074
rect 7750 50022 7802 50074
rect 7814 50022 7866 50074
rect 7878 50022 7930 50074
rect 7942 50022 7994 50074
rect 8006 50022 8058 50074
rect 9350 50022 9402 50074
rect 9414 50022 9466 50074
rect 9478 50022 9530 50074
rect 9542 50022 9594 50074
rect 9606 50022 9658 50074
rect 2320 49852 2372 49904
rect 3792 49852 3844 49904
rect 1032 49784 1084 49836
rect 4436 49920 4488 49972
rect 5080 49920 5132 49972
rect 4712 49852 4764 49904
rect 5540 49852 5592 49904
rect 3332 49716 3384 49768
rect 4344 49716 4396 49768
rect 4344 49580 4396 49632
rect 7656 49920 7708 49972
rect 6736 49784 6788 49836
rect 8300 49827 8352 49836
rect 8300 49793 8309 49827
rect 8309 49793 8343 49827
rect 8343 49793 8352 49827
rect 8300 49784 8352 49793
rect 4896 49580 4948 49632
rect 8300 49580 8352 49632
rect 3610 49478 3662 49530
rect 3674 49478 3726 49530
rect 3738 49478 3790 49530
rect 3802 49478 3854 49530
rect 3866 49478 3918 49530
rect 5210 49478 5262 49530
rect 5274 49478 5326 49530
rect 5338 49478 5390 49530
rect 5402 49478 5454 49530
rect 5466 49478 5518 49530
rect 6810 49478 6862 49530
rect 6874 49478 6926 49530
rect 6938 49478 6990 49530
rect 7002 49478 7054 49530
rect 7066 49478 7118 49530
rect 8410 49478 8462 49530
rect 8474 49478 8526 49530
rect 8538 49478 8590 49530
rect 8602 49478 8654 49530
rect 8666 49478 8718 49530
rect 2228 49376 2280 49428
rect 4712 49376 4764 49428
rect 5172 49376 5224 49428
rect 6644 49376 6696 49428
rect 8116 49376 8168 49428
rect 9220 49376 9272 49428
rect 6736 49215 6788 49224
rect 6736 49181 6745 49215
rect 6745 49181 6779 49215
rect 6779 49181 6788 49215
rect 6736 49172 6788 49181
rect 7472 49172 7524 49224
rect 8576 49240 8628 49292
rect 9128 49240 9180 49292
rect 11336 49172 11388 49224
rect 7656 49104 7708 49156
rect 940 49036 992 49088
rect 6644 49079 6696 49088
rect 6644 49045 6653 49079
rect 6653 49045 6687 49079
rect 6687 49045 6696 49079
rect 6644 49036 6696 49045
rect 8116 49079 8168 49088
rect 8116 49045 8125 49079
rect 8125 49045 8159 49079
rect 8159 49045 8168 49079
rect 8116 49036 8168 49045
rect 8760 49036 8812 49088
rect 2950 48934 3002 48986
rect 3014 48934 3066 48986
rect 3078 48934 3130 48986
rect 3142 48934 3194 48986
rect 3206 48934 3258 48986
rect 4550 48934 4602 48986
rect 4614 48934 4666 48986
rect 4678 48934 4730 48986
rect 4742 48934 4794 48986
rect 4806 48934 4858 48986
rect 6150 48934 6202 48986
rect 6214 48934 6266 48986
rect 6278 48934 6330 48986
rect 6342 48934 6394 48986
rect 6406 48934 6458 48986
rect 7750 48934 7802 48986
rect 7814 48934 7866 48986
rect 7878 48934 7930 48986
rect 7942 48934 7994 48986
rect 8006 48934 8058 48986
rect 9350 48934 9402 48986
rect 9414 48934 9466 48986
rect 9478 48934 9530 48986
rect 9542 48934 9594 48986
rect 9606 48934 9658 48986
rect 4160 48832 4212 48884
rect 4804 48832 4856 48884
rect 4896 48832 4948 48884
rect 2872 48764 2924 48816
rect 6092 48696 6144 48748
rect 6736 48696 6788 48748
rect 8208 48764 8260 48816
rect 8668 48696 8720 48748
rect 9128 48696 9180 48748
rect 4712 48560 4764 48612
rect 5172 48560 5224 48612
rect 1584 48535 1636 48544
rect 1584 48501 1593 48535
rect 1593 48501 1627 48535
rect 1627 48501 1636 48535
rect 1584 48492 1636 48501
rect 4252 48492 4304 48544
rect 8208 48492 8260 48544
rect 8576 48492 8628 48544
rect 8944 48492 8996 48544
rect 3610 48390 3662 48442
rect 3674 48390 3726 48442
rect 3738 48390 3790 48442
rect 3802 48390 3854 48442
rect 3866 48390 3918 48442
rect 5210 48390 5262 48442
rect 5274 48390 5326 48442
rect 5338 48390 5390 48442
rect 5402 48390 5454 48442
rect 5466 48390 5518 48442
rect 6810 48390 6862 48442
rect 6874 48390 6926 48442
rect 6938 48390 6990 48442
rect 7002 48390 7054 48442
rect 7066 48390 7118 48442
rect 8410 48390 8462 48442
rect 8474 48390 8526 48442
rect 8538 48390 8590 48442
rect 8602 48390 8654 48442
rect 8666 48390 8718 48442
rect 4712 48288 4764 48340
rect 5172 48288 5224 48340
rect 6736 48084 6788 48136
rect 7196 48084 7248 48136
rect 7472 48084 7524 48136
rect 6092 47948 6144 48000
rect 6828 47948 6880 48000
rect 7196 47948 7248 48000
rect 7472 47948 7524 48000
rect 2950 47846 3002 47898
rect 3014 47846 3066 47898
rect 3078 47846 3130 47898
rect 3142 47846 3194 47898
rect 3206 47846 3258 47898
rect 4550 47846 4602 47898
rect 4614 47846 4666 47898
rect 4678 47846 4730 47898
rect 4742 47846 4794 47898
rect 4806 47846 4858 47898
rect 6150 47846 6202 47898
rect 6214 47846 6266 47898
rect 6278 47846 6330 47898
rect 6342 47846 6394 47898
rect 6406 47846 6458 47898
rect 7750 47846 7802 47898
rect 7814 47846 7866 47898
rect 7878 47846 7930 47898
rect 7942 47846 7994 47898
rect 8006 47846 8058 47898
rect 9350 47846 9402 47898
rect 9414 47846 9466 47898
rect 9478 47846 9530 47898
rect 9542 47846 9594 47898
rect 9606 47846 9658 47898
rect 2688 47676 2740 47728
rect 6460 47608 6512 47660
rect 6828 47608 6880 47660
rect 4896 47472 4948 47524
rect 9036 47472 9088 47524
rect 9312 47472 9364 47524
rect 940 47404 992 47456
rect 2872 47404 2924 47456
rect 5172 47404 5224 47456
rect 7288 47404 7340 47456
rect 3610 47302 3662 47354
rect 3674 47302 3726 47354
rect 3738 47302 3790 47354
rect 3802 47302 3854 47354
rect 3866 47302 3918 47354
rect 5210 47302 5262 47354
rect 5274 47302 5326 47354
rect 5338 47302 5390 47354
rect 5402 47302 5454 47354
rect 5466 47302 5518 47354
rect 6810 47302 6862 47354
rect 6874 47302 6926 47354
rect 6938 47302 6990 47354
rect 7002 47302 7054 47354
rect 7066 47302 7118 47354
rect 8410 47302 8462 47354
rect 8474 47302 8526 47354
rect 8538 47302 8590 47354
rect 8602 47302 8654 47354
rect 8666 47302 8718 47354
rect 1584 47064 1636 47116
rect 3332 47064 3384 47116
rect 8852 47064 8904 47116
rect 9036 47064 9088 47116
rect 9220 47064 9272 47116
rect 6828 46996 6880 47048
rect 2780 46928 2832 46980
rect 3332 46928 3384 46980
rect 4252 46928 4304 46980
rect 5540 46928 5592 46980
rect 6460 46928 6512 46980
rect 7104 46928 7156 46980
rect 5172 46903 5224 46912
rect 5172 46869 5181 46903
rect 5181 46869 5215 46903
rect 5215 46869 5224 46903
rect 5172 46860 5224 46869
rect 5724 46860 5776 46912
rect 6736 46860 6788 46912
rect 8852 46860 8904 46912
rect 2950 46758 3002 46810
rect 3014 46758 3066 46810
rect 3078 46758 3130 46810
rect 3142 46758 3194 46810
rect 3206 46758 3258 46810
rect 4550 46758 4602 46810
rect 4614 46758 4666 46810
rect 4678 46758 4730 46810
rect 4742 46758 4794 46810
rect 4806 46758 4858 46810
rect 6150 46758 6202 46810
rect 6214 46758 6266 46810
rect 6278 46758 6330 46810
rect 6342 46758 6394 46810
rect 6406 46758 6458 46810
rect 7750 46758 7802 46810
rect 7814 46758 7866 46810
rect 7878 46758 7930 46810
rect 7942 46758 7994 46810
rect 8006 46758 8058 46810
rect 9350 46758 9402 46810
rect 9414 46758 9466 46810
rect 9478 46758 9530 46810
rect 9542 46758 9594 46810
rect 9606 46758 9658 46810
rect 5724 46656 5776 46708
rect 5908 46656 5960 46708
rect 6828 46656 6880 46708
rect 2412 46588 2464 46640
rect 6460 46588 6512 46640
rect 6736 46588 6788 46640
rect 7196 46588 7248 46640
rect 11152 46588 11204 46640
rect 5540 46520 5592 46572
rect 6000 46452 6052 46504
rect 6368 46495 6420 46504
rect 6368 46461 6377 46495
rect 6377 46461 6411 46495
rect 6411 46461 6420 46495
rect 6368 46452 6420 46461
rect 9956 46520 10008 46572
rect 940 46316 992 46368
rect 4344 46316 4396 46368
rect 5172 46316 5224 46368
rect 6092 46384 6144 46436
rect 5908 46316 5960 46368
rect 6276 46316 6328 46368
rect 3610 46214 3662 46266
rect 3674 46214 3726 46266
rect 3738 46214 3790 46266
rect 3802 46214 3854 46266
rect 3866 46214 3918 46266
rect 5210 46214 5262 46266
rect 5274 46214 5326 46266
rect 5338 46214 5390 46266
rect 5402 46214 5454 46266
rect 5466 46214 5518 46266
rect 6810 46214 6862 46266
rect 6874 46214 6926 46266
rect 6938 46214 6990 46266
rect 7002 46214 7054 46266
rect 7066 46214 7118 46266
rect 8410 46214 8462 46266
rect 8474 46214 8526 46266
rect 8538 46214 8590 46266
rect 8602 46214 8654 46266
rect 8666 46214 8718 46266
rect 2504 46112 2556 46164
rect 2872 46112 2924 46164
rect 7012 46112 7064 46164
rect 7288 46112 7340 46164
rect 6368 45976 6420 46028
rect 6644 46019 6696 46028
rect 6644 45985 6653 46019
rect 6653 45985 6687 46019
rect 6687 45985 6696 46019
rect 6644 45976 6696 45985
rect 4528 45908 4580 45960
rect 5172 45908 5224 45960
rect 6460 45908 6512 45960
rect 8208 46112 8260 46164
rect 8300 46155 8352 46164
rect 8300 46121 8309 46155
rect 8309 46121 8343 46155
rect 8343 46121 8352 46155
rect 8300 46112 8352 46121
rect 8668 46112 8720 46164
rect 8944 46112 8996 46164
rect 5540 45840 5592 45892
rect 8392 45840 8444 45892
rect 9312 45840 9364 45892
rect 2504 45772 2556 45824
rect 4160 45772 4212 45824
rect 7380 45772 7432 45824
rect 8300 45772 8352 45824
rect 8944 45772 8996 45824
rect 2950 45670 3002 45722
rect 3014 45670 3066 45722
rect 3078 45670 3130 45722
rect 3142 45670 3194 45722
rect 3206 45670 3258 45722
rect 4550 45670 4602 45722
rect 4614 45670 4666 45722
rect 4678 45670 4730 45722
rect 4742 45670 4794 45722
rect 4806 45670 4858 45722
rect 6150 45670 6202 45722
rect 6214 45670 6266 45722
rect 6278 45670 6330 45722
rect 6342 45670 6394 45722
rect 6406 45670 6458 45722
rect 7750 45670 7802 45722
rect 7814 45670 7866 45722
rect 7878 45670 7930 45722
rect 7942 45670 7994 45722
rect 8006 45670 8058 45722
rect 9350 45670 9402 45722
rect 9414 45670 9466 45722
rect 9478 45670 9530 45722
rect 9542 45670 9594 45722
rect 9606 45670 9658 45722
rect 7840 45568 7892 45620
rect 8392 45568 8444 45620
rect 1492 45543 1544 45552
rect 1492 45509 1501 45543
rect 1501 45509 1535 45543
rect 1535 45509 1544 45543
rect 1492 45500 1544 45509
rect 4252 45432 4304 45484
rect 4620 45475 4672 45484
rect 4620 45441 4629 45475
rect 4629 45441 4663 45475
rect 4663 45441 4672 45475
rect 4620 45432 4672 45441
rect 9128 45500 9180 45552
rect 4988 45432 5040 45484
rect 5448 45432 5500 45484
rect 7012 45432 7064 45484
rect 940 45228 992 45280
rect 4160 45228 4212 45280
rect 4252 45228 4304 45280
rect 4988 45296 5040 45348
rect 8760 45432 8812 45484
rect 7472 45271 7524 45280
rect 7472 45237 7481 45271
rect 7481 45237 7515 45271
rect 7515 45237 7524 45271
rect 7472 45228 7524 45237
rect 7656 45271 7708 45280
rect 7656 45237 7665 45271
rect 7665 45237 7699 45271
rect 7699 45237 7708 45271
rect 7656 45228 7708 45237
rect 9128 45296 9180 45348
rect 9220 45228 9272 45280
rect 3610 45126 3662 45178
rect 3674 45126 3726 45178
rect 3738 45126 3790 45178
rect 3802 45126 3854 45178
rect 3866 45126 3918 45178
rect 5210 45126 5262 45178
rect 5274 45126 5326 45178
rect 5338 45126 5390 45178
rect 5402 45126 5454 45178
rect 5466 45126 5518 45178
rect 6810 45126 6862 45178
rect 6874 45126 6926 45178
rect 6938 45126 6990 45178
rect 7002 45126 7054 45178
rect 7066 45126 7118 45178
rect 8410 45126 8462 45178
rect 8474 45126 8526 45178
rect 8538 45126 8590 45178
rect 8602 45126 8654 45178
rect 8666 45126 8718 45178
rect 4344 45067 4396 45076
rect 4344 45033 4353 45067
rect 4353 45033 4387 45067
rect 4387 45033 4396 45067
rect 4344 45024 4396 45033
rect 4620 45024 4672 45076
rect 2320 44956 2372 45008
rect 5632 44956 5684 45008
rect 9220 44956 9272 45008
rect 9588 44956 9640 45008
rect 2044 44888 2096 44940
rect 4528 44888 4580 44940
rect 940 44820 992 44872
rect 4620 44863 4672 44872
rect 4620 44829 4629 44863
rect 4629 44829 4663 44863
rect 4663 44829 4672 44863
rect 4620 44820 4672 44829
rect 5264 44863 5316 44872
rect 5264 44829 5273 44863
rect 5273 44829 5307 44863
rect 5307 44829 5316 44863
rect 5264 44820 5316 44829
rect 7840 44888 7892 44940
rect 8116 44888 8168 44940
rect 5448 44863 5500 44872
rect 5448 44829 5457 44863
rect 5457 44829 5491 44863
rect 5491 44829 5500 44863
rect 5448 44820 5500 44829
rect 5908 44820 5960 44872
rect 2688 44684 2740 44736
rect 3516 44684 3568 44736
rect 7748 44752 7800 44804
rect 5908 44684 5960 44736
rect 6092 44684 6144 44736
rect 2950 44582 3002 44634
rect 3014 44582 3066 44634
rect 3078 44582 3130 44634
rect 3142 44582 3194 44634
rect 3206 44582 3258 44634
rect 4550 44582 4602 44634
rect 4614 44582 4666 44634
rect 4678 44582 4730 44634
rect 4742 44582 4794 44634
rect 4806 44582 4858 44634
rect 6150 44582 6202 44634
rect 6214 44582 6266 44634
rect 6278 44582 6330 44634
rect 6342 44582 6394 44634
rect 6406 44582 6458 44634
rect 7750 44582 7802 44634
rect 7814 44582 7866 44634
rect 7878 44582 7930 44634
rect 7942 44582 7994 44634
rect 8006 44582 8058 44634
rect 9350 44582 9402 44634
rect 9414 44582 9466 44634
rect 9478 44582 9530 44634
rect 9542 44582 9594 44634
rect 9606 44582 9658 44634
rect 4712 44480 4764 44532
rect 5264 44480 5316 44532
rect 7656 44480 7708 44532
rect 7748 44480 7800 44532
rect 8208 44480 8260 44532
rect 2872 44344 2924 44396
rect 4344 44387 4396 44396
rect 4344 44353 4377 44387
rect 4377 44353 4396 44387
rect 4344 44344 4396 44353
rect 4712 44344 4764 44396
rect 5080 44387 5132 44396
rect 5080 44353 5089 44387
rect 5089 44353 5123 44387
rect 5123 44353 5132 44387
rect 5080 44344 5132 44353
rect 5172 44387 5224 44396
rect 5172 44353 5181 44387
rect 5181 44353 5215 44387
rect 5215 44353 5224 44387
rect 5172 44344 5224 44353
rect 6644 44344 6696 44396
rect 7564 44344 7616 44396
rect 8116 44344 8168 44396
rect 4896 44276 4948 44328
rect 4712 44208 4764 44260
rect 6736 44208 6788 44260
rect 4344 44140 4396 44192
rect 8116 44183 8168 44192
rect 8116 44149 8125 44183
rect 8125 44149 8159 44183
rect 8159 44149 8168 44183
rect 8116 44140 8168 44149
rect 8208 44140 8260 44192
rect 3610 44038 3662 44090
rect 3674 44038 3726 44090
rect 3738 44038 3790 44090
rect 3802 44038 3854 44090
rect 3866 44038 3918 44090
rect 5210 44038 5262 44090
rect 5274 44038 5326 44090
rect 5338 44038 5390 44090
rect 5402 44038 5454 44090
rect 5466 44038 5518 44090
rect 6810 44038 6862 44090
rect 6874 44038 6926 44090
rect 6938 44038 6990 44090
rect 7002 44038 7054 44090
rect 7066 44038 7118 44090
rect 8410 44038 8462 44090
rect 8474 44038 8526 44090
rect 8538 44038 8590 44090
rect 8602 44038 8654 44090
rect 8666 44038 8718 44090
rect 4068 43936 4120 43988
rect 940 43732 992 43784
rect 8208 43936 8260 43988
rect 6644 43800 6696 43852
rect 8760 43732 8812 43784
rect 9036 43732 9088 43784
rect 4896 43596 4948 43648
rect 7196 43596 7248 43648
rect 9036 43596 9088 43648
rect 2950 43494 3002 43546
rect 3014 43494 3066 43546
rect 3078 43494 3130 43546
rect 3142 43494 3194 43546
rect 3206 43494 3258 43546
rect 4550 43494 4602 43546
rect 4614 43494 4666 43546
rect 4678 43494 4730 43546
rect 4742 43494 4794 43546
rect 4806 43494 4858 43546
rect 6150 43494 6202 43546
rect 6214 43494 6266 43546
rect 6278 43494 6330 43546
rect 6342 43494 6394 43546
rect 6406 43494 6458 43546
rect 7750 43494 7802 43546
rect 7814 43494 7866 43546
rect 7878 43494 7930 43546
rect 7942 43494 7994 43546
rect 8006 43494 8058 43546
rect 9350 43494 9402 43546
rect 9414 43494 9466 43546
rect 9478 43494 9530 43546
rect 9542 43494 9594 43546
rect 9606 43494 9658 43546
rect 7748 43392 7800 43444
rect 8208 43392 8260 43444
rect 7656 43324 7708 43376
rect 8668 43324 8720 43376
rect 6644 43256 6696 43308
rect 8116 43095 8168 43104
rect 8116 43061 8125 43095
rect 8125 43061 8159 43095
rect 8159 43061 8168 43095
rect 8116 43052 8168 43061
rect 3610 42950 3662 43002
rect 3674 42950 3726 43002
rect 3738 42950 3790 43002
rect 3802 42950 3854 43002
rect 3866 42950 3918 43002
rect 5210 42950 5262 43002
rect 5274 42950 5326 43002
rect 5338 42950 5390 43002
rect 5402 42950 5454 43002
rect 5466 42950 5518 43002
rect 6810 42950 6862 43002
rect 6874 42950 6926 43002
rect 6938 42950 6990 43002
rect 7002 42950 7054 43002
rect 7066 42950 7118 43002
rect 8410 42950 8462 43002
rect 8474 42950 8526 43002
rect 8538 42950 8590 43002
rect 8602 42950 8654 43002
rect 8666 42950 8718 43002
rect 3976 42780 4028 42832
rect 3332 42712 3384 42764
rect 1952 42644 2004 42696
rect 2596 42644 2648 42696
rect 4528 42712 4580 42764
rect 940 42576 992 42628
rect 5264 42644 5316 42696
rect 5908 42848 5960 42900
rect 7196 42780 7248 42832
rect 8668 42780 8720 42832
rect 5724 42712 5776 42764
rect 7748 42712 7800 42764
rect 5448 42687 5500 42696
rect 5448 42653 5457 42687
rect 5457 42653 5491 42687
rect 5491 42653 5500 42687
rect 5448 42644 5500 42653
rect 8300 42644 8352 42696
rect 8576 42644 8628 42696
rect 8852 42644 8904 42696
rect 3884 42508 3936 42560
rect 4068 42508 4120 42560
rect 4344 42508 4396 42560
rect 5540 42576 5592 42628
rect 5080 42508 5132 42560
rect 5172 42551 5224 42560
rect 5172 42517 5181 42551
rect 5181 42517 5215 42551
rect 5215 42517 5224 42551
rect 5172 42508 5224 42517
rect 5264 42508 5316 42560
rect 7380 42508 7432 42560
rect 7748 42508 7800 42560
rect 8300 42508 8352 42560
rect 2950 42406 3002 42458
rect 3014 42406 3066 42458
rect 3078 42406 3130 42458
rect 3142 42406 3194 42458
rect 3206 42406 3258 42458
rect 4550 42406 4602 42458
rect 4614 42406 4666 42458
rect 4678 42406 4730 42458
rect 4742 42406 4794 42458
rect 4806 42406 4858 42458
rect 6150 42406 6202 42458
rect 6214 42406 6266 42458
rect 6278 42406 6330 42458
rect 6342 42406 6394 42458
rect 6406 42406 6458 42458
rect 7750 42406 7802 42458
rect 7814 42406 7866 42458
rect 7878 42406 7930 42458
rect 7942 42406 7994 42458
rect 8006 42406 8058 42458
rect 9350 42406 9402 42458
rect 9414 42406 9466 42458
rect 9478 42406 9530 42458
rect 9542 42406 9594 42458
rect 9606 42406 9658 42458
rect 2504 42304 2556 42356
rect 3976 42304 4028 42356
rect 5264 42304 5316 42356
rect 7748 42304 7800 42356
rect 9956 42304 10008 42356
rect 5448 42236 5500 42288
rect 7288 42236 7340 42288
rect 2596 42168 2648 42220
rect 6644 42168 6696 42220
rect 10048 42168 10100 42220
rect 1584 42032 1636 42084
rect 3332 42032 3384 42084
rect 3884 42032 3936 42084
rect 1952 41964 2004 42016
rect 5172 41964 5224 42016
rect 5540 41964 5592 42016
rect 7380 41964 7432 42016
rect 8576 41964 8628 42016
rect 8852 41964 8904 42016
rect 3610 41862 3662 41914
rect 3674 41862 3726 41914
rect 3738 41862 3790 41914
rect 3802 41862 3854 41914
rect 3866 41862 3918 41914
rect 5210 41862 5262 41914
rect 5274 41862 5326 41914
rect 5338 41862 5390 41914
rect 5402 41862 5454 41914
rect 5466 41862 5518 41914
rect 6810 41862 6862 41914
rect 6874 41862 6926 41914
rect 6938 41862 6990 41914
rect 7002 41862 7054 41914
rect 7066 41862 7118 41914
rect 8410 41862 8462 41914
rect 8474 41862 8526 41914
rect 8538 41862 8590 41914
rect 8602 41862 8654 41914
rect 8666 41862 8718 41914
rect 4160 41760 4212 41812
rect 2780 41692 2832 41744
rect 4528 41556 4580 41608
rect 4896 41556 4948 41608
rect 7288 41556 7340 41608
rect 7656 41556 7708 41608
rect 940 41488 992 41540
rect 2136 41488 2188 41540
rect 2504 41420 2556 41472
rect 2950 41318 3002 41370
rect 3014 41318 3066 41370
rect 3078 41318 3130 41370
rect 3142 41318 3194 41370
rect 3206 41318 3258 41370
rect 4550 41318 4602 41370
rect 4614 41318 4666 41370
rect 4678 41318 4730 41370
rect 4742 41318 4794 41370
rect 4806 41318 4858 41370
rect 6150 41318 6202 41370
rect 6214 41318 6266 41370
rect 6278 41318 6330 41370
rect 6342 41318 6394 41370
rect 6406 41318 6458 41370
rect 7750 41318 7802 41370
rect 7814 41318 7866 41370
rect 7878 41318 7930 41370
rect 7942 41318 7994 41370
rect 8006 41318 8058 41370
rect 9350 41318 9402 41370
rect 9414 41318 9466 41370
rect 9478 41318 9530 41370
rect 9542 41318 9594 41370
rect 9606 41318 9658 41370
rect 1032 41080 1084 41132
rect 4068 40876 4120 40928
rect 3610 40774 3662 40826
rect 3674 40774 3726 40826
rect 3738 40774 3790 40826
rect 3802 40774 3854 40826
rect 3866 40774 3918 40826
rect 5210 40774 5262 40826
rect 5274 40774 5326 40826
rect 5338 40774 5390 40826
rect 5402 40774 5454 40826
rect 5466 40774 5518 40826
rect 6810 40774 6862 40826
rect 6874 40774 6926 40826
rect 6938 40774 6990 40826
rect 7002 40774 7054 40826
rect 7066 40774 7118 40826
rect 8410 40774 8462 40826
rect 8474 40774 8526 40826
rect 8538 40774 8590 40826
rect 8602 40774 8654 40826
rect 8666 40774 8718 40826
rect 5632 40672 5684 40724
rect 6828 40672 6880 40724
rect 4344 40536 4396 40588
rect 4804 40536 4856 40588
rect 572 40468 624 40520
rect 2596 40468 2648 40520
rect 7564 40604 7616 40656
rect 9128 40672 9180 40724
rect 8024 40604 8076 40656
rect 4344 40400 4396 40452
rect 5908 40400 5960 40452
rect 6000 40400 6052 40452
rect 7104 40400 7156 40452
rect 4804 40332 4856 40384
rect 4988 40332 5040 40384
rect 5632 40332 5684 40384
rect 7564 40468 7616 40520
rect 8852 40536 8904 40588
rect 8392 40332 8444 40384
rect 2950 40230 3002 40282
rect 3014 40230 3066 40282
rect 3078 40230 3130 40282
rect 3142 40230 3194 40282
rect 3206 40230 3258 40282
rect 4550 40230 4602 40282
rect 4614 40230 4666 40282
rect 4678 40230 4730 40282
rect 4742 40230 4794 40282
rect 4806 40230 4858 40282
rect 6150 40230 6202 40282
rect 6214 40230 6266 40282
rect 6278 40230 6330 40282
rect 6342 40230 6394 40282
rect 6406 40230 6458 40282
rect 7750 40230 7802 40282
rect 7814 40230 7866 40282
rect 7878 40230 7930 40282
rect 7942 40230 7994 40282
rect 8006 40230 8058 40282
rect 9350 40230 9402 40282
rect 9414 40230 9466 40282
rect 9478 40230 9530 40282
rect 9542 40230 9594 40282
rect 9606 40230 9658 40282
rect 4804 40128 4856 40180
rect 5172 40128 5224 40180
rect 5816 40128 5868 40180
rect 7104 40128 7156 40180
rect 7472 40128 7524 40180
rect 1492 40103 1544 40112
rect 1492 40069 1501 40103
rect 1501 40069 1535 40103
rect 1535 40069 1544 40103
rect 1492 40060 1544 40069
rect 7656 40060 7708 40112
rect 8944 40171 8996 40180
rect 8944 40137 8953 40171
rect 8953 40137 8987 40171
rect 8987 40137 8996 40171
rect 8944 40128 8996 40137
rect 9956 40060 10008 40112
rect 7472 39924 7524 39976
rect 8024 39924 8076 39976
rect 8116 39924 8168 39976
rect 8300 39967 8352 39976
rect 8300 39933 8309 39967
rect 8309 39933 8343 39967
rect 8343 39933 8352 39967
rect 8300 39924 8352 39933
rect 9036 40035 9088 40044
rect 9036 40001 9045 40035
rect 9045 40001 9079 40035
rect 9079 40001 9088 40035
rect 9036 39992 9088 40001
rect 9128 39992 9180 40044
rect 6828 39856 6880 39908
rect 2688 39788 2740 39840
rect 8852 39788 8904 39840
rect 3610 39686 3662 39738
rect 3674 39686 3726 39738
rect 3738 39686 3790 39738
rect 3802 39686 3854 39738
rect 3866 39686 3918 39738
rect 5210 39686 5262 39738
rect 5274 39686 5326 39738
rect 5338 39686 5390 39738
rect 5402 39686 5454 39738
rect 5466 39686 5518 39738
rect 6810 39686 6862 39738
rect 6874 39686 6926 39738
rect 6938 39686 6990 39738
rect 7002 39686 7054 39738
rect 7066 39686 7118 39738
rect 8410 39686 8462 39738
rect 8474 39686 8526 39738
rect 8538 39686 8590 39738
rect 8602 39686 8654 39738
rect 8666 39686 8718 39738
rect 4344 39584 4396 39636
rect 5540 39584 5592 39636
rect 6920 39584 6972 39636
rect 5448 39516 5500 39568
rect 7472 39516 7524 39568
rect 7564 39448 7616 39500
rect 7656 39448 7708 39500
rect 7840 39491 7892 39500
rect 7840 39457 7849 39491
rect 7849 39457 7883 39491
rect 7883 39457 7892 39491
rect 7840 39448 7892 39457
rect 664 39380 716 39432
rect 5540 39380 5592 39432
rect 7288 39380 7340 39432
rect 4160 39244 4212 39296
rect 6000 39244 6052 39296
rect 6920 39244 6972 39296
rect 7564 39244 7616 39296
rect 2950 39142 3002 39194
rect 3014 39142 3066 39194
rect 3078 39142 3130 39194
rect 3142 39142 3194 39194
rect 3206 39142 3258 39194
rect 4550 39142 4602 39194
rect 4614 39142 4666 39194
rect 4678 39142 4730 39194
rect 4742 39142 4794 39194
rect 4806 39142 4858 39194
rect 6150 39142 6202 39194
rect 6214 39142 6266 39194
rect 6278 39142 6330 39194
rect 6342 39142 6394 39194
rect 6406 39142 6458 39194
rect 7750 39142 7802 39194
rect 7814 39142 7866 39194
rect 7878 39142 7930 39194
rect 7942 39142 7994 39194
rect 8006 39142 8058 39194
rect 9350 39142 9402 39194
rect 9414 39142 9466 39194
rect 9478 39142 9530 39194
rect 9542 39142 9594 39194
rect 9606 39142 9658 39194
rect 1308 39040 1360 39092
rect 4068 38972 4120 39024
rect 1032 38904 1084 38956
rect 5540 38904 5592 38956
rect 6736 38972 6788 39024
rect 7288 38904 7340 38956
rect 2780 38700 2832 38752
rect 7656 38879 7708 38888
rect 7656 38845 7665 38879
rect 7665 38845 7699 38879
rect 7699 38845 7708 38879
rect 7656 38836 7708 38845
rect 6828 38768 6880 38820
rect 6644 38700 6696 38752
rect 9128 38700 9180 38752
rect 11704 38700 11756 38752
rect 3610 38598 3662 38650
rect 3674 38598 3726 38650
rect 3738 38598 3790 38650
rect 3802 38598 3854 38650
rect 3866 38598 3918 38650
rect 5210 38598 5262 38650
rect 5274 38598 5326 38650
rect 5338 38598 5390 38650
rect 5402 38598 5454 38650
rect 5466 38598 5518 38650
rect 6810 38598 6862 38650
rect 6874 38598 6926 38650
rect 6938 38598 6990 38650
rect 7002 38598 7054 38650
rect 7066 38598 7118 38650
rect 8410 38598 8462 38650
rect 8474 38598 8526 38650
rect 8538 38598 8590 38650
rect 8602 38598 8654 38650
rect 8666 38598 8718 38650
rect 1860 38496 1912 38548
rect 2872 38496 2924 38548
rect 11520 38428 11572 38480
rect 7104 38224 7156 38276
rect 7656 38224 7708 38276
rect 8116 38156 8168 38208
rect 2950 38054 3002 38106
rect 3014 38054 3066 38106
rect 3078 38054 3130 38106
rect 3142 38054 3194 38106
rect 3206 38054 3258 38106
rect 4550 38054 4602 38106
rect 4614 38054 4666 38106
rect 4678 38054 4730 38106
rect 4742 38054 4794 38106
rect 4806 38054 4858 38106
rect 6150 38054 6202 38106
rect 6214 38054 6266 38106
rect 6278 38054 6330 38106
rect 6342 38054 6394 38106
rect 6406 38054 6458 38106
rect 7750 38054 7802 38106
rect 7814 38054 7866 38106
rect 7878 38054 7930 38106
rect 7942 38054 7994 38106
rect 8006 38054 8058 38106
rect 9350 38054 9402 38106
rect 9414 38054 9466 38106
rect 9478 38054 9530 38106
rect 9542 38054 9594 38106
rect 9606 38054 9658 38106
rect 7196 37952 7248 38004
rect 7380 37952 7432 38004
rect 8208 37952 8260 38004
rect 1032 37816 1084 37868
rect 7472 37748 7524 37800
rect 8116 37791 8168 37800
rect 8116 37757 8125 37791
rect 8125 37757 8159 37791
rect 8159 37757 8168 37791
rect 8116 37748 8168 37757
rect 2320 37612 2372 37664
rect 4344 37612 4396 37664
rect 7472 37612 7524 37664
rect 11980 37612 12032 37664
rect 3610 37510 3662 37562
rect 3674 37510 3726 37562
rect 3738 37510 3790 37562
rect 3802 37510 3854 37562
rect 3866 37510 3918 37562
rect 5210 37510 5262 37562
rect 5274 37510 5326 37562
rect 5338 37510 5390 37562
rect 5402 37510 5454 37562
rect 5466 37510 5518 37562
rect 6810 37510 6862 37562
rect 6874 37510 6926 37562
rect 6938 37510 6990 37562
rect 7002 37510 7054 37562
rect 7066 37510 7118 37562
rect 8410 37510 8462 37562
rect 8474 37510 8526 37562
rect 8538 37510 8590 37562
rect 8602 37510 8654 37562
rect 8666 37510 8718 37562
rect 2688 37408 2740 37460
rect 7380 37408 7432 37460
rect 8852 37340 8904 37392
rect 6920 37315 6972 37324
rect 6920 37281 6929 37315
rect 6929 37281 6963 37315
rect 6963 37281 6972 37315
rect 6920 37272 6972 37281
rect 7748 37315 7800 37324
rect 7748 37281 7757 37315
rect 7757 37281 7791 37315
rect 7791 37281 7800 37315
rect 7748 37272 7800 37281
rect 1032 37204 1084 37256
rect 1860 37204 1912 37256
rect 4988 37204 5040 37256
rect 5540 37204 5592 37256
rect 2412 37136 2464 37188
rect 480 37068 532 37120
rect 7104 37068 7156 37120
rect 9772 37204 9824 37256
rect 7380 37068 7432 37120
rect 2950 36966 3002 37018
rect 3014 36966 3066 37018
rect 3078 36966 3130 37018
rect 3142 36966 3194 37018
rect 3206 36966 3258 37018
rect 4550 36966 4602 37018
rect 4614 36966 4666 37018
rect 4678 36966 4730 37018
rect 4742 36966 4794 37018
rect 4806 36966 4858 37018
rect 6150 36966 6202 37018
rect 6214 36966 6266 37018
rect 6278 36966 6330 37018
rect 6342 36966 6394 37018
rect 6406 36966 6458 37018
rect 7750 36966 7802 37018
rect 7814 36966 7866 37018
rect 7878 36966 7930 37018
rect 7942 36966 7994 37018
rect 8006 36966 8058 37018
rect 9350 36966 9402 37018
rect 9414 36966 9466 37018
rect 9478 36966 9530 37018
rect 9542 36966 9594 37018
rect 9606 36966 9658 37018
rect 7104 36796 7156 36848
rect 8300 36864 8352 36916
rect 11612 36864 11664 36916
rect 4988 36592 5040 36644
rect 5448 36592 5500 36644
rect 6460 36592 6512 36644
rect 6644 36592 6696 36644
rect 8852 36660 8904 36712
rect 9220 36592 9272 36644
rect 848 36524 900 36576
rect 3610 36422 3662 36474
rect 3674 36422 3726 36474
rect 3738 36422 3790 36474
rect 3802 36422 3854 36474
rect 3866 36422 3918 36474
rect 5210 36422 5262 36474
rect 5274 36422 5326 36474
rect 5338 36422 5390 36474
rect 5402 36422 5454 36474
rect 5466 36422 5518 36474
rect 6810 36422 6862 36474
rect 6874 36422 6926 36474
rect 6938 36422 6990 36474
rect 7002 36422 7054 36474
rect 7066 36422 7118 36474
rect 8410 36422 8462 36474
rect 8474 36422 8526 36474
rect 8538 36422 8590 36474
rect 8602 36422 8654 36474
rect 8666 36422 8718 36474
rect 1676 36184 1728 36236
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 1216 36048 1268 36100
rect 8852 36184 8904 36236
rect 9128 36116 9180 36168
rect 6552 35980 6604 36032
rect 7196 35980 7248 36032
rect 7656 35980 7708 36032
rect 8852 36048 8904 36100
rect 2950 35878 3002 35930
rect 3014 35878 3066 35930
rect 3078 35878 3130 35930
rect 3142 35878 3194 35930
rect 3206 35878 3258 35930
rect 4550 35878 4602 35930
rect 4614 35878 4666 35930
rect 4678 35878 4730 35930
rect 4742 35878 4794 35930
rect 4806 35878 4858 35930
rect 6150 35878 6202 35930
rect 6214 35878 6266 35930
rect 6278 35878 6330 35930
rect 6342 35878 6394 35930
rect 6406 35878 6458 35930
rect 7750 35878 7802 35930
rect 7814 35878 7866 35930
rect 7878 35878 7930 35930
rect 7942 35878 7994 35930
rect 8006 35878 8058 35930
rect 9350 35878 9402 35930
rect 9414 35878 9466 35930
rect 9478 35878 9530 35930
rect 9542 35878 9594 35930
rect 9606 35878 9658 35930
rect 2228 35776 2280 35828
rect 7196 35776 7248 35828
rect 1124 35708 1176 35760
rect 8300 35708 8352 35760
rect 4068 35640 4120 35692
rect 4896 35640 4948 35692
rect 3610 35334 3662 35386
rect 3674 35334 3726 35386
rect 3738 35334 3790 35386
rect 3802 35334 3854 35386
rect 3866 35334 3918 35386
rect 5210 35334 5262 35386
rect 5274 35334 5326 35386
rect 5338 35334 5390 35386
rect 5402 35334 5454 35386
rect 5466 35334 5518 35386
rect 6810 35334 6862 35386
rect 6874 35334 6926 35386
rect 6938 35334 6990 35386
rect 7002 35334 7054 35386
rect 7066 35334 7118 35386
rect 8410 35334 8462 35386
rect 8474 35334 8526 35386
rect 8538 35334 8590 35386
rect 8602 35334 8654 35386
rect 8666 35334 8718 35386
rect 848 35232 900 35284
rect 1308 35232 1360 35284
rect 2688 35096 2740 35148
rect 3332 35096 3384 35148
rect 940 35028 992 35080
rect 2872 34892 2924 34944
rect 2950 34790 3002 34842
rect 3014 34790 3066 34842
rect 3078 34790 3130 34842
rect 3142 34790 3194 34842
rect 3206 34790 3258 34842
rect 4550 34790 4602 34842
rect 4614 34790 4666 34842
rect 4678 34790 4730 34842
rect 4742 34790 4794 34842
rect 4806 34790 4858 34842
rect 6150 34790 6202 34842
rect 6214 34790 6266 34842
rect 6278 34790 6330 34842
rect 6342 34790 6394 34842
rect 6406 34790 6458 34842
rect 7750 34790 7802 34842
rect 7814 34790 7866 34842
rect 7878 34790 7930 34842
rect 7942 34790 7994 34842
rect 8006 34790 8058 34842
rect 9350 34790 9402 34842
rect 9414 34790 9466 34842
rect 9478 34790 9530 34842
rect 9542 34790 9594 34842
rect 9606 34790 9658 34842
rect 10692 34688 10744 34740
rect 1768 34620 1820 34672
rect 9036 34552 9088 34604
rect 8852 34484 8904 34536
rect 3610 34246 3662 34298
rect 3674 34246 3726 34298
rect 3738 34246 3790 34298
rect 3802 34246 3854 34298
rect 3866 34246 3918 34298
rect 5210 34246 5262 34298
rect 5274 34246 5326 34298
rect 5338 34246 5390 34298
rect 5402 34246 5454 34298
rect 5466 34246 5518 34298
rect 6810 34246 6862 34298
rect 6874 34246 6926 34298
rect 6938 34246 6990 34298
rect 7002 34246 7054 34298
rect 7066 34246 7118 34298
rect 8410 34246 8462 34298
rect 8474 34246 8526 34298
rect 8538 34246 8590 34298
rect 8602 34246 8654 34298
rect 8666 34246 8718 34298
rect 3332 34144 3384 34196
rect 3884 34144 3936 34196
rect 11888 34076 11940 34128
rect 8576 34051 8628 34060
rect 8576 34017 8585 34051
rect 8585 34017 8619 34051
rect 8619 34017 8628 34051
rect 8576 34008 8628 34017
rect 940 33940 992 33992
rect 7196 33872 7248 33924
rect 8668 33915 8720 33924
rect 8668 33881 8677 33915
rect 8677 33881 8711 33915
rect 8711 33881 8720 33915
rect 8668 33872 8720 33881
rect 8852 33872 8904 33924
rect 3332 33804 3384 33856
rect 8484 33804 8536 33856
rect 8944 33804 8996 33856
rect 2950 33702 3002 33754
rect 3014 33702 3066 33754
rect 3078 33702 3130 33754
rect 3142 33702 3194 33754
rect 3206 33702 3258 33754
rect 4550 33702 4602 33754
rect 4614 33702 4666 33754
rect 4678 33702 4730 33754
rect 4742 33702 4794 33754
rect 4806 33702 4858 33754
rect 6150 33702 6202 33754
rect 6214 33702 6266 33754
rect 6278 33702 6330 33754
rect 6342 33702 6394 33754
rect 6406 33702 6458 33754
rect 7750 33702 7802 33754
rect 7814 33702 7866 33754
rect 7878 33702 7930 33754
rect 7942 33702 7994 33754
rect 8006 33702 8058 33754
rect 9350 33702 9402 33754
rect 9414 33702 9466 33754
rect 9478 33702 9530 33754
rect 9542 33702 9594 33754
rect 9606 33702 9658 33754
rect 3884 33600 3936 33652
rect 8668 33600 8720 33652
rect 9312 33600 9364 33652
rect 8116 33532 8168 33584
rect 1492 33507 1544 33516
rect 1492 33473 1501 33507
rect 1501 33473 1535 33507
rect 1535 33473 1544 33507
rect 1492 33464 1544 33473
rect 8392 33507 8444 33516
rect 8392 33473 8401 33507
rect 8401 33473 8435 33507
rect 8435 33473 8444 33507
rect 8392 33464 8444 33473
rect 8944 33464 8996 33516
rect 7288 33396 7340 33448
rect 8484 33396 8536 33448
rect 1124 33328 1176 33380
rect 7472 33260 7524 33312
rect 3610 33158 3662 33210
rect 3674 33158 3726 33210
rect 3738 33158 3790 33210
rect 3802 33158 3854 33210
rect 3866 33158 3918 33210
rect 5210 33158 5262 33210
rect 5274 33158 5326 33210
rect 5338 33158 5390 33210
rect 5402 33158 5454 33210
rect 5466 33158 5518 33210
rect 6810 33158 6862 33210
rect 6874 33158 6926 33210
rect 6938 33158 6990 33210
rect 7002 33158 7054 33210
rect 7066 33158 7118 33210
rect 8410 33158 8462 33210
rect 8474 33158 8526 33210
rect 8538 33158 8590 33210
rect 8602 33158 8654 33210
rect 8666 33158 8718 33210
rect 6552 33056 6604 33108
rect 7104 33056 7156 33108
rect 8668 33056 8720 33108
rect 9312 33056 9364 33108
rect 10508 32988 10560 33040
rect 8944 32920 8996 32972
rect 2136 32852 2188 32904
rect 8116 32852 8168 32904
rect 6644 32784 6696 32836
rect 9864 32784 9916 32836
rect 2950 32614 3002 32666
rect 3014 32614 3066 32666
rect 3078 32614 3130 32666
rect 3142 32614 3194 32666
rect 3206 32614 3258 32666
rect 4550 32614 4602 32666
rect 4614 32614 4666 32666
rect 4678 32614 4730 32666
rect 4742 32614 4794 32666
rect 4806 32614 4858 32666
rect 6150 32614 6202 32666
rect 6214 32614 6266 32666
rect 6278 32614 6330 32666
rect 6342 32614 6394 32666
rect 6406 32614 6458 32666
rect 7750 32614 7802 32666
rect 7814 32614 7866 32666
rect 7878 32614 7930 32666
rect 7942 32614 7994 32666
rect 8006 32614 8058 32666
rect 9350 32614 9402 32666
rect 9414 32614 9466 32666
rect 9478 32614 9530 32666
rect 9542 32614 9594 32666
rect 9606 32614 9658 32666
rect 8208 32512 8260 32564
rect 8668 32512 8720 32564
rect 9312 32512 9364 32564
rect 6552 32444 6604 32496
rect 8024 32444 8076 32496
rect 940 32376 992 32428
rect 7196 32376 7248 32428
rect 7472 32376 7524 32428
rect 7748 32308 7800 32360
rect 8208 32308 8260 32360
rect 8852 32308 8904 32360
rect 10600 32308 10652 32360
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 4896 32172 4948 32224
rect 7288 32172 7340 32224
rect 7840 32172 7892 32224
rect 10784 32172 10836 32224
rect 3610 32070 3662 32122
rect 3674 32070 3726 32122
rect 3738 32070 3790 32122
rect 3802 32070 3854 32122
rect 3866 32070 3918 32122
rect 5210 32070 5262 32122
rect 5274 32070 5326 32122
rect 5338 32070 5390 32122
rect 5402 32070 5454 32122
rect 5466 32070 5518 32122
rect 6810 32070 6862 32122
rect 6874 32070 6926 32122
rect 6938 32070 6990 32122
rect 7002 32070 7054 32122
rect 7066 32070 7118 32122
rect 8410 32070 8462 32122
rect 8474 32070 8526 32122
rect 8538 32070 8590 32122
rect 8602 32070 8654 32122
rect 8666 32070 8718 32122
rect 1032 31968 1084 32020
rect 8116 31968 8168 32020
rect 5448 31900 5500 31952
rect 5908 31900 5960 31952
rect 7472 31900 7524 31952
rect 7656 31900 7708 31952
rect 9220 31968 9272 32020
rect 10140 31968 10192 32020
rect 1768 31832 1820 31884
rect 7748 31832 7800 31884
rect 8116 31832 8168 31884
rect 7196 31764 7248 31816
rect 7840 31764 7892 31816
rect 9588 31900 9640 31952
rect 8208 31696 8260 31748
rect 10048 31696 10100 31748
rect 7564 31628 7616 31680
rect 7748 31628 7800 31680
rect 2950 31526 3002 31578
rect 3014 31526 3066 31578
rect 3078 31526 3130 31578
rect 3142 31526 3194 31578
rect 3206 31526 3258 31578
rect 4550 31526 4602 31578
rect 4614 31526 4666 31578
rect 4678 31526 4730 31578
rect 4742 31526 4794 31578
rect 4806 31526 4858 31578
rect 6150 31526 6202 31578
rect 6214 31526 6266 31578
rect 6278 31526 6330 31578
rect 6342 31526 6394 31578
rect 6406 31526 6458 31578
rect 7750 31526 7802 31578
rect 7814 31526 7866 31578
rect 7878 31526 7930 31578
rect 7942 31526 7994 31578
rect 8006 31526 8058 31578
rect 9350 31526 9402 31578
rect 9414 31526 9466 31578
rect 9478 31526 9530 31578
rect 9542 31526 9594 31578
rect 9606 31526 9658 31578
rect 7380 31424 7432 31476
rect 8116 31424 8168 31476
rect 5908 31356 5960 31408
rect 7012 31356 7064 31408
rect 940 31288 992 31340
rect 5448 31288 5500 31340
rect 6092 31288 6144 31340
rect 7564 31288 7616 31340
rect 1584 31152 1636 31204
rect 2688 31152 2740 31204
rect 7380 31152 7432 31204
rect 7472 31084 7524 31136
rect 3610 30982 3662 31034
rect 3674 30982 3726 31034
rect 3738 30982 3790 31034
rect 3802 30982 3854 31034
rect 3866 30982 3918 31034
rect 5210 30982 5262 31034
rect 5274 30982 5326 31034
rect 5338 30982 5390 31034
rect 5402 30982 5454 31034
rect 5466 30982 5518 31034
rect 6810 30982 6862 31034
rect 6874 30982 6926 31034
rect 6938 30982 6990 31034
rect 7002 30982 7054 31034
rect 7066 30982 7118 31034
rect 8410 30982 8462 31034
rect 8474 30982 8526 31034
rect 8538 30982 8590 31034
rect 8602 30982 8654 31034
rect 8666 30982 8718 31034
rect 2950 30438 3002 30490
rect 3014 30438 3066 30490
rect 3078 30438 3130 30490
rect 3142 30438 3194 30490
rect 3206 30438 3258 30490
rect 4550 30438 4602 30490
rect 4614 30438 4666 30490
rect 4678 30438 4730 30490
rect 4742 30438 4794 30490
rect 4806 30438 4858 30490
rect 6150 30438 6202 30490
rect 6214 30438 6266 30490
rect 6278 30438 6330 30490
rect 6342 30438 6394 30490
rect 6406 30438 6458 30490
rect 7750 30438 7802 30490
rect 7814 30438 7866 30490
rect 7878 30438 7930 30490
rect 7942 30438 7994 30490
rect 8006 30438 8058 30490
rect 9350 30438 9402 30490
rect 9414 30438 9466 30490
rect 9478 30438 9530 30490
rect 9542 30438 9594 30490
rect 9606 30438 9658 30490
rect 4160 30268 4212 30320
rect 4804 30268 4856 30320
rect 9220 30268 9272 30320
rect 940 30200 992 30252
rect 7288 30200 7340 30252
rect 4160 30132 4212 30184
rect 4988 30132 5040 30184
rect 4988 29996 5040 30048
rect 3610 29894 3662 29946
rect 3674 29894 3726 29946
rect 3738 29894 3790 29946
rect 3802 29894 3854 29946
rect 3866 29894 3918 29946
rect 5210 29894 5262 29946
rect 5274 29894 5326 29946
rect 5338 29894 5390 29946
rect 5402 29894 5454 29946
rect 5466 29894 5518 29946
rect 6810 29894 6862 29946
rect 6874 29894 6926 29946
rect 6938 29894 6990 29946
rect 7002 29894 7054 29946
rect 7066 29894 7118 29946
rect 8410 29894 8462 29946
rect 8474 29894 8526 29946
rect 8538 29894 8590 29946
rect 8602 29894 8654 29946
rect 8666 29894 8718 29946
rect 5632 29656 5684 29708
rect 5724 29656 5776 29708
rect 6828 29656 6880 29708
rect 940 29588 992 29640
rect 4804 29520 4856 29572
rect 5172 29520 5224 29572
rect 5540 29452 5592 29504
rect 5632 29452 5684 29504
rect 2950 29350 3002 29402
rect 3014 29350 3066 29402
rect 3078 29350 3130 29402
rect 3142 29350 3194 29402
rect 3206 29350 3258 29402
rect 4550 29350 4602 29402
rect 4614 29350 4666 29402
rect 4678 29350 4730 29402
rect 4742 29350 4794 29402
rect 4806 29350 4858 29402
rect 6150 29350 6202 29402
rect 6214 29350 6266 29402
rect 6278 29350 6330 29402
rect 6342 29350 6394 29402
rect 6406 29350 6458 29402
rect 7750 29350 7802 29402
rect 7814 29350 7866 29402
rect 7878 29350 7930 29402
rect 7942 29350 7994 29402
rect 8006 29350 8058 29402
rect 9350 29350 9402 29402
rect 9414 29350 9466 29402
rect 9478 29350 9530 29402
rect 9542 29350 9594 29402
rect 9606 29350 9658 29402
rect 6736 29248 6788 29300
rect 8852 29223 8904 29232
rect 8852 29189 8861 29223
rect 8861 29189 8895 29223
rect 8895 29189 8904 29223
rect 8852 29180 8904 29189
rect 8944 29180 8996 29232
rect 9864 29180 9916 29232
rect 7288 29155 7340 29164
rect 7288 29121 7297 29155
rect 7297 29121 7331 29155
rect 7331 29121 7340 29155
rect 7288 29112 7340 29121
rect 11888 29112 11940 29164
rect 4804 28908 4856 28960
rect 5172 28908 5224 28960
rect 6828 28908 6880 28960
rect 7840 28908 7892 28960
rect 9036 28908 9088 28960
rect 3610 28806 3662 28858
rect 3674 28806 3726 28858
rect 3738 28806 3790 28858
rect 3802 28806 3854 28858
rect 3866 28806 3918 28858
rect 5210 28806 5262 28858
rect 5274 28806 5326 28858
rect 5338 28806 5390 28858
rect 5402 28806 5454 28858
rect 5466 28806 5518 28858
rect 6810 28806 6862 28858
rect 6874 28806 6926 28858
rect 6938 28806 6990 28858
rect 7002 28806 7054 28858
rect 7066 28806 7118 28858
rect 8410 28806 8462 28858
rect 8474 28806 8526 28858
rect 8538 28806 8590 28858
rect 8602 28806 8654 28858
rect 8666 28806 8718 28858
rect 6092 28704 6144 28756
rect 7012 28704 7064 28756
rect 9220 28704 9272 28756
rect 7196 28636 7248 28688
rect 7656 28611 7708 28620
rect 7656 28577 7665 28611
rect 7665 28577 7699 28611
rect 7699 28577 7708 28611
rect 7656 28568 7708 28577
rect 940 28500 992 28552
rect 6092 28500 6144 28552
rect 6828 28500 6880 28552
rect 7472 28543 7524 28552
rect 7472 28509 7481 28543
rect 7481 28509 7515 28543
rect 7515 28509 7524 28543
rect 7472 28500 7524 28509
rect 7840 28636 7892 28688
rect 10324 28636 10376 28688
rect 1400 28407 1452 28416
rect 1400 28373 1409 28407
rect 1409 28373 1443 28407
rect 1443 28373 1452 28407
rect 1400 28364 1452 28373
rect 4804 28364 4856 28416
rect 5448 28364 5500 28416
rect 5816 28364 5868 28416
rect 6000 28364 6052 28416
rect 7196 28364 7248 28416
rect 7748 28364 7800 28416
rect 8208 28568 8260 28620
rect 8484 28568 8536 28620
rect 8852 28568 8904 28620
rect 8760 28500 8812 28552
rect 8116 28364 8168 28416
rect 2950 28262 3002 28314
rect 3014 28262 3066 28314
rect 3078 28262 3130 28314
rect 3142 28262 3194 28314
rect 3206 28262 3258 28314
rect 4550 28262 4602 28314
rect 4614 28262 4666 28314
rect 4678 28262 4730 28314
rect 4742 28262 4794 28314
rect 4806 28262 4858 28314
rect 6150 28262 6202 28314
rect 6214 28262 6266 28314
rect 6278 28262 6330 28314
rect 6342 28262 6394 28314
rect 6406 28262 6458 28314
rect 7750 28262 7802 28314
rect 7814 28262 7866 28314
rect 7878 28262 7930 28314
rect 7942 28262 7994 28314
rect 8006 28262 8058 28314
rect 9350 28262 9402 28314
rect 9414 28262 9466 28314
rect 9478 28262 9530 28314
rect 9542 28262 9594 28314
rect 9606 28262 9658 28314
rect 1400 28160 1452 28212
rect 5816 28160 5868 28212
rect 2596 27820 2648 27872
rect 3332 27820 3384 27872
rect 3610 27718 3662 27770
rect 3674 27718 3726 27770
rect 3738 27718 3790 27770
rect 3802 27718 3854 27770
rect 3866 27718 3918 27770
rect 5210 27718 5262 27770
rect 5274 27718 5326 27770
rect 5338 27718 5390 27770
rect 5402 27718 5454 27770
rect 5466 27718 5518 27770
rect 6810 27718 6862 27770
rect 6874 27718 6926 27770
rect 6938 27718 6990 27770
rect 7002 27718 7054 27770
rect 7066 27718 7118 27770
rect 8410 27718 8462 27770
rect 8474 27718 8526 27770
rect 8538 27718 8590 27770
rect 8602 27718 8654 27770
rect 8666 27718 8718 27770
rect 3332 27616 3384 27668
rect 4160 27616 4212 27668
rect 7656 27616 7708 27668
rect 940 27412 992 27464
rect 1676 27387 1728 27396
rect 1676 27353 1685 27387
rect 1685 27353 1719 27387
rect 1719 27353 1728 27387
rect 1676 27344 1728 27353
rect 6920 27344 6972 27396
rect 7380 27344 7432 27396
rect 2950 27174 3002 27226
rect 3014 27174 3066 27226
rect 3078 27174 3130 27226
rect 3142 27174 3194 27226
rect 3206 27174 3258 27226
rect 4550 27174 4602 27226
rect 4614 27174 4666 27226
rect 4678 27174 4730 27226
rect 4742 27174 4794 27226
rect 4806 27174 4858 27226
rect 6150 27174 6202 27226
rect 6214 27174 6266 27226
rect 6278 27174 6330 27226
rect 6342 27174 6394 27226
rect 6406 27174 6458 27226
rect 7750 27174 7802 27226
rect 7814 27174 7866 27226
rect 7878 27174 7930 27226
rect 7942 27174 7994 27226
rect 8006 27174 8058 27226
rect 9350 27174 9402 27226
rect 9414 27174 9466 27226
rect 9478 27174 9530 27226
rect 9542 27174 9594 27226
rect 9606 27174 9658 27226
rect 5540 27072 5592 27124
rect 8208 27072 8260 27124
rect 11612 27072 11664 27124
rect 6460 26936 6512 26988
rect 7104 26936 7156 26988
rect 6092 26868 6144 26920
rect 6920 26868 6972 26920
rect 7656 26868 7708 26920
rect 756 26800 808 26852
rect 9496 26800 9548 26852
rect 6644 26732 6696 26784
rect 6828 26732 6880 26784
rect 8208 26732 8260 26784
rect 8944 26732 8996 26784
rect 10048 26732 10100 26784
rect 3610 26630 3662 26682
rect 3674 26630 3726 26682
rect 3738 26630 3790 26682
rect 3802 26630 3854 26682
rect 3866 26630 3918 26682
rect 5210 26630 5262 26682
rect 5274 26630 5326 26682
rect 5338 26630 5390 26682
rect 5402 26630 5454 26682
rect 5466 26630 5518 26682
rect 6810 26630 6862 26682
rect 6874 26630 6926 26682
rect 6938 26630 6990 26682
rect 7002 26630 7054 26682
rect 7066 26630 7118 26682
rect 8410 26630 8462 26682
rect 8474 26630 8526 26682
rect 8538 26630 8590 26682
rect 8602 26630 8654 26682
rect 8666 26630 8718 26682
rect 7380 26528 7432 26580
rect 7564 26528 7616 26580
rect 5356 26460 5408 26512
rect 6460 26460 6512 26512
rect 8944 26460 8996 26512
rect 940 26324 992 26376
rect 7104 26392 7156 26444
rect 7472 26392 7524 26444
rect 7656 26392 7708 26444
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 4988 26324 5040 26376
rect 5540 26324 5592 26376
rect 6552 26324 6604 26376
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 7012 26367 7064 26376
rect 7012 26333 7021 26367
rect 7021 26333 7055 26367
rect 7055 26333 7064 26367
rect 7012 26324 7064 26333
rect 7196 26367 7248 26376
rect 7196 26333 7205 26367
rect 7205 26333 7239 26367
rect 7239 26333 7248 26367
rect 7196 26324 7248 26333
rect 9496 26571 9548 26580
rect 9496 26537 9505 26571
rect 9505 26537 9539 26571
rect 9539 26537 9548 26571
rect 9496 26528 9548 26537
rect 10140 26528 10192 26580
rect 2872 26188 2924 26240
rect 4160 26231 4212 26240
rect 4160 26197 4169 26231
rect 4169 26197 4203 26231
rect 4203 26197 4212 26231
rect 4160 26188 4212 26197
rect 9588 26256 9640 26308
rect 10416 26256 10468 26308
rect 8392 26188 8444 26240
rect 2950 26086 3002 26138
rect 3014 26086 3066 26138
rect 3078 26086 3130 26138
rect 3142 26086 3194 26138
rect 3206 26086 3258 26138
rect 4550 26086 4602 26138
rect 4614 26086 4666 26138
rect 4678 26086 4730 26138
rect 4742 26086 4794 26138
rect 4806 26086 4858 26138
rect 6150 26086 6202 26138
rect 6214 26086 6266 26138
rect 6278 26086 6330 26138
rect 6342 26086 6394 26138
rect 6406 26086 6458 26138
rect 7750 26086 7802 26138
rect 7814 26086 7866 26138
rect 7878 26086 7930 26138
rect 7942 26086 7994 26138
rect 8006 26086 8058 26138
rect 9350 26086 9402 26138
rect 9414 26086 9466 26138
rect 9478 26086 9530 26138
rect 9542 26086 9594 26138
rect 9606 26086 9658 26138
rect 1584 26027 1636 26036
rect 1584 25993 1593 26027
rect 1593 25993 1627 26027
rect 1627 25993 1636 26027
rect 1584 25984 1636 25993
rect 4988 25984 5040 26036
rect 5356 25984 5408 26036
rect 5816 25984 5868 26036
rect 7656 25984 7708 26036
rect 8392 26027 8444 26036
rect 8392 25993 8401 26027
rect 8401 25993 8435 26027
rect 8435 25993 8444 26027
rect 8392 25984 8444 25993
rect 9128 26027 9180 26036
rect 9128 25993 9137 26027
rect 9137 25993 9171 26027
rect 9171 25993 9180 26027
rect 9128 25984 9180 25993
rect 940 25848 992 25900
rect 5908 25916 5960 25968
rect 6920 25916 6972 25968
rect 5540 25848 5592 25900
rect 5816 25891 5868 25900
rect 5816 25857 5825 25891
rect 5825 25857 5859 25891
rect 5859 25857 5868 25891
rect 5816 25848 5868 25857
rect 6184 25848 6236 25900
rect 7012 25848 7064 25900
rect 7564 25848 7616 25900
rect 8116 25916 8168 25968
rect 5908 25780 5960 25832
rect 7104 25780 7156 25832
rect 7656 25823 7708 25832
rect 7656 25789 7665 25823
rect 7665 25789 7699 25823
rect 7699 25789 7708 25823
rect 7656 25780 7708 25789
rect 8024 25848 8076 25900
rect 7288 25712 7340 25764
rect 7840 25780 7892 25832
rect 8760 25780 8812 25832
rect 1768 25644 1820 25696
rect 7656 25644 7708 25696
rect 8760 25644 8812 25696
rect 3610 25542 3662 25594
rect 3674 25542 3726 25594
rect 3738 25542 3790 25594
rect 3802 25542 3854 25594
rect 3866 25542 3918 25594
rect 5210 25542 5262 25594
rect 5274 25542 5326 25594
rect 5338 25542 5390 25594
rect 5402 25542 5454 25594
rect 5466 25542 5518 25594
rect 6810 25542 6862 25594
rect 6874 25542 6926 25594
rect 6938 25542 6990 25594
rect 7002 25542 7054 25594
rect 7066 25542 7118 25594
rect 8410 25542 8462 25594
rect 8474 25542 8526 25594
rect 8538 25542 8590 25594
rect 8602 25542 8654 25594
rect 8666 25542 8718 25594
rect 2780 25440 2832 25492
rect 7196 25440 7248 25492
rect 7840 25372 7892 25424
rect 9588 25372 9640 25424
rect 1584 25304 1636 25356
rect 6184 25304 6236 25356
rect 4988 25100 5040 25152
rect 7288 25100 7340 25152
rect 2950 24998 3002 25050
rect 3014 24998 3066 25050
rect 3078 24998 3130 25050
rect 3142 24998 3194 25050
rect 3206 24998 3258 25050
rect 4550 24998 4602 25050
rect 4614 24998 4666 25050
rect 4678 24998 4730 25050
rect 4742 24998 4794 25050
rect 4806 24998 4858 25050
rect 6150 24998 6202 25050
rect 6214 24998 6266 25050
rect 6278 24998 6330 25050
rect 6342 24998 6394 25050
rect 6406 24998 6458 25050
rect 7750 24998 7802 25050
rect 7814 24998 7866 25050
rect 7878 24998 7930 25050
rect 7942 24998 7994 25050
rect 8006 24998 8058 25050
rect 9350 24998 9402 25050
rect 9414 24998 9466 25050
rect 9478 24998 9530 25050
rect 9542 24998 9594 25050
rect 9606 24998 9658 25050
rect 5540 24896 5592 24948
rect 7932 24896 7984 24948
rect 940 24760 992 24812
rect 6644 24760 6696 24812
rect 11060 24760 11112 24812
rect 2320 24692 2372 24744
rect 7748 24692 7800 24744
rect 8116 24692 8168 24744
rect 9312 24692 9364 24744
rect 848 24556 900 24608
rect 3610 24454 3662 24506
rect 3674 24454 3726 24506
rect 3738 24454 3790 24506
rect 3802 24454 3854 24506
rect 3866 24454 3918 24506
rect 5210 24454 5262 24506
rect 5274 24454 5326 24506
rect 5338 24454 5390 24506
rect 5402 24454 5454 24506
rect 5466 24454 5518 24506
rect 6810 24454 6862 24506
rect 6874 24454 6926 24506
rect 6938 24454 6990 24506
rect 7002 24454 7054 24506
rect 7066 24454 7118 24506
rect 8410 24454 8462 24506
rect 8474 24454 8526 24506
rect 8538 24454 8590 24506
rect 8602 24454 8654 24506
rect 8666 24454 8718 24506
rect 7380 24352 7432 24404
rect 7840 24352 7892 24404
rect 8300 24352 8352 24404
rect 10876 24352 10928 24404
rect 7472 24284 7524 24336
rect 8116 24327 8168 24336
rect 8116 24293 8125 24327
rect 8125 24293 8159 24327
rect 8159 24293 8168 24327
rect 8116 24284 8168 24293
rect 9220 24284 9272 24336
rect 2596 24148 2648 24200
rect 5724 24148 5776 24200
rect 2872 24080 2924 24132
rect 5816 24080 5868 24132
rect 2228 24012 2280 24064
rect 4988 24012 5040 24064
rect 5724 24012 5776 24064
rect 7288 24148 7340 24200
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 7932 24216 7984 24268
rect 7840 24080 7892 24132
rect 7748 24012 7800 24064
rect 8392 24012 8444 24064
rect 2950 23910 3002 23962
rect 3014 23910 3066 23962
rect 3078 23910 3130 23962
rect 3142 23910 3194 23962
rect 3206 23910 3258 23962
rect 4550 23910 4602 23962
rect 4614 23910 4666 23962
rect 4678 23910 4730 23962
rect 4742 23910 4794 23962
rect 4806 23910 4858 23962
rect 6150 23910 6202 23962
rect 6214 23910 6266 23962
rect 6278 23910 6330 23962
rect 6342 23910 6394 23962
rect 6406 23910 6458 23962
rect 7750 23910 7802 23962
rect 7814 23910 7866 23962
rect 7878 23910 7930 23962
rect 7942 23910 7994 23962
rect 8006 23910 8058 23962
rect 9350 23910 9402 23962
rect 9414 23910 9466 23962
rect 9478 23910 9530 23962
rect 9542 23910 9594 23962
rect 9606 23910 9658 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 7472 23808 7524 23860
rect 8300 23808 8352 23860
rect 940 23672 992 23724
rect 5632 23672 5684 23724
rect 8392 23604 8444 23656
rect 9312 23604 9364 23656
rect 2412 23536 2464 23588
rect 4988 23536 5040 23588
rect 3332 23468 3384 23520
rect 3610 23366 3662 23418
rect 3674 23366 3726 23418
rect 3738 23366 3790 23418
rect 3802 23366 3854 23418
rect 3866 23366 3918 23418
rect 5210 23366 5262 23418
rect 5274 23366 5326 23418
rect 5338 23366 5390 23418
rect 5402 23366 5454 23418
rect 5466 23366 5518 23418
rect 6810 23366 6862 23418
rect 6874 23366 6926 23418
rect 6938 23366 6990 23418
rect 7002 23366 7054 23418
rect 7066 23366 7118 23418
rect 8410 23366 8462 23418
rect 8474 23366 8526 23418
rect 8538 23366 8590 23418
rect 8602 23366 8654 23418
rect 8666 23366 8718 23418
rect 3240 23264 3292 23316
rect 3608 23264 3660 23316
rect 9220 23264 9272 23316
rect 11428 23264 11480 23316
rect 5816 23196 5868 23248
rect 10048 23196 10100 23248
rect 6000 23060 6052 23112
rect 8208 23060 8260 23112
rect 8944 23060 8996 23112
rect 9588 22992 9640 23044
rect 2320 22924 2372 22976
rect 7380 22924 7432 22976
rect 8208 22924 8260 22976
rect 8944 22924 8996 22976
rect 2950 22822 3002 22874
rect 3014 22822 3066 22874
rect 3078 22822 3130 22874
rect 3142 22822 3194 22874
rect 3206 22822 3258 22874
rect 4550 22822 4602 22874
rect 4614 22822 4666 22874
rect 4678 22822 4730 22874
rect 4742 22822 4794 22874
rect 4806 22822 4858 22874
rect 6150 22822 6202 22874
rect 6214 22822 6266 22874
rect 6278 22822 6330 22874
rect 6342 22822 6394 22874
rect 6406 22822 6458 22874
rect 7750 22822 7802 22874
rect 7814 22822 7866 22874
rect 7878 22822 7930 22874
rect 7942 22822 7994 22874
rect 8006 22822 8058 22874
rect 9350 22822 9402 22874
rect 9414 22822 9466 22874
rect 9478 22822 9530 22874
rect 9542 22822 9594 22874
rect 9606 22822 9658 22874
rect 3056 22720 3108 22772
rect 3516 22720 3568 22772
rect 4252 22720 4304 22772
rect 4528 22720 4580 22772
rect 2872 22652 2924 22704
rect 940 22584 992 22636
rect 6552 22652 6604 22704
rect 7196 22652 7248 22704
rect 9956 22584 10008 22636
rect 3976 22380 4028 22432
rect 4620 22380 4672 22432
rect 7840 22423 7892 22432
rect 7840 22389 7849 22423
rect 7849 22389 7883 22423
rect 7883 22389 7892 22423
rect 7840 22380 7892 22389
rect 3610 22278 3662 22330
rect 3674 22278 3726 22330
rect 3738 22278 3790 22330
rect 3802 22278 3854 22330
rect 3866 22278 3918 22330
rect 5210 22278 5262 22330
rect 5274 22278 5326 22330
rect 5338 22278 5390 22330
rect 5402 22278 5454 22330
rect 5466 22278 5518 22330
rect 6810 22278 6862 22330
rect 6874 22278 6926 22330
rect 6938 22278 6990 22330
rect 7002 22278 7054 22330
rect 7066 22278 7118 22330
rect 8410 22278 8462 22330
rect 8474 22278 8526 22330
rect 8538 22278 8590 22330
rect 8602 22278 8654 22330
rect 8666 22278 8718 22330
rect 4252 22108 4304 22160
rect 4620 22108 4672 22160
rect 7656 22040 7708 22092
rect 940 21972 992 22024
rect 4528 21972 4580 22024
rect 5908 21904 5960 21956
rect 2136 21836 2188 21888
rect 6736 21836 6788 21888
rect 2950 21734 3002 21786
rect 3014 21734 3066 21786
rect 3078 21734 3130 21786
rect 3142 21734 3194 21786
rect 3206 21734 3258 21786
rect 4550 21734 4602 21786
rect 4614 21734 4666 21786
rect 4678 21734 4730 21786
rect 4742 21734 4794 21786
rect 4806 21734 4858 21786
rect 6150 21734 6202 21786
rect 6214 21734 6266 21786
rect 6278 21734 6330 21786
rect 6342 21734 6394 21786
rect 6406 21734 6458 21786
rect 7750 21734 7802 21786
rect 7814 21734 7866 21786
rect 7878 21734 7930 21786
rect 7942 21734 7994 21786
rect 8006 21734 8058 21786
rect 9350 21734 9402 21786
rect 9414 21734 9466 21786
rect 9478 21734 9530 21786
rect 9542 21734 9594 21786
rect 9606 21734 9658 21786
rect 5724 21496 5776 21548
rect 7288 21496 7340 21548
rect 7472 21428 7524 21480
rect 7564 21335 7616 21344
rect 7564 21301 7573 21335
rect 7573 21301 7607 21335
rect 7607 21301 7616 21335
rect 7564 21292 7616 21301
rect 3610 21190 3662 21242
rect 3674 21190 3726 21242
rect 3738 21190 3790 21242
rect 3802 21190 3854 21242
rect 3866 21190 3918 21242
rect 5210 21190 5262 21242
rect 5274 21190 5326 21242
rect 5338 21190 5390 21242
rect 5402 21190 5454 21242
rect 5466 21190 5518 21242
rect 6810 21190 6862 21242
rect 6874 21190 6926 21242
rect 6938 21190 6990 21242
rect 7002 21190 7054 21242
rect 7066 21190 7118 21242
rect 8410 21190 8462 21242
rect 8474 21190 8526 21242
rect 8538 21190 8590 21242
rect 8602 21190 8654 21242
rect 8666 21190 8718 21242
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 6000 20816 6052 20868
rect 6736 20748 6788 20800
rect 7380 20748 7432 20800
rect 2950 20646 3002 20698
rect 3014 20646 3066 20698
rect 3078 20646 3130 20698
rect 3142 20646 3194 20698
rect 3206 20646 3258 20698
rect 4550 20646 4602 20698
rect 4614 20646 4666 20698
rect 4678 20646 4730 20698
rect 4742 20646 4794 20698
rect 4806 20646 4858 20698
rect 6150 20646 6202 20698
rect 6214 20646 6266 20698
rect 6278 20646 6330 20698
rect 6342 20646 6394 20698
rect 6406 20646 6458 20698
rect 7750 20646 7802 20698
rect 7814 20646 7866 20698
rect 7878 20646 7930 20698
rect 7942 20646 7994 20698
rect 8006 20646 8058 20698
rect 9350 20646 9402 20698
rect 9414 20646 9466 20698
rect 9478 20646 9530 20698
rect 9542 20646 9594 20698
rect 9606 20646 9658 20698
rect 8760 20408 8812 20460
rect 8852 20204 8904 20256
rect 9588 20204 9640 20256
rect 3610 20102 3662 20154
rect 3674 20102 3726 20154
rect 3738 20102 3790 20154
rect 3802 20102 3854 20154
rect 3866 20102 3918 20154
rect 5210 20102 5262 20154
rect 5274 20102 5326 20154
rect 5338 20102 5390 20154
rect 5402 20102 5454 20154
rect 5466 20102 5518 20154
rect 6810 20102 6862 20154
rect 6874 20102 6926 20154
rect 6938 20102 6990 20154
rect 7002 20102 7054 20154
rect 7066 20102 7118 20154
rect 8410 20102 8462 20154
rect 8474 20102 8526 20154
rect 8538 20102 8590 20154
rect 8602 20102 8654 20154
rect 8666 20102 8718 20154
rect 940 19796 992 19848
rect 8300 19796 8352 19848
rect 5724 19728 5776 19780
rect 9036 19660 9088 19712
rect 2950 19558 3002 19610
rect 3014 19558 3066 19610
rect 3078 19558 3130 19610
rect 3142 19558 3194 19610
rect 3206 19558 3258 19610
rect 4550 19558 4602 19610
rect 4614 19558 4666 19610
rect 4678 19558 4730 19610
rect 4742 19558 4794 19610
rect 4806 19558 4858 19610
rect 6150 19558 6202 19610
rect 6214 19558 6266 19610
rect 6278 19558 6330 19610
rect 6342 19558 6394 19610
rect 6406 19558 6458 19610
rect 7750 19558 7802 19610
rect 7814 19558 7866 19610
rect 7878 19558 7930 19610
rect 7942 19558 7994 19610
rect 8006 19558 8058 19610
rect 9350 19558 9402 19610
rect 9414 19558 9466 19610
rect 9478 19558 9530 19610
rect 9542 19558 9594 19610
rect 9606 19558 9658 19610
rect 3610 19014 3662 19066
rect 3674 19014 3726 19066
rect 3738 19014 3790 19066
rect 3802 19014 3854 19066
rect 3866 19014 3918 19066
rect 5210 19014 5262 19066
rect 5274 19014 5326 19066
rect 5338 19014 5390 19066
rect 5402 19014 5454 19066
rect 5466 19014 5518 19066
rect 6810 19014 6862 19066
rect 6874 19014 6926 19066
rect 6938 19014 6990 19066
rect 7002 19014 7054 19066
rect 7066 19014 7118 19066
rect 8410 19014 8462 19066
rect 8474 19014 8526 19066
rect 8538 19014 8590 19066
rect 8602 19014 8654 19066
rect 8666 19014 8718 19066
rect 7288 18912 7340 18964
rect 7656 18912 7708 18964
rect 7196 18844 7248 18896
rect 7748 18844 7800 18896
rect 3424 18776 3476 18828
rect 7288 18776 7340 18828
rect 4896 18708 4948 18760
rect 940 18640 992 18692
rect 7288 18640 7340 18692
rect 8208 18708 8260 18760
rect 6736 18572 6788 18624
rect 2950 18470 3002 18522
rect 3014 18470 3066 18522
rect 3078 18470 3130 18522
rect 3142 18470 3194 18522
rect 3206 18470 3258 18522
rect 4550 18470 4602 18522
rect 4614 18470 4666 18522
rect 4678 18470 4730 18522
rect 4742 18470 4794 18522
rect 4806 18470 4858 18522
rect 6150 18470 6202 18522
rect 6214 18470 6266 18522
rect 6278 18470 6330 18522
rect 6342 18470 6394 18522
rect 6406 18470 6458 18522
rect 7750 18470 7802 18522
rect 7814 18470 7866 18522
rect 7878 18470 7930 18522
rect 7942 18470 7994 18522
rect 8006 18470 8058 18522
rect 9350 18470 9402 18522
rect 9414 18470 9466 18522
rect 9478 18470 9530 18522
rect 9542 18470 9594 18522
rect 9606 18470 9658 18522
rect 2596 18300 2648 18352
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3610 17926 3662 17978
rect 3674 17926 3726 17978
rect 3738 17926 3790 17978
rect 3802 17926 3854 17978
rect 3866 17926 3918 17978
rect 5210 17926 5262 17978
rect 5274 17926 5326 17978
rect 5338 17926 5390 17978
rect 5402 17926 5454 17978
rect 5466 17926 5518 17978
rect 6810 17926 6862 17978
rect 6874 17926 6926 17978
rect 6938 17926 6990 17978
rect 7002 17926 7054 17978
rect 7066 17926 7118 17978
rect 8410 17926 8462 17978
rect 8474 17926 8526 17978
rect 8538 17926 8590 17978
rect 8602 17926 8654 17978
rect 8666 17926 8718 17978
rect 7288 17688 7340 17740
rect 7472 17688 7524 17740
rect 8300 17484 8352 17536
rect 2950 17382 3002 17434
rect 3014 17382 3066 17434
rect 3078 17382 3130 17434
rect 3142 17382 3194 17434
rect 3206 17382 3258 17434
rect 4550 17382 4602 17434
rect 4614 17382 4666 17434
rect 4678 17382 4730 17434
rect 4742 17382 4794 17434
rect 4806 17382 4858 17434
rect 6150 17382 6202 17434
rect 6214 17382 6266 17434
rect 6278 17382 6330 17434
rect 6342 17382 6394 17434
rect 6406 17382 6458 17434
rect 7750 17382 7802 17434
rect 7814 17382 7866 17434
rect 7878 17382 7930 17434
rect 7942 17382 7994 17434
rect 8006 17382 8058 17434
rect 9350 17382 9402 17434
rect 9414 17382 9466 17434
rect 9478 17382 9530 17434
rect 9542 17382 9594 17434
rect 9606 17382 9658 17434
rect 7564 17280 7616 17332
rect 2044 17212 2096 17264
rect 940 16940 992 16992
rect 7564 16940 7616 16992
rect 3610 16838 3662 16890
rect 3674 16838 3726 16890
rect 3738 16838 3790 16890
rect 3802 16838 3854 16890
rect 3866 16838 3918 16890
rect 5210 16838 5262 16890
rect 5274 16838 5326 16890
rect 5338 16838 5390 16890
rect 5402 16838 5454 16890
rect 5466 16838 5518 16890
rect 6810 16838 6862 16890
rect 6874 16838 6926 16890
rect 6938 16838 6990 16890
rect 7002 16838 7054 16890
rect 7066 16838 7118 16890
rect 8410 16838 8462 16890
rect 8474 16838 8526 16890
rect 8538 16838 8590 16890
rect 8602 16838 8654 16890
rect 8666 16838 8718 16890
rect 7196 16736 7248 16788
rect 8208 16711 8260 16720
rect 8208 16677 8217 16711
rect 8217 16677 8251 16711
rect 8251 16677 8260 16711
rect 8208 16668 8260 16677
rect 7656 16532 7708 16584
rect 8300 16575 8352 16584
rect 8300 16541 8309 16575
rect 8309 16541 8343 16575
rect 8343 16541 8352 16575
rect 8300 16532 8352 16541
rect 9864 16532 9916 16584
rect 7288 16396 7340 16448
rect 7472 16439 7524 16448
rect 7472 16405 7481 16439
rect 7481 16405 7515 16439
rect 7515 16405 7524 16439
rect 7472 16396 7524 16405
rect 8852 16464 8904 16516
rect 8300 16396 8352 16448
rect 2950 16294 3002 16346
rect 3014 16294 3066 16346
rect 3078 16294 3130 16346
rect 3142 16294 3194 16346
rect 3206 16294 3258 16346
rect 4550 16294 4602 16346
rect 4614 16294 4666 16346
rect 4678 16294 4730 16346
rect 4742 16294 4794 16346
rect 4806 16294 4858 16346
rect 6150 16294 6202 16346
rect 6214 16294 6266 16346
rect 6278 16294 6330 16346
rect 6342 16294 6394 16346
rect 6406 16294 6458 16346
rect 7750 16294 7802 16346
rect 7814 16294 7866 16346
rect 7878 16294 7930 16346
rect 7942 16294 7994 16346
rect 8006 16294 8058 16346
rect 9350 16294 9402 16346
rect 9414 16294 9466 16346
rect 9478 16294 9530 16346
rect 9542 16294 9594 16346
rect 9606 16294 9658 16346
rect 7656 16192 7708 16244
rect 4344 16124 4396 16176
rect 8760 16124 8812 16176
rect 9864 16192 9916 16244
rect 8208 15988 8260 16040
rect 940 15852 992 15904
rect 5632 15852 5684 15904
rect 3610 15750 3662 15802
rect 3674 15750 3726 15802
rect 3738 15750 3790 15802
rect 3802 15750 3854 15802
rect 3866 15750 3918 15802
rect 5210 15750 5262 15802
rect 5274 15750 5326 15802
rect 5338 15750 5390 15802
rect 5402 15750 5454 15802
rect 5466 15750 5518 15802
rect 6810 15750 6862 15802
rect 6874 15750 6926 15802
rect 6938 15750 6990 15802
rect 7002 15750 7054 15802
rect 7066 15750 7118 15802
rect 8410 15750 8462 15802
rect 8474 15750 8526 15802
rect 8538 15750 8590 15802
rect 8602 15750 8654 15802
rect 8666 15750 8718 15802
rect 9036 15512 9088 15564
rect 9220 15512 9272 15564
rect 3516 15444 3568 15496
rect 9220 15308 9272 15360
rect 2950 15206 3002 15258
rect 3014 15206 3066 15258
rect 3078 15206 3130 15258
rect 3142 15206 3194 15258
rect 3206 15206 3258 15258
rect 4550 15206 4602 15258
rect 4614 15206 4666 15258
rect 4678 15206 4730 15258
rect 4742 15206 4794 15258
rect 4806 15206 4858 15258
rect 6150 15206 6202 15258
rect 6214 15206 6266 15258
rect 6278 15206 6330 15258
rect 6342 15206 6394 15258
rect 6406 15206 6458 15258
rect 7750 15206 7802 15258
rect 7814 15206 7866 15258
rect 7878 15206 7930 15258
rect 7942 15206 7994 15258
rect 8006 15206 8058 15258
rect 9350 15206 9402 15258
rect 9414 15206 9466 15258
rect 9478 15206 9530 15258
rect 9542 15206 9594 15258
rect 9606 15206 9658 15258
rect 4436 15036 4488 15088
rect 940 14764 992 14816
rect 3610 14662 3662 14714
rect 3674 14662 3726 14714
rect 3738 14662 3790 14714
rect 3802 14662 3854 14714
rect 3866 14662 3918 14714
rect 5210 14662 5262 14714
rect 5274 14662 5326 14714
rect 5338 14662 5390 14714
rect 5402 14662 5454 14714
rect 5466 14662 5518 14714
rect 6810 14662 6862 14714
rect 6874 14662 6926 14714
rect 6938 14662 6990 14714
rect 7002 14662 7054 14714
rect 7066 14662 7118 14714
rect 8410 14662 8462 14714
rect 8474 14662 8526 14714
rect 8538 14662 8590 14714
rect 8602 14662 8654 14714
rect 8666 14662 8718 14714
rect 7656 14492 7708 14544
rect 8208 14424 8260 14476
rect 8760 14424 8812 14476
rect 9036 14424 9088 14476
rect 4068 14356 4120 14408
rect 9772 14356 9824 14408
rect 7288 14288 7340 14340
rect 940 14220 992 14272
rect 9036 14220 9088 14272
rect 2950 14118 3002 14170
rect 3014 14118 3066 14170
rect 3078 14118 3130 14170
rect 3142 14118 3194 14170
rect 3206 14118 3258 14170
rect 4550 14118 4602 14170
rect 4614 14118 4666 14170
rect 4678 14118 4730 14170
rect 4742 14118 4794 14170
rect 4806 14118 4858 14170
rect 6150 14118 6202 14170
rect 6214 14118 6266 14170
rect 6278 14118 6330 14170
rect 6342 14118 6394 14170
rect 6406 14118 6458 14170
rect 7750 14118 7802 14170
rect 7814 14118 7866 14170
rect 7878 14118 7930 14170
rect 7942 14118 7994 14170
rect 8006 14118 8058 14170
rect 9350 14118 9402 14170
rect 9414 14118 9466 14170
rect 9478 14118 9530 14170
rect 9542 14118 9594 14170
rect 9606 14118 9658 14170
rect 3610 13574 3662 13626
rect 3674 13574 3726 13626
rect 3738 13574 3790 13626
rect 3802 13574 3854 13626
rect 3866 13574 3918 13626
rect 5210 13574 5262 13626
rect 5274 13574 5326 13626
rect 5338 13574 5390 13626
rect 5402 13574 5454 13626
rect 5466 13574 5518 13626
rect 6810 13574 6862 13626
rect 6874 13574 6926 13626
rect 6938 13574 6990 13626
rect 7002 13574 7054 13626
rect 7066 13574 7118 13626
rect 8410 13574 8462 13626
rect 8474 13574 8526 13626
rect 8538 13574 8590 13626
rect 8602 13574 8654 13626
rect 8666 13574 8718 13626
rect 7380 13336 7432 13388
rect 7564 13336 7616 13388
rect 1860 13268 1912 13320
rect 8024 13311 8076 13320
rect 8024 13277 8033 13311
rect 8033 13277 8067 13311
rect 8067 13277 8076 13311
rect 8024 13268 8076 13277
rect 7288 13200 7340 13252
rect 7564 13200 7616 13252
rect 940 13132 992 13184
rect 10968 13132 11020 13184
rect 2950 13030 3002 13082
rect 3014 13030 3066 13082
rect 3078 13030 3130 13082
rect 3142 13030 3194 13082
rect 3206 13030 3258 13082
rect 4550 13030 4602 13082
rect 4614 13030 4666 13082
rect 4678 13030 4730 13082
rect 4742 13030 4794 13082
rect 4806 13030 4858 13082
rect 6150 13030 6202 13082
rect 6214 13030 6266 13082
rect 6278 13030 6330 13082
rect 6342 13030 6394 13082
rect 6406 13030 6458 13082
rect 7750 13030 7802 13082
rect 7814 13030 7866 13082
rect 7878 13030 7930 13082
rect 7942 13030 7994 13082
rect 8006 13030 8058 13082
rect 9350 13030 9402 13082
rect 9414 13030 9466 13082
rect 9478 13030 9530 13082
rect 9542 13030 9594 13082
rect 9606 13030 9658 13082
rect 8944 12724 8996 12776
rect 9220 12724 9272 12776
rect 8944 12588 8996 12640
rect 9680 12588 9732 12640
rect 3610 12486 3662 12538
rect 3674 12486 3726 12538
rect 3738 12486 3790 12538
rect 3802 12486 3854 12538
rect 3866 12486 3918 12538
rect 5210 12486 5262 12538
rect 5274 12486 5326 12538
rect 5338 12486 5390 12538
rect 5402 12486 5454 12538
rect 5466 12486 5518 12538
rect 6810 12486 6862 12538
rect 6874 12486 6926 12538
rect 6938 12486 6990 12538
rect 7002 12486 7054 12538
rect 7066 12486 7118 12538
rect 8410 12486 8462 12538
rect 8474 12486 8526 12538
rect 8538 12486 8590 12538
rect 8602 12486 8654 12538
rect 8666 12486 8718 12538
rect 1952 12180 2004 12232
rect 940 12044 992 12096
rect 2950 11942 3002 11994
rect 3014 11942 3066 11994
rect 3078 11942 3130 11994
rect 3142 11942 3194 11994
rect 3206 11942 3258 11994
rect 4550 11942 4602 11994
rect 4614 11942 4666 11994
rect 4678 11942 4730 11994
rect 4742 11942 4794 11994
rect 4806 11942 4858 11994
rect 6150 11942 6202 11994
rect 6214 11942 6266 11994
rect 6278 11942 6330 11994
rect 6342 11942 6394 11994
rect 6406 11942 6458 11994
rect 7750 11942 7802 11994
rect 7814 11942 7866 11994
rect 7878 11942 7930 11994
rect 7942 11942 7994 11994
rect 8006 11942 8058 11994
rect 9350 11942 9402 11994
rect 9414 11942 9466 11994
rect 9478 11942 9530 11994
rect 9542 11942 9594 11994
rect 9606 11942 9658 11994
rect 6736 11840 6788 11892
rect 7380 11704 7432 11756
rect 8116 11500 8168 11552
rect 3610 11398 3662 11450
rect 3674 11398 3726 11450
rect 3738 11398 3790 11450
rect 3802 11398 3854 11450
rect 3866 11398 3918 11450
rect 5210 11398 5262 11450
rect 5274 11398 5326 11450
rect 5338 11398 5390 11450
rect 5402 11398 5454 11450
rect 5466 11398 5518 11450
rect 6810 11398 6862 11450
rect 6874 11398 6926 11450
rect 6938 11398 6990 11450
rect 7002 11398 7054 11450
rect 7066 11398 7118 11450
rect 8410 11398 8462 11450
rect 8474 11398 8526 11450
rect 8538 11398 8590 11450
rect 8602 11398 8654 11450
rect 8666 11398 8718 11450
rect 940 11296 992 11348
rect 5540 11296 5592 11348
rect 9588 11296 9640 11348
rect 10232 11228 10284 11280
rect 7380 11160 7432 11212
rect 2504 11092 2556 11144
rect 7472 11024 7524 11076
rect 2950 10854 3002 10906
rect 3014 10854 3066 10906
rect 3078 10854 3130 10906
rect 3142 10854 3194 10906
rect 3206 10854 3258 10906
rect 4550 10854 4602 10906
rect 4614 10854 4666 10906
rect 4678 10854 4730 10906
rect 4742 10854 4794 10906
rect 4806 10854 4858 10906
rect 6150 10854 6202 10906
rect 6214 10854 6266 10906
rect 6278 10854 6330 10906
rect 6342 10854 6394 10906
rect 6406 10854 6458 10906
rect 7750 10854 7802 10906
rect 7814 10854 7866 10906
rect 7878 10854 7930 10906
rect 7942 10854 7994 10906
rect 8006 10854 8058 10906
rect 9350 10854 9402 10906
rect 9414 10854 9466 10906
rect 9478 10854 9530 10906
rect 9542 10854 9594 10906
rect 9606 10854 9658 10906
rect 2228 10684 2280 10736
rect 940 10412 992 10464
rect 3610 10310 3662 10362
rect 3674 10310 3726 10362
rect 3738 10310 3790 10362
rect 3802 10310 3854 10362
rect 3866 10310 3918 10362
rect 5210 10310 5262 10362
rect 5274 10310 5326 10362
rect 5338 10310 5390 10362
rect 5402 10310 5454 10362
rect 5466 10310 5518 10362
rect 6810 10310 6862 10362
rect 6874 10310 6926 10362
rect 6938 10310 6990 10362
rect 7002 10310 7054 10362
rect 7066 10310 7118 10362
rect 8410 10310 8462 10362
rect 8474 10310 8526 10362
rect 8538 10310 8590 10362
rect 8602 10310 8654 10362
rect 8666 10310 8718 10362
rect 2950 9766 3002 9818
rect 3014 9766 3066 9818
rect 3078 9766 3130 9818
rect 3142 9766 3194 9818
rect 3206 9766 3258 9818
rect 4550 9766 4602 9818
rect 4614 9766 4666 9818
rect 4678 9766 4730 9818
rect 4742 9766 4794 9818
rect 4806 9766 4858 9818
rect 6150 9766 6202 9818
rect 6214 9766 6266 9818
rect 6278 9766 6330 9818
rect 6342 9766 6394 9818
rect 6406 9766 6458 9818
rect 7750 9766 7802 9818
rect 7814 9766 7866 9818
rect 7878 9766 7930 9818
rect 7942 9766 7994 9818
rect 8006 9766 8058 9818
rect 9350 9766 9402 9818
rect 9414 9766 9466 9818
rect 9478 9766 9530 9818
rect 9542 9766 9594 9818
rect 9606 9766 9658 9818
rect 4160 9596 4212 9648
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 7380 9460 7432 9512
rect 940 9324 992 9376
rect 8208 9324 8260 9376
rect 3610 9222 3662 9274
rect 3674 9222 3726 9274
rect 3738 9222 3790 9274
rect 3802 9222 3854 9274
rect 3866 9222 3918 9274
rect 5210 9222 5262 9274
rect 5274 9222 5326 9274
rect 5338 9222 5390 9274
rect 5402 9222 5454 9274
rect 5466 9222 5518 9274
rect 6810 9222 6862 9274
rect 6874 9222 6926 9274
rect 6938 9222 6990 9274
rect 7002 9222 7054 9274
rect 7066 9222 7118 9274
rect 8410 9222 8462 9274
rect 8474 9222 8526 9274
rect 8538 9222 8590 9274
rect 8602 9222 8654 9274
rect 8666 9222 8718 9274
rect 8300 8916 8352 8968
rect 9588 8916 9640 8968
rect 2950 8678 3002 8730
rect 3014 8678 3066 8730
rect 3078 8678 3130 8730
rect 3142 8678 3194 8730
rect 3206 8678 3258 8730
rect 4550 8678 4602 8730
rect 4614 8678 4666 8730
rect 4678 8678 4730 8730
rect 4742 8678 4794 8730
rect 4806 8678 4858 8730
rect 6150 8678 6202 8730
rect 6214 8678 6266 8730
rect 6278 8678 6330 8730
rect 6342 8678 6394 8730
rect 6406 8678 6458 8730
rect 7750 8678 7802 8730
rect 7814 8678 7866 8730
rect 7878 8678 7930 8730
rect 7942 8678 7994 8730
rect 8006 8678 8058 8730
rect 9350 8678 9402 8730
rect 9414 8678 9466 8730
rect 9478 8678 9530 8730
rect 9542 8678 9594 8730
rect 9606 8678 9658 8730
rect 1768 8508 1820 8560
rect 1400 8304 1452 8356
rect 3610 8134 3662 8186
rect 3674 8134 3726 8186
rect 3738 8134 3790 8186
rect 3802 8134 3854 8186
rect 3866 8134 3918 8186
rect 5210 8134 5262 8186
rect 5274 8134 5326 8186
rect 5338 8134 5390 8186
rect 5402 8134 5454 8186
rect 5466 8134 5518 8186
rect 6810 8134 6862 8186
rect 6874 8134 6926 8186
rect 6938 8134 6990 8186
rect 7002 8134 7054 8186
rect 7066 8134 7118 8186
rect 8410 8134 8462 8186
rect 8474 8134 8526 8186
rect 8538 8134 8590 8186
rect 8602 8134 8654 8186
rect 8666 8134 8718 8186
rect 2950 7590 3002 7642
rect 3014 7590 3066 7642
rect 3078 7590 3130 7642
rect 3142 7590 3194 7642
rect 3206 7590 3258 7642
rect 4550 7590 4602 7642
rect 4614 7590 4666 7642
rect 4678 7590 4730 7642
rect 4742 7590 4794 7642
rect 4806 7590 4858 7642
rect 6150 7590 6202 7642
rect 6214 7590 6266 7642
rect 6278 7590 6330 7642
rect 6342 7590 6394 7642
rect 6406 7590 6458 7642
rect 7750 7590 7802 7642
rect 7814 7590 7866 7642
rect 7878 7590 7930 7642
rect 7942 7590 7994 7642
rect 8006 7590 8058 7642
rect 9350 7590 9402 7642
rect 9414 7590 9466 7642
rect 9478 7590 9530 7642
rect 9542 7590 9594 7642
rect 9606 7590 9658 7642
rect 3332 7420 3384 7472
rect 940 7148 992 7200
rect 3610 7046 3662 7098
rect 3674 7046 3726 7098
rect 3738 7046 3790 7098
rect 3802 7046 3854 7098
rect 3866 7046 3918 7098
rect 5210 7046 5262 7098
rect 5274 7046 5326 7098
rect 5338 7046 5390 7098
rect 5402 7046 5454 7098
rect 5466 7046 5518 7098
rect 6810 7046 6862 7098
rect 6874 7046 6926 7098
rect 6938 7046 6990 7098
rect 7002 7046 7054 7098
rect 7066 7046 7118 7098
rect 8410 7046 8462 7098
rect 8474 7046 8526 7098
rect 8538 7046 8590 7098
rect 8602 7046 8654 7098
rect 8666 7046 8718 7098
rect 2136 6740 2188 6792
rect 940 6604 992 6656
rect 2950 6502 3002 6554
rect 3014 6502 3066 6554
rect 3078 6502 3130 6554
rect 3142 6502 3194 6554
rect 3206 6502 3258 6554
rect 4550 6502 4602 6554
rect 4614 6502 4666 6554
rect 4678 6502 4730 6554
rect 4742 6502 4794 6554
rect 4806 6502 4858 6554
rect 6150 6502 6202 6554
rect 6214 6502 6266 6554
rect 6278 6502 6330 6554
rect 6342 6502 6394 6554
rect 6406 6502 6458 6554
rect 7750 6502 7802 6554
rect 7814 6502 7866 6554
rect 7878 6502 7930 6554
rect 7942 6502 7994 6554
rect 8006 6502 8058 6554
rect 9350 6502 9402 6554
rect 9414 6502 9466 6554
rect 9478 6502 9530 6554
rect 9542 6502 9594 6554
rect 9606 6502 9658 6554
rect 3610 5958 3662 6010
rect 3674 5958 3726 6010
rect 3738 5958 3790 6010
rect 3802 5958 3854 6010
rect 3866 5958 3918 6010
rect 5210 5958 5262 6010
rect 5274 5958 5326 6010
rect 5338 5958 5390 6010
rect 5402 5958 5454 6010
rect 5466 5958 5518 6010
rect 6810 5958 6862 6010
rect 6874 5958 6926 6010
rect 6938 5958 6990 6010
rect 7002 5958 7054 6010
rect 7066 5958 7118 6010
rect 8410 5958 8462 6010
rect 8474 5958 8526 6010
rect 8538 5958 8590 6010
rect 8602 5958 8654 6010
rect 8666 5958 8718 6010
rect 3976 5652 4028 5704
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 2950 5414 3002 5466
rect 3014 5414 3066 5466
rect 3078 5414 3130 5466
rect 3142 5414 3194 5466
rect 3206 5414 3258 5466
rect 4550 5414 4602 5466
rect 4614 5414 4666 5466
rect 4678 5414 4730 5466
rect 4742 5414 4794 5466
rect 4806 5414 4858 5466
rect 6150 5414 6202 5466
rect 6214 5414 6266 5466
rect 6278 5414 6330 5466
rect 6342 5414 6394 5466
rect 6406 5414 6458 5466
rect 7750 5414 7802 5466
rect 7814 5414 7866 5466
rect 7878 5414 7930 5466
rect 7942 5414 7994 5466
rect 8006 5414 8058 5466
rect 9350 5414 9402 5466
rect 9414 5414 9466 5466
rect 9478 5414 9530 5466
rect 9542 5414 9594 5466
rect 9606 5414 9658 5466
rect 3610 4870 3662 4922
rect 3674 4870 3726 4922
rect 3738 4870 3790 4922
rect 3802 4870 3854 4922
rect 3866 4870 3918 4922
rect 5210 4870 5262 4922
rect 5274 4870 5326 4922
rect 5338 4870 5390 4922
rect 5402 4870 5454 4922
rect 5466 4870 5518 4922
rect 6810 4870 6862 4922
rect 6874 4870 6926 4922
rect 6938 4870 6990 4922
rect 7002 4870 7054 4922
rect 7066 4870 7118 4922
rect 8410 4870 8462 4922
rect 8474 4870 8526 4922
rect 8538 4870 8590 4922
rect 8602 4870 8654 4922
rect 8666 4870 8718 4922
rect 4252 4564 4304 4616
rect 940 4428 992 4480
rect 2950 4326 3002 4378
rect 3014 4326 3066 4378
rect 3078 4326 3130 4378
rect 3142 4326 3194 4378
rect 3206 4326 3258 4378
rect 4550 4326 4602 4378
rect 4614 4326 4666 4378
rect 4678 4326 4730 4378
rect 4742 4326 4794 4378
rect 4806 4326 4858 4378
rect 6150 4326 6202 4378
rect 6214 4326 6266 4378
rect 6278 4326 6330 4378
rect 6342 4326 6394 4378
rect 6406 4326 6458 4378
rect 7750 4326 7802 4378
rect 7814 4326 7866 4378
rect 7878 4326 7930 4378
rect 7942 4326 7994 4378
rect 8006 4326 8058 4378
rect 9350 4326 9402 4378
rect 9414 4326 9466 4378
rect 9478 4326 9530 4378
rect 9542 4326 9594 4378
rect 9606 4326 9658 4378
rect 11704 3952 11756 4004
rect 17868 3952 17920 4004
rect 9036 3884 9088 3936
rect 54392 3884 54444 3936
rect 3610 3782 3662 3834
rect 3674 3782 3726 3834
rect 3738 3782 3790 3834
rect 3802 3782 3854 3834
rect 3866 3782 3918 3834
rect 5210 3782 5262 3834
rect 5274 3782 5326 3834
rect 5338 3782 5390 3834
rect 5402 3782 5454 3834
rect 5466 3782 5518 3834
rect 6810 3782 6862 3834
rect 6874 3782 6926 3834
rect 6938 3782 6990 3834
rect 7002 3782 7054 3834
rect 7066 3782 7118 3834
rect 8410 3782 8462 3834
rect 8474 3782 8526 3834
rect 8538 3782 8590 3834
rect 8602 3782 8654 3834
rect 8666 3782 8718 3834
rect 11428 3816 11480 3868
rect 46112 3816 46164 3868
rect 10784 3748 10836 3800
rect 40316 3748 40368 3800
rect 9128 3680 9180 3732
rect 50896 3680 50948 3732
rect 7564 3612 7616 3664
rect 45008 3612 45060 3664
rect 5080 3544 5132 3596
rect 39212 3544 39264 3596
rect 2320 3476 2372 3528
rect 10968 3476 11020 3528
rect 29828 3476 29880 3528
rect 6644 3408 6696 3460
rect 54576 3408 54628 3460
rect 940 3340 992 3392
rect 10232 3340 10284 3392
rect 28724 3340 28776 3392
rect 2950 3238 3002 3290
rect 3014 3238 3066 3290
rect 3078 3238 3130 3290
rect 3142 3238 3194 3290
rect 3206 3238 3258 3290
rect 4550 3238 4602 3290
rect 4614 3238 4666 3290
rect 4678 3238 4730 3290
rect 4742 3238 4794 3290
rect 4806 3238 4858 3290
rect 6150 3238 6202 3290
rect 6214 3238 6266 3290
rect 6278 3238 6330 3290
rect 6342 3238 6394 3290
rect 6406 3238 6458 3290
rect 7750 3238 7802 3290
rect 7814 3238 7866 3290
rect 7878 3238 7930 3290
rect 7942 3238 7994 3290
rect 8006 3238 8058 3290
rect 9350 3238 9402 3290
rect 9414 3238 9466 3290
rect 9478 3238 9530 3290
rect 9542 3238 9594 3290
rect 9606 3238 9658 3290
rect 10324 3272 10376 3324
rect 32128 3272 32180 3324
rect 5816 3136 5868 3188
rect 47492 3136 47544 3188
rect 3610 2694 3662 2746
rect 3674 2694 3726 2746
rect 3738 2694 3790 2746
rect 3802 2694 3854 2746
rect 3866 2694 3918 2746
rect 5210 2694 5262 2746
rect 5274 2694 5326 2746
rect 5338 2694 5390 2746
rect 5402 2694 5454 2746
rect 5466 2694 5518 2746
rect 6810 2694 6862 2746
rect 6874 2694 6926 2746
rect 6938 2694 6990 2746
rect 7002 2694 7054 2746
rect 7066 2694 7118 2746
rect 8410 2694 8462 2746
rect 8474 2694 8526 2746
rect 8538 2694 8590 2746
rect 8602 2694 8654 2746
rect 8666 2694 8718 2746
rect 11888 2728 11940 2780
rect 27528 2728 27580 2780
rect 11796 2660 11848 2712
rect 34704 2660 34756 2712
rect 6000 2592 6052 2644
rect 107936 2592 107988 2644
rect 8116 2524 8168 2576
rect 32036 2524 32088 2576
rect 8944 2456 8996 2508
rect 43812 2456 43864 2508
rect 8760 2388 8812 2440
rect 55404 2388 55456 2440
rect 8300 2320 8352 2372
rect 57980 2320 58032 2372
rect 848 2252 900 2304
rect 49700 2252 49752 2304
rect 2950 2150 3002 2202
rect 3014 2150 3066 2202
rect 3078 2150 3130 2202
rect 3142 2150 3194 2202
rect 3206 2150 3258 2202
rect 4550 2150 4602 2202
rect 4614 2150 4666 2202
rect 4678 2150 4730 2202
rect 4742 2150 4794 2202
rect 4806 2150 4858 2202
rect 6150 2150 6202 2202
rect 6214 2150 6266 2202
rect 6278 2150 6330 2202
rect 6342 2150 6394 2202
rect 6406 2150 6458 2202
rect 7750 2150 7802 2202
rect 7814 2150 7866 2202
rect 7878 2150 7930 2202
rect 7942 2150 7994 2202
rect 8006 2150 8058 2202
rect 9350 2150 9402 2202
rect 9414 2150 9466 2202
rect 9478 2150 9530 2202
rect 9542 2150 9594 2202
rect 9606 2150 9658 2202
rect 11612 2184 11664 2236
rect 37004 2184 37056 2236
rect 10876 2116 10928 2168
rect 48596 2116 48648 2168
rect 6552 2048 6604 2100
rect 94964 2048 95016 2100
rect 9220 1980 9272 2032
rect 42800 1980 42852 2032
rect 3610 1606 3662 1658
rect 3674 1606 3726 1658
rect 3738 1606 3790 1658
rect 3802 1606 3854 1658
rect 3866 1606 3918 1658
rect 5210 1606 5262 1658
rect 5274 1606 5326 1658
rect 5338 1606 5390 1658
rect 5402 1606 5454 1658
rect 5466 1606 5518 1658
rect 6810 1606 6862 1658
rect 6874 1606 6926 1658
rect 6938 1606 6990 1658
rect 7002 1606 7054 1658
rect 7066 1606 7118 1658
rect 8410 1606 8462 1658
rect 8474 1606 8526 1658
rect 8538 1606 8590 1658
rect 8602 1606 8654 1658
rect 8666 1606 8718 1658
rect 10010 1606 10062 1658
rect 10074 1606 10126 1658
rect 10138 1606 10190 1658
rect 10202 1606 10254 1658
rect 10266 1606 10318 1658
rect 11610 1606 11662 1658
rect 11674 1606 11726 1658
rect 11738 1606 11790 1658
rect 11802 1606 11854 1658
rect 11866 1606 11918 1658
rect 13210 1606 13262 1658
rect 13274 1606 13326 1658
rect 13338 1606 13390 1658
rect 13402 1606 13454 1658
rect 13466 1606 13518 1658
rect 14810 1606 14862 1658
rect 14874 1606 14926 1658
rect 14938 1606 14990 1658
rect 15002 1606 15054 1658
rect 15066 1606 15118 1658
rect 16410 1606 16462 1658
rect 16474 1606 16526 1658
rect 16538 1606 16590 1658
rect 16602 1606 16654 1658
rect 16666 1606 16718 1658
rect 18010 1606 18062 1658
rect 18074 1606 18126 1658
rect 18138 1606 18190 1658
rect 18202 1606 18254 1658
rect 18266 1606 18318 1658
rect 19610 1606 19662 1658
rect 19674 1606 19726 1658
rect 19738 1606 19790 1658
rect 19802 1606 19854 1658
rect 19866 1606 19918 1658
rect 21210 1606 21262 1658
rect 21274 1606 21326 1658
rect 21338 1606 21390 1658
rect 21402 1606 21454 1658
rect 21466 1606 21518 1658
rect 22810 1606 22862 1658
rect 22874 1606 22926 1658
rect 22938 1606 22990 1658
rect 23002 1606 23054 1658
rect 23066 1606 23118 1658
rect 24410 1606 24462 1658
rect 24474 1606 24526 1658
rect 24538 1606 24590 1658
rect 24602 1606 24654 1658
rect 24666 1606 24718 1658
rect 26010 1606 26062 1658
rect 26074 1606 26126 1658
rect 26138 1606 26190 1658
rect 26202 1606 26254 1658
rect 26266 1606 26318 1658
rect 27610 1606 27662 1658
rect 27674 1606 27726 1658
rect 27738 1606 27790 1658
rect 27802 1606 27854 1658
rect 27866 1606 27918 1658
rect 29210 1606 29262 1658
rect 29274 1606 29326 1658
rect 29338 1606 29390 1658
rect 29402 1606 29454 1658
rect 29466 1606 29518 1658
rect 30810 1606 30862 1658
rect 30874 1606 30926 1658
rect 30938 1606 30990 1658
rect 31002 1606 31054 1658
rect 31066 1606 31118 1658
rect 32410 1606 32462 1658
rect 32474 1606 32526 1658
rect 32538 1606 32590 1658
rect 32602 1606 32654 1658
rect 32666 1606 32718 1658
rect 34010 1606 34062 1658
rect 34074 1606 34126 1658
rect 34138 1606 34190 1658
rect 34202 1606 34254 1658
rect 34266 1606 34318 1658
rect 35610 1606 35662 1658
rect 35674 1606 35726 1658
rect 35738 1606 35790 1658
rect 35802 1606 35854 1658
rect 35866 1606 35918 1658
rect 37210 1606 37262 1658
rect 37274 1606 37326 1658
rect 37338 1606 37390 1658
rect 37402 1606 37454 1658
rect 37466 1606 37518 1658
rect 38810 1606 38862 1658
rect 38874 1606 38926 1658
rect 38938 1606 38990 1658
rect 39002 1606 39054 1658
rect 39066 1606 39118 1658
rect 40410 1606 40462 1658
rect 40474 1606 40526 1658
rect 40538 1606 40590 1658
rect 40602 1606 40654 1658
rect 40666 1606 40718 1658
rect 42010 1606 42062 1658
rect 42074 1606 42126 1658
rect 42138 1606 42190 1658
rect 42202 1606 42254 1658
rect 42266 1606 42318 1658
rect 43610 1606 43662 1658
rect 43674 1606 43726 1658
rect 43738 1606 43790 1658
rect 43802 1606 43854 1658
rect 43866 1606 43918 1658
rect 45210 1606 45262 1658
rect 45274 1606 45326 1658
rect 45338 1606 45390 1658
rect 45402 1606 45454 1658
rect 45466 1606 45518 1658
rect 46810 1606 46862 1658
rect 46874 1606 46926 1658
rect 46938 1606 46990 1658
rect 47002 1606 47054 1658
rect 47066 1606 47118 1658
rect 48410 1606 48462 1658
rect 48474 1606 48526 1658
rect 48538 1606 48590 1658
rect 48602 1606 48654 1658
rect 48666 1606 48718 1658
rect 50010 1606 50062 1658
rect 50074 1606 50126 1658
rect 50138 1606 50190 1658
rect 50202 1606 50254 1658
rect 50266 1606 50318 1658
rect 51610 1606 51662 1658
rect 51674 1606 51726 1658
rect 51738 1606 51790 1658
rect 51802 1606 51854 1658
rect 51866 1606 51918 1658
rect 53210 1606 53262 1658
rect 53274 1606 53326 1658
rect 53338 1606 53390 1658
rect 53402 1606 53454 1658
rect 53466 1606 53518 1658
rect 54810 1606 54862 1658
rect 54874 1606 54926 1658
rect 54938 1606 54990 1658
rect 55002 1606 55054 1658
rect 55066 1606 55118 1658
rect 56410 1606 56462 1658
rect 56474 1606 56526 1658
rect 56538 1606 56590 1658
rect 56602 1606 56654 1658
rect 56666 1606 56718 1658
rect 58010 1606 58062 1658
rect 58074 1606 58126 1658
rect 58138 1606 58190 1658
rect 58202 1606 58254 1658
rect 58266 1606 58318 1658
rect 59610 1606 59662 1658
rect 59674 1606 59726 1658
rect 59738 1606 59790 1658
rect 59802 1606 59854 1658
rect 59866 1606 59918 1658
rect 61210 1606 61262 1658
rect 61274 1606 61326 1658
rect 61338 1606 61390 1658
rect 61402 1606 61454 1658
rect 61466 1606 61518 1658
rect 62810 1606 62862 1658
rect 62874 1606 62926 1658
rect 62938 1606 62990 1658
rect 63002 1606 63054 1658
rect 63066 1606 63118 1658
rect 64410 1606 64462 1658
rect 64474 1606 64526 1658
rect 64538 1606 64590 1658
rect 64602 1606 64654 1658
rect 64666 1606 64718 1658
rect 66010 1606 66062 1658
rect 66074 1606 66126 1658
rect 66138 1606 66190 1658
rect 66202 1606 66254 1658
rect 66266 1606 66318 1658
rect 67610 1606 67662 1658
rect 67674 1606 67726 1658
rect 67738 1606 67790 1658
rect 67802 1606 67854 1658
rect 67866 1606 67918 1658
rect 69210 1606 69262 1658
rect 69274 1606 69326 1658
rect 69338 1606 69390 1658
rect 69402 1606 69454 1658
rect 69466 1606 69518 1658
rect 70810 1606 70862 1658
rect 70874 1606 70926 1658
rect 70938 1606 70990 1658
rect 71002 1606 71054 1658
rect 71066 1606 71118 1658
rect 72410 1606 72462 1658
rect 72474 1606 72526 1658
rect 72538 1606 72590 1658
rect 72602 1606 72654 1658
rect 72666 1606 72718 1658
rect 74010 1606 74062 1658
rect 74074 1606 74126 1658
rect 74138 1606 74190 1658
rect 74202 1606 74254 1658
rect 74266 1606 74318 1658
rect 75610 1606 75662 1658
rect 75674 1606 75726 1658
rect 75738 1606 75790 1658
rect 75802 1606 75854 1658
rect 75866 1606 75918 1658
rect 77210 1606 77262 1658
rect 77274 1606 77326 1658
rect 77338 1606 77390 1658
rect 77402 1606 77454 1658
rect 77466 1606 77518 1658
rect 78810 1606 78862 1658
rect 78874 1606 78926 1658
rect 78938 1606 78990 1658
rect 79002 1606 79054 1658
rect 79066 1606 79118 1658
rect 80410 1606 80462 1658
rect 80474 1606 80526 1658
rect 80538 1606 80590 1658
rect 80602 1606 80654 1658
rect 80666 1606 80718 1658
rect 82010 1606 82062 1658
rect 82074 1606 82126 1658
rect 82138 1606 82190 1658
rect 82202 1606 82254 1658
rect 82266 1606 82318 1658
rect 83610 1606 83662 1658
rect 83674 1606 83726 1658
rect 83738 1606 83790 1658
rect 83802 1606 83854 1658
rect 83866 1606 83918 1658
rect 85210 1606 85262 1658
rect 85274 1606 85326 1658
rect 85338 1606 85390 1658
rect 85402 1606 85454 1658
rect 85466 1606 85518 1658
rect 86810 1606 86862 1658
rect 86874 1606 86926 1658
rect 86938 1606 86990 1658
rect 87002 1606 87054 1658
rect 87066 1606 87118 1658
rect 88410 1606 88462 1658
rect 88474 1606 88526 1658
rect 88538 1606 88590 1658
rect 88602 1606 88654 1658
rect 88666 1606 88718 1658
rect 90010 1606 90062 1658
rect 90074 1606 90126 1658
rect 90138 1606 90190 1658
rect 90202 1606 90254 1658
rect 90266 1606 90318 1658
rect 91610 1606 91662 1658
rect 91674 1606 91726 1658
rect 91738 1606 91790 1658
rect 91802 1606 91854 1658
rect 91866 1606 91918 1658
rect 93210 1606 93262 1658
rect 93274 1606 93326 1658
rect 93338 1606 93390 1658
rect 93402 1606 93454 1658
rect 93466 1606 93518 1658
rect 94810 1606 94862 1658
rect 94874 1606 94926 1658
rect 94938 1606 94990 1658
rect 95002 1606 95054 1658
rect 95066 1606 95118 1658
rect 96410 1606 96462 1658
rect 96474 1606 96526 1658
rect 96538 1606 96590 1658
rect 96602 1606 96654 1658
rect 96666 1606 96718 1658
rect 98010 1606 98062 1658
rect 98074 1606 98126 1658
rect 98138 1606 98190 1658
rect 98202 1606 98254 1658
rect 98266 1606 98318 1658
rect 99610 1606 99662 1658
rect 99674 1606 99726 1658
rect 99738 1606 99790 1658
rect 99802 1606 99854 1658
rect 99866 1606 99918 1658
rect 101210 1606 101262 1658
rect 101274 1606 101326 1658
rect 101338 1606 101390 1658
rect 101402 1606 101454 1658
rect 101466 1606 101518 1658
rect 102810 1606 102862 1658
rect 102874 1606 102926 1658
rect 102938 1606 102990 1658
rect 103002 1606 103054 1658
rect 103066 1606 103118 1658
rect 104410 1606 104462 1658
rect 104474 1606 104526 1658
rect 104538 1606 104590 1658
rect 104602 1606 104654 1658
rect 104666 1606 104718 1658
rect 106010 1606 106062 1658
rect 106074 1606 106126 1658
rect 106138 1606 106190 1658
rect 106202 1606 106254 1658
rect 106266 1606 106318 1658
rect 107610 1606 107662 1658
rect 107674 1606 107726 1658
rect 107738 1606 107790 1658
rect 107802 1606 107854 1658
rect 107866 1606 107918 1658
rect 23664 1436 23716 1488
rect 11520 1300 11572 1352
rect 1032 1232 1084 1284
rect 23204 1368 23256 1420
rect 24124 1300 24176 1352
rect 1124 1164 1176 1216
rect 17224 1164 17276 1216
rect 22928 1207 22980 1216
rect 22928 1173 22937 1207
rect 22937 1173 22971 1207
rect 22971 1173 22980 1207
rect 22928 1164 22980 1173
rect 23480 1232 23532 1284
rect 27528 1411 27580 1420
rect 27528 1377 27537 1411
rect 27537 1377 27571 1411
rect 27571 1377 27580 1411
rect 27528 1368 27580 1377
rect 27804 1343 27856 1352
rect 27804 1309 27813 1343
rect 27813 1309 27847 1343
rect 27847 1309 27856 1343
rect 27804 1300 27856 1309
rect 34704 1411 34756 1420
rect 34704 1377 34713 1411
rect 34713 1377 34747 1411
rect 34747 1377 34756 1411
rect 34704 1368 34756 1377
rect 29644 1343 29696 1352
rect 29644 1309 29653 1343
rect 29653 1309 29687 1343
rect 29687 1309 29696 1343
rect 29644 1300 29696 1309
rect 26240 1164 26292 1216
rect 26332 1207 26384 1216
rect 26332 1173 26341 1207
rect 26341 1173 26375 1207
rect 26375 1173 26384 1207
rect 26332 1164 26384 1173
rect 27344 1232 27396 1284
rect 32128 1343 32180 1352
rect 32128 1309 32137 1343
rect 32137 1309 32171 1343
rect 32171 1309 32180 1343
rect 32128 1300 32180 1309
rect 32404 1343 32456 1352
rect 32404 1309 32413 1343
rect 32413 1309 32447 1343
rect 32447 1309 32456 1343
rect 32404 1300 32456 1309
rect 33140 1300 33192 1352
rect 33876 1343 33928 1352
rect 33876 1309 33885 1343
rect 33885 1309 33919 1343
rect 33919 1309 33928 1343
rect 33876 1300 33928 1309
rect 37372 1300 37424 1352
rect 37556 1300 37608 1352
rect 37740 1343 37792 1352
rect 37740 1309 37749 1343
rect 37749 1309 37783 1343
rect 37783 1309 37792 1343
rect 37740 1300 37792 1309
rect 29460 1164 29512 1216
rect 29736 1207 29788 1216
rect 29736 1173 29745 1207
rect 29745 1173 29779 1207
rect 29779 1173 29788 1207
rect 29736 1164 29788 1173
rect 29828 1164 29880 1216
rect 59360 1232 59412 1284
rect 30656 1207 30708 1216
rect 30656 1173 30665 1207
rect 30665 1173 30699 1207
rect 30699 1173 30708 1207
rect 30656 1164 30708 1173
rect 32312 1164 32364 1216
rect 37280 1164 37332 1216
rect 37556 1164 37608 1216
rect 2950 1062 3002 1114
rect 3014 1062 3066 1114
rect 3078 1062 3130 1114
rect 3142 1062 3194 1114
rect 3206 1062 3258 1114
rect 4550 1062 4602 1114
rect 4614 1062 4666 1114
rect 4678 1062 4730 1114
rect 4742 1062 4794 1114
rect 4806 1062 4858 1114
rect 6150 1062 6202 1114
rect 6214 1062 6266 1114
rect 6278 1062 6330 1114
rect 6342 1062 6394 1114
rect 6406 1062 6458 1114
rect 7750 1062 7802 1114
rect 7814 1062 7866 1114
rect 7878 1062 7930 1114
rect 7942 1062 7994 1114
rect 8006 1062 8058 1114
rect 9350 1062 9402 1114
rect 9414 1062 9466 1114
rect 9478 1062 9530 1114
rect 9542 1062 9594 1114
rect 9606 1062 9658 1114
rect 10950 1062 11002 1114
rect 11014 1062 11066 1114
rect 11078 1062 11130 1114
rect 11142 1062 11194 1114
rect 11206 1062 11258 1114
rect 12550 1062 12602 1114
rect 12614 1062 12666 1114
rect 12678 1062 12730 1114
rect 12742 1062 12794 1114
rect 12806 1062 12858 1114
rect 14150 1062 14202 1114
rect 14214 1062 14266 1114
rect 14278 1062 14330 1114
rect 14342 1062 14394 1114
rect 14406 1062 14458 1114
rect 15750 1062 15802 1114
rect 15814 1062 15866 1114
rect 15878 1062 15930 1114
rect 15942 1062 15994 1114
rect 16006 1062 16058 1114
rect 17350 1062 17402 1114
rect 17414 1062 17466 1114
rect 17478 1062 17530 1114
rect 17542 1062 17594 1114
rect 17606 1062 17658 1114
rect 18950 1062 19002 1114
rect 19014 1062 19066 1114
rect 19078 1062 19130 1114
rect 19142 1062 19194 1114
rect 19206 1062 19258 1114
rect 20550 1062 20602 1114
rect 20614 1062 20666 1114
rect 20678 1062 20730 1114
rect 20742 1062 20794 1114
rect 20806 1062 20858 1114
rect 22150 1062 22202 1114
rect 22214 1062 22266 1114
rect 22278 1062 22330 1114
rect 22342 1062 22394 1114
rect 22406 1062 22458 1114
rect 23750 1062 23802 1114
rect 23814 1062 23866 1114
rect 23878 1062 23930 1114
rect 23942 1062 23994 1114
rect 24006 1062 24058 1114
rect 25350 1062 25402 1114
rect 25414 1062 25466 1114
rect 25478 1062 25530 1114
rect 25542 1062 25594 1114
rect 25606 1062 25658 1114
rect 26950 1062 27002 1114
rect 27014 1062 27066 1114
rect 27078 1062 27130 1114
rect 27142 1062 27194 1114
rect 27206 1062 27258 1114
rect 28550 1062 28602 1114
rect 28614 1062 28666 1114
rect 28678 1062 28730 1114
rect 28742 1062 28794 1114
rect 28806 1062 28858 1114
rect 30150 1062 30202 1114
rect 30214 1062 30266 1114
rect 30278 1062 30330 1114
rect 30342 1062 30394 1114
rect 30406 1062 30458 1114
rect 31750 1062 31802 1114
rect 31814 1062 31866 1114
rect 31878 1062 31930 1114
rect 31942 1062 31994 1114
rect 32006 1062 32058 1114
rect 33350 1062 33402 1114
rect 33414 1062 33466 1114
rect 33478 1062 33530 1114
rect 33542 1062 33594 1114
rect 33606 1062 33658 1114
rect 34950 1062 35002 1114
rect 35014 1062 35066 1114
rect 35078 1062 35130 1114
rect 35142 1062 35194 1114
rect 35206 1062 35258 1114
rect 36550 1062 36602 1114
rect 36614 1062 36666 1114
rect 36678 1062 36730 1114
rect 36742 1062 36794 1114
rect 36806 1062 36858 1114
rect 38150 1062 38202 1114
rect 38214 1062 38266 1114
rect 38278 1062 38330 1114
rect 38342 1062 38394 1114
rect 38406 1062 38458 1114
rect 39750 1062 39802 1114
rect 39814 1062 39866 1114
rect 39878 1062 39930 1114
rect 39942 1062 39994 1114
rect 40006 1062 40058 1114
rect 41350 1062 41402 1114
rect 41414 1062 41466 1114
rect 41478 1062 41530 1114
rect 41542 1062 41594 1114
rect 41606 1062 41658 1114
rect 42950 1062 43002 1114
rect 43014 1062 43066 1114
rect 43078 1062 43130 1114
rect 43142 1062 43194 1114
rect 43206 1062 43258 1114
rect 44550 1062 44602 1114
rect 44614 1062 44666 1114
rect 44678 1062 44730 1114
rect 44742 1062 44794 1114
rect 44806 1062 44858 1114
rect 46150 1062 46202 1114
rect 46214 1062 46266 1114
rect 46278 1062 46330 1114
rect 46342 1062 46394 1114
rect 46406 1062 46458 1114
rect 47750 1062 47802 1114
rect 47814 1062 47866 1114
rect 47878 1062 47930 1114
rect 47942 1062 47994 1114
rect 48006 1062 48058 1114
rect 49350 1062 49402 1114
rect 49414 1062 49466 1114
rect 49478 1062 49530 1114
rect 49542 1062 49594 1114
rect 49606 1062 49658 1114
rect 50950 1062 51002 1114
rect 51014 1062 51066 1114
rect 51078 1062 51130 1114
rect 51142 1062 51194 1114
rect 51206 1062 51258 1114
rect 52550 1062 52602 1114
rect 52614 1062 52666 1114
rect 52678 1062 52730 1114
rect 52742 1062 52794 1114
rect 52806 1062 52858 1114
rect 54150 1062 54202 1114
rect 54214 1062 54266 1114
rect 54278 1062 54330 1114
rect 54342 1062 54394 1114
rect 54406 1062 54458 1114
rect 55750 1062 55802 1114
rect 55814 1062 55866 1114
rect 55878 1062 55930 1114
rect 55942 1062 55994 1114
rect 56006 1062 56058 1114
rect 57350 1062 57402 1114
rect 57414 1062 57466 1114
rect 57478 1062 57530 1114
rect 57542 1062 57594 1114
rect 57606 1062 57658 1114
rect 58950 1062 59002 1114
rect 59014 1062 59066 1114
rect 59078 1062 59130 1114
rect 59142 1062 59194 1114
rect 59206 1062 59258 1114
rect 60550 1062 60602 1114
rect 60614 1062 60666 1114
rect 60678 1062 60730 1114
rect 60742 1062 60794 1114
rect 60806 1062 60858 1114
rect 62150 1062 62202 1114
rect 62214 1062 62266 1114
rect 62278 1062 62330 1114
rect 62342 1062 62394 1114
rect 62406 1062 62458 1114
rect 63750 1062 63802 1114
rect 63814 1062 63866 1114
rect 63878 1062 63930 1114
rect 63942 1062 63994 1114
rect 64006 1062 64058 1114
rect 65350 1062 65402 1114
rect 65414 1062 65466 1114
rect 65478 1062 65530 1114
rect 65542 1062 65594 1114
rect 65606 1062 65658 1114
rect 66950 1062 67002 1114
rect 67014 1062 67066 1114
rect 67078 1062 67130 1114
rect 67142 1062 67194 1114
rect 67206 1062 67258 1114
rect 68550 1062 68602 1114
rect 68614 1062 68666 1114
rect 68678 1062 68730 1114
rect 68742 1062 68794 1114
rect 68806 1062 68858 1114
rect 70150 1062 70202 1114
rect 70214 1062 70266 1114
rect 70278 1062 70330 1114
rect 70342 1062 70394 1114
rect 70406 1062 70458 1114
rect 71750 1062 71802 1114
rect 71814 1062 71866 1114
rect 71878 1062 71930 1114
rect 71942 1062 71994 1114
rect 72006 1062 72058 1114
rect 73350 1062 73402 1114
rect 73414 1062 73466 1114
rect 73478 1062 73530 1114
rect 73542 1062 73594 1114
rect 73606 1062 73658 1114
rect 74950 1062 75002 1114
rect 75014 1062 75066 1114
rect 75078 1062 75130 1114
rect 75142 1062 75194 1114
rect 75206 1062 75258 1114
rect 76550 1062 76602 1114
rect 76614 1062 76666 1114
rect 76678 1062 76730 1114
rect 76742 1062 76794 1114
rect 76806 1062 76858 1114
rect 78150 1062 78202 1114
rect 78214 1062 78266 1114
rect 78278 1062 78330 1114
rect 78342 1062 78394 1114
rect 78406 1062 78458 1114
rect 79750 1062 79802 1114
rect 79814 1062 79866 1114
rect 79878 1062 79930 1114
rect 79942 1062 79994 1114
rect 80006 1062 80058 1114
rect 81350 1062 81402 1114
rect 81414 1062 81466 1114
rect 81478 1062 81530 1114
rect 81542 1062 81594 1114
rect 81606 1062 81658 1114
rect 82950 1062 83002 1114
rect 83014 1062 83066 1114
rect 83078 1062 83130 1114
rect 83142 1062 83194 1114
rect 83206 1062 83258 1114
rect 84550 1062 84602 1114
rect 84614 1062 84666 1114
rect 84678 1062 84730 1114
rect 84742 1062 84794 1114
rect 84806 1062 84858 1114
rect 86150 1062 86202 1114
rect 86214 1062 86266 1114
rect 86278 1062 86330 1114
rect 86342 1062 86394 1114
rect 86406 1062 86458 1114
rect 87750 1062 87802 1114
rect 87814 1062 87866 1114
rect 87878 1062 87930 1114
rect 87942 1062 87994 1114
rect 88006 1062 88058 1114
rect 89350 1062 89402 1114
rect 89414 1062 89466 1114
rect 89478 1062 89530 1114
rect 89542 1062 89594 1114
rect 89606 1062 89658 1114
rect 90950 1062 91002 1114
rect 91014 1062 91066 1114
rect 91078 1062 91130 1114
rect 91142 1062 91194 1114
rect 91206 1062 91258 1114
rect 92550 1062 92602 1114
rect 92614 1062 92666 1114
rect 92678 1062 92730 1114
rect 92742 1062 92794 1114
rect 92806 1062 92858 1114
rect 94150 1062 94202 1114
rect 94214 1062 94266 1114
rect 94278 1062 94330 1114
rect 94342 1062 94394 1114
rect 94406 1062 94458 1114
rect 95750 1062 95802 1114
rect 95814 1062 95866 1114
rect 95878 1062 95930 1114
rect 95942 1062 95994 1114
rect 96006 1062 96058 1114
rect 97350 1062 97402 1114
rect 97414 1062 97466 1114
rect 97478 1062 97530 1114
rect 97542 1062 97594 1114
rect 97606 1062 97658 1114
rect 98950 1062 99002 1114
rect 99014 1062 99066 1114
rect 99078 1062 99130 1114
rect 99142 1062 99194 1114
rect 99206 1062 99258 1114
rect 100550 1062 100602 1114
rect 100614 1062 100666 1114
rect 100678 1062 100730 1114
rect 100742 1062 100794 1114
rect 100806 1062 100858 1114
rect 102150 1062 102202 1114
rect 102214 1062 102266 1114
rect 102278 1062 102330 1114
rect 102342 1062 102394 1114
rect 102406 1062 102458 1114
rect 103750 1062 103802 1114
rect 103814 1062 103866 1114
rect 103878 1062 103930 1114
rect 103942 1062 103994 1114
rect 104006 1062 104058 1114
rect 105350 1062 105402 1114
rect 105414 1062 105466 1114
rect 105478 1062 105530 1114
rect 105542 1062 105594 1114
rect 105606 1062 105658 1114
rect 106950 1062 107002 1114
rect 107014 1062 107066 1114
rect 107078 1062 107130 1114
rect 107142 1062 107194 1114
rect 107206 1062 107258 1114
rect 108550 1062 108602 1114
rect 108614 1062 108666 1114
rect 108678 1062 108730 1114
rect 108742 1062 108794 1114
rect 108806 1062 108858 1114
rect 5632 960 5684 1012
rect 17224 960 17276 1012
rect 24124 892 24176 944
rect 8208 756 8260 808
rect 24400 756 24452 808
rect 26240 960 26292 1012
rect 29736 960 29788 1012
rect 65156 960 65208 1012
rect 33876 892 33928 944
rect 67640 892 67692 944
rect 56600 824 56652 876
rect 29552 756 29604 808
rect 30656 756 30708 808
rect 64880 756 64932 808
rect 11980 688 12032 740
rect 23480 688 23532 740
rect 10416 620 10468 672
rect 29460 688 29512 740
rect 32220 688 32272 740
rect 32312 688 32364 740
rect 8852 552 8904 604
rect 7656 484 7708 536
rect 23664 484 23716 536
rect 10508 416 10560 468
rect 23204 416 23256 468
rect 9864 280 9916 332
rect 27344 552 27396 604
rect 27804 552 27856 604
rect 60924 688 60976 740
rect 37740 620 37792 672
rect 69020 620 69072 672
rect 37372 552 37424 604
rect 66260 552 66312 604
rect 32404 484 32456 536
rect 62488 484 62540 536
rect 63500 348 63552 400
rect 33232 280 33284 332
rect 34520 280 34572 332
rect 24400 212 24452 264
rect 30564 212 30616 264
rect 22928 76 22980 128
rect 57980 212 58032 264
<< metal2 >>
rect 36544 87644 36596 87650
rect 36544 87586 36596 87592
rect 47308 87644 47360 87650
rect 47308 87586 47360 87592
rect 27528 87576 27580 87582
rect 27528 87518 27580 87524
rect 3424 87372 3476 87378
rect 3424 87314 3476 87320
rect 1308 87236 1360 87242
rect 1308 87178 1360 87184
rect 1032 85536 1084 85542
rect 1032 85478 1084 85484
rect 940 84652 992 84658
rect 940 84594 992 84600
rect 952 84425 980 84594
rect 938 84416 994 84425
rect 938 84351 994 84360
rect 940 83564 992 83570
rect 940 83506 992 83512
rect 952 83473 980 83506
rect 938 83464 994 83473
rect 938 83399 994 83408
rect 940 81796 992 81802
rect 940 81738 992 81744
rect 952 81569 980 81738
rect 938 81560 994 81569
rect 938 81495 994 81504
rect 940 80708 992 80714
rect 940 80650 992 80656
rect 952 80617 980 80650
rect 938 80608 994 80617
rect 938 80543 994 80552
rect 938 79656 994 79665
rect 938 79591 940 79600
rect 992 79591 994 79600
rect 940 79562 992 79568
rect 940 79212 992 79218
rect 940 79154 992 79160
rect 952 78713 980 79154
rect 938 78704 994 78713
rect 938 78639 994 78648
rect 940 78124 992 78130
rect 940 78066 992 78072
rect 952 77761 980 78066
rect 938 77752 994 77761
rect 938 77687 994 77696
rect 940 77036 992 77042
rect 940 76978 992 76984
rect 952 76809 980 76978
rect 938 76800 994 76809
rect 938 76735 994 76744
rect 940 75268 992 75274
rect 940 75210 992 75216
rect 952 74905 980 75210
rect 938 74896 994 74905
rect 938 74831 994 74840
rect 940 74248 992 74254
rect 940 74190 992 74196
rect 952 73953 980 74190
rect 938 73944 994 73953
rect 938 73879 994 73888
rect 940 73092 992 73098
rect 940 73034 992 73040
rect 952 73001 980 73034
rect 938 72992 994 73001
rect 938 72927 994 72936
rect 938 72040 994 72049
rect 938 71975 940 71984
rect 992 71975 994 71984
rect 940 71946 992 71952
rect 664 71664 716 71670
rect 492 71624 664 71652
rect 296 68128 348 68134
rect 296 68070 348 68076
rect 308 67674 336 68070
rect 308 67646 428 67674
rect 296 65408 348 65414
rect 296 65350 348 65356
rect 308 59022 336 65350
rect 400 60734 428 67646
rect 492 60858 520 71624
rect 664 71606 716 71612
rect 940 71596 992 71602
rect 940 71538 992 71544
rect 572 71392 624 71398
rect 572 71334 624 71340
rect 480 60852 532 60858
rect 480 60794 532 60800
rect 400 60706 520 60734
rect 296 59016 348 59022
rect 296 58958 348 58964
rect 492 37126 520 60706
rect 584 40526 612 71334
rect 952 71097 980 71538
rect 938 71088 994 71097
rect 938 71023 994 71032
rect 664 70644 716 70650
rect 664 70586 716 70592
rect 572 40520 624 40526
rect 572 40462 624 40468
rect 676 39438 704 70586
rect 940 69420 992 69426
rect 940 69362 992 69368
rect 952 69193 980 69362
rect 938 69184 994 69193
rect 938 69119 994 69128
rect 940 68332 992 68338
rect 940 68274 992 68280
rect 952 68241 980 68274
rect 938 68232 994 68241
rect 848 68196 900 68202
rect 938 68167 994 68176
rect 848 68138 900 68144
rect 756 67788 808 67794
rect 756 67730 808 67736
rect 768 53106 796 67730
rect 860 67634 888 68138
rect 860 67606 980 67634
rect 952 66722 980 67606
rect 1044 66842 1072 85478
rect 1216 79008 1268 79014
rect 1216 78950 1268 78956
rect 1124 76288 1176 76294
rect 1124 76230 1176 76236
rect 1136 71670 1164 76230
rect 1124 71664 1176 71670
rect 1124 71606 1176 71612
rect 1124 71528 1176 71534
rect 1124 71470 1176 71476
rect 1032 66836 1084 66842
rect 1032 66778 1084 66784
rect 860 66694 980 66722
rect 860 63050 888 66694
rect 940 66564 992 66570
rect 940 66506 992 66512
rect 952 66337 980 66506
rect 938 66328 994 66337
rect 938 66263 994 66272
rect 940 65476 992 65482
rect 940 65418 992 65424
rect 952 65385 980 65418
rect 938 65376 994 65385
rect 938 65311 994 65320
rect 1136 65226 1164 71470
rect 1228 65414 1256 78950
rect 1320 71534 1348 87178
rect 2950 85980 3258 85989
rect 2950 85978 2956 85980
rect 3012 85978 3036 85980
rect 3092 85978 3116 85980
rect 3172 85978 3196 85980
rect 3252 85978 3258 85980
rect 3012 85926 3014 85978
rect 3194 85926 3196 85978
rect 2950 85924 2956 85926
rect 3012 85924 3036 85926
rect 3092 85924 3116 85926
rect 3172 85924 3196 85926
rect 3252 85924 3258 85926
rect 2950 85915 3258 85924
rect 2950 84892 3258 84901
rect 2950 84890 2956 84892
rect 3012 84890 3036 84892
rect 3092 84890 3116 84892
rect 3172 84890 3196 84892
rect 3252 84890 3258 84892
rect 3012 84838 3014 84890
rect 3194 84838 3196 84890
rect 2950 84836 2956 84838
rect 3012 84836 3036 84838
rect 3092 84836 3116 84838
rect 3172 84836 3196 84838
rect 3252 84836 3258 84838
rect 2950 84827 3258 84836
rect 1676 84516 1728 84522
rect 1676 84458 1728 84464
rect 1492 82884 1544 82890
rect 1492 82826 1544 82832
rect 1504 82793 1532 82826
rect 1490 82784 1546 82793
rect 1490 82719 1546 82728
rect 1492 75948 1544 75954
rect 1492 75890 1544 75896
rect 1504 75857 1532 75890
rect 1490 75848 1546 75857
rect 1490 75783 1546 75792
rect 1584 73024 1636 73030
rect 1504 72984 1584 73012
rect 1308 71528 1360 71534
rect 1308 71470 1360 71476
rect 1400 70508 1452 70514
rect 1400 70450 1452 70456
rect 1412 70417 1440 70450
rect 1398 70408 1454 70417
rect 1398 70343 1454 70352
rect 1308 70304 1360 70310
rect 1308 70246 1360 70252
rect 1216 65408 1268 65414
rect 1216 65350 1268 65356
rect 1136 65198 1256 65226
rect 1122 65104 1178 65113
rect 1044 65062 1122 65090
rect 938 64424 994 64433
rect 938 64359 940 64368
rect 992 64359 994 64368
rect 940 64330 992 64336
rect 1044 63186 1072 65062
rect 1122 65039 1178 65048
rect 1228 63442 1256 65198
rect 1216 63436 1268 63442
rect 1216 63378 1268 63384
rect 1044 63158 1256 63186
rect 860 63022 1164 63050
rect 1032 62960 1084 62966
rect 1032 62902 1084 62908
rect 940 62892 992 62898
rect 940 62834 992 62840
rect 952 62529 980 62834
rect 938 62520 994 62529
rect 938 62455 994 62464
rect 940 61804 992 61810
rect 940 61746 992 61752
rect 952 61577 980 61746
rect 938 61568 994 61577
rect 938 61503 994 61512
rect 940 60716 992 60722
rect 940 60658 992 60664
rect 952 60625 980 60658
rect 938 60616 994 60625
rect 938 60551 994 60560
rect 940 59968 992 59974
rect 940 59910 992 59916
rect 952 59673 980 59910
rect 938 59664 994 59673
rect 938 59599 994 59608
rect 940 58880 992 58886
rect 940 58822 992 58828
rect 952 58721 980 58822
rect 938 58712 994 58721
rect 938 58647 994 58656
rect 938 56808 994 56817
rect 938 56743 994 56752
rect 952 56710 980 56743
rect 940 56704 992 56710
rect 940 56646 992 56652
rect 940 56160 992 56166
rect 940 56102 992 56108
rect 952 55865 980 56102
rect 938 55856 994 55865
rect 938 55791 994 55800
rect 940 55072 992 55078
rect 940 55014 992 55020
rect 952 54913 980 55014
rect 938 54904 994 54913
rect 938 54839 994 54848
rect 940 53984 992 53990
rect 938 53952 940 53961
rect 992 53952 994 53961
rect 938 53887 994 53896
rect 756 53100 808 53106
rect 756 53042 808 53048
rect 938 53000 994 53009
rect 938 52935 994 52944
rect 952 52902 980 52935
rect 940 52896 992 52902
rect 940 52838 992 52844
rect 940 51264 992 51270
rect 940 51206 992 51212
rect 952 51105 980 51206
rect 938 51096 994 51105
rect 1044 51074 1072 62902
rect 1136 53038 1164 63022
rect 1228 59702 1256 63158
rect 1216 59696 1268 59702
rect 1216 59638 1268 59644
rect 1320 59514 1348 70246
rect 1504 67810 1532 72984
rect 1584 72966 1636 72972
rect 1584 71936 1636 71942
rect 1582 71904 1584 71913
rect 1636 71904 1638 71913
rect 1582 71839 1638 71848
rect 1584 69420 1636 69426
rect 1584 69362 1636 69368
rect 1228 59486 1348 59514
rect 1412 67782 1532 67810
rect 1228 55962 1256 59486
rect 1412 57974 1440 67782
rect 1492 67652 1544 67658
rect 1492 67594 1544 67600
rect 1504 67561 1532 67594
rect 1490 67552 1546 67561
rect 1490 67487 1546 67496
rect 1596 65113 1624 69362
rect 1582 65104 1638 65113
rect 1582 65039 1638 65048
rect 1584 64320 1636 64326
rect 1584 64262 1636 64268
rect 1596 64122 1624 64262
rect 1584 64116 1636 64122
rect 1584 64058 1636 64064
rect 1492 63980 1544 63986
rect 1492 63922 1544 63928
rect 1504 63481 1532 63922
rect 1584 63776 1636 63782
rect 1584 63718 1636 63724
rect 1596 63578 1624 63718
rect 1584 63572 1636 63578
rect 1584 63514 1636 63520
rect 1490 63472 1546 63481
rect 1490 63407 1546 63416
rect 1584 62144 1636 62150
rect 1584 62086 1636 62092
rect 1492 60036 1544 60042
rect 1492 59978 1544 59984
rect 1504 59770 1532 59978
rect 1492 59764 1544 59770
rect 1492 59706 1544 59712
rect 1320 57946 1440 57974
rect 1216 55956 1268 55962
rect 1216 55898 1268 55904
rect 1124 53032 1176 53038
rect 1124 52974 1176 52980
rect 1044 51046 1164 51074
rect 938 51031 994 51040
rect 940 50176 992 50182
rect 938 50144 940 50153
rect 992 50144 994 50153
rect 938 50079 994 50088
rect 1032 49836 1084 49842
rect 1032 49778 1084 49784
rect 938 49192 994 49201
rect 938 49127 994 49136
rect 952 49094 980 49127
rect 940 49088 992 49094
rect 940 49030 992 49036
rect 940 47456 992 47462
rect 940 47398 992 47404
rect 952 47297 980 47398
rect 938 47288 994 47297
rect 938 47223 994 47232
rect 940 46368 992 46374
rect 938 46336 940 46345
rect 992 46336 994 46345
rect 938 46271 994 46280
rect 938 45384 994 45393
rect 938 45319 994 45328
rect 952 45286 980 45319
rect 940 45280 992 45286
rect 940 45222 992 45228
rect 940 44872 992 44878
rect 940 44814 992 44820
rect 952 44441 980 44814
rect 938 44432 994 44441
rect 938 44367 994 44376
rect 940 43784 992 43790
rect 940 43726 992 43732
rect 952 43489 980 43726
rect 938 43480 994 43489
rect 938 43415 994 43424
rect 940 42628 992 42634
rect 940 42570 992 42576
rect 952 42537 980 42570
rect 938 42528 994 42537
rect 938 42463 994 42472
rect 938 41576 994 41585
rect 938 41511 940 41520
rect 992 41511 994 41520
rect 940 41482 992 41488
rect 1044 41414 1072 49778
rect 952 41386 1072 41414
rect 664 39432 716 39438
rect 664 39374 716 39380
rect 480 37120 532 37126
rect 480 37062 532 37068
rect 848 36576 900 36582
rect 848 36518 900 36524
rect 860 35290 888 36518
rect 848 35284 900 35290
rect 848 35226 900 35232
rect 952 35170 980 41386
rect 1032 41132 1084 41138
rect 1032 41074 1084 41080
rect 1044 40633 1072 41074
rect 1030 40624 1086 40633
rect 1030 40559 1086 40568
rect 1032 38956 1084 38962
rect 1032 38898 1084 38904
rect 1044 38729 1072 38898
rect 1030 38720 1086 38729
rect 1030 38655 1086 38664
rect 1032 37868 1084 37874
rect 1032 37810 1084 37816
rect 1044 37777 1072 37810
rect 1030 37768 1086 37777
rect 1030 37703 1086 37712
rect 1032 37256 1084 37262
rect 1032 37198 1084 37204
rect 1044 36825 1072 37198
rect 1030 36816 1086 36825
rect 1030 36751 1086 36760
rect 1136 35766 1164 51046
rect 1320 39098 1348 57946
rect 1596 57882 1624 62086
rect 1412 57854 1624 57882
rect 1412 54262 1440 57854
rect 1584 57792 1636 57798
rect 1582 57760 1584 57769
rect 1636 57760 1638 57769
rect 1582 57695 1638 57704
rect 1492 56228 1544 56234
rect 1492 56170 1544 56176
rect 1400 54256 1452 54262
rect 1400 54198 1452 54204
rect 1504 51406 1532 56170
rect 1584 52352 1636 52358
rect 1582 52320 1584 52329
rect 1636 52320 1638 52329
rect 1582 52255 1638 52264
rect 1584 51808 1636 51814
rect 1584 51750 1636 51756
rect 1492 51400 1544 51406
rect 1492 51342 1544 51348
rect 1596 51074 1624 51750
rect 1504 51046 1624 51074
rect 1504 45558 1532 51046
rect 1584 48544 1636 48550
rect 1584 48486 1636 48492
rect 1596 48249 1624 48486
rect 1582 48240 1638 48249
rect 1582 48175 1638 48184
rect 1584 47116 1636 47122
rect 1584 47058 1636 47064
rect 1492 45552 1544 45558
rect 1492 45494 1544 45500
rect 1596 42090 1624 47058
rect 1584 42084 1636 42090
rect 1584 42026 1636 42032
rect 1492 40112 1544 40118
rect 1492 40054 1544 40060
rect 1504 39953 1532 40054
rect 1490 39944 1546 39953
rect 1490 39879 1546 39888
rect 1308 39092 1360 39098
rect 1308 39034 1360 39040
rect 1688 36242 1716 84458
rect 2950 83804 3258 83813
rect 2950 83802 2956 83804
rect 3012 83802 3036 83804
rect 3092 83802 3116 83804
rect 3172 83802 3196 83804
rect 3252 83802 3258 83804
rect 3012 83750 3014 83802
rect 3194 83750 3196 83802
rect 2950 83748 2956 83750
rect 3012 83748 3036 83750
rect 3092 83748 3116 83750
rect 3172 83748 3196 83750
rect 3252 83748 3258 83750
rect 2950 83739 3258 83748
rect 2228 82884 2280 82890
rect 2228 82826 2280 82832
rect 1768 81796 1820 81802
rect 1768 81738 1820 81744
rect 1676 36236 1728 36242
rect 1676 36178 1728 36184
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1216 36100 1268 36106
rect 1216 36042 1268 36048
rect 1124 35760 1176 35766
rect 1124 35702 1176 35708
rect 860 35142 980 35170
rect 756 26852 808 26858
rect 756 26794 808 26800
rect 768 16574 796 26794
rect 860 24614 888 35142
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34921 980 35022
rect 938 34912 994 34921
rect 938 34847 994 34856
rect 940 33992 992 33998
rect 938 33960 940 33969
rect 992 33960 994 33969
rect 938 33895 994 33904
rect 1124 33380 1176 33386
rect 1124 33322 1176 33328
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 952 32065 980 32370
rect 938 32056 994 32065
rect 938 31991 994 32000
rect 1032 32020 1084 32026
rect 1032 31962 1084 31968
rect 940 31340 992 31346
rect 940 31282 992 31288
rect 952 31113 980 31282
rect 938 31104 994 31113
rect 938 31039 994 31048
rect 940 30252 992 30258
rect 940 30194 992 30200
rect 952 30161 980 30194
rect 938 30152 994 30161
rect 938 30087 994 30096
rect 940 29640 992 29646
rect 940 29582 992 29588
rect 952 29209 980 29582
rect 938 29200 994 29209
rect 938 29135 994 29144
rect 940 28552 992 28558
rect 940 28494 992 28500
rect 952 28257 980 28494
rect 938 28248 994 28257
rect 938 28183 994 28192
rect 940 27464 992 27470
rect 940 27406 992 27412
rect 952 27305 980 27406
rect 938 27296 994 27305
rect 938 27231 994 27240
rect 940 26376 992 26382
rect 938 26344 940 26353
rect 992 26344 994 26353
rect 938 26279 994 26288
rect 940 25900 992 25906
rect 940 25842 992 25848
rect 952 25401 980 25842
rect 938 25392 994 25401
rect 938 25327 994 25336
rect 940 24812 992 24818
rect 940 24754 992 24760
rect 848 24608 900 24614
rect 848 24550 900 24556
rect 952 24449 980 24754
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 940 23724 992 23730
rect 940 23666 992 23672
rect 952 23497 980 23666
rect 938 23488 994 23497
rect 938 23423 994 23432
rect 940 22636 992 22642
rect 940 22578 992 22584
rect 952 22545 980 22578
rect 938 22536 994 22545
rect 938 22471 994 22480
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 952 19689 980 19790
rect 938 19680 994 19689
rect 938 19615 994 19624
rect 938 18728 994 18737
rect 938 18663 940 18672
rect 992 18663 994 18672
rect 940 18634 992 18640
rect 940 16992 992 16998
rect 940 16934 992 16940
rect 952 16833 980 16934
rect 938 16824 994 16833
rect 938 16759 994 16768
rect 768 16546 888 16574
rect 860 2310 888 16546
rect 940 15904 992 15910
rect 938 15872 940 15881
rect 992 15872 994 15881
rect 938 15807 994 15816
rect 938 14920 994 14929
rect 938 14855 994 14864
rect 952 14822 980 14855
rect 940 14816 992 14822
rect 940 14758 992 14764
rect 940 14272 992 14278
rect 940 14214 992 14220
rect 952 13977 980 14214
rect 938 13968 994 13977
rect 938 13903 994 13912
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 952 13025 980 13126
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 940 12096 992 12102
rect 938 12064 940 12073
rect 992 12064 994 12073
rect 938 11999 994 12008
rect 940 11348 992 11354
rect 940 11290 992 11296
rect 952 11121 980 11290
rect 938 11112 994 11121
rect 938 11047 994 11056
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10169 980 10406
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 952 9217 980 9318
rect 938 9208 994 9217
rect 938 9143 994 9152
rect 938 7304 994 7313
rect 938 7239 994 7248
rect 952 7206 980 7239
rect 940 7200 992 7206
rect 940 7142 992 7148
rect 940 6656 992 6662
rect 940 6598 992 6604
rect 952 6361 980 6598
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 940 4480 992 4486
rect 938 4448 940 4457
rect 992 4448 994 4457
rect 938 4383 994 4392
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 3398 980 3431
rect 940 3392 992 3398
rect 940 3334 992 3340
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 1044 1290 1072 31962
rect 1032 1284 1084 1290
rect 1032 1226 1084 1232
rect 1136 1222 1164 33322
rect 1228 2553 1256 36042
rect 1412 35873 1440 36110
rect 1398 35864 1454 35873
rect 1398 35799 1454 35808
rect 1308 35284 1360 35290
rect 1308 35226 1360 35232
rect 1214 2544 1270 2553
rect 1214 2479 1270 2488
rect 1124 1216 1176 1222
rect 1124 1158 1176 1164
rect 1320 377 1348 35226
rect 1780 34678 1808 81738
rect 1860 80708 1912 80714
rect 1860 80650 1912 80656
rect 1872 38554 1900 80650
rect 2044 79620 2096 79626
rect 2044 79562 2096 79568
rect 2056 74534 2084 79562
rect 2056 74506 2176 74534
rect 1952 74112 2004 74118
rect 1952 74054 2004 74060
rect 1964 42702 1992 74054
rect 2044 72684 2096 72690
rect 2044 72626 2096 72632
rect 2056 70514 2084 72626
rect 2044 70508 2096 70514
rect 2044 70450 2096 70456
rect 2148 70394 2176 74506
rect 2056 70366 2176 70394
rect 2056 60734 2084 70366
rect 2134 69320 2190 69329
rect 2134 69255 2136 69264
rect 2188 69255 2190 69264
rect 2136 69226 2188 69232
rect 2136 65476 2188 65482
rect 2136 65418 2188 65424
rect 2148 65113 2176 65418
rect 2134 65104 2190 65113
rect 2134 65039 2190 65048
rect 2136 65000 2188 65006
rect 2136 64942 2188 64948
rect 2148 63510 2176 64942
rect 2136 63504 2188 63510
rect 2136 63446 2188 63452
rect 2056 60706 2176 60734
rect 2148 55894 2176 60706
rect 2136 55888 2188 55894
rect 2136 55830 2188 55836
rect 2240 55214 2268 82826
rect 2950 82716 3258 82725
rect 2950 82714 2956 82716
rect 3012 82714 3036 82716
rect 3092 82714 3116 82716
rect 3172 82714 3196 82716
rect 3252 82714 3258 82716
rect 3012 82662 3014 82714
rect 3194 82662 3196 82714
rect 2950 82660 2956 82662
rect 3012 82660 3036 82662
rect 3092 82660 3116 82662
rect 3172 82660 3196 82662
rect 3252 82660 3258 82662
rect 2950 82651 3258 82660
rect 2950 81628 3258 81637
rect 2950 81626 2956 81628
rect 3012 81626 3036 81628
rect 3092 81626 3116 81628
rect 3172 81626 3196 81628
rect 3252 81626 3258 81628
rect 3012 81574 3014 81626
rect 3194 81574 3196 81626
rect 2950 81572 2956 81574
rect 3012 81572 3036 81574
rect 3092 81572 3116 81574
rect 3172 81572 3196 81574
rect 3252 81572 3258 81574
rect 2950 81563 3258 81572
rect 2950 80540 3258 80549
rect 2950 80538 2956 80540
rect 3012 80538 3036 80540
rect 3092 80538 3116 80540
rect 3172 80538 3196 80540
rect 3252 80538 3258 80540
rect 3012 80486 3014 80538
rect 3194 80486 3196 80538
rect 2950 80484 2956 80486
rect 3012 80484 3036 80486
rect 3092 80484 3116 80486
rect 3172 80484 3196 80486
rect 3252 80484 3258 80486
rect 2950 80475 3258 80484
rect 2950 79452 3258 79461
rect 2950 79450 2956 79452
rect 3012 79450 3036 79452
rect 3092 79450 3116 79452
rect 3172 79450 3196 79452
rect 3252 79450 3258 79452
rect 3012 79398 3014 79450
rect 3194 79398 3196 79450
rect 2950 79396 2956 79398
rect 3012 79396 3036 79398
rect 3092 79396 3116 79398
rect 3172 79396 3196 79398
rect 3252 79396 3258 79398
rect 2950 79387 3258 79396
rect 2950 78364 3258 78373
rect 2950 78362 2956 78364
rect 3012 78362 3036 78364
rect 3092 78362 3116 78364
rect 3172 78362 3196 78364
rect 3252 78362 3258 78364
rect 3012 78310 3014 78362
rect 3194 78310 3196 78362
rect 2950 78308 2956 78310
rect 3012 78308 3036 78310
rect 3092 78308 3116 78310
rect 3172 78308 3196 78310
rect 3252 78308 3258 78310
rect 2950 78299 3258 78308
rect 3332 77920 3384 77926
rect 3332 77862 3384 77868
rect 2950 77276 3258 77285
rect 2950 77274 2956 77276
rect 3012 77274 3036 77276
rect 3092 77274 3116 77276
rect 3172 77274 3196 77276
rect 3252 77274 3258 77276
rect 3012 77222 3014 77274
rect 3194 77222 3196 77274
rect 2950 77220 2956 77222
rect 3012 77220 3036 77222
rect 3092 77220 3116 77222
rect 3172 77220 3196 77222
rect 3252 77220 3258 77222
rect 2950 77211 3258 77220
rect 2596 76900 2648 76906
rect 2596 76842 2648 76848
rect 2504 76832 2556 76838
rect 2504 76774 2556 76780
rect 2412 70848 2464 70854
rect 2412 70790 2464 70796
rect 2320 67652 2372 67658
rect 2320 67594 2372 67600
rect 2332 62966 2360 67594
rect 2424 65686 2452 70790
rect 2516 68218 2544 76774
rect 2608 69873 2636 76842
rect 2950 76188 3258 76197
rect 2950 76186 2956 76188
rect 3012 76186 3036 76188
rect 3092 76186 3116 76188
rect 3172 76186 3196 76188
rect 3252 76186 3258 76188
rect 3012 76134 3014 76186
rect 3194 76134 3196 76186
rect 2950 76132 2956 76134
rect 3012 76132 3036 76134
rect 3092 76132 3116 76134
rect 3172 76132 3196 76134
rect 3252 76132 3258 76134
rect 2950 76123 3258 76132
rect 2688 75268 2740 75274
rect 2688 75210 2740 75216
rect 2700 70009 2728 75210
rect 2950 75100 3258 75109
rect 2950 75098 2956 75100
rect 3012 75098 3036 75100
rect 3092 75098 3116 75100
rect 3172 75098 3196 75100
rect 3252 75098 3258 75100
rect 3012 75046 3014 75098
rect 3194 75046 3196 75098
rect 2950 75044 2956 75046
rect 3012 75044 3036 75046
rect 3092 75044 3116 75046
rect 3172 75044 3196 75046
rect 3252 75044 3258 75046
rect 2950 75035 3258 75044
rect 2950 74012 3258 74021
rect 2950 74010 2956 74012
rect 3012 74010 3036 74012
rect 3092 74010 3116 74012
rect 3172 74010 3196 74012
rect 3252 74010 3258 74012
rect 3012 73958 3014 74010
rect 3194 73958 3196 74010
rect 2950 73956 2956 73958
rect 3012 73956 3036 73958
rect 3092 73956 3116 73958
rect 3172 73956 3196 73958
rect 3252 73956 3258 73958
rect 2950 73947 3258 73956
rect 2950 72924 3258 72933
rect 2950 72922 2956 72924
rect 3012 72922 3036 72924
rect 3092 72922 3116 72924
rect 3172 72922 3196 72924
rect 3252 72922 3258 72924
rect 3012 72870 3014 72922
rect 3194 72870 3196 72922
rect 2950 72868 2956 72870
rect 3012 72868 3036 72870
rect 3092 72868 3116 72870
rect 3172 72868 3196 72870
rect 3252 72868 3258 72870
rect 2950 72859 3258 72868
rect 2950 71836 3258 71845
rect 2950 71834 2956 71836
rect 3012 71834 3036 71836
rect 3092 71834 3116 71836
rect 3172 71834 3196 71836
rect 3252 71834 3258 71836
rect 3012 71782 3014 71834
rect 3194 71782 3196 71834
rect 2950 71780 2956 71782
rect 3012 71780 3036 71782
rect 3092 71780 3116 71782
rect 3172 71780 3196 71782
rect 3252 71780 3258 71782
rect 2950 71771 3258 71780
rect 2870 71496 2926 71505
rect 2870 71431 2926 71440
rect 2780 70916 2832 70922
rect 2780 70858 2832 70864
rect 2686 70000 2742 70009
rect 2686 69935 2742 69944
rect 2594 69864 2650 69873
rect 2594 69799 2650 69808
rect 2792 68932 2820 70858
rect 2700 68904 2820 68932
rect 2516 68190 2636 68218
rect 2504 68128 2556 68134
rect 2504 68070 2556 68076
rect 2412 65680 2464 65686
rect 2412 65622 2464 65628
rect 2412 65544 2464 65550
rect 2412 65486 2464 65492
rect 2424 64920 2452 65486
rect 2516 65142 2544 68070
rect 2504 65136 2556 65142
rect 2504 65078 2556 65084
rect 2608 65074 2636 68190
rect 2700 65634 2728 68904
rect 2778 68232 2834 68241
rect 2778 68167 2834 68176
rect 2792 65793 2820 68167
rect 2884 68134 2912 71431
rect 2950 70748 3258 70757
rect 2950 70746 2956 70748
rect 3012 70746 3036 70748
rect 3092 70746 3116 70748
rect 3172 70746 3196 70748
rect 3252 70746 3258 70748
rect 3012 70694 3014 70746
rect 3194 70694 3196 70746
rect 2950 70692 2956 70694
rect 3012 70692 3036 70694
rect 3092 70692 3116 70694
rect 3172 70692 3196 70694
rect 3252 70692 3258 70694
rect 2950 70683 3258 70692
rect 2950 69660 3258 69669
rect 2950 69658 2956 69660
rect 3012 69658 3036 69660
rect 3092 69658 3116 69660
rect 3172 69658 3196 69660
rect 3252 69658 3258 69660
rect 3012 69606 3014 69658
rect 3194 69606 3196 69658
rect 2950 69604 2956 69606
rect 3012 69604 3036 69606
rect 3092 69604 3116 69606
rect 3172 69604 3196 69606
rect 3252 69604 3258 69606
rect 2950 69595 3258 69604
rect 2950 68572 3258 68581
rect 2950 68570 2956 68572
rect 3012 68570 3036 68572
rect 3092 68570 3116 68572
rect 3172 68570 3196 68572
rect 3252 68570 3258 68572
rect 3012 68518 3014 68570
rect 3194 68518 3196 68570
rect 2950 68516 2956 68518
rect 3012 68516 3036 68518
rect 3092 68516 3116 68518
rect 3172 68516 3196 68518
rect 3252 68516 3258 68518
rect 2950 68507 3258 68516
rect 2872 68128 2924 68134
rect 2872 68070 2924 68076
rect 2950 67484 3258 67493
rect 2950 67482 2956 67484
rect 3012 67482 3036 67484
rect 3092 67482 3116 67484
rect 3172 67482 3196 67484
rect 3252 67482 3258 67484
rect 3012 67430 3014 67482
rect 3194 67430 3196 67482
rect 2950 67428 2956 67430
rect 3012 67428 3036 67430
rect 3092 67428 3116 67430
rect 3172 67428 3196 67430
rect 3252 67428 3258 67430
rect 2950 67419 3258 67428
rect 2950 66396 3258 66405
rect 2950 66394 2956 66396
rect 3012 66394 3036 66396
rect 3092 66394 3116 66396
rect 3172 66394 3196 66396
rect 3252 66394 3258 66396
rect 3012 66342 3014 66394
rect 3194 66342 3196 66394
rect 2950 66340 2956 66342
rect 3012 66340 3036 66342
rect 3092 66340 3116 66342
rect 3172 66340 3196 66342
rect 3252 66340 3258 66342
rect 2950 66331 3258 66340
rect 2778 65784 2834 65793
rect 3344 65754 3372 77862
rect 2778 65719 2834 65728
rect 3332 65748 3384 65754
rect 3332 65690 3384 65696
rect 2700 65606 2820 65634
rect 2688 65544 2740 65550
rect 2688 65486 2740 65492
rect 2596 65068 2648 65074
rect 2596 65010 2648 65016
rect 2424 64892 2544 64920
rect 2412 64660 2464 64666
rect 2412 64602 2464 64608
rect 2320 62960 2372 62966
rect 2320 62902 2372 62908
rect 2320 62824 2372 62830
rect 2320 62766 2372 62772
rect 2056 55186 2268 55214
rect 2056 46186 2084 55186
rect 2136 53576 2188 53582
rect 2136 53518 2188 53524
rect 2148 48314 2176 53518
rect 2228 51060 2280 51066
rect 2228 51002 2280 51008
rect 2240 49434 2268 51002
rect 2332 49910 2360 62766
rect 2424 55350 2452 64602
rect 2516 63594 2544 64892
rect 2700 64546 2728 65486
rect 2792 65482 2820 65606
rect 2780 65476 2832 65482
rect 2780 65418 2832 65424
rect 3332 65476 3384 65482
rect 3332 65418 3384 65424
rect 2778 65376 2834 65385
rect 2778 65311 2834 65320
rect 2792 64666 2820 65311
rect 2950 65308 3258 65317
rect 2950 65306 2956 65308
rect 3012 65306 3036 65308
rect 3092 65306 3116 65308
rect 3172 65306 3196 65308
rect 3252 65306 3258 65308
rect 3012 65254 3014 65306
rect 3194 65254 3196 65306
rect 2950 65252 2956 65254
rect 3012 65252 3036 65254
rect 3092 65252 3116 65254
rect 3172 65252 3196 65254
rect 3252 65252 3258 65254
rect 2950 65243 3258 65252
rect 3240 65000 3292 65006
rect 3240 64942 3292 64948
rect 2872 64864 2924 64870
rect 2872 64806 2924 64812
rect 2780 64660 2832 64666
rect 2780 64602 2832 64608
rect 2700 64518 2820 64546
rect 2688 64456 2740 64462
rect 2688 64398 2740 64404
rect 2516 63566 2636 63594
rect 2504 63504 2556 63510
rect 2504 63446 2556 63452
rect 2516 62218 2544 63446
rect 2504 62212 2556 62218
rect 2504 62154 2556 62160
rect 2608 57594 2636 63566
rect 2700 60722 2728 64398
rect 2688 60716 2740 60722
rect 2688 60658 2740 60664
rect 2792 60602 2820 64518
rect 2700 60574 2820 60602
rect 2700 57934 2728 60574
rect 2780 60512 2832 60518
rect 2780 60454 2832 60460
rect 2792 60178 2820 60454
rect 2780 60172 2832 60178
rect 2780 60114 2832 60120
rect 2780 59424 2832 59430
rect 2780 59366 2832 59372
rect 2688 57928 2740 57934
rect 2688 57870 2740 57876
rect 2596 57588 2648 57594
rect 2596 57530 2648 57536
rect 2688 56160 2740 56166
rect 2688 56102 2740 56108
rect 2412 55344 2464 55350
rect 2412 55286 2464 55292
rect 2700 55214 2728 56102
rect 2516 55186 2728 55214
rect 2412 52896 2464 52902
rect 2412 52838 2464 52844
rect 2424 50998 2452 52838
rect 2516 51066 2544 55186
rect 2596 54052 2648 54058
rect 2596 53994 2648 54000
rect 2608 51066 2636 53994
rect 2688 53984 2740 53990
rect 2688 53926 2740 53932
rect 2504 51060 2556 51066
rect 2504 51002 2556 51008
rect 2596 51060 2648 51066
rect 2596 51002 2648 51008
rect 2412 50992 2464 50998
rect 2412 50934 2464 50940
rect 2412 50788 2464 50794
rect 2412 50730 2464 50736
rect 2320 49904 2372 49910
rect 2320 49846 2372 49852
rect 2228 49428 2280 49434
rect 2228 49370 2280 49376
rect 2148 48286 2360 48314
rect 2056 46158 2268 46186
rect 2044 44940 2096 44946
rect 2044 44882 2096 44888
rect 1952 42696 2004 42702
rect 1952 42638 2004 42644
rect 1952 42016 2004 42022
rect 1952 41958 2004 41964
rect 1860 38548 1912 38554
rect 1860 38490 1912 38496
rect 1860 37256 1912 37262
rect 1860 37198 1912 37204
rect 1768 34672 1820 34678
rect 1768 34614 1820 34620
rect 1492 33516 1544 33522
rect 1492 33458 1544 33464
rect 1504 33153 1532 33458
rect 1490 33144 1546 33153
rect 1490 33079 1546 33088
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 31890 1808 32166
rect 1768 31884 1820 31890
rect 1768 31826 1820 31832
rect 1584 31204 1636 31210
rect 1584 31146 1636 31152
rect 1400 28416 1452 28422
rect 1400 28358 1452 28364
rect 1412 28218 1440 28358
rect 1400 28212 1452 28218
rect 1400 28154 1452 28160
rect 1596 26042 1624 31146
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1596 23866 1624 25298
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20641 1440 20878
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17785 1624 18022
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 1688 2009 1716 27338
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1780 8566 1808 25638
rect 1872 13326 1900 37198
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1964 12238 1992 41958
rect 2056 17270 2084 44882
rect 2136 41540 2188 41546
rect 2136 41482 2188 41488
rect 2148 32910 2176 41482
rect 2240 35834 2268 46158
rect 2332 45014 2360 48286
rect 2424 46646 2452 50730
rect 2504 50720 2556 50726
rect 2504 50662 2556 50668
rect 2412 46640 2464 46646
rect 2412 46582 2464 46588
rect 2516 46170 2544 50662
rect 2700 47734 2728 53926
rect 2792 53174 2820 59366
rect 2884 59022 2912 64806
rect 3252 64462 3280 64942
rect 3240 64456 3292 64462
rect 3240 64398 3292 64404
rect 2950 64220 3258 64229
rect 2950 64218 2956 64220
rect 3012 64218 3036 64220
rect 3092 64218 3116 64220
rect 3172 64218 3196 64220
rect 3252 64218 3258 64220
rect 3012 64166 3014 64218
rect 3194 64166 3196 64218
rect 2950 64164 2956 64166
rect 3012 64164 3036 64166
rect 3092 64164 3116 64166
rect 3172 64164 3196 64166
rect 3252 64164 3258 64166
rect 2950 64155 3258 64164
rect 2950 63132 3258 63141
rect 2950 63130 2956 63132
rect 3012 63130 3036 63132
rect 3092 63130 3116 63132
rect 3172 63130 3196 63132
rect 3252 63130 3258 63132
rect 3012 63078 3014 63130
rect 3194 63078 3196 63130
rect 2950 63076 2956 63078
rect 3012 63076 3036 63078
rect 3092 63076 3116 63078
rect 3172 63076 3196 63078
rect 3252 63076 3258 63078
rect 2950 63067 3258 63076
rect 2950 62044 3258 62053
rect 2950 62042 2956 62044
rect 3012 62042 3036 62044
rect 3092 62042 3116 62044
rect 3172 62042 3196 62044
rect 3252 62042 3258 62044
rect 3012 61990 3014 62042
rect 3194 61990 3196 62042
rect 2950 61988 2956 61990
rect 3012 61988 3036 61990
rect 3092 61988 3116 61990
rect 3172 61988 3196 61990
rect 3252 61988 3258 61990
rect 2950 61979 3258 61988
rect 2950 60956 3258 60965
rect 2950 60954 2956 60956
rect 3012 60954 3036 60956
rect 3092 60954 3116 60956
rect 3172 60954 3196 60956
rect 3252 60954 3258 60956
rect 3012 60902 3014 60954
rect 3194 60902 3196 60954
rect 2950 60900 2956 60902
rect 3012 60900 3036 60902
rect 3092 60900 3116 60902
rect 3172 60900 3196 60902
rect 3252 60900 3258 60902
rect 2950 60891 3258 60900
rect 2950 59868 3258 59877
rect 2950 59866 2956 59868
rect 3012 59866 3036 59868
rect 3092 59866 3116 59868
rect 3172 59866 3196 59868
rect 3252 59866 3258 59868
rect 3012 59814 3014 59866
rect 3194 59814 3196 59866
rect 2950 59812 2956 59814
rect 3012 59812 3036 59814
rect 3092 59812 3116 59814
rect 3172 59812 3196 59814
rect 3252 59812 3258 59814
rect 2950 59803 3258 59812
rect 2872 59016 2924 59022
rect 2872 58958 2924 58964
rect 2950 58780 3258 58789
rect 2950 58778 2956 58780
rect 3012 58778 3036 58780
rect 3092 58778 3116 58780
rect 3172 58778 3196 58780
rect 3252 58778 3258 58780
rect 3012 58726 3014 58778
rect 3194 58726 3196 58778
rect 2950 58724 2956 58726
rect 3012 58724 3036 58726
rect 3092 58724 3116 58726
rect 3172 58724 3196 58726
rect 3252 58724 3258 58726
rect 2950 58715 3258 58724
rect 2950 57692 3258 57701
rect 2950 57690 2956 57692
rect 3012 57690 3036 57692
rect 3092 57690 3116 57692
rect 3172 57690 3196 57692
rect 3252 57690 3258 57692
rect 3012 57638 3014 57690
rect 3194 57638 3196 57690
rect 2950 57636 2956 57638
rect 3012 57636 3036 57638
rect 3092 57636 3116 57638
rect 3172 57636 3196 57638
rect 3252 57636 3258 57638
rect 2950 57627 3258 57636
rect 2950 56604 3258 56613
rect 2950 56602 2956 56604
rect 3012 56602 3036 56604
rect 3092 56602 3116 56604
rect 3172 56602 3196 56604
rect 3252 56602 3258 56604
rect 3012 56550 3014 56602
rect 3194 56550 3196 56602
rect 2950 56548 2956 56550
rect 3012 56548 3036 56550
rect 3092 56548 3116 56550
rect 3172 56548 3196 56550
rect 3252 56548 3258 56550
rect 2950 56539 3258 56548
rect 3344 56438 3372 65418
rect 3332 56432 3384 56438
rect 3332 56374 3384 56380
rect 3332 56296 3384 56302
rect 3332 56238 3384 56244
rect 2950 55516 3258 55525
rect 2950 55514 2956 55516
rect 3012 55514 3036 55516
rect 3092 55514 3116 55516
rect 3172 55514 3196 55516
rect 3252 55514 3258 55516
rect 3012 55462 3014 55514
rect 3194 55462 3196 55514
rect 2950 55460 2956 55462
rect 3012 55460 3036 55462
rect 3092 55460 3116 55462
rect 3172 55460 3196 55462
rect 3252 55460 3258 55462
rect 2950 55451 3258 55460
rect 2872 54528 2924 54534
rect 2872 54470 2924 54476
rect 2780 53168 2832 53174
rect 2780 53110 2832 53116
rect 2780 52964 2832 52970
rect 2780 52906 2832 52912
rect 2688 47728 2740 47734
rect 2688 47670 2740 47676
rect 2792 46986 2820 52906
rect 2884 48822 2912 54470
rect 2950 54428 3258 54437
rect 2950 54426 2956 54428
rect 3012 54426 3036 54428
rect 3092 54426 3116 54428
rect 3172 54426 3196 54428
rect 3252 54426 3258 54428
rect 3012 54374 3014 54426
rect 3194 54374 3196 54426
rect 2950 54372 2956 54374
rect 3012 54372 3036 54374
rect 3092 54372 3116 54374
rect 3172 54372 3196 54374
rect 3252 54372 3258 54374
rect 2950 54363 3258 54372
rect 2950 53340 3258 53349
rect 2950 53338 2956 53340
rect 3012 53338 3036 53340
rect 3092 53338 3116 53340
rect 3172 53338 3196 53340
rect 3252 53338 3258 53340
rect 3012 53286 3014 53338
rect 3194 53286 3196 53338
rect 2950 53284 2956 53286
rect 3012 53284 3036 53286
rect 3092 53284 3116 53286
rect 3172 53284 3196 53286
rect 3252 53284 3258 53286
rect 2950 53275 3258 53284
rect 2950 52252 3258 52261
rect 2950 52250 2956 52252
rect 3012 52250 3036 52252
rect 3092 52250 3116 52252
rect 3172 52250 3196 52252
rect 3252 52250 3258 52252
rect 3012 52198 3014 52250
rect 3194 52198 3196 52250
rect 2950 52196 2956 52198
rect 3012 52196 3036 52198
rect 3092 52196 3116 52198
rect 3172 52196 3196 52198
rect 3252 52196 3258 52198
rect 2950 52187 3258 52196
rect 2950 51164 3258 51173
rect 2950 51162 2956 51164
rect 3012 51162 3036 51164
rect 3092 51162 3116 51164
rect 3172 51162 3196 51164
rect 3252 51162 3258 51164
rect 3012 51110 3014 51162
rect 3194 51110 3196 51162
rect 2950 51108 2956 51110
rect 3012 51108 3036 51110
rect 3092 51108 3116 51110
rect 3172 51108 3196 51110
rect 3252 51108 3258 51110
rect 2950 51099 3258 51108
rect 3344 50318 3372 56238
rect 3332 50312 3384 50318
rect 3332 50254 3384 50260
rect 2950 50076 3258 50085
rect 2950 50074 2956 50076
rect 3012 50074 3036 50076
rect 3092 50074 3116 50076
rect 3172 50074 3196 50076
rect 3252 50074 3258 50076
rect 3012 50022 3014 50074
rect 3194 50022 3196 50074
rect 2950 50020 2956 50022
rect 3012 50020 3036 50022
rect 3092 50020 3116 50022
rect 3172 50020 3196 50022
rect 3252 50020 3258 50022
rect 2950 50011 3258 50020
rect 3332 49768 3384 49774
rect 3332 49710 3384 49716
rect 2950 48988 3258 48997
rect 2950 48986 2956 48988
rect 3012 48986 3036 48988
rect 3092 48986 3116 48988
rect 3172 48986 3196 48988
rect 3252 48986 3258 48988
rect 3012 48934 3014 48986
rect 3194 48934 3196 48986
rect 2950 48932 2956 48934
rect 3012 48932 3036 48934
rect 3092 48932 3116 48934
rect 3172 48932 3196 48934
rect 3252 48932 3258 48934
rect 2950 48923 3258 48932
rect 2872 48816 2924 48822
rect 2872 48758 2924 48764
rect 2950 47900 3258 47909
rect 2950 47898 2956 47900
rect 3012 47898 3036 47900
rect 3092 47898 3116 47900
rect 3172 47898 3196 47900
rect 3252 47898 3258 47900
rect 3012 47846 3014 47898
rect 3194 47846 3196 47898
rect 2950 47844 2956 47846
rect 3012 47844 3036 47846
rect 3092 47844 3116 47846
rect 3172 47844 3196 47846
rect 3252 47844 3258 47846
rect 2950 47835 3258 47844
rect 2872 47456 2924 47462
rect 2872 47398 2924 47404
rect 2780 46980 2832 46986
rect 2780 46922 2832 46928
rect 2884 46322 2912 47398
rect 3344 47122 3372 49710
rect 3332 47116 3384 47122
rect 3332 47058 3384 47064
rect 3332 46980 3384 46986
rect 3332 46922 3384 46928
rect 2950 46812 3258 46821
rect 2950 46810 2956 46812
rect 3012 46810 3036 46812
rect 3092 46810 3116 46812
rect 3172 46810 3196 46812
rect 3252 46810 3258 46812
rect 3012 46758 3014 46810
rect 3194 46758 3196 46810
rect 2950 46756 2956 46758
rect 3012 46756 3036 46758
rect 3092 46756 3116 46758
rect 3172 46756 3196 46758
rect 3252 46756 3258 46758
rect 2950 46747 3258 46756
rect 2792 46294 2912 46322
rect 2504 46164 2556 46170
rect 2504 46106 2556 46112
rect 2504 45824 2556 45830
rect 2504 45766 2556 45772
rect 2320 45008 2372 45014
rect 2320 44950 2372 44956
rect 2516 42362 2544 45766
rect 2688 44736 2740 44742
rect 2688 44678 2740 44684
rect 2596 42696 2648 42702
rect 2596 42638 2648 42644
rect 2504 42356 2556 42362
rect 2504 42298 2556 42304
rect 2608 42226 2636 42638
rect 2596 42220 2648 42226
rect 2596 42162 2648 42168
rect 2504 41472 2556 41478
rect 2504 41414 2556 41420
rect 2700 41414 2728 44678
rect 2792 41750 2820 46294
rect 2872 46164 2924 46170
rect 2872 46106 2924 46112
rect 2884 44402 2912 46106
rect 2950 45724 3258 45733
rect 2950 45722 2956 45724
rect 3012 45722 3036 45724
rect 3092 45722 3116 45724
rect 3172 45722 3196 45724
rect 3252 45722 3258 45724
rect 3012 45670 3014 45722
rect 3194 45670 3196 45722
rect 2950 45668 2956 45670
rect 3012 45668 3036 45670
rect 3092 45668 3116 45670
rect 3172 45668 3196 45670
rect 3252 45668 3258 45670
rect 2950 45659 3258 45668
rect 2950 44636 3258 44645
rect 2950 44634 2956 44636
rect 3012 44634 3036 44636
rect 3092 44634 3116 44636
rect 3172 44634 3196 44636
rect 3252 44634 3258 44636
rect 3012 44582 3014 44634
rect 3194 44582 3196 44634
rect 2950 44580 2956 44582
rect 3012 44580 3036 44582
rect 3092 44580 3116 44582
rect 3172 44580 3196 44582
rect 3252 44580 3258 44582
rect 2950 44571 3258 44580
rect 2872 44396 2924 44402
rect 2872 44338 2924 44344
rect 2950 43548 3258 43557
rect 2950 43546 2956 43548
rect 3012 43546 3036 43548
rect 3092 43546 3116 43548
rect 3172 43546 3196 43548
rect 3252 43546 3258 43548
rect 3012 43494 3014 43546
rect 3194 43494 3196 43546
rect 2950 43492 2956 43494
rect 3012 43492 3036 43494
rect 3092 43492 3116 43494
rect 3172 43492 3196 43494
rect 3252 43492 3258 43494
rect 2950 43483 3258 43492
rect 3344 42770 3372 46922
rect 3332 42764 3384 42770
rect 3332 42706 3384 42712
rect 2950 42460 3258 42469
rect 2950 42458 2956 42460
rect 3012 42458 3036 42460
rect 3092 42458 3116 42460
rect 3172 42458 3196 42460
rect 3252 42458 3258 42460
rect 3012 42406 3014 42458
rect 3194 42406 3196 42458
rect 2950 42404 2956 42406
rect 3012 42404 3036 42406
rect 3092 42404 3116 42406
rect 3172 42404 3196 42406
rect 3252 42404 3258 42406
rect 2950 42395 3258 42404
rect 3332 42084 3384 42090
rect 3332 42026 3384 42032
rect 2780 41744 2832 41750
rect 2780 41686 2832 41692
rect 2320 37664 2372 37670
rect 2320 37606 2372 37612
rect 2228 35828 2280 35834
rect 2228 35770 2280 35776
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2332 24750 2360 37606
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2320 24744 2372 24750
rect 2320 24686 2372 24692
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 2148 6798 2176 21830
rect 2240 10742 2268 24006
rect 2424 23594 2452 37130
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2332 3534 2360 22918
rect 2516 11150 2544 41414
rect 2608 41386 2728 41414
rect 2608 40526 2636 41386
rect 2950 41372 3258 41381
rect 2950 41370 2956 41372
rect 3012 41370 3036 41372
rect 3092 41370 3116 41372
rect 3172 41370 3196 41372
rect 3252 41370 3258 41372
rect 3012 41318 3014 41370
rect 3194 41318 3196 41370
rect 2950 41316 2956 41318
rect 3012 41316 3036 41318
rect 3092 41316 3116 41318
rect 3172 41316 3196 41318
rect 3252 41316 3258 41318
rect 2950 41307 3258 41316
rect 2596 40520 2648 40526
rect 2596 40462 2648 40468
rect 2950 40284 3258 40293
rect 2950 40282 2956 40284
rect 3012 40282 3036 40284
rect 3092 40282 3116 40284
rect 3172 40282 3196 40284
rect 3252 40282 3258 40284
rect 3012 40230 3014 40282
rect 3194 40230 3196 40282
rect 2950 40228 2956 40230
rect 3012 40228 3036 40230
rect 3092 40228 3116 40230
rect 3172 40228 3196 40230
rect 3252 40228 3258 40230
rect 2950 40219 3258 40228
rect 2688 39840 2740 39846
rect 2688 39782 2740 39788
rect 2700 37466 2728 39782
rect 2950 39196 3258 39205
rect 2950 39194 2956 39196
rect 3012 39194 3036 39196
rect 3092 39194 3116 39196
rect 3172 39194 3196 39196
rect 3252 39194 3258 39196
rect 3012 39142 3014 39194
rect 3194 39142 3196 39194
rect 2950 39140 2956 39142
rect 3012 39140 3036 39142
rect 3092 39140 3116 39142
rect 3172 39140 3196 39142
rect 3252 39140 3258 39142
rect 2950 39131 3258 39140
rect 2780 38752 2832 38758
rect 2780 38694 2832 38700
rect 2688 37460 2740 37466
rect 2688 37402 2740 37408
rect 2688 35148 2740 35154
rect 2688 35090 2740 35096
rect 2700 31210 2728 35090
rect 2688 31204 2740 31210
rect 2688 31146 2740 31152
rect 2596 27872 2648 27878
rect 2596 27814 2648 27820
rect 2608 24206 2636 27814
rect 2792 26466 2820 38694
rect 2872 38548 2924 38554
rect 2872 38490 2924 38496
rect 2884 35196 2912 38490
rect 2950 38108 3258 38117
rect 2950 38106 2956 38108
rect 3012 38106 3036 38108
rect 3092 38106 3116 38108
rect 3172 38106 3196 38108
rect 3252 38106 3258 38108
rect 3012 38054 3014 38106
rect 3194 38054 3196 38106
rect 2950 38052 2956 38054
rect 3012 38052 3036 38054
rect 3092 38052 3116 38054
rect 3172 38052 3196 38054
rect 3252 38052 3258 38054
rect 2950 38043 3258 38052
rect 2950 37020 3258 37029
rect 2950 37018 2956 37020
rect 3012 37018 3036 37020
rect 3092 37018 3116 37020
rect 3172 37018 3196 37020
rect 3252 37018 3258 37020
rect 3012 36966 3014 37018
rect 3194 36966 3196 37018
rect 2950 36964 2956 36966
rect 3012 36964 3036 36966
rect 3092 36964 3116 36966
rect 3172 36964 3196 36966
rect 3252 36964 3258 36966
rect 2950 36955 3258 36964
rect 2950 35932 3258 35941
rect 2950 35930 2956 35932
rect 3012 35930 3036 35932
rect 3092 35930 3116 35932
rect 3172 35930 3196 35932
rect 3252 35930 3258 35932
rect 3012 35878 3014 35930
rect 3194 35878 3196 35930
rect 2950 35876 2956 35878
rect 3012 35876 3036 35878
rect 3092 35876 3116 35878
rect 3172 35876 3196 35878
rect 3252 35876 3258 35878
rect 2950 35867 3258 35876
rect 2884 35168 3280 35196
rect 3252 35034 3280 35168
rect 3344 35154 3372 42026
rect 3332 35148 3384 35154
rect 3332 35090 3384 35096
rect 3252 35006 3372 35034
rect 2872 34944 2924 34950
rect 2872 34886 2924 34892
rect 2700 26438 2820 26466
rect 2700 25650 2728 26438
rect 2884 26246 2912 34886
rect 2950 34844 3258 34853
rect 2950 34842 2956 34844
rect 3012 34842 3036 34844
rect 3092 34842 3116 34844
rect 3172 34842 3196 34844
rect 3252 34842 3258 34844
rect 3012 34790 3014 34842
rect 3194 34790 3196 34842
rect 2950 34788 2956 34790
rect 3012 34788 3036 34790
rect 3092 34788 3116 34790
rect 3172 34788 3196 34790
rect 3252 34788 3258 34790
rect 2950 34779 3258 34788
rect 3344 34202 3372 35006
rect 3332 34196 3384 34202
rect 3332 34138 3384 34144
rect 3332 33856 3384 33862
rect 3332 33798 3384 33804
rect 2950 33756 3258 33765
rect 2950 33754 2956 33756
rect 3012 33754 3036 33756
rect 3092 33754 3116 33756
rect 3172 33754 3196 33756
rect 3252 33754 3258 33756
rect 3012 33702 3014 33754
rect 3194 33702 3196 33754
rect 2950 33700 2956 33702
rect 3012 33700 3036 33702
rect 3092 33700 3116 33702
rect 3172 33700 3196 33702
rect 3252 33700 3258 33702
rect 2950 33691 3258 33700
rect 2950 32668 3258 32677
rect 2950 32666 2956 32668
rect 3012 32666 3036 32668
rect 3092 32666 3116 32668
rect 3172 32666 3196 32668
rect 3252 32666 3258 32668
rect 3012 32614 3014 32666
rect 3194 32614 3196 32666
rect 2950 32612 2956 32614
rect 3012 32612 3036 32614
rect 3092 32612 3116 32614
rect 3172 32612 3196 32614
rect 3252 32612 3258 32614
rect 2950 32603 3258 32612
rect 2950 31580 3258 31589
rect 2950 31578 2956 31580
rect 3012 31578 3036 31580
rect 3092 31578 3116 31580
rect 3172 31578 3196 31580
rect 3252 31578 3258 31580
rect 3012 31526 3014 31578
rect 3194 31526 3196 31578
rect 2950 31524 2956 31526
rect 3012 31524 3036 31526
rect 3092 31524 3116 31526
rect 3172 31524 3196 31526
rect 3252 31524 3258 31526
rect 2950 31515 3258 31524
rect 2950 30492 3258 30501
rect 2950 30490 2956 30492
rect 3012 30490 3036 30492
rect 3092 30490 3116 30492
rect 3172 30490 3196 30492
rect 3252 30490 3258 30492
rect 3012 30438 3014 30490
rect 3194 30438 3196 30490
rect 2950 30436 2956 30438
rect 3012 30436 3036 30438
rect 3092 30436 3116 30438
rect 3172 30436 3196 30438
rect 3252 30436 3258 30438
rect 2950 30427 3258 30436
rect 2950 29404 3258 29413
rect 2950 29402 2956 29404
rect 3012 29402 3036 29404
rect 3092 29402 3116 29404
rect 3172 29402 3196 29404
rect 3252 29402 3258 29404
rect 3012 29350 3014 29402
rect 3194 29350 3196 29402
rect 2950 29348 2956 29350
rect 3012 29348 3036 29350
rect 3092 29348 3116 29350
rect 3172 29348 3196 29350
rect 3252 29348 3258 29350
rect 2950 29339 3258 29348
rect 2950 28316 3258 28325
rect 2950 28314 2956 28316
rect 3012 28314 3036 28316
rect 3092 28314 3116 28316
rect 3172 28314 3196 28316
rect 3252 28314 3258 28316
rect 3012 28262 3014 28314
rect 3194 28262 3196 28314
rect 2950 28260 2956 28262
rect 3012 28260 3036 28262
rect 3092 28260 3116 28262
rect 3172 28260 3196 28262
rect 3252 28260 3258 28262
rect 2950 28251 3258 28260
rect 3344 27878 3372 33798
rect 3332 27872 3384 27878
rect 3332 27814 3384 27820
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 2950 27228 3258 27237
rect 2950 27226 2956 27228
rect 3012 27226 3036 27228
rect 3092 27226 3116 27228
rect 3172 27226 3196 27228
rect 3252 27226 3258 27228
rect 3012 27174 3014 27226
rect 3194 27174 3196 27226
rect 2950 27172 2956 27174
rect 3012 27172 3036 27174
rect 3092 27172 3116 27174
rect 3172 27172 3196 27174
rect 3252 27172 3258 27174
rect 2950 27163 3258 27172
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2950 26140 3258 26149
rect 2950 26138 2956 26140
rect 3012 26138 3036 26140
rect 3092 26138 3116 26140
rect 3172 26138 3196 26140
rect 3252 26138 3258 26140
rect 3012 26086 3014 26138
rect 3194 26086 3196 26138
rect 2950 26084 2956 26086
rect 3012 26084 3036 26086
rect 3092 26084 3116 26086
rect 3172 26084 3196 26086
rect 3252 26084 3258 26086
rect 2950 26075 3258 26084
rect 2700 25622 2820 25650
rect 2792 25498 2820 25622
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2950 25052 3258 25061
rect 2950 25050 2956 25052
rect 3012 25050 3036 25052
rect 3092 25050 3116 25052
rect 3172 25050 3196 25052
rect 3252 25050 3258 25052
rect 3012 24998 3014 25050
rect 3194 24998 3196 25050
rect 2950 24996 2956 24998
rect 3012 24996 3036 24998
rect 3092 24996 3116 24998
rect 3172 24996 3196 24998
rect 3252 24996 3258 24998
rect 2950 24987 3258 24996
rect 2596 24200 2648 24206
rect 2596 24142 2648 24148
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2884 22710 2912 24074
rect 2950 23964 3258 23973
rect 2950 23962 2956 23964
rect 3012 23962 3036 23964
rect 3092 23962 3116 23964
rect 3172 23962 3196 23964
rect 3252 23962 3258 23964
rect 3012 23910 3014 23962
rect 3194 23910 3196 23962
rect 2950 23908 2956 23910
rect 3012 23908 3036 23910
rect 3092 23908 3116 23910
rect 3172 23908 3196 23910
rect 3252 23908 3258 23910
rect 2950 23899 3258 23908
rect 3344 23610 3372 27610
rect 3252 23582 3372 23610
rect 3252 23322 3280 23582
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 2950 22876 3258 22885
rect 2950 22874 2956 22876
rect 3012 22874 3036 22876
rect 3092 22874 3116 22876
rect 3172 22874 3196 22876
rect 3252 22874 3258 22876
rect 3012 22822 3014 22874
rect 3194 22822 3196 22874
rect 2950 22820 2956 22822
rect 3012 22820 3036 22822
rect 3092 22820 3116 22822
rect 3172 22820 3196 22822
rect 3252 22820 3258 22822
rect 2950 22811 3258 22820
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 3068 22094 3096 22714
rect 2884 22066 3096 22094
rect 2884 21978 2912 22066
rect 2608 21950 2912 21978
rect 2608 18358 2636 21950
rect 2950 21788 3258 21797
rect 2950 21786 2956 21788
rect 3012 21786 3036 21788
rect 3092 21786 3116 21788
rect 3172 21786 3196 21788
rect 3252 21786 3258 21788
rect 3012 21734 3014 21786
rect 3194 21734 3196 21786
rect 2950 21732 2956 21734
rect 3012 21732 3036 21734
rect 3092 21732 3116 21734
rect 3172 21732 3196 21734
rect 3252 21732 3258 21734
rect 2950 21723 3258 21732
rect 2950 20700 3258 20709
rect 2950 20698 2956 20700
rect 3012 20698 3036 20700
rect 3092 20698 3116 20700
rect 3172 20698 3196 20700
rect 3252 20698 3258 20700
rect 3012 20646 3014 20698
rect 3194 20646 3196 20698
rect 2950 20644 2956 20646
rect 3012 20644 3036 20646
rect 3092 20644 3116 20646
rect 3172 20644 3196 20646
rect 3252 20644 3258 20646
rect 2950 20635 3258 20644
rect 2950 19612 3258 19621
rect 2950 19610 2956 19612
rect 3012 19610 3036 19612
rect 3092 19610 3116 19612
rect 3172 19610 3196 19612
rect 3252 19610 3258 19612
rect 3012 19558 3014 19610
rect 3194 19558 3196 19610
rect 2950 19556 2956 19558
rect 3012 19556 3036 19558
rect 3092 19556 3116 19558
rect 3172 19556 3196 19558
rect 3252 19556 3258 19558
rect 2950 19547 3258 19556
rect 2950 18524 3258 18533
rect 2950 18522 2956 18524
rect 3012 18522 3036 18524
rect 3092 18522 3116 18524
rect 3172 18522 3196 18524
rect 3252 18522 3258 18524
rect 3012 18470 3014 18522
rect 3194 18470 3196 18522
rect 2950 18468 2956 18470
rect 3012 18468 3036 18470
rect 3092 18468 3116 18470
rect 3172 18468 3196 18470
rect 3252 18468 3258 18470
rect 2950 18459 3258 18468
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2950 17436 3258 17445
rect 2950 17434 2956 17436
rect 3012 17434 3036 17436
rect 3092 17434 3116 17436
rect 3172 17434 3196 17436
rect 3252 17434 3258 17436
rect 3012 17382 3014 17434
rect 3194 17382 3196 17434
rect 2950 17380 2956 17382
rect 3012 17380 3036 17382
rect 3092 17380 3116 17382
rect 3172 17380 3196 17382
rect 3252 17380 3258 17382
rect 2950 17371 3258 17380
rect 2950 16348 3258 16357
rect 2950 16346 2956 16348
rect 3012 16346 3036 16348
rect 3092 16346 3116 16348
rect 3172 16346 3196 16348
rect 3252 16346 3258 16348
rect 3012 16294 3014 16346
rect 3194 16294 3196 16346
rect 2950 16292 2956 16294
rect 3012 16292 3036 16294
rect 3092 16292 3116 16294
rect 3172 16292 3196 16294
rect 3252 16292 3258 16294
rect 2950 16283 3258 16292
rect 2950 15260 3258 15269
rect 2950 15258 2956 15260
rect 3012 15258 3036 15260
rect 3092 15258 3116 15260
rect 3172 15258 3196 15260
rect 3252 15258 3258 15260
rect 3012 15206 3014 15258
rect 3194 15206 3196 15258
rect 2950 15204 2956 15206
rect 3012 15204 3036 15206
rect 3092 15204 3116 15206
rect 3172 15204 3196 15206
rect 3252 15204 3258 15206
rect 2950 15195 3258 15204
rect 2950 14172 3258 14181
rect 2950 14170 2956 14172
rect 3012 14170 3036 14172
rect 3092 14170 3116 14172
rect 3172 14170 3196 14172
rect 3252 14170 3258 14172
rect 3012 14118 3014 14170
rect 3194 14118 3196 14170
rect 2950 14116 2956 14118
rect 3012 14116 3036 14118
rect 3092 14116 3116 14118
rect 3172 14116 3196 14118
rect 3252 14116 3258 14118
rect 2950 14107 3258 14116
rect 2950 13084 3258 13093
rect 2950 13082 2956 13084
rect 3012 13082 3036 13084
rect 3092 13082 3116 13084
rect 3172 13082 3196 13084
rect 3252 13082 3258 13084
rect 3012 13030 3014 13082
rect 3194 13030 3196 13082
rect 2950 13028 2956 13030
rect 3012 13028 3036 13030
rect 3092 13028 3116 13030
rect 3172 13028 3196 13030
rect 3252 13028 3258 13030
rect 2950 13019 3258 13028
rect 2950 11996 3258 12005
rect 2950 11994 2956 11996
rect 3012 11994 3036 11996
rect 3092 11994 3116 11996
rect 3172 11994 3196 11996
rect 3252 11994 3258 11996
rect 3012 11942 3014 11994
rect 3194 11942 3196 11994
rect 2950 11940 2956 11942
rect 3012 11940 3036 11942
rect 3092 11940 3116 11942
rect 3172 11940 3196 11942
rect 3252 11940 3258 11942
rect 2950 11931 3258 11940
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2950 10908 3258 10917
rect 2950 10906 2956 10908
rect 3012 10906 3036 10908
rect 3092 10906 3116 10908
rect 3172 10906 3196 10908
rect 3252 10906 3258 10908
rect 3012 10854 3014 10906
rect 3194 10854 3196 10906
rect 2950 10852 2956 10854
rect 3012 10852 3036 10854
rect 3092 10852 3116 10854
rect 3172 10852 3196 10854
rect 3252 10852 3258 10854
rect 2950 10843 3258 10852
rect 2950 9820 3258 9829
rect 2950 9818 2956 9820
rect 3012 9818 3036 9820
rect 3092 9818 3116 9820
rect 3172 9818 3196 9820
rect 3252 9818 3258 9820
rect 3012 9766 3014 9818
rect 3194 9766 3196 9818
rect 2950 9764 2956 9766
rect 3012 9764 3036 9766
rect 3092 9764 3116 9766
rect 3172 9764 3196 9766
rect 3252 9764 3258 9766
rect 2950 9755 3258 9764
rect 2950 8732 3258 8741
rect 2950 8730 2956 8732
rect 3012 8730 3036 8732
rect 3092 8730 3116 8732
rect 3172 8730 3196 8732
rect 3252 8730 3258 8732
rect 3012 8678 3014 8730
rect 3194 8678 3196 8730
rect 2950 8676 2956 8678
rect 3012 8676 3036 8678
rect 3092 8676 3116 8678
rect 3172 8676 3196 8678
rect 3252 8676 3258 8678
rect 2950 8667 3258 8676
rect 2950 7644 3258 7653
rect 2950 7642 2956 7644
rect 3012 7642 3036 7644
rect 3092 7642 3116 7644
rect 3172 7642 3196 7644
rect 3252 7642 3258 7644
rect 3012 7590 3014 7642
rect 3194 7590 3196 7642
rect 2950 7588 2956 7590
rect 3012 7588 3036 7590
rect 3092 7588 3116 7590
rect 3172 7588 3196 7590
rect 3252 7588 3258 7590
rect 2950 7579 3258 7588
rect 3344 7478 3372 23462
rect 3436 18834 3464 87314
rect 11336 87304 11388 87310
rect 11336 87246 11388 87252
rect 9036 87168 9088 87174
rect 9036 87110 9088 87116
rect 4896 86828 4948 86834
rect 4896 86770 4948 86776
rect 3610 86524 3918 86533
rect 3610 86522 3616 86524
rect 3672 86522 3696 86524
rect 3752 86522 3776 86524
rect 3832 86522 3856 86524
rect 3912 86522 3918 86524
rect 3672 86470 3674 86522
rect 3854 86470 3856 86522
rect 3610 86468 3616 86470
rect 3672 86468 3696 86470
rect 3752 86468 3776 86470
rect 3832 86468 3856 86470
rect 3912 86468 3918 86470
rect 3610 86459 3918 86468
rect 4344 86284 4396 86290
rect 4344 86226 4396 86232
rect 3610 85436 3918 85445
rect 3610 85434 3616 85436
rect 3672 85434 3696 85436
rect 3752 85434 3776 85436
rect 3832 85434 3856 85436
rect 3912 85434 3918 85436
rect 3672 85382 3674 85434
rect 3854 85382 3856 85434
rect 3610 85380 3616 85382
rect 3672 85380 3696 85382
rect 3752 85380 3776 85382
rect 3832 85380 3856 85382
rect 3912 85380 3918 85382
rect 3610 85371 3918 85380
rect 4160 84652 4212 84658
rect 4160 84594 4212 84600
rect 3610 84348 3918 84357
rect 3610 84346 3616 84348
rect 3672 84346 3696 84348
rect 3752 84346 3776 84348
rect 3832 84346 3856 84348
rect 3912 84346 3918 84348
rect 3672 84294 3674 84346
rect 3854 84294 3856 84346
rect 3610 84292 3616 84294
rect 3672 84292 3696 84294
rect 3752 84292 3776 84294
rect 3832 84292 3856 84294
rect 3912 84292 3918 84294
rect 3610 84283 3918 84292
rect 3976 83428 4028 83434
rect 3976 83370 4028 83376
rect 3610 83260 3918 83269
rect 3610 83258 3616 83260
rect 3672 83258 3696 83260
rect 3752 83258 3776 83260
rect 3832 83258 3856 83260
rect 3912 83258 3918 83260
rect 3672 83206 3674 83258
rect 3854 83206 3856 83258
rect 3610 83204 3616 83206
rect 3672 83204 3696 83206
rect 3752 83204 3776 83206
rect 3832 83204 3856 83206
rect 3912 83204 3918 83206
rect 3610 83195 3918 83204
rect 3610 82172 3918 82181
rect 3610 82170 3616 82172
rect 3672 82170 3696 82172
rect 3752 82170 3776 82172
rect 3832 82170 3856 82172
rect 3912 82170 3918 82172
rect 3672 82118 3674 82170
rect 3854 82118 3856 82170
rect 3610 82116 3616 82118
rect 3672 82116 3696 82118
rect 3752 82116 3776 82118
rect 3832 82116 3856 82118
rect 3912 82116 3918 82118
rect 3610 82107 3918 82116
rect 3610 81084 3918 81093
rect 3610 81082 3616 81084
rect 3672 81082 3696 81084
rect 3752 81082 3776 81084
rect 3832 81082 3856 81084
rect 3912 81082 3918 81084
rect 3672 81030 3674 81082
rect 3854 81030 3856 81082
rect 3610 81028 3616 81030
rect 3672 81028 3696 81030
rect 3752 81028 3776 81030
rect 3832 81028 3856 81030
rect 3912 81028 3918 81030
rect 3610 81019 3918 81028
rect 3610 79996 3918 80005
rect 3610 79994 3616 79996
rect 3672 79994 3696 79996
rect 3752 79994 3776 79996
rect 3832 79994 3856 79996
rect 3912 79994 3918 79996
rect 3672 79942 3674 79994
rect 3854 79942 3856 79994
rect 3610 79940 3616 79942
rect 3672 79940 3696 79942
rect 3752 79940 3776 79942
rect 3832 79940 3856 79942
rect 3912 79940 3918 79942
rect 3610 79931 3918 79940
rect 3610 78908 3918 78917
rect 3610 78906 3616 78908
rect 3672 78906 3696 78908
rect 3752 78906 3776 78908
rect 3832 78906 3856 78908
rect 3912 78906 3918 78908
rect 3672 78854 3674 78906
rect 3854 78854 3856 78906
rect 3610 78852 3616 78854
rect 3672 78852 3696 78854
rect 3752 78852 3776 78854
rect 3832 78852 3856 78854
rect 3912 78852 3918 78854
rect 3610 78843 3918 78852
rect 3610 77820 3918 77829
rect 3610 77818 3616 77820
rect 3672 77818 3696 77820
rect 3752 77818 3776 77820
rect 3832 77818 3856 77820
rect 3912 77818 3918 77820
rect 3672 77766 3674 77818
rect 3854 77766 3856 77818
rect 3610 77764 3616 77766
rect 3672 77764 3696 77766
rect 3752 77764 3776 77766
rect 3832 77764 3856 77766
rect 3912 77764 3918 77766
rect 3610 77755 3918 77764
rect 3610 76732 3918 76741
rect 3610 76730 3616 76732
rect 3672 76730 3696 76732
rect 3752 76730 3776 76732
rect 3832 76730 3856 76732
rect 3912 76730 3918 76732
rect 3672 76678 3674 76730
rect 3854 76678 3856 76730
rect 3610 76676 3616 76678
rect 3672 76676 3696 76678
rect 3752 76676 3776 76678
rect 3832 76676 3856 76678
rect 3912 76676 3918 76678
rect 3610 76667 3918 76676
rect 3610 75644 3918 75653
rect 3610 75642 3616 75644
rect 3672 75642 3696 75644
rect 3752 75642 3776 75644
rect 3832 75642 3856 75644
rect 3912 75642 3918 75644
rect 3672 75590 3674 75642
rect 3854 75590 3856 75642
rect 3610 75588 3616 75590
rect 3672 75588 3696 75590
rect 3752 75588 3776 75590
rect 3832 75588 3856 75590
rect 3912 75588 3918 75590
rect 3610 75579 3918 75588
rect 3610 74556 3918 74565
rect 3610 74554 3616 74556
rect 3672 74554 3696 74556
rect 3752 74554 3776 74556
rect 3832 74554 3856 74556
rect 3912 74554 3918 74556
rect 3672 74502 3674 74554
rect 3854 74502 3856 74554
rect 3610 74500 3616 74502
rect 3672 74500 3696 74502
rect 3752 74500 3776 74502
rect 3832 74500 3856 74502
rect 3912 74500 3918 74502
rect 3610 74491 3918 74500
rect 3516 73908 3568 73914
rect 3516 73850 3568 73856
rect 3528 70854 3556 73850
rect 3610 73468 3918 73477
rect 3610 73466 3616 73468
rect 3672 73466 3696 73468
rect 3752 73466 3776 73468
rect 3832 73466 3856 73468
rect 3912 73466 3918 73468
rect 3672 73414 3674 73466
rect 3854 73414 3856 73466
rect 3610 73412 3616 73414
rect 3672 73412 3696 73414
rect 3752 73412 3776 73414
rect 3832 73412 3856 73414
rect 3912 73412 3918 73414
rect 3610 73403 3918 73412
rect 3610 72380 3918 72389
rect 3610 72378 3616 72380
rect 3672 72378 3696 72380
rect 3752 72378 3776 72380
rect 3832 72378 3856 72380
rect 3912 72378 3918 72380
rect 3672 72326 3674 72378
rect 3854 72326 3856 72378
rect 3610 72324 3616 72326
rect 3672 72324 3696 72326
rect 3752 72324 3776 72326
rect 3832 72324 3856 72326
rect 3912 72324 3918 72326
rect 3610 72315 3918 72324
rect 3610 71292 3918 71301
rect 3610 71290 3616 71292
rect 3672 71290 3696 71292
rect 3752 71290 3776 71292
rect 3832 71290 3856 71292
rect 3912 71290 3918 71292
rect 3672 71238 3674 71290
rect 3854 71238 3856 71290
rect 3610 71236 3616 71238
rect 3672 71236 3696 71238
rect 3752 71236 3776 71238
rect 3832 71236 3856 71238
rect 3912 71236 3918 71238
rect 3610 71227 3918 71236
rect 3516 70848 3568 70854
rect 3516 70790 3568 70796
rect 3516 70508 3568 70514
rect 3516 70450 3568 70456
rect 3528 65550 3556 70450
rect 3610 70204 3918 70213
rect 3610 70202 3616 70204
rect 3672 70202 3696 70204
rect 3752 70202 3776 70204
rect 3832 70202 3856 70204
rect 3912 70202 3918 70204
rect 3672 70150 3674 70202
rect 3854 70150 3856 70202
rect 3610 70148 3616 70150
rect 3672 70148 3696 70150
rect 3752 70148 3776 70150
rect 3832 70148 3856 70150
rect 3912 70148 3918 70150
rect 3610 70139 3918 70148
rect 3610 69116 3918 69125
rect 3610 69114 3616 69116
rect 3672 69114 3696 69116
rect 3752 69114 3776 69116
rect 3832 69114 3856 69116
rect 3912 69114 3918 69116
rect 3672 69062 3674 69114
rect 3854 69062 3856 69114
rect 3610 69060 3616 69062
rect 3672 69060 3696 69062
rect 3752 69060 3776 69062
rect 3832 69060 3856 69062
rect 3912 69060 3918 69062
rect 3610 69051 3918 69060
rect 3884 68876 3936 68882
rect 3884 68818 3936 68824
rect 3896 68134 3924 68818
rect 3884 68128 3936 68134
rect 3884 68070 3936 68076
rect 3610 68028 3918 68037
rect 3610 68026 3616 68028
rect 3672 68026 3696 68028
rect 3752 68026 3776 68028
rect 3832 68026 3856 68028
rect 3912 68026 3918 68028
rect 3672 67974 3674 68026
rect 3854 67974 3856 68026
rect 3610 67972 3616 67974
rect 3672 67972 3696 67974
rect 3752 67972 3776 67974
rect 3832 67972 3856 67974
rect 3912 67972 3918 67974
rect 3610 67963 3918 67972
rect 3882 67824 3938 67833
rect 3882 67759 3938 67768
rect 3896 67250 3924 67759
rect 3884 67244 3936 67250
rect 3884 67186 3936 67192
rect 3610 66940 3918 66949
rect 3610 66938 3616 66940
rect 3672 66938 3696 66940
rect 3752 66938 3776 66940
rect 3832 66938 3856 66940
rect 3912 66938 3918 66940
rect 3672 66886 3674 66938
rect 3854 66886 3856 66938
rect 3610 66884 3616 66886
rect 3672 66884 3696 66886
rect 3752 66884 3776 66886
rect 3832 66884 3856 66886
rect 3912 66884 3918 66886
rect 3610 66875 3918 66884
rect 3988 66638 4016 83370
rect 4172 80054 4200 84594
rect 4172 80026 4292 80054
rect 4160 79552 4212 79558
rect 4160 79494 4212 79500
rect 4068 75812 4120 75818
rect 4068 75754 4120 75760
rect 3976 66632 4028 66638
rect 3976 66574 4028 66580
rect 3976 66020 4028 66026
rect 3976 65962 4028 65968
rect 3610 65852 3918 65861
rect 3610 65850 3616 65852
rect 3672 65850 3696 65852
rect 3752 65850 3776 65852
rect 3832 65850 3856 65852
rect 3912 65850 3918 65852
rect 3672 65798 3674 65850
rect 3854 65798 3856 65850
rect 3610 65796 3616 65798
rect 3672 65796 3696 65798
rect 3752 65796 3776 65798
rect 3832 65796 3856 65798
rect 3912 65796 3918 65798
rect 3610 65787 3918 65796
rect 3608 65680 3660 65686
rect 3608 65622 3660 65628
rect 3516 65544 3568 65550
rect 3516 65486 3568 65492
rect 3620 65362 3648 65622
rect 3528 65334 3648 65362
rect 3528 56846 3556 65334
rect 3610 64764 3918 64773
rect 3610 64762 3616 64764
rect 3672 64762 3696 64764
rect 3752 64762 3776 64764
rect 3832 64762 3856 64764
rect 3912 64762 3918 64764
rect 3672 64710 3674 64762
rect 3854 64710 3856 64762
rect 3610 64708 3616 64710
rect 3672 64708 3696 64710
rect 3752 64708 3776 64710
rect 3832 64708 3856 64710
rect 3912 64708 3918 64710
rect 3610 64699 3918 64708
rect 3610 63676 3918 63685
rect 3610 63674 3616 63676
rect 3672 63674 3696 63676
rect 3752 63674 3776 63676
rect 3832 63674 3856 63676
rect 3912 63674 3918 63676
rect 3672 63622 3674 63674
rect 3854 63622 3856 63674
rect 3610 63620 3616 63622
rect 3672 63620 3696 63622
rect 3752 63620 3776 63622
rect 3832 63620 3856 63622
rect 3912 63620 3918 63622
rect 3610 63611 3918 63620
rect 3608 63436 3660 63442
rect 3608 63378 3660 63384
rect 3620 62937 3648 63378
rect 3606 62928 3662 62937
rect 3606 62863 3662 62872
rect 3610 62588 3918 62597
rect 3610 62586 3616 62588
rect 3672 62586 3696 62588
rect 3752 62586 3776 62588
rect 3832 62586 3856 62588
rect 3912 62586 3918 62588
rect 3672 62534 3674 62586
rect 3854 62534 3856 62586
rect 3610 62532 3616 62534
rect 3672 62532 3696 62534
rect 3752 62532 3776 62534
rect 3832 62532 3856 62534
rect 3912 62532 3918 62534
rect 3610 62523 3918 62532
rect 3610 61500 3918 61509
rect 3610 61498 3616 61500
rect 3672 61498 3696 61500
rect 3752 61498 3776 61500
rect 3832 61498 3856 61500
rect 3912 61498 3918 61500
rect 3672 61446 3674 61498
rect 3854 61446 3856 61498
rect 3610 61444 3616 61446
rect 3672 61444 3696 61446
rect 3752 61444 3776 61446
rect 3832 61444 3856 61446
rect 3912 61444 3918 61446
rect 3610 61435 3918 61444
rect 3610 60412 3918 60421
rect 3610 60410 3616 60412
rect 3672 60410 3696 60412
rect 3752 60410 3776 60412
rect 3832 60410 3856 60412
rect 3912 60410 3918 60412
rect 3672 60358 3674 60410
rect 3854 60358 3856 60410
rect 3610 60356 3616 60358
rect 3672 60356 3696 60358
rect 3752 60356 3776 60358
rect 3832 60356 3856 60358
rect 3912 60356 3918 60358
rect 3610 60347 3918 60356
rect 3884 60172 3936 60178
rect 3884 60114 3936 60120
rect 3896 59514 3924 60114
rect 3988 59634 4016 65962
rect 3976 59628 4028 59634
rect 3976 59570 4028 59576
rect 3896 59486 4016 59514
rect 3610 59324 3918 59333
rect 3610 59322 3616 59324
rect 3672 59322 3696 59324
rect 3752 59322 3776 59324
rect 3832 59322 3856 59324
rect 3912 59322 3918 59324
rect 3672 59270 3674 59322
rect 3854 59270 3856 59322
rect 3610 59268 3616 59270
rect 3672 59268 3696 59270
rect 3752 59268 3776 59270
rect 3832 59268 3856 59270
rect 3912 59268 3918 59270
rect 3610 59259 3918 59268
rect 3610 58236 3918 58245
rect 3610 58234 3616 58236
rect 3672 58234 3696 58236
rect 3752 58234 3776 58236
rect 3832 58234 3856 58236
rect 3912 58234 3918 58236
rect 3672 58182 3674 58234
rect 3854 58182 3856 58234
rect 3610 58180 3616 58182
rect 3672 58180 3696 58182
rect 3752 58180 3776 58182
rect 3832 58180 3856 58182
rect 3912 58180 3918 58182
rect 3610 58171 3918 58180
rect 3610 57148 3918 57157
rect 3610 57146 3616 57148
rect 3672 57146 3696 57148
rect 3752 57146 3776 57148
rect 3832 57146 3856 57148
rect 3912 57146 3918 57148
rect 3672 57094 3674 57146
rect 3854 57094 3856 57146
rect 3610 57092 3616 57094
rect 3672 57092 3696 57094
rect 3752 57092 3776 57094
rect 3832 57092 3856 57094
rect 3912 57092 3918 57094
rect 3610 57083 3918 57092
rect 3516 56840 3568 56846
rect 3516 56782 3568 56788
rect 3516 56704 3568 56710
rect 3516 56646 3568 56652
rect 3528 56302 3556 56646
rect 3516 56296 3568 56302
rect 3516 56238 3568 56244
rect 3610 56060 3918 56069
rect 3610 56058 3616 56060
rect 3672 56058 3696 56060
rect 3752 56058 3776 56060
rect 3832 56058 3856 56060
rect 3912 56058 3918 56060
rect 3672 56006 3674 56058
rect 3854 56006 3856 56058
rect 3610 56004 3616 56006
rect 3672 56004 3696 56006
rect 3752 56004 3776 56006
rect 3832 56004 3856 56006
rect 3912 56004 3918 56006
rect 3610 55995 3918 56004
rect 3610 54972 3918 54981
rect 3610 54970 3616 54972
rect 3672 54970 3696 54972
rect 3752 54970 3776 54972
rect 3832 54970 3856 54972
rect 3912 54970 3918 54972
rect 3672 54918 3674 54970
rect 3854 54918 3856 54970
rect 3610 54916 3616 54918
rect 3672 54916 3696 54918
rect 3752 54916 3776 54918
rect 3832 54916 3856 54918
rect 3912 54916 3918 54918
rect 3610 54907 3918 54916
rect 3610 53884 3918 53893
rect 3610 53882 3616 53884
rect 3672 53882 3696 53884
rect 3752 53882 3776 53884
rect 3832 53882 3856 53884
rect 3912 53882 3918 53884
rect 3672 53830 3674 53882
rect 3854 53830 3856 53882
rect 3610 53828 3616 53830
rect 3672 53828 3696 53830
rect 3752 53828 3776 53830
rect 3832 53828 3856 53830
rect 3912 53828 3918 53830
rect 3610 53819 3918 53828
rect 3988 53666 4016 59486
rect 3804 53638 4016 53666
rect 3516 53440 3568 53446
rect 3516 53382 3568 53388
rect 3528 44826 3556 53382
rect 3804 52970 3832 53638
rect 3976 53508 4028 53514
rect 3976 53450 4028 53456
rect 3792 52964 3844 52970
rect 3792 52906 3844 52912
rect 3610 52796 3918 52805
rect 3610 52794 3616 52796
rect 3672 52794 3696 52796
rect 3752 52794 3776 52796
rect 3832 52794 3856 52796
rect 3912 52794 3918 52796
rect 3672 52742 3674 52794
rect 3854 52742 3856 52794
rect 3610 52740 3616 52742
rect 3672 52740 3696 52742
rect 3752 52740 3776 52742
rect 3832 52740 3856 52742
rect 3912 52740 3918 52742
rect 3610 52731 3918 52740
rect 3610 51708 3918 51717
rect 3610 51706 3616 51708
rect 3672 51706 3696 51708
rect 3752 51706 3776 51708
rect 3832 51706 3856 51708
rect 3912 51706 3918 51708
rect 3672 51654 3674 51706
rect 3854 51654 3856 51706
rect 3610 51652 3616 51654
rect 3672 51652 3696 51654
rect 3752 51652 3776 51654
rect 3832 51652 3856 51654
rect 3912 51652 3918 51654
rect 3610 51643 3918 51652
rect 3610 50620 3918 50629
rect 3610 50618 3616 50620
rect 3672 50618 3696 50620
rect 3752 50618 3776 50620
rect 3832 50618 3856 50620
rect 3912 50618 3918 50620
rect 3672 50566 3674 50618
rect 3854 50566 3856 50618
rect 3610 50564 3616 50566
rect 3672 50564 3696 50566
rect 3752 50564 3776 50566
rect 3832 50564 3856 50566
rect 3912 50564 3918 50566
rect 3610 50555 3918 50564
rect 3792 50244 3844 50250
rect 3792 50186 3844 50192
rect 3804 49910 3832 50186
rect 3792 49904 3844 49910
rect 3792 49846 3844 49852
rect 3610 49532 3918 49541
rect 3610 49530 3616 49532
rect 3672 49530 3696 49532
rect 3752 49530 3776 49532
rect 3832 49530 3856 49532
rect 3912 49530 3918 49532
rect 3672 49478 3674 49530
rect 3854 49478 3856 49530
rect 3610 49476 3616 49478
rect 3672 49476 3696 49478
rect 3752 49476 3776 49478
rect 3832 49476 3856 49478
rect 3912 49476 3918 49478
rect 3610 49467 3918 49476
rect 3610 48444 3918 48453
rect 3610 48442 3616 48444
rect 3672 48442 3696 48444
rect 3752 48442 3776 48444
rect 3832 48442 3856 48444
rect 3912 48442 3918 48444
rect 3672 48390 3674 48442
rect 3854 48390 3856 48442
rect 3610 48388 3616 48390
rect 3672 48388 3696 48390
rect 3752 48388 3776 48390
rect 3832 48388 3856 48390
rect 3912 48388 3918 48390
rect 3610 48379 3918 48388
rect 3610 47356 3918 47365
rect 3610 47354 3616 47356
rect 3672 47354 3696 47356
rect 3752 47354 3776 47356
rect 3832 47354 3856 47356
rect 3912 47354 3918 47356
rect 3672 47302 3674 47354
rect 3854 47302 3856 47354
rect 3610 47300 3616 47302
rect 3672 47300 3696 47302
rect 3752 47300 3776 47302
rect 3832 47300 3856 47302
rect 3912 47300 3918 47302
rect 3610 47291 3918 47300
rect 3610 46268 3918 46277
rect 3610 46266 3616 46268
rect 3672 46266 3696 46268
rect 3752 46266 3776 46268
rect 3832 46266 3856 46268
rect 3912 46266 3918 46268
rect 3672 46214 3674 46266
rect 3854 46214 3856 46266
rect 3610 46212 3616 46214
rect 3672 46212 3696 46214
rect 3752 46212 3776 46214
rect 3832 46212 3856 46214
rect 3912 46212 3918 46214
rect 3610 46203 3918 46212
rect 3610 45180 3918 45189
rect 3610 45178 3616 45180
rect 3672 45178 3696 45180
rect 3752 45178 3776 45180
rect 3832 45178 3856 45180
rect 3912 45178 3918 45180
rect 3672 45126 3674 45178
rect 3854 45126 3856 45178
rect 3610 45124 3616 45126
rect 3672 45124 3696 45126
rect 3752 45124 3776 45126
rect 3832 45124 3856 45126
rect 3912 45124 3918 45126
rect 3610 45115 3918 45124
rect 3988 44985 4016 53450
rect 4080 45529 4108 75754
rect 4172 68921 4200 79494
rect 4264 75002 4292 80026
rect 4252 74996 4304 75002
rect 4252 74938 4304 74944
rect 4356 73098 4384 86226
rect 4550 85980 4858 85989
rect 4550 85978 4556 85980
rect 4612 85978 4636 85980
rect 4692 85978 4716 85980
rect 4772 85978 4796 85980
rect 4852 85978 4858 85980
rect 4612 85926 4614 85978
rect 4794 85926 4796 85978
rect 4550 85924 4556 85926
rect 4612 85924 4636 85926
rect 4692 85924 4716 85926
rect 4772 85924 4796 85926
rect 4852 85924 4858 85926
rect 4550 85915 4858 85924
rect 4436 85876 4488 85882
rect 4436 85818 4488 85824
rect 4448 75410 4476 85818
rect 4550 84892 4858 84901
rect 4550 84890 4556 84892
rect 4612 84890 4636 84892
rect 4692 84890 4716 84892
rect 4772 84890 4796 84892
rect 4852 84890 4858 84892
rect 4612 84838 4614 84890
rect 4794 84838 4796 84890
rect 4550 84836 4556 84838
rect 4612 84836 4636 84838
rect 4692 84836 4716 84838
rect 4772 84836 4796 84838
rect 4852 84836 4858 84838
rect 4550 84827 4858 84836
rect 4550 83804 4858 83813
rect 4550 83802 4556 83804
rect 4612 83802 4636 83804
rect 4692 83802 4716 83804
rect 4772 83802 4796 83804
rect 4852 83802 4858 83804
rect 4612 83750 4614 83802
rect 4794 83750 4796 83802
rect 4550 83748 4556 83750
rect 4612 83748 4636 83750
rect 4692 83748 4716 83750
rect 4772 83748 4796 83750
rect 4852 83748 4858 83750
rect 4550 83739 4858 83748
rect 4550 82716 4858 82725
rect 4550 82714 4556 82716
rect 4612 82714 4636 82716
rect 4692 82714 4716 82716
rect 4772 82714 4796 82716
rect 4852 82714 4858 82716
rect 4612 82662 4614 82714
rect 4794 82662 4796 82714
rect 4550 82660 4556 82662
rect 4612 82660 4636 82662
rect 4692 82660 4716 82662
rect 4772 82660 4796 82662
rect 4852 82660 4858 82662
rect 4550 82651 4858 82660
rect 4550 81628 4858 81637
rect 4550 81626 4556 81628
rect 4612 81626 4636 81628
rect 4692 81626 4716 81628
rect 4772 81626 4796 81628
rect 4852 81626 4858 81628
rect 4612 81574 4614 81626
rect 4794 81574 4796 81626
rect 4550 81572 4556 81574
rect 4612 81572 4636 81574
rect 4692 81572 4716 81574
rect 4772 81572 4796 81574
rect 4852 81572 4858 81574
rect 4550 81563 4858 81572
rect 4550 80540 4858 80549
rect 4550 80538 4556 80540
rect 4612 80538 4636 80540
rect 4692 80538 4716 80540
rect 4772 80538 4796 80540
rect 4852 80538 4858 80540
rect 4612 80486 4614 80538
rect 4794 80486 4796 80538
rect 4550 80484 4556 80486
rect 4612 80484 4636 80486
rect 4692 80484 4716 80486
rect 4772 80484 4796 80486
rect 4852 80484 4858 80486
rect 4550 80475 4858 80484
rect 4550 79452 4858 79461
rect 4550 79450 4556 79452
rect 4612 79450 4636 79452
rect 4692 79450 4716 79452
rect 4772 79450 4796 79452
rect 4852 79450 4858 79452
rect 4612 79398 4614 79450
rect 4794 79398 4796 79450
rect 4550 79396 4556 79398
rect 4612 79396 4636 79398
rect 4692 79396 4716 79398
rect 4772 79396 4796 79398
rect 4852 79396 4858 79398
rect 4550 79387 4858 79396
rect 4550 78364 4858 78373
rect 4550 78362 4556 78364
rect 4612 78362 4636 78364
rect 4692 78362 4716 78364
rect 4772 78362 4796 78364
rect 4852 78362 4858 78364
rect 4612 78310 4614 78362
rect 4794 78310 4796 78362
rect 4550 78308 4556 78310
rect 4612 78308 4636 78310
rect 4692 78308 4716 78310
rect 4772 78308 4796 78310
rect 4852 78308 4858 78310
rect 4550 78299 4858 78308
rect 4550 77276 4858 77285
rect 4550 77274 4556 77276
rect 4612 77274 4636 77276
rect 4692 77274 4716 77276
rect 4772 77274 4796 77276
rect 4852 77274 4858 77276
rect 4612 77222 4614 77274
rect 4794 77222 4796 77274
rect 4550 77220 4556 77222
rect 4612 77220 4636 77222
rect 4692 77220 4716 77222
rect 4772 77220 4796 77222
rect 4852 77220 4858 77222
rect 4550 77211 4858 77220
rect 4550 76188 4858 76197
rect 4550 76186 4556 76188
rect 4612 76186 4636 76188
rect 4692 76186 4716 76188
rect 4772 76186 4796 76188
rect 4852 76186 4858 76188
rect 4612 76134 4614 76186
rect 4794 76134 4796 76186
rect 4550 76132 4556 76134
rect 4612 76132 4636 76134
rect 4692 76132 4716 76134
rect 4772 76132 4796 76134
rect 4852 76132 4858 76134
rect 4550 76123 4858 76132
rect 4436 75404 4488 75410
rect 4436 75346 4488 75352
rect 4908 75206 4936 86770
rect 5540 86760 5592 86766
rect 5540 86702 5592 86708
rect 5210 86524 5518 86533
rect 5210 86522 5216 86524
rect 5272 86522 5296 86524
rect 5352 86522 5376 86524
rect 5432 86522 5456 86524
rect 5512 86522 5518 86524
rect 5272 86470 5274 86522
rect 5454 86470 5456 86522
rect 5210 86468 5216 86470
rect 5272 86468 5296 86470
rect 5352 86468 5376 86470
rect 5432 86468 5456 86470
rect 5512 86468 5518 86470
rect 5210 86459 5518 86468
rect 4988 86216 5040 86222
rect 4988 86158 5040 86164
rect 5000 79558 5028 86158
rect 5210 85436 5518 85445
rect 5210 85434 5216 85436
rect 5272 85434 5296 85436
rect 5352 85434 5376 85436
rect 5432 85434 5456 85436
rect 5512 85434 5518 85436
rect 5272 85382 5274 85434
rect 5454 85382 5456 85434
rect 5210 85380 5216 85382
rect 5272 85380 5296 85382
rect 5352 85380 5376 85382
rect 5432 85380 5456 85382
rect 5512 85380 5518 85382
rect 5210 85371 5518 85380
rect 5078 85096 5134 85105
rect 5078 85031 5134 85040
rect 4988 79552 5040 79558
rect 4988 79494 5040 79500
rect 4436 75200 4488 75206
rect 4436 75142 4488 75148
rect 4896 75200 4948 75206
rect 4896 75142 4948 75148
rect 4344 73092 4396 73098
rect 4344 73034 4396 73040
rect 4252 72684 4304 72690
rect 4252 72626 4304 72632
rect 4264 69834 4292 72626
rect 4344 71732 4396 71738
rect 4344 71674 4396 71680
rect 4356 70514 4384 71674
rect 4344 70508 4396 70514
rect 4344 70450 4396 70456
rect 4448 70394 4476 75142
rect 4550 75100 4858 75109
rect 4550 75098 4556 75100
rect 4612 75098 4636 75100
rect 4692 75098 4716 75100
rect 4772 75098 4796 75100
rect 4852 75098 4858 75100
rect 4612 75046 4614 75098
rect 4794 75046 4796 75098
rect 4550 75044 4556 75046
rect 4612 75044 4636 75046
rect 4692 75044 4716 75046
rect 4772 75044 4796 75046
rect 4852 75044 4858 75046
rect 4550 75035 4858 75044
rect 4896 74996 4948 75002
rect 4896 74938 4948 74944
rect 4550 74012 4858 74021
rect 4550 74010 4556 74012
rect 4612 74010 4636 74012
rect 4692 74010 4716 74012
rect 4772 74010 4796 74012
rect 4852 74010 4858 74012
rect 4612 73958 4614 74010
rect 4794 73958 4796 74010
rect 4550 73956 4556 73958
rect 4612 73956 4636 73958
rect 4692 73956 4716 73958
rect 4772 73956 4796 73958
rect 4852 73956 4858 73958
rect 4550 73947 4858 73956
rect 4550 72924 4858 72933
rect 4550 72922 4556 72924
rect 4612 72922 4636 72924
rect 4692 72922 4716 72924
rect 4772 72922 4796 72924
rect 4852 72922 4858 72924
rect 4612 72870 4614 72922
rect 4794 72870 4796 72922
rect 4550 72868 4556 72870
rect 4612 72868 4636 72870
rect 4692 72868 4716 72870
rect 4772 72868 4796 72870
rect 4852 72868 4858 72870
rect 4550 72859 4858 72868
rect 4908 72554 4936 74938
rect 4988 73364 5040 73370
rect 4988 73306 5040 73312
rect 4896 72548 4948 72554
rect 4896 72490 4948 72496
rect 4550 71836 4858 71845
rect 4550 71834 4556 71836
rect 4612 71834 4636 71836
rect 4692 71834 4716 71836
rect 4772 71834 4796 71836
rect 4852 71834 4858 71836
rect 4612 71782 4614 71834
rect 4794 71782 4796 71834
rect 4550 71780 4556 71782
rect 4612 71780 4636 71782
rect 4692 71780 4716 71782
rect 4772 71780 4796 71782
rect 4852 71780 4858 71782
rect 4550 71771 4858 71780
rect 4896 71664 4948 71670
rect 4896 71606 4948 71612
rect 4550 70748 4858 70757
rect 4550 70746 4556 70748
rect 4612 70746 4636 70748
rect 4692 70746 4716 70748
rect 4772 70746 4796 70748
rect 4852 70746 4858 70748
rect 4612 70694 4614 70746
rect 4794 70694 4796 70746
rect 4550 70692 4556 70694
rect 4612 70692 4636 70694
rect 4692 70692 4716 70694
rect 4772 70692 4796 70694
rect 4852 70692 4858 70694
rect 4550 70683 4858 70692
rect 4710 70408 4766 70417
rect 4356 70366 4476 70394
rect 4632 70366 4710 70394
rect 4252 69828 4304 69834
rect 4252 69770 4304 69776
rect 4264 69018 4292 69770
rect 4356 69562 4384 70366
rect 4436 70304 4488 70310
rect 4436 70246 4488 70252
rect 4344 69556 4396 69562
rect 4344 69498 4396 69504
rect 4252 69012 4304 69018
rect 4252 68954 4304 68960
rect 4344 69012 4396 69018
rect 4344 68954 4396 68960
rect 4158 68912 4214 68921
rect 4356 68898 4384 68954
rect 4158 68847 4214 68856
rect 4264 68870 4384 68898
rect 4264 68762 4292 68870
rect 4172 68734 4292 68762
rect 4344 68808 4396 68814
rect 4344 68750 4396 68756
rect 4172 64870 4200 68734
rect 4252 68672 4304 68678
rect 4252 68614 4304 68620
rect 4264 67862 4292 68614
rect 4252 67856 4304 67862
rect 4356 67833 4384 68750
rect 4448 68270 4476 70246
rect 4632 69970 4660 70366
rect 4710 70343 4766 70352
rect 4712 70304 4764 70310
rect 4712 70246 4764 70252
rect 4620 69964 4672 69970
rect 4620 69906 4672 69912
rect 4724 69834 4752 70246
rect 4712 69828 4764 69834
rect 4712 69770 4764 69776
rect 4550 69660 4858 69669
rect 4550 69658 4556 69660
rect 4612 69658 4636 69660
rect 4692 69658 4716 69660
rect 4772 69658 4796 69660
rect 4852 69658 4858 69660
rect 4612 69606 4614 69658
rect 4794 69606 4796 69658
rect 4550 69604 4556 69606
rect 4612 69604 4636 69606
rect 4692 69604 4716 69606
rect 4772 69604 4796 69606
rect 4852 69604 4858 69606
rect 4550 69595 4858 69604
rect 4804 69556 4856 69562
rect 4804 69498 4856 69504
rect 4620 69216 4672 69222
rect 4620 69158 4672 69164
rect 4712 69216 4764 69222
rect 4712 69158 4764 69164
rect 4632 68678 4660 69158
rect 4724 68746 4752 69158
rect 4816 68746 4844 69498
rect 4712 68740 4764 68746
rect 4712 68682 4764 68688
rect 4804 68740 4856 68746
rect 4804 68682 4856 68688
rect 4620 68672 4672 68678
rect 4620 68614 4672 68620
rect 4550 68572 4858 68581
rect 4550 68570 4556 68572
rect 4612 68570 4636 68572
rect 4692 68570 4716 68572
rect 4772 68570 4796 68572
rect 4852 68570 4858 68572
rect 4612 68518 4614 68570
rect 4794 68518 4796 68570
rect 4550 68516 4556 68518
rect 4612 68516 4636 68518
rect 4692 68516 4716 68518
rect 4772 68516 4796 68518
rect 4852 68516 4858 68518
rect 4550 68507 4858 68516
rect 4528 68332 4580 68338
rect 4528 68274 4580 68280
rect 4804 68332 4856 68338
rect 4804 68274 4856 68280
rect 4436 68264 4488 68270
rect 4436 68206 4488 68212
rect 4436 68128 4488 68134
rect 4436 68070 4488 68076
rect 4252 67798 4304 67804
rect 4342 67824 4398 67833
rect 4264 67182 4292 67798
rect 4342 67759 4398 67768
rect 4344 67312 4396 67318
rect 4342 67280 4344 67289
rect 4396 67280 4398 67289
rect 4342 67215 4398 67224
rect 4252 67176 4304 67182
rect 4252 67118 4304 67124
rect 4264 66570 4292 67118
rect 4252 66564 4304 66570
rect 4252 66506 4304 66512
rect 4160 64864 4212 64870
rect 4160 64806 4212 64812
rect 4160 64524 4212 64530
rect 4160 64466 4212 64472
rect 4172 57594 4200 64466
rect 4264 59226 4292 66506
rect 4356 66473 4384 67215
rect 4448 66502 4476 68070
rect 4540 67697 4568 68274
rect 4618 67824 4674 67833
rect 4618 67759 4620 67768
rect 4672 67759 4674 67768
rect 4620 67730 4672 67736
rect 4526 67688 4582 67697
rect 4816 67658 4844 68274
rect 4908 68082 4936 71606
rect 5000 70106 5028 73306
rect 4988 70100 5040 70106
rect 4988 70042 5040 70048
rect 4988 69828 5040 69834
rect 4988 69770 5040 69776
rect 5000 68474 5028 69770
rect 4988 68468 5040 68474
rect 4988 68410 5040 68416
rect 5092 68406 5120 85031
rect 5210 84348 5518 84357
rect 5210 84346 5216 84348
rect 5272 84346 5296 84348
rect 5352 84346 5376 84348
rect 5432 84346 5456 84348
rect 5512 84346 5518 84348
rect 5272 84294 5274 84346
rect 5454 84294 5456 84346
rect 5210 84292 5216 84294
rect 5272 84292 5296 84294
rect 5352 84292 5376 84294
rect 5432 84292 5456 84294
rect 5512 84292 5518 84294
rect 5210 84283 5518 84292
rect 5210 83260 5518 83269
rect 5210 83258 5216 83260
rect 5272 83258 5296 83260
rect 5352 83258 5376 83260
rect 5432 83258 5456 83260
rect 5512 83258 5518 83260
rect 5272 83206 5274 83258
rect 5454 83206 5456 83258
rect 5210 83204 5216 83206
rect 5272 83204 5296 83206
rect 5352 83204 5376 83206
rect 5432 83204 5456 83206
rect 5512 83204 5518 83206
rect 5210 83195 5518 83204
rect 5210 82172 5518 82181
rect 5210 82170 5216 82172
rect 5272 82170 5296 82172
rect 5352 82170 5376 82172
rect 5432 82170 5456 82172
rect 5512 82170 5518 82172
rect 5272 82118 5274 82170
rect 5454 82118 5456 82170
rect 5210 82116 5216 82118
rect 5272 82116 5296 82118
rect 5352 82116 5376 82118
rect 5432 82116 5456 82118
rect 5512 82116 5518 82118
rect 5210 82107 5518 82116
rect 5210 81084 5518 81093
rect 5210 81082 5216 81084
rect 5272 81082 5296 81084
rect 5352 81082 5376 81084
rect 5432 81082 5456 81084
rect 5512 81082 5518 81084
rect 5272 81030 5274 81082
rect 5454 81030 5456 81082
rect 5210 81028 5216 81030
rect 5272 81028 5296 81030
rect 5352 81028 5376 81030
rect 5432 81028 5456 81030
rect 5512 81028 5518 81030
rect 5210 81019 5518 81028
rect 5210 79996 5518 80005
rect 5210 79994 5216 79996
rect 5272 79994 5296 79996
rect 5352 79994 5376 79996
rect 5432 79994 5456 79996
rect 5512 79994 5518 79996
rect 5272 79942 5274 79994
rect 5454 79942 5456 79994
rect 5210 79940 5216 79942
rect 5272 79940 5296 79942
rect 5352 79940 5376 79942
rect 5432 79940 5456 79942
rect 5512 79940 5518 79942
rect 5210 79931 5518 79940
rect 5210 78908 5518 78917
rect 5210 78906 5216 78908
rect 5272 78906 5296 78908
rect 5352 78906 5376 78908
rect 5432 78906 5456 78908
rect 5512 78906 5518 78908
rect 5272 78854 5274 78906
rect 5454 78854 5456 78906
rect 5210 78852 5216 78854
rect 5272 78852 5296 78854
rect 5352 78852 5376 78854
rect 5432 78852 5456 78854
rect 5512 78852 5518 78854
rect 5210 78843 5518 78852
rect 5210 77820 5518 77829
rect 5210 77818 5216 77820
rect 5272 77818 5296 77820
rect 5352 77818 5376 77820
rect 5432 77818 5456 77820
rect 5512 77818 5518 77820
rect 5272 77766 5274 77818
rect 5454 77766 5456 77818
rect 5210 77764 5216 77766
rect 5272 77764 5296 77766
rect 5352 77764 5376 77766
rect 5432 77764 5456 77766
rect 5512 77764 5518 77766
rect 5210 77755 5518 77764
rect 5210 76732 5518 76741
rect 5210 76730 5216 76732
rect 5272 76730 5296 76732
rect 5352 76730 5376 76732
rect 5432 76730 5456 76732
rect 5512 76730 5518 76732
rect 5272 76678 5274 76730
rect 5454 76678 5456 76730
rect 5210 76676 5216 76678
rect 5272 76676 5296 76678
rect 5352 76676 5376 76678
rect 5432 76676 5456 76678
rect 5512 76676 5518 76678
rect 5210 76667 5518 76676
rect 5210 75644 5518 75653
rect 5210 75642 5216 75644
rect 5272 75642 5296 75644
rect 5352 75642 5376 75644
rect 5432 75642 5456 75644
rect 5512 75642 5518 75644
rect 5272 75590 5274 75642
rect 5454 75590 5456 75642
rect 5210 75588 5216 75590
rect 5272 75588 5296 75590
rect 5352 75588 5376 75590
rect 5432 75588 5456 75590
rect 5512 75588 5518 75590
rect 5210 75579 5518 75588
rect 5210 74556 5518 74565
rect 5210 74554 5216 74556
rect 5272 74554 5296 74556
rect 5352 74554 5376 74556
rect 5432 74554 5456 74556
rect 5512 74554 5518 74556
rect 5272 74502 5274 74554
rect 5454 74502 5456 74554
rect 5210 74500 5216 74502
rect 5272 74500 5296 74502
rect 5352 74500 5376 74502
rect 5432 74500 5456 74502
rect 5512 74500 5518 74502
rect 5210 74491 5518 74500
rect 5210 73468 5518 73477
rect 5210 73466 5216 73468
rect 5272 73466 5296 73468
rect 5352 73466 5376 73468
rect 5432 73466 5456 73468
rect 5512 73466 5518 73468
rect 5272 73414 5274 73466
rect 5454 73414 5456 73466
rect 5210 73412 5216 73414
rect 5272 73412 5296 73414
rect 5352 73412 5376 73414
rect 5432 73412 5456 73414
rect 5512 73412 5518 73414
rect 5210 73403 5518 73412
rect 5210 72380 5518 72389
rect 5210 72378 5216 72380
rect 5272 72378 5296 72380
rect 5352 72378 5376 72380
rect 5432 72378 5456 72380
rect 5512 72378 5518 72380
rect 5272 72326 5274 72378
rect 5454 72326 5456 72378
rect 5210 72324 5216 72326
rect 5272 72324 5296 72326
rect 5352 72324 5376 72326
rect 5432 72324 5456 72326
rect 5512 72324 5518 72326
rect 5210 72315 5518 72324
rect 5552 72282 5580 86702
rect 6810 86524 7118 86533
rect 6810 86522 6816 86524
rect 6872 86522 6896 86524
rect 6952 86522 6976 86524
rect 7032 86522 7056 86524
rect 7112 86522 7118 86524
rect 6872 86470 6874 86522
rect 7054 86470 7056 86522
rect 6810 86468 6816 86470
rect 6872 86468 6896 86470
rect 6952 86468 6976 86470
rect 7032 86468 7056 86470
rect 7112 86468 7118 86470
rect 6810 86459 7118 86468
rect 8410 86524 8718 86533
rect 8410 86522 8416 86524
rect 8472 86522 8496 86524
rect 8552 86522 8576 86524
rect 8632 86522 8656 86524
rect 8712 86522 8718 86524
rect 8472 86470 8474 86522
rect 8654 86470 8656 86522
rect 8410 86468 8416 86470
rect 8472 86468 8496 86470
rect 8552 86468 8576 86470
rect 8632 86468 8656 86470
rect 8712 86468 8718 86470
rect 8410 86459 8718 86468
rect 6000 86420 6052 86426
rect 6000 86362 6052 86368
rect 5908 86352 5960 86358
rect 5908 86294 5960 86300
rect 5920 80054 5948 86294
rect 5828 80026 5948 80054
rect 5724 75404 5776 75410
rect 5724 75346 5776 75352
rect 5632 75200 5684 75206
rect 5632 75142 5684 75148
rect 5540 72276 5592 72282
rect 5540 72218 5592 72224
rect 5540 72072 5592 72078
rect 5540 72014 5592 72020
rect 5552 71398 5580 72014
rect 5540 71392 5592 71398
rect 5540 71334 5592 71340
rect 5210 71292 5518 71301
rect 5210 71290 5216 71292
rect 5272 71290 5296 71292
rect 5352 71290 5376 71292
rect 5432 71290 5456 71292
rect 5512 71290 5518 71292
rect 5272 71238 5274 71290
rect 5454 71238 5456 71290
rect 5210 71236 5216 71238
rect 5272 71236 5296 71238
rect 5352 71236 5376 71238
rect 5432 71236 5456 71238
rect 5512 71236 5518 71238
rect 5210 71227 5518 71236
rect 5540 70984 5592 70990
rect 5540 70926 5592 70932
rect 5210 70204 5518 70213
rect 5210 70202 5216 70204
rect 5272 70202 5296 70204
rect 5352 70202 5376 70204
rect 5432 70202 5456 70204
rect 5512 70202 5518 70204
rect 5272 70150 5274 70202
rect 5454 70150 5456 70202
rect 5210 70148 5216 70150
rect 5272 70148 5296 70150
rect 5352 70148 5376 70150
rect 5432 70148 5456 70150
rect 5512 70148 5518 70150
rect 5210 70139 5518 70148
rect 5172 70100 5224 70106
rect 5172 70042 5224 70048
rect 5184 69562 5212 70042
rect 5354 70000 5410 70009
rect 5354 69935 5410 69944
rect 5172 69556 5224 69562
rect 5172 69498 5224 69504
rect 5368 69465 5396 69935
rect 5448 69896 5500 69902
rect 5448 69838 5500 69844
rect 5460 69766 5488 69838
rect 5448 69760 5500 69766
rect 5448 69702 5500 69708
rect 5354 69456 5410 69465
rect 5354 69391 5410 69400
rect 5460 69222 5488 69702
rect 5448 69216 5500 69222
rect 5448 69158 5500 69164
rect 5210 69116 5518 69125
rect 5210 69114 5216 69116
rect 5272 69114 5296 69116
rect 5352 69114 5376 69116
rect 5432 69114 5456 69116
rect 5512 69114 5518 69116
rect 5272 69062 5274 69114
rect 5454 69062 5456 69114
rect 5210 69060 5216 69062
rect 5272 69060 5296 69062
rect 5352 69060 5376 69062
rect 5432 69060 5456 69062
rect 5512 69060 5518 69062
rect 5210 69051 5518 69060
rect 5552 69000 5580 70926
rect 5460 68972 5580 69000
rect 5356 68944 5408 68950
rect 5356 68886 5408 68892
rect 5264 68740 5316 68746
rect 5264 68682 5316 68688
rect 5172 68672 5224 68678
rect 5172 68614 5224 68620
rect 5080 68400 5132 68406
rect 5080 68342 5132 68348
rect 5184 68252 5212 68614
rect 5276 68474 5304 68682
rect 5264 68468 5316 68474
rect 5264 68410 5316 68416
rect 5092 68224 5212 68252
rect 4908 68054 5028 68082
rect 4896 67924 4948 67930
rect 4896 67866 4948 67872
rect 4526 67623 4582 67632
rect 4804 67652 4856 67658
rect 4804 67594 4856 67600
rect 4550 67484 4858 67493
rect 4550 67482 4556 67484
rect 4612 67482 4636 67484
rect 4692 67482 4716 67484
rect 4772 67482 4796 67484
rect 4852 67482 4858 67484
rect 4612 67430 4614 67482
rect 4794 67430 4796 67482
rect 4550 67428 4556 67430
rect 4612 67428 4636 67430
rect 4692 67428 4716 67430
rect 4772 67428 4796 67430
rect 4852 67428 4858 67430
rect 4550 67419 4858 67428
rect 4620 67244 4672 67250
rect 4620 67186 4672 67192
rect 4526 66736 4582 66745
rect 4526 66671 4528 66680
rect 4580 66671 4582 66680
rect 4528 66642 4580 66648
rect 4436 66496 4488 66502
rect 4342 66464 4398 66473
rect 4632 66484 4660 67186
rect 4712 67176 4764 67182
rect 4712 67118 4764 67124
rect 4724 66609 4752 67118
rect 4908 66774 4936 67866
rect 4896 66768 4948 66774
rect 4896 66710 4948 66716
rect 4710 66600 4766 66609
rect 4710 66535 4766 66544
rect 4632 66456 4936 66484
rect 4436 66438 4488 66444
rect 4342 66399 4398 66408
rect 4344 66292 4396 66298
rect 4344 66234 4396 66240
rect 4356 62422 4384 66234
rect 4344 62416 4396 62422
rect 4344 62358 4396 62364
rect 4344 62212 4396 62218
rect 4344 62154 4396 62160
rect 4252 59220 4304 59226
rect 4252 59162 4304 59168
rect 4356 59090 4384 62154
rect 4448 60722 4476 66438
rect 4550 66396 4858 66405
rect 4550 66394 4556 66396
rect 4612 66394 4636 66396
rect 4692 66394 4716 66396
rect 4772 66394 4796 66396
rect 4852 66394 4858 66396
rect 4612 66342 4614 66394
rect 4794 66342 4796 66394
rect 4550 66340 4556 66342
rect 4612 66340 4636 66342
rect 4692 66340 4716 66342
rect 4772 66340 4796 66342
rect 4852 66340 4858 66342
rect 4550 66331 4858 66340
rect 4618 66192 4674 66201
rect 4618 66127 4674 66136
rect 4632 65414 4660 66127
rect 4908 65618 4936 66456
rect 5000 66230 5028 68054
rect 5092 67930 5120 68224
rect 5368 68202 5396 68886
rect 5356 68196 5408 68202
rect 5460 68184 5488 68972
rect 5540 68672 5592 68678
rect 5540 68614 5592 68620
rect 5552 68252 5580 68614
rect 5644 68406 5672 75142
rect 5736 72185 5764 75346
rect 5722 72176 5778 72185
rect 5722 72111 5778 72120
rect 5724 72072 5776 72078
rect 5724 72014 5776 72020
rect 5736 71058 5764 72014
rect 5724 71052 5776 71058
rect 5724 70994 5776 71000
rect 5736 70378 5764 70994
rect 5828 70553 5856 80026
rect 5908 74656 5960 74662
rect 5908 74598 5960 74604
rect 5814 70544 5870 70553
rect 5814 70479 5870 70488
rect 5724 70372 5776 70378
rect 5724 70314 5776 70320
rect 5816 70372 5868 70378
rect 5816 70314 5868 70320
rect 5724 70100 5776 70106
rect 5724 70042 5776 70048
rect 5736 68785 5764 70042
rect 5828 68814 5856 70314
rect 5920 68950 5948 74598
rect 6012 72758 6040 86362
rect 8760 86080 8812 86086
rect 8760 86022 8812 86028
rect 6150 85980 6458 85989
rect 6150 85978 6156 85980
rect 6212 85978 6236 85980
rect 6292 85978 6316 85980
rect 6372 85978 6396 85980
rect 6452 85978 6458 85980
rect 6212 85926 6214 85978
rect 6394 85926 6396 85978
rect 6150 85924 6156 85926
rect 6212 85924 6236 85926
rect 6292 85924 6316 85926
rect 6372 85924 6396 85926
rect 6452 85924 6458 85926
rect 6150 85915 6458 85924
rect 7750 85980 8058 85989
rect 7750 85978 7756 85980
rect 7812 85978 7836 85980
rect 7892 85978 7916 85980
rect 7972 85978 7996 85980
rect 8052 85978 8058 85980
rect 7812 85926 7814 85978
rect 7994 85926 7996 85978
rect 7750 85924 7756 85926
rect 7812 85924 7836 85926
rect 7892 85924 7916 85926
rect 7972 85924 7996 85926
rect 8052 85924 8058 85926
rect 7750 85915 8058 85924
rect 6810 85436 7118 85445
rect 6810 85434 6816 85436
rect 6872 85434 6896 85436
rect 6952 85434 6976 85436
rect 7032 85434 7056 85436
rect 7112 85434 7118 85436
rect 6872 85382 6874 85434
rect 7054 85382 7056 85434
rect 6810 85380 6816 85382
rect 6872 85380 6896 85382
rect 6952 85380 6976 85382
rect 7032 85380 7056 85382
rect 7112 85380 7118 85382
rect 6810 85371 7118 85380
rect 8410 85436 8718 85445
rect 8410 85434 8416 85436
rect 8472 85434 8496 85436
rect 8552 85434 8576 85436
rect 8632 85434 8656 85436
rect 8712 85434 8718 85436
rect 8472 85382 8474 85434
rect 8654 85382 8656 85434
rect 8410 85380 8416 85382
rect 8472 85380 8496 85382
rect 8552 85380 8576 85382
rect 8632 85380 8656 85382
rect 8712 85380 8718 85382
rect 8410 85371 8718 85380
rect 8208 85264 8260 85270
rect 8208 85206 8260 85212
rect 8116 85196 8168 85202
rect 8116 85138 8168 85144
rect 7472 85128 7524 85134
rect 7472 85070 7524 85076
rect 7196 85060 7248 85066
rect 7196 85002 7248 85008
rect 6552 84992 6604 84998
rect 6552 84934 6604 84940
rect 6150 84892 6458 84901
rect 6150 84890 6156 84892
rect 6212 84890 6236 84892
rect 6292 84890 6316 84892
rect 6372 84890 6396 84892
rect 6452 84890 6458 84892
rect 6212 84838 6214 84890
rect 6394 84838 6396 84890
rect 6150 84836 6156 84838
rect 6212 84836 6236 84838
rect 6292 84836 6316 84838
rect 6372 84836 6396 84838
rect 6452 84836 6458 84838
rect 6150 84827 6458 84836
rect 6150 83804 6458 83813
rect 6150 83802 6156 83804
rect 6212 83802 6236 83804
rect 6292 83802 6316 83804
rect 6372 83802 6396 83804
rect 6452 83802 6458 83804
rect 6212 83750 6214 83802
rect 6394 83750 6396 83802
rect 6150 83748 6156 83750
rect 6212 83748 6236 83750
rect 6292 83748 6316 83750
rect 6372 83748 6396 83750
rect 6452 83748 6458 83750
rect 6150 83739 6458 83748
rect 6150 82716 6458 82725
rect 6150 82714 6156 82716
rect 6212 82714 6236 82716
rect 6292 82714 6316 82716
rect 6372 82714 6396 82716
rect 6452 82714 6458 82716
rect 6212 82662 6214 82714
rect 6394 82662 6396 82714
rect 6150 82660 6156 82662
rect 6212 82660 6236 82662
rect 6292 82660 6316 82662
rect 6372 82660 6396 82662
rect 6452 82660 6458 82662
rect 6150 82651 6458 82660
rect 6150 81628 6458 81637
rect 6150 81626 6156 81628
rect 6212 81626 6236 81628
rect 6292 81626 6316 81628
rect 6372 81626 6396 81628
rect 6452 81626 6458 81628
rect 6212 81574 6214 81626
rect 6394 81574 6396 81626
rect 6150 81572 6156 81574
rect 6212 81572 6236 81574
rect 6292 81572 6316 81574
rect 6372 81572 6396 81574
rect 6452 81572 6458 81574
rect 6150 81563 6458 81572
rect 6150 80540 6458 80549
rect 6150 80538 6156 80540
rect 6212 80538 6236 80540
rect 6292 80538 6316 80540
rect 6372 80538 6396 80540
rect 6452 80538 6458 80540
rect 6212 80486 6214 80538
rect 6394 80486 6396 80538
rect 6150 80484 6156 80486
rect 6212 80484 6236 80486
rect 6292 80484 6316 80486
rect 6372 80484 6396 80486
rect 6452 80484 6458 80486
rect 6150 80475 6458 80484
rect 6150 79452 6458 79461
rect 6150 79450 6156 79452
rect 6212 79450 6236 79452
rect 6292 79450 6316 79452
rect 6372 79450 6396 79452
rect 6452 79450 6458 79452
rect 6212 79398 6214 79450
rect 6394 79398 6396 79450
rect 6150 79396 6156 79398
rect 6212 79396 6236 79398
rect 6292 79396 6316 79398
rect 6372 79396 6396 79398
rect 6452 79396 6458 79398
rect 6150 79387 6458 79396
rect 6150 78364 6458 78373
rect 6150 78362 6156 78364
rect 6212 78362 6236 78364
rect 6292 78362 6316 78364
rect 6372 78362 6396 78364
rect 6452 78362 6458 78364
rect 6212 78310 6214 78362
rect 6394 78310 6396 78362
rect 6150 78308 6156 78310
rect 6212 78308 6236 78310
rect 6292 78308 6316 78310
rect 6372 78308 6396 78310
rect 6452 78308 6458 78310
rect 6150 78299 6458 78308
rect 6150 77276 6458 77285
rect 6150 77274 6156 77276
rect 6212 77274 6236 77276
rect 6292 77274 6316 77276
rect 6372 77274 6396 77276
rect 6452 77274 6458 77276
rect 6212 77222 6214 77274
rect 6394 77222 6396 77274
rect 6150 77220 6156 77222
rect 6212 77220 6236 77222
rect 6292 77220 6316 77222
rect 6372 77220 6396 77222
rect 6452 77220 6458 77222
rect 6150 77211 6458 77220
rect 6150 76188 6458 76197
rect 6150 76186 6156 76188
rect 6212 76186 6236 76188
rect 6292 76186 6316 76188
rect 6372 76186 6396 76188
rect 6452 76186 6458 76188
rect 6212 76134 6214 76186
rect 6394 76134 6396 76186
rect 6150 76132 6156 76134
rect 6212 76132 6236 76134
rect 6292 76132 6316 76134
rect 6372 76132 6396 76134
rect 6452 76132 6458 76134
rect 6150 76123 6458 76132
rect 6150 75100 6458 75109
rect 6150 75098 6156 75100
rect 6212 75098 6236 75100
rect 6292 75098 6316 75100
rect 6372 75098 6396 75100
rect 6452 75098 6458 75100
rect 6212 75046 6214 75098
rect 6394 75046 6396 75098
rect 6150 75044 6156 75046
rect 6212 75044 6236 75046
rect 6292 75044 6316 75046
rect 6372 75044 6396 75046
rect 6452 75044 6458 75046
rect 6150 75035 6458 75044
rect 6150 74012 6458 74021
rect 6150 74010 6156 74012
rect 6212 74010 6236 74012
rect 6292 74010 6316 74012
rect 6372 74010 6396 74012
rect 6452 74010 6458 74012
rect 6212 73958 6214 74010
rect 6394 73958 6396 74010
rect 6150 73956 6156 73958
rect 6212 73956 6236 73958
rect 6292 73956 6316 73958
rect 6372 73956 6396 73958
rect 6452 73956 6458 73958
rect 6150 73947 6458 73956
rect 6460 73704 6512 73710
rect 6460 73646 6512 73652
rect 6472 73166 6500 73646
rect 6460 73160 6512 73166
rect 6460 73102 6512 73108
rect 6150 72924 6458 72933
rect 6150 72922 6156 72924
rect 6212 72922 6236 72924
rect 6292 72922 6316 72924
rect 6372 72922 6396 72924
rect 6452 72922 6458 72924
rect 6212 72870 6214 72922
rect 6394 72870 6396 72922
rect 6150 72868 6156 72870
rect 6212 72868 6236 72870
rect 6292 72868 6316 72870
rect 6372 72868 6396 72870
rect 6452 72868 6458 72870
rect 6150 72859 6458 72868
rect 6000 72752 6052 72758
rect 6000 72694 6052 72700
rect 6274 72720 6330 72729
rect 6274 72655 6330 72664
rect 6460 72684 6512 72690
rect 6000 72616 6052 72622
rect 6000 72558 6052 72564
rect 6012 71942 6040 72558
rect 6288 72010 6316 72655
rect 6460 72626 6512 72632
rect 6472 72146 6500 72626
rect 6460 72140 6512 72146
rect 6460 72082 6512 72088
rect 6276 72004 6328 72010
rect 6276 71946 6328 71952
rect 6000 71936 6052 71942
rect 6000 71878 6052 71884
rect 6012 70632 6040 71878
rect 6150 71836 6458 71845
rect 6150 71834 6156 71836
rect 6212 71834 6236 71836
rect 6292 71834 6316 71836
rect 6372 71834 6396 71836
rect 6452 71834 6458 71836
rect 6212 71782 6214 71834
rect 6394 71782 6396 71834
rect 6150 71780 6156 71782
rect 6212 71780 6236 71782
rect 6292 71780 6316 71782
rect 6372 71780 6396 71782
rect 6452 71780 6458 71782
rect 6150 71771 6458 71780
rect 6564 71720 6592 84934
rect 6810 84348 7118 84357
rect 6810 84346 6816 84348
rect 6872 84346 6896 84348
rect 6952 84346 6976 84348
rect 7032 84346 7056 84348
rect 7112 84346 7118 84348
rect 6872 84294 6874 84346
rect 7054 84294 7056 84346
rect 6810 84292 6816 84294
rect 6872 84292 6896 84294
rect 6952 84292 6976 84294
rect 7032 84292 7056 84294
rect 7112 84292 7118 84294
rect 6810 84283 7118 84292
rect 6644 83904 6696 83910
rect 6644 83846 6696 83852
rect 6656 74338 6684 83846
rect 6810 83260 7118 83269
rect 6810 83258 6816 83260
rect 6872 83258 6896 83260
rect 6952 83258 6976 83260
rect 7032 83258 7056 83260
rect 7112 83258 7118 83260
rect 6872 83206 6874 83258
rect 7054 83206 7056 83258
rect 6810 83204 6816 83206
rect 6872 83204 6896 83206
rect 6952 83204 6976 83206
rect 7032 83204 7056 83206
rect 7112 83204 7118 83206
rect 6810 83195 7118 83204
rect 6810 82172 7118 82181
rect 6810 82170 6816 82172
rect 6872 82170 6896 82172
rect 6952 82170 6976 82172
rect 7032 82170 7056 82172
rect 7112 82170 7118 82172
rect 6872 82118 6874 82170
rect 7054 82118 7056 82170
rect 6810 82116 6816 82118
rect 6872 82116 6896 82118
rect 6952 82116 6976 82118
rect 7032 82116 7056 82118
rect 7112 82116 7118 82118
rect 6810 82107 7118 82116
rect 6810 81084 7118 81093
rect 6810 81082 6816 81084
rect 6872 81082 6896 81084
rect 6952 81082 6976 81084
rect 7032 81082 7056 81084
rect 7112 81082 7118 81084
rect 6872 81030 6874 81082
rect 7054 81030 7056 81082
rect 6810 81028 6816 81030
rect 6872 81028 6896 81030
rect 6952 81028 6976 81030
rect 7032 81028 7056 81030
rect 7112 81028 7118 81030
rect 6810 81019 7118 81028
rect 6810 79996 7118 80005
rect 6810 79994 6816 79996
rect 6872 79994 6896 79996
rect 6952 79994 6976 79996
rect 7032 79994 7056 79996
rect 7112 79994 7118 79996
rect 6872 79942 6874 79994
rect 7054 79942 7056 79994
rect 6810 79940 6816 79942
rect 6872 79940 6896 79942
rect 6952 79940 6976 79942
rect 7032 79940 7056 79942
rect 7112 79940 7118 79942
rect 6810 79931 7118 79940
rect 6810 78908 7118 78917
rect 6810 78906 6816 78908
rect 6872 78906 6896 78908
rect 6952 78906 6976 78908
rect 7032 78906 7056 78908
rect 7112 78906 7118 78908
rect 6872 78854 6874 78906
rect 7054 78854 7056 78906
rect 6810 78852 6816 78854
rect 6872 78852 6896 78854
rect 6952 78852 6976 78854
rect 7032 78852 7056 78854
rect 7112 78852 7118 78854
rect 6810 78843 7118 78852
rect 6810 77820 7118 77829
rect 6810 77818 6816 77820
rect 6872 77818 6896 77820
rect 6952 77818 6976 77820
rect 7032 77818 7056 77820
rect 7112 77818 7118 77820
rect 6872 77766 6874 77818
rect 7054 77766 7056 77818
rect 6810 77764 6816 77766
rect 6872 77764 6896 77766
rect 6952 77764 6976 77766
rect 7032 77764 7056 77766
rect 7112 77764 7118 77766
rect 6810 77755 7118 77764
rect 7208 77294 7236 85002
rect 7380 83700 7432 83706
rect 7380 83642 7432 83648
rect 7208 77266 7328 77294
rect 6810 76732 7118 76741
rect 6810 76730 6816 76732
rect 6872 76730 6896 76732
rect 6952 76730 6976 76732
rect 7032 76730 7056 76732
rect 7112 76730 7118 76732
rect 6872 76678 6874 76730
rect 7054 76678 7056 76730
rect 6810 76676 6816 76678
rect 6872 76676 6896 76678
rect 6952 76676 6976 76678
rect 7032 76676 7056 76678
rect 7112 76676 7118 76678
rect 6810 76667 7118 76676
rect 6810 75644 7118 75653
rect 6810 75642 6816 75644
rect 6872 75642 6896 75644
rect 6952 75642 6976 75644
rect 7032 75642 7056 75644
rect 7112 75642 7118 75644
rect 6872 75590 6874 75642
rect 7054 75590 7056 75642
rect 6810 75588 6816 75590
rect 6872 75588 6896 75590
rect 6952 75588 6976 75590
rect 7032 75588 7056 75590
rect 7112 75588 7118 75590
rect 6810 75579 7118 75588
rect 7196 75268 7248 75274
rect 7196 75210 7248 75216
rect 6810 74556 7118 74565
rect 6810 74554 6816 74556
rect 6872 74554 6896 74556
rect 6952 74554 6976 74556
rect 7032 74554 7056 74556
rect 7112 74554 7118 74556
rect 6872 74502 6874 74554
rect 7054 74502 7056 74554
rect 6810 74500 6816 74502
rect 6872 74500 6896 74502
rect 6952 74500 6976 74502
rect 7032 74500 7056 74502
rect 7112 74500 7118 74502
rect 6810 74491 7118 74500
rect 6656 74310 6868 74338
rect 6840 73846 6868 74310
rect 7208 74254 7236 75210
rect 7300 74633 7328 77266
rect 7286 74624 7342 74633
rect 7286 74559 7342 74568
rect 7288 74452 7340 74458
rect 7288 74394 7340 74400
rect 6920 74248 6972 74254
rect 6920 74190 6972 74196
rect 7196 74248 7248 74254
rect 7196 74190 7248 74196
rect 6828 73840 6880 73846
rect 6828 73782 6880 73788
rect 6736 73772 6788 73778
rect 6736 73714 6788 73720
rect 6748 73352 6776 73714
rect 6932 73574 6960 74190
rect 7196 73704 7248 73710
rect 7196 73646 7248 73652
rect 6920 73568 6972 73574
rect 6920 73510 6972 73516
rect 6810 73468 7118 73477
rect 6810 73466 6816 73468
rect 6872 73466 6896 73468
rect 6952 73466 6976 73468
rect 7032 73466 7056 73468
rect 7112 73466 7118 73468
rect 6872 73414 6874 73466
rect 7054 73414 7056 73466
rect 6810 73412 6816 73414
rect 6872 73412 6896 73414
rect 6952 73412 6976 73414
rect 7032 73412 7056 73414
rect 7112 73412 7118 73414
rect 6810 73403 7118 73412
rect 6748 73324 6868 73352
rect 6644 73228 6696 73234
rect 6644 73170 6696 73176
rect 6380 71692 6592 71720
rect 6380 71602 6408 71692
rect 6656 71652 6684 73170
rect 6840 73166 6868 73324
rect 7010 73264 7066 73273
rect 6920 73228 6972 73234
rect 7010 73199 7066 73208
rect 6920 73170 6972 73176
rect 6828 73160 6880 73166
rect 6734 73128 6790 73137
rect 6828 73102 6880 73108
rect 6734 73063 6790 73072
rect 6564 71624 6684 71652
rect 6368 71596 6420 71602
rect 6368 71538 6420 71544
rect 6460 71596 6512 71602
rect 6460 71538 6512 71544
rect 6472 71194 6500 71538
rect 6460 71188 6512 71194
rect 6460 71130 6512 71136
rect 6564 71074 6592 71624
rect 6748 71584 6776 73063
rect 6840 72690 6868 73102
rect 6828 72684 6880 72690
rect 6828 72626 6880 72632
rect 6932 72622 6960 73170
rect 6920 72616 6972 72622
rect 6826 72584 6882 72593
rect 6920 72558 6972 72564
rect 6826 72519 6882 72528
rect 6840 72486 6868 72519
rect 7024 72486 7052 73199
rect 7104 73092 7156 73098
rect 7104 73034 7156 73040
rect 7116 72622 7144 73034
rect 7208 72865 7236 73646
rect 7194 72856 7250 72865
rect 7194 72791 7250 72800
rect 7196 72684 7248 72690
rect 7196 72626 7248 72632
rect 7104 72616 7156 72622
rect 7104 72558 7156 72564
rect 6828 72480 6880 72486
rect 6828 72422 6880 72428
rect 7012 72480 7064 72486
rect 7012 72422 7064 72428
rect 6810 72380 7118 72389
rect 6810 72378 6816 72380
rect 6872 72378 6896 72380
rect 6952 72378 6976 72380
rect 7032 72378 7056 72380
rect 7112 72378 7118 72380
rect 6872 72326 6874 72378
rect 7054 72326 7056 72378
rect 6810 72324 6816 72326
rect 6872 72324 6896 72326
rect 6952 72324 6976 72326
rect 7032 72324 7056 72326
rect 7112 72324 7118 72326
rect 6810 72315 7118 72324
rect 7208 72264 7236 72626
rect 7300 72604 7328 74394
rect 7392 73370 7420 83642
rect 7484 73710 7512 85070
rect 7750 84892 8058 84901
rect 7750 84890 7756 84892
rect 7812 84890 7836 84892
rect 7892 84890 7916 84892
rect 7972 84890 7996 84892
rect 8052 84890 8058 84892
rect 7812 84838 7814 84890
rect 7994 84838 7996 84890
rect 7750 84836 7756 84838
rect 7812 84836 7836 84838
rect 7892 84836 7916 84838
rect 7972 84836 7996 84838
rect 8052 84836 8058 84838
rect 7750 84827 8058 84836
rect 7750 83804 8058 83813
rect 7750 83802 7756 83804
rect 7812 83802 7836 83804
rect 7892 83802 7916 83804
rect 7972 83802 7996 83804
rect 8052 83802 8058 83804
rect 7812 83750 7814 83802
rect 7994 83750 7996 83802
rect 7750 83748 7756 83750
rect 7812 83748 7836 83750
rect 7892 83748 7916 83750
rect 7972 83748 7996 83750
rect 8052 83748 8058 83750
rect 7750 83739 8058 83748
rect 7750 82716 8058 82725
rect 7750 82714 7756 82716
rect 7812 82714 7836 82716
rect 7892 82714 7916 82716
rect 7972 82714 7996 82716
rect 8052 82714 8058 82716
rect 7812 82662 7814 82714
rect 7994 82662 7996 82714
rect 7750 82660 7756 82662
rect 7812 82660 7836 82662
rect 7892 82660 7916 82662
rect 7972 82660 7996 82662
rect 8052 82660 8058 82662
rect 7750 82651 8058 82660
rect 7750 81628 8058 81637
rect 7750 81626 7756 81628
rect 7812 81626 7836 81628
rect 7892 81626 7916 81628
rect 7972 81626 7996 81628
rect 8052 81626 8058 81628
rect 7812 81574 7814 81626
rect 7994 81574 7996 81626
rect 7750 81572 7756 81574
rect 7812 81572 7836 81574
rect 7892 81572 7916 81574
rect 7972 81572 7996 81574
rect 8052 81572 8058 81574
rect 7750 81563 8058 81572
rect 7750 80540 8058 80549
rect 7750 80538 7756 80540
rect 7812 80538 7836 80540
rect 7892 80538 7916 80540
rect 7972 80538 7996 80540
rect 8052 80538 8058 80540
rect 7812 80486 7814 80538
rect 7994 80486 7996 80538
rect 7750 80484 7756 80486
rect 7812 80484 7836 80486
rect 7892 80484 7916 80486
rect 7972 80484 7996 80486
rect 8052 80484 8058 80486
rect 7750 80475 8058 80484
rect 7750 79452 8058 79461
rect 7750 79450 7756 79452
rect 7812 79450 7836 79452
rect 7892 79450 7916 79452
rect 7972 79450 7996 79452
rect 8052 79450 8058 79452
rect 7812 79398 7814 79450
rect 7994 79398 7996 79450
rect 7750 79396 7756 79398
rect 7812 79396 7836 79398
rect 7892 79396 7916 79398
rect 7972 79396 7996 79398
rect 8052 79396 8058 79398
rect 7750 79387 8058 79396
rect 7750 78364 8058 78373
rect 7750 78362 7756 78364
rect 7812 78362 7836 78364
rect 7892 78362 7916 78364
rect 7972 78362 7996 78364
rect 8052 78362 8058 78364
rect 7812 78310 7814 78362
rect 7994 78310 7996 78362
rect 7750 78308 7756 78310
rect 7812 78308 7836 78310
rect 7892 78308 7916 78310
rect 7972 78308 7996 78310
rect 8052 78308 8058 78310
rect 7750 78299 8058 78308
rect 7750 77276 8058 77285
rect 7750 77274 7756 77276
rect 7812 77274 7836 77276
rect 7892 77274 7916 77276
rect 7972 77274 7996 77276
rect 8052 77274 8058 77276
rect 7812 77222 7814 77274
rect 7994 77222 7996 77274
rect 7750 77220 7756 77222
rect 7812 77220 7836 77222
rect 7892 77220 7916 77222
rect 7972 77220 7996 77222
rect 8052 77220 8058 77222
rect 7750 77211 8058 77220
rect 7656 77036 7708 77042
rect 7656 76978 7708 76984
rect 7564 74792 7616 74798
rect 7564 74734 7616 74740
rect 7472 73704 7524 73710
rect 7472 73646 7524 73652
rect 7470 73536 7526 73545
rect 7470 73471 7526 73480
rect 7380 73364 7432 73370
rect 7380 73306 7432 73312
rect 7484 73216 7512 73471
rect 7392 73188 7512 73216
rect 7392 72690 7420 73188
rect 7576 73166 7604 74734
rect 7564 73160 7616 73166
rect 7564 73102 7616 73108
rect 7668 73098 7696 76978
rect 7750 76188 8058 76197
rect 7750 76186 7756 76188
rect 7812 76186 7836 76188
rect 7892 76186 7916 76188
rect 7972 76186 7996 76188
rect 8052 76186 8058 76188
rect 7812 76134 7814 76186
rect 7994 76134 7996 76186
rect 7750 76132 7756 76134
rect 7812 76132 7836 76134
rect 7892 76132 7916 76134
rect 7972 76132 7996 76134
rect 8052 76132 8058 76134
rect 7750 76123 8058 76132
rect 7750 75100 8058 75109
rect 7750 75098 7756 75100
rect 7812 75098 7836 75100
rect 7892 75098 7916 75100
rect 7972 75098 7996 75100
rect 8052 75098 8058 75100
rect 7812 75046 7814 75098
rect 7994 75046 7996 75098
rect 7750 75044 7756 75046
rect 7812 75044 7836 75046
rect 7892 75044 7916 75046
rect 7972 75044 7996 75046
rect 8052 75044 8058 75046
rect 7750 75035 8058 75044
rect 7750 74012 8058 74021
rect 7750 74010 7756 74012
rect 7812 74010 7836 74012
rect 7892 74010 7916 74012
rect 7972 74010 7996 74012
rect 8052 74010 8058 74012
rect 7812 73958 7814 74010
rect 7994 73958 7996 74010
rect 7750 73956 7756 73958
rect 7812 73956 7836 73958
rect 7892 73956 7916 73958
rect 7972 73956 7996 73958
rect 8052 73956 8058 73958
rect 7750 73947 8058 73956
rect 8128 73896 8156 85138
rect 8220 76430 8248 85206
rect 8410 84348 8718 84357
rect 8410 84346 8416 84348
rect 8472 84346 8496 84348
rect 8552 84346 8576 84348
rect 8632 84346 8656 84348
rect 8712 84346 8718 84348
rect 8472 84294 8474 84346
rect 8654 84294 8656 84346
rect 8410 84292 8416 84294
rect 8472 84292 8496 84294
rect 8552 84292 8576 84294
rect 8632 84292 8656 84294
rect 8712 84292 8718 84294
rect 8410 84283 8718 84292
rect 8300 83632 8352 83638
rect 8300 83574 8352 83580
rect 8208 76424 8260 76430
rect 8208 76366 8260 76372
rect 8312 74730 8340 83574
rect 8410 83260 8718 83269
rect 8410 83258 8416 83260
rect 8472 83258 8496 83260
rect 8552 83258 8576 83260
rect 8632 83258 8656 83260
rect 8712 83258 8718 83260
rect 8472 83206 8474 83258
rect 8654 83206 8656 83258
rect 8410 83204 8416 83206
rect 8472 83204 8496 83206
rect 8552 83204 8576 83206
rect 8632 83204 8656 83206
rect 8712 83204 8718 83206
rect 8410 83195 8718 83204
rect 8410 82172 8718 82181
rect 8410 82170 8416 82172
rect 8472 82170 8496 82172
rect 8552 82170 8576 82172
rect 8632 82170 8656 82172
rect 8712 82170 8718 82172
rect 8472 82118 8474 82170
rect 8654 82118 8656 82170
rect 8410 82116 8416 82118
rect 8472 82116 8496 82118
rect 8552 82116 8576 82118
rect 8632 82116 8656 82118
rect 8712 82116 8718 82118
rect 8410 82107 8718 82116
rect 8410 81084 8718 81093
rect 8410 81082 8416 81084
rect 8472 81082 8496 81084
rect 8552 81082 8576 81084
rect 8632 81082 8656 81084
rect 8712 81082 8718 81084
rect 8472 81030 8474 81082
rect 8654 81030 8656 81082
rect 8410 81028 8416 81030
rect 8472 81028 8496 81030
rect 8552 81028 8576 81030
rect 8632 81028 8656 81030
rect 8712 81028 8718 81030
rect 8410 81019 8718 81028
rect 8410 79996 8718 80005
rect 8410 79994 8416 79996
rect 8472 79994 8496 79996
rect 8552 79994 8576 79996
rect 8632 79994 8656 79996
rect 8712 79994 8718 79996
rect 8472 79942 8474 79994
rect 8654 79942 8656 79994
rect 8410 79940 8416 79942
rect 8472 79940 8496 79942
rect 8552 79940 8576 79942
rect 8632 79940 8656 79942
rect 8712 79940 8718 79942
rect 8410 79931 8718 79940
rect 8410 78908 8718 78917
rect 8410 78906 8416 78908
rect 8472 78906 8496 78908
rect 8552 78906 8576 78908
rect 8632 78906 8656 78908
rect 8712 78906 8718 78908
rect 8472 78854 8474 78906
rect 8654 78854 8656 78906
rect 8410 78852 8416 78854
rect 8472 78852 8496 78854
rect 8552 78852 8576 78854
rect 8632 78852 8656 78854
rect 8712 78852 8718 78854
rect 8410 78843 8718 78852
rect 8410 77820 8718 77829
rect 8410 77818 8416 77820
rect 8472 77818 8496 77820
rect 8552 77818 8576 77820
rect 8632 77818 8656 77820
rect 8712 77818 8718 77820
rect 8472 77766 8474 77818
rect 8654 77766 8656 77818
rect 8410 77764 8416 77766
rect 8472 77764 8496 77766
rect 8552 77764 8576 77766
rect 8632 77764 8656 77766
rect 8712 77764 8718 77766
rect 8410 77755 8718 77764
rect 8410 76732 8718 76741
rect 8410 76730 8416 76732
rect 8472 76730 8496 76732
rect 8552 76730 8576 76732
rect 8632 76730 8656 76732
rect 8712 76730 8718 76732
rect 8472 76678 8474 76730
rect 8654 76678 8656 76730
rect 8410 76676 8416 76678
rect 8472 76676 8496 76678
rect 8552 76676 8576 76678
rect 8632 76676 8656 76678
rect 8712 76676 8718 76678
rect 8410 76667 8718 76676
rect 8772 76498 8800 86022
rect 8944 85740 8996 85746
rect 8944 85682 8996 85688
rect 8956 76974 8984 85682
rect 9048 77178 9076 87110
rect 10784 87100 10836 87106
rect 10784 87042 10836 87048
rect 10416 87032 10468 87038
rect 10416 86974 10468 86980
rect 10010 86524 10318 86533
rect 10010 86522 10016 86524
rect 10072 86522 10096 86524
rect 10152 86522 10176 86524
rect 10232 86522 10256 86524
rect 10312 86522 10318 86524
rect 10072 86470 10074 86522
rect 10254 86470 10256 86522
rect 10010 86468 10016 86470
rect 10072 86468 10096 86470
rect 10152 86468 10176 86470
rect 10232 86468 10256 86470
rect 10312 86468 10318 86470
rect 10010 86459 10318 86468
rect 9350 85980 9658 85989
rect 9350 85978 9356 85980
rect 9412 85978 9436 85980
rect 9492 85978 9516 85980
rect 9572 85978 9596 85980
rect 9652 85978 9658 85980
rect 9412 85926 9414 85978
rect 9594 85926 9596 85978
rect 9350 85924 9356 85926
rect 9412 85924 9436 85926
rect 9492 85924 9516 85926
rect 9572 85924 9596 85926
rect 9652 85924 9658 85926
rect 9350 85915 9658 85924
rect 9220 85808 9272 85814
rect 9220 85750 9272 85756
rect 9128 85604 9180 85610
rect 9128 85546 9180 85552
rect 9036 77172 9088 77178
rect 9036 77114 9088 77120
rect 8944 76968 8996 76974
rect 8944 76910 8996 76916
rect 8956 76498 8984 76910
rect 8760 76492 8812 76498
rect 8760 76434 8812 76440
rect 8944 76492 8996 76498
rect 8944 76434 8996 76440
rect 8410 75644 8718 75653
rect 8410 75642 8416 75644
rect 8472 75642 8496 75644
rect 8552 75642 8576 75644
rect 8632 75642 8656 75644
rect 8712 75642 8718 75644
rect 8472 75590 8474 75642
rect 8654 75590 8656 75642
rect 8410 75588 8416 75590
rect 8472 75588 8496 75590
rect 8552 75588 8576 75590
rect 8632 75588 8656 75590
rect 8712 75588 8718 75590
rect 8410 75579 8718 75588
rect 8484 75404 8536 75410
rect 8484 75346 8536 75352
rect 8496 74866 8524 75346
rect 8772 75002 8800 76434
rect 8852 76356 8904 76362
rect 8852 76298 8904 76304
rect 8760 74996 8812 75002
rect 8760 74938 8812 74944
rect 8484 74860 8536 74866
rect 8484 74802 8536 74808
rect 8300 74724 8352 74730
rect 8300 74666 8352 74672
rect 8496 74662 8524 74802
rect 8760 74724 8812 74730
rect 8760 74666 8812 74672
rect 8208 74656 8260 74662
rect 8208 74598 8260 74604
rect 8484 74656 8536 74662
rect 8484 74598 8536 74604
rect 8220 74254 8248 74598
rect 8410 74556 8718 74565
rect 8410 74554 8416 74556
rect 8472 74554 8496 74556
rect 8552 74554 8576 74556
rect 8632 74554 8656 74556
rect 8712 74554 8718 74556
rect 8472 74502 8474 74554
rect 8654 74502 8656 74554
rect 8410 74500 8416 74502
rect 8472 74500 8496 74502
rect 8552 74500 8576 74502
rect 8632 74500 8656 74502
rect 8712 74500 8718 74502
rect 8410 74491 8718 74500
rect 8208 74248 8260 74254
rect 8208 74190 8260 74196
rect 8036 73868 8156 73896
rect 8036 73778 8064 73868
rect 7840 73772 7892 73778
rect 7840 73714 7892 73720
rect 8024 73772 8076 73778
rect 8024 73714 8076 73720
rect 8116 73772 8168 73778
rect 8116 73714 8168 73720
rect 7746 73536 7802 73545
rect 7746 73471 7802 73480
rect 7760 73234 7788 73471
rect 7852 73302 7880 73714
rect 7840 73296 7892 73302
rect 7840 73238 7892 73244
rect 8036 73250 8064 73714
rect 8128 73370 8156 73714
rect 8220 73545 8248 74190
rect 8392 73772 8444 73778
rect 8392 73714 8444 73720
rect 8404 73574 8432 73714
rect 8300 73568 8352 73574
rect 8206 73536 8262 73545
rect 8300 73510 8352 73516
rect 8392 73568 8444 73574
rect 8392 73510 8444 73516
rect 8206 73471 8262 73480
rect 8116 73364 8168 73370
rect 8116 73306 8168 73312
rect 8208 73296 8260 73302
rect 8114 73264 8170 73273
rect 7748 73228 7800 73234
rect 7748 73170 7800 73176
rect 7932 73228 7984 73234
rect 8036 73222 8114 73250
rect 8208 73238 8260 73244
rect 8114 73199 8170 73208
rect 7932 73170 7984 73176
rect 7944 73114 7972 73170
rect 7472 73092 7524 73098
rect 7472 73034 7524 73040
rect 7656 73092 7708 73098
rect 7944 73086 8156 73114
rect 7656 73034 7708 73040
rect 7484 72690 7512 73034
rect 7750 72924 8058 72933
rect 7750 72922 7756 72924
rect 7812 72922 7836 72924
rect 7892 72922 7916 72924
rect 7972 72922 7996 72924
rect 8052 72922 8058 72924
rect 7812 72870 7814 72922
rect 7994 72870 7996 72922
rect 7750 72868 7756 72870
rect 7812 72868 7836 72870
rect 7892 72868 7916 72870
rect 7972 72868 7996 72870
rect 8052 72868 8058 72870
rect 7562 72856 7618 72865
rect 7750 72859 8058 72868
rect 7562 72791 7618 72800
rect 7380 72684 7432 72690
rect 7380 72626 7432 72632
rect 7472 72684 7524 72690
rect 7472 72626 7524 72632
rect 7300 72576 7333 72604
rect 7116 72236 7236 72264
rect 6826 72040 6882 72049
rect 6826 71975 6882 71984
rect 6840 71738 6868 71975
rect 6828 71732 6880 71738
rect 6828 71674 6880 71680
rect 7116 71602 7144 72236
rect 7194 72176 7250 72185
rect 7305 72128 7333 72576
rect 7484 72570 7512 72626
rect 7194 72111 7196 72120
rect 7248 72111 7250 72120
rect 7196 72082 7248 72088
rect 7300 72100 7333 72128
rect 7392 72542 7512 72570
rect 7208 71602 7236 72082
rect 7300 71738 7328 72100
rect 7288 71732 7340 71738
rect 7288 71674 7340 71680
rect 7392 71618 7420 72542
rect 7472 72480 7524 72486
rect 7472 72422 7524 72428
rect 6472 71046 6592 71074
rect 6656 71556 6776 71584
rect 7104 71596 7156 71602
rect 6472 70836 6500 71046
rect 6552 70984 6604 70990
rect 6550 70952 6552 70961
rect 6604 70952 6606 70961
rect 6550 70887 6606 70896
rect 6472 70808 6592 70836
rect 6150 70748 6458 70757
rect 6150 70746 6156 70748
rect 6212 70746 6236 70748
rect 6292 70746 6316 70748
rect 6372 70746 6396 70748
rect 6452 70746 6458 70748
rect 6212 70694 6214 70746
rect 6394 70694 6396 70746
rect 6150 70692 6156 70694
rect 6212 70692 6236 70694
rect 6292 70692 6316 70694
rect 6372 70692 6396 70694
rect 6452 70692 6458 70694
rect 6150 70683 6458 70692
rect 6368 70644 6420 70650
rect 6012 70604 6132 70632
rect 6000 70440 6052 70446
rect 6000 70382 6052 70388
rect 5908 68944 5960 68950
rect 5908 68886 5960 68892
rect 5816 68808 5868 68814
rect 5722 68776 5778 68785
rect 5816 68750 5868 68756
rect 5906 68776 5962 68785
rect 5722 68711 5778 68720
rect 5632 68400 5684 68406
rect 5632 68342 5684 68348
rect 5552 68224 5672 68252
rect 5460 68156 5580 68184
rect 5356 68138 5408 68144
rect 5210 68028 5518 68037
rect 5210 68026 5216 68028
rect 5272 68026 5296 68028
rect 5352 68026 5376 68028
rect 5432 68026 5456 68028
rect 5512 68026 5518 68028
rect 5272 67974 5274 68026
rect 5454 67974 5456 68026
rect 5210 67972 5216 67974
rect 5272 67972 5296 67974
rect 5352 67972 5376 67974
rect 5432 67972 5456 67974
rect 5512 67972 5518 67974
rect 5210 67963 5518 67972
rect 5080 67924 5132 67930
rect 5080 67866 5132 67872
rect 5264 67924 5316 67930
rect 5264 67866 5316 67872
rect 5356 67924 5408 67930
rect 5552 67912 5580 68156
rect 5356 67866 5408 67872
rect 5460 67884 5580 67912
rect 5080 67652 5132 67658
rect 5080 67594 5132 67600
rect 5092 67046 5120 67594
rect 5276 67386 5304 67866
rect 5368 67538 5396 67866
rect 5460 67658 5488 67884
rect 5540 67720 5592 67726
rect 5540 67662 5592 67668
rect 5448 67652 5500 67658
rect 5448 67594 5500 67600
rect 5368 67510 5488 67538
rect 5264 67380 5316 67386
rect 5264 67322 5316 67328
rect 5356 67244 5408 67250
rect 5356 67186 5408 67192
rect 5368 67153 5396 67186
rect 5354 67144 5410 67153
rect 5354 67079 5410 67088
rect 5460 67046 5488 67510
rect 5080 67040 5132 67046
rect 5080 66982 5132 66988
rect 5448 67040 5500 67046
rect 5448 66982 5500 66988
rect 4988 66224 5040 66230
rect 4988 66166 5040 66172
rect 4988 66088 5040 66094
rect 4988 66030 5040 66036
rect 4896 65612 4948 65618
rect 4896 65554 4948 65560
rect 5000 65498 5028 66030
rect 4908 65470 5028 65498
rect 5092 65482 5120 66982
rect 5210 66940 5518 66949
rect 5210 66938 5216 66940
rect 5272 66938 5296 66940
rect 5352 66938 5376 66940
rect 5432 66938 5456 66940
rect 5512 66938 5518 66940
rect 5272 66886 5274 66938
rect 5454 66886 5456 66938
rect 5210 66884 5216 66886
rect 5272 66884 5296 66886
rect 5352 66884 5376 66886
rect 5432 66884 5456 66886
rect 5512 66884 5518 66886
rect 5210 66875 5518 66884
rect 5172 66768 5224 66774
rect 5172 66710 5224 66716
rect 5356 66768 5408 66774
rect 5356 66710 5408 66716
rect 5184 66162 5212 66710
rect 5264 66564 5316 66570
rect 5264 66506 5316 66512
rect 5172 66156 5224 66162
rect 5172 66098 5224 66104
rect 5276 66094 5304 66506
rect 5368 66162 5396 66710
rect 5552 66450 5580 67662
rect 5460 66422 5580 66450
rect 5356 66156 5408 66162
rect 5356 66098 5408 66104
rect 5264 66088 5316 66094
rect 5264 66030 5316 66036
rect 5368 65940 5396 66098
rect 5460 66008 5488 66422
rect 5540 66292 5592 66298
rect 5644 66280 5672 68224
rect 5724 68196 5776 68202
rect 5724 68138 5776 68144
rect 5592 66252 5672 66280
rect 5540 66234 5592 66240
rect 5736 66230 5764 68138
rect 5724 66224 5776 66230
rect 5724 66166 5776 66172
rect 5828 66162 5856 68750
rect 5906 68711 5962 68720
rect 5920 67862 5948 68711
rect 5908 67856 5960 67862
rect 5908 67798 5960 67804
rect 6012 67640 6040 70382
rect 6104 70310 6132 70604
rect 6368 70586 6420 70592
rect 6092 70304 6144 70310
rect 6092 70246 6144 70252
rect 6184 70304 6236 70310
rect 6184 70246 6236 70252
rect 6104 69952 6132 70246
rect 6196 70106 6224 70246
rect 6380 70106 6408 70586
rect 6564 70582 6592 70808
rect 6552 70576 6604 70582
rect 6552 70518 6604 70524
rect 6460 70508 6512 70514
rect 6460 70450 6512 70456
rect 6472 70394 6500 70450
rect 6472 70366 6592 70394
rect 6184 70100 6236 70106
rect 6184 70042 6236 70048
rect 6368 70100 6420 70106
rect 6368 70042 6420 70048
rect 6184 69964 6236 69970
rect 6104 69924 6184 69952
rect 6184 69906 6236 69912
rect 6092 69760 6144 69766
rect 6276 69760 6328 69766
rect 6144 69720 6276 69748
rect 6092 69702 6144 69708
rect 6276 69702 6328 69708
rect 6150 69660 6458 69669
rect 6150 69658 6156 69660
rect 6212 69658 6236 69660
rect 6292 69658 6316 69660
rect 6372 69658 6396 69660
rect 6452 69658 6458 69660
rect 6212 69606 6214 69658
rect 6394 69606 6396 69658
rect 6150 69604 6156 69606
rect 6212 69604 6236 69606
rect 6292 69604 6316 69606
rect 6372 69604 6396 69606
rect 6452 69604 6458 69606
rect 6150 69595 6458 69604
rect 6564 69562 6592 70366
rect 6552 69556 6604 69562
rect 6552 69498 6604 69504
rect 6368 69420 6420 69426
rect 6368 69362 6420 69368
rect 6380 69306 6408 69362
rect 6380 69290 6592 69306
rect 6380 69284 6604 69290
rect 6380 69278 6552 69284
rect 6552 69226 6604 69232
rect 6092 69216 6144 69222
rect 6092 69158 6144 69164
rect 6460 69216 6512 69222
rect 6460 69158 6512 69164
rect 6104 68678 6132 69158
rect 6472 68898 6500 69158
rect 6656 69000 6684 71556
rect 7104 71538 7156 71544
rect 7196 71596 7248 71602
rect 7196 71538 7248 71544
rect 7300 71590 7420 71618
rect 6736 71392 6788 71398
rect 6736 71334 6788 71340
rect 7104 71392 7156 71398
rect 7156 71352 7236 71380
rect 7104 71334 7156 71340
rect 6748 69834 6776 71334
rect 6810 71292 7118 71301
rect 6810 71290 6816 71292
rect 6872 71290 6896 71292
rect 6952 71290 6976 71292
rect 7032 71290 7056 71292
rect 7112 71290 7118 71292
rect 6872 71238 6874 71290
rect 7054 71238 7056 71290
rect 6810 71236 6816 71238
rect 6872 71236 6896 71238
rect 6952 71236 6976 71238
rect 7032 71236 7056 71238
rect 7112 71236 7118 71238
rect 6810 71227 7118 71236
rect 6920 71188 6972 71194
rect 6920 71130 6972 71136
rect 7012 71188 7064 71194
rect 7012 71130 7064 71136
rect 6828 71120 6880 71126
rect 6828 71062 6880 71068
rect 6840 70650 6868 71062
rect 6828 70644 6880 70650
rect 6828 70586 6880 70592
rect 6932 70553 6960 71130
rect 7024 70990 7052 71130
rect 7012 70984 7064 70990
rect 7012 70926 7064 70932
rect 7104 70984 7156 70990
rect 7208 70972 7236 71352
rect 7300 71194 7328 71590
rect 7380 71528 7432 71534
rect 7380 71470 7432 71476
rect 7288 71188 7340 71194
rect 7288 71130 7340 71136
rect 7208 70944 7328 70972
rect 7104 70926 7156 70932
rect 7024 70582 7052 70926
rect 7012 70576 7064 70582
rect 6918 70544 6974 70553
rect 7012 70518 7064 70524
rect 7116 70514 7144 70926
rect 7196 70848 7248 70854
rect 7196 70790 7248 70796
rect 6918 70479 6920 70488
rect 6972 70479 6974 70488
rect 7104 70508 7156 70514
rect 6920 70450 6972 70456
rect 7104 70450 7156 70456
rect 6810 70204 7118 70213
rect 6810 70202 6816 70204
rect 6872 70202 6896 70204
rect 6952 70202 6976 70204
rect 7032 70202 7056 70204
rect 7112 70202 7118 70204
rect 6872 70150 6874 70202
rect 7054 70150 7056 70202
rect 6810 70148 6816 70150
rect 6872 70148 6896 70150
rect 6952 70148 6976 70150
rect 7032 70148 7056 70150
rect 7112 70148 7118 70150
rect 6810 70139 7118 70148
rect 6920 70100 6972 70106
rect 6920 70042 6972 70048
rect 6828 69964 6880 69970
rect 6828 69906 6880 69912
rect 6736 69828 6788 69834
rect 6736 69770 6788 69776
rect 6840 69562 6868 69906
rect 6932 69562 6960 70042
rect 7208 70038 7236 70790
rect 7300 70038 7328 70944
rect 7392 70854 7420 71470
rect 7380 70848 7432 70854
rect 7380 70790 7432 70796
rect 7380 70508 7432 70514
rect 7380 70450 7432 70456
rect 7196 70032 7248 70038
rect 7196 69974 7248 69980
rect 7288 70032 7340 70038
rect 7288 69974 7340 69980
rect 7392 69902 7420 70450
rect 7196 69896 7248 69902
rect 7196 69838 7248 69844
rect 7288 69896 7340 69902
rect 7288 69838 7340 69844
rect 7380 69896 7432 69902
rect 7380 69838 7432 69844
rect 7104 69760 7156 69766
rect 7104 69702 7156 69708
rect 6828 69556 6880 69562
rect 6828 69498 6880 69504
rect 6920 69556 6972 69562
rect 6920 69498 6972 69504
rect 7116 69426 7144 69702
rect 7104 69420 7156 69426
rect 7104 69362 7156 69368
rect 6920 69352 6972 69358
rect 6920 69294 6972 69300
rect 6932 69222 6960 69294
rect 6920 69216 6972 69222
rect 6920 69158 6972 69164
rect 6810 69116 7118 69125
rect 6810 69114 6816 69116
rect 6872 69114 6896 69116
rect 6952 69114 6976 69116
rect 7032 69114 7056 69116
rect 7112 69114 7118 69116
rect 6872 69062 6874 69114
rect 7054 69062 7056 69114
rect 6810 69060 6816 69062
rect 6872 69060 6896 69062
rect 6952 69060 6976 69062
rect 7032 69060 7056 69062
rect 7112 69060 7118 69062
rect 6810 69051 7118 69060
rect 6656 68972 6868 69000
rect 6840 68932 6868 68972
rect 7012 68944 7064 68950
rect 6840 68904 7012 68932
rect 6472 68870 6679 68898
rect 7012 68886 7064 68892
rect 7104 68944 7156 68950
rect 7104 68886 7156 68892
rect 6460 68808 6512 68814
rect 6651 68806 6679 68870
rect 6736 68808 6788 68814
rect 6651 68778 6684 68806
rect 6512 68756 6592 68762
rect 6460 68750 6592 68756
rect 6472 68734 6592 68750
rect 6092 68672 6144 68678
rect 6092 68614 6144 68620
rect 6150 68572 6458 68581
rect 6150 68570 6156 68572
rect 6212 68570 6236 68572
rect 6292 68570 6316 68572
rect 6372 68570 6396 68572
rect 6452 68570 6458 68572
rect 6212 68518 6214 68570
rect 6394 68518 6396 68570
rect 6150 68516 6156 68518
rect 6212 68516 6236 68518
rect 6292 68516 6316 68518
rect 6372 68516 6396 68518
rect 6452 68516 6458 68518
rect 6150 68507 6458 68516
rect 6276 68468 6328 68474
rect 6276 68410 6328 68416
rect 6090 68368 6146 68377
rect 6090 68303 6146 68312
rect 6104 67726 6132 68303
rect 6184 68264 6236 68270
rect 6184 68206 6236 68212
rect 6092 67720 6144 67726
rect 6196 67697 6224 68206
rect 6092 67662 6144 67668
rect 6182 67688 6238 67697
rect 5920 67612 6040 67640
rect 6182 67623 6238 67632
rect 5920 67386 5948 67612
rect 6288 67572 6316 68410
rect 6460 68332 6512 68338
rect 6460 68274 6512 68280
rect 6012 67544 6316 67572
rect 6472 67572 6500 68274
rect 6564 68202 6592 68734
rect 6552 68196 6604 68202
rect 6552 68138 6604 68144
rect 6564 67794 6592 68138
rect 6552 67788 6604 67794
rect 6552 67730 6604 67736
rect 6656 67634 6684 68778
rect 7012 68808 7064 68814
rect 6788 68768 6868 68796
rect 6736 68750 6788 68756
rect 6736 68672 6788 68678
rect 6736 68614 6788 68620
rect 6748 68474 6776 68614
rect 6736 68468 6788 68474
rect 6736 68410 6788 68416
rect 6840 68202 6868 68768
rect 6932 68768 7012 68796
rect 6932 68241 6960 68768
rect 7012 68750 7064 68756
rect 7012 68400 7064 68406
rect 7116 68388 7144 68886
rect 7064 68360 7144 68388
rect 7012 68342 7064 68348
rect 6918 68232 6974 68241
rect 6828 68196 6880 68202
rect 6748 68156 6828 68184
rect 6748 67844 6776 68156
rect 6918 68167 6974 68176
rect 6828 68138 6880 68144
rect 6810 68028 7118 68037
rect 6810 68026 6816 68028
rect 6872 68026 6896 68028
rect 6952 68026 6976 68028
rect 7032 68026 7056 68028
rect 7112 68026 7118 68028
rect 6872 67974 6874 68026
rect 7054 67974 7056 68026
rect 6810 67972 6816 67974
rect 6872 67972 6896 67974
rect 6952 67972 6976 67974
rect 7032 67972 7056 67974
rect 7112 67972 7118 67974
rect 6810 67963 7118 67972
rect 6840 67884 7144 67912
rect 6840 67844 6868 67884
rect 6748 67816 6868 67844
rect 7116 67658 7144 67884
rect 6920 67652 6972 67658
rect 6656 67606 6776 67634
rect 6472 67544 6684 67572
rect 5908 67380 5960 67386
rect 6012 67368 6040 67544
rect 6150 67484 6458 67493
rect 6150 67482 6156 67484
rect 6212 67482 6236 67484
rect 6292 67482 6316 67484
rect 6372 67482 6396 67484
rect 6452 67482 6458 67484
rect 6212 67430 6214 67482
rect 6394 67430 6396 67482
rect 6150 67428 6156 67430
rect 6212 67428 6236 67430
rect 6292 67428 6316 67430
rect 6372 67428 6396 67430
rect 6452 67428 6458 67430
rect 6150 67419 6458 67428
rect 6460 67380 6512 67386
rect 6012 67340 6224 67368
rect 5908 67322 5960 67328
rect 6092 67176 6144 67182
rect 6092 67118 6144 67124
rect 6000 67108 6052 67114
rect 6000 67050 6052 67056
rect 5908 67040 5960 67046
rect 5908 66982 5960 66988
rect 5920 66774 5948 66982
rect 5908 66768 5960 66774
rect 5908 66710 5960 66716
rect 5908 66632 5960 66638
rect 5908 66574 5960 66580
rect 5816 66156 5868 66162
rect 5816 66098 5868 66104
rect 5816 66020 5868 66026
rect 5460 65980 5672 66008
rect 5368 65912 5580 65940
rect 5210 65852 5518 65861
rect 5210 65850 5216 65852
rect 5272 65850 5296 65852
rect 5352 65850 5376 65852
rect 5432 65850 5456 65852
rect 5512 65850 5518 65852
rect 5272 65798 5274 65850
rect 5454 65798 5456 65850
rect 5210 65796 5216 65798
rect 5272 65796 5296 65798
rect 5352 65796 5376 65798
rect 5432 65796 5456 65798
rect 5512 65796 5518 65798
rect 5210 65787 5518 65796
rect 5354 65648 5410 65657
rect 5354 65583 5410 65592
rect 5080 65476 5132 65482
rect 4620 65408 4672 65414
rect 4620 65350 4672 65356
rect 4550 65308 4858 65317
rect 4550 65306 4556 65308
rect 4612 65306 4636 65308
rect 4692 65306 4716 65308
rect 4772 65306 4796 65308
rect 4852 65306 4858 65308
rect 4612 65254 4614 65306
rect 4794 65254 4796 65306
rect 4550 65252 4556 65254
rect 4612 65252 4636 65254
rect 4692 65252 4716 65254
rect 4772 65252 4796 65254
rect 4852 65252 4858 65254
rect 4550 65243 4858 65252
rect 4908 65090 4936 65470
rect 5080 65418 5132 65424
rect 5172 65408 5224 65414
rect 5172 65350 5224 65356
rect 5080 65204 5132 65210
rect 4712 65068 4764 65074
rect 4712 65010 4764 65016
rect 4816 65062 4936 65090
rect 5000 65164 5080 65192
rect 4724 64326 4752 65010
rect 4816 64666 4844 65062
rect 4896 64864 4948 64870
rect 4896 64806 4948 64812
rect 4804 64660 4856 64666
rect 4804 64602 4856 64608
rect 4712 64320 4764 64326
rect 4712 64262 4764 64268
rect 4550 64220 4858 64229
rect 4550 64218 4556 64220
rect 4612 64218 4636 64220
rect 4692 64218 4716 64220
rect 4772 64218 4796 64220
rect 4852 64218 4858 64220
rect 4612 64166 4614 64218
rect 4794 64166 4796 64218
rect 4550 64164 4556 64166
rect 4612 64164 4636 64166
rect 4692 64164 4716 64166
rect 4772 64164 4796 64166
rect 4852 64164 4858 64166
rect 4550 64155 4858 64164
rect 4804 64116 4856 64122
rect 4804 64058 4856 64064
rect 4816 63510 4844 64058
rect 4804 63504 4856 63510
rect 4804 63446 4856 63452
rect 4550 63132 4858 63141
rect 4550 63130 4556 63132
rect 4612 63130 4636 63132
rect 4692 63130 4716 63132
rect 4772 63130 4796 63132
rect 4852 63130 4858 63132
rect 4612 63078 4614 63130
rect 4794 63078 4796 63130
rect 4550 63076 4556 63078
rect 4612 63076 4636 63078
rect 4692 63076 4716 63078
rect 4772 63076 4796 63078
rect 4852 63076 4858 63078
rect 4550 63067 4858 63076
rect 4908 63016 4936 64806
rect 4724 62988 4936 63016
rect 4724 62218 4752 62988
rect 4804 62892 4856 62898
rect 4804 62834 4856 62840
rect 4816 62268 4844 62834
rect 4816 62240 4936 62268
rect 4712 62212 4764 62218
rect 4712 62154 4764 62160
rect 4550 62044 4858 62053
rect 4550 62042 4556 62044
rect 4612 62042 4636 62044
rect 4692 62042 4716 62044
rect 4772 62042 4796 62044
rect 4852 62042 4858 62044
rect 4612 61990 4614 62042
rect 4794 61990 4796 62042
rect 4550 61988 4556 61990
rect 4612 61988 4636 61990
rect 4692 61988 4716 61990
rect 4772 61988 4796 61990
rect 4852 61988 4858 61990
rect 4550 61979 4858 61988
rect 4550 60956 4858 60965
rect 4550 60954 4556 60956
rect 4612 60954 4636 60956
rect 4692 60954 4716 60956
rect 4772 60954 4796 60956
rect 4852 60954 4858 60956
rect 4612 60902 4614 60954
rect 4794 60902 4796 60954
rect 4550 60900 4556 60902
rect 4612 60900 4636 60902
rect 4692 60900 4716 60902
rect 4772 60900 4796 60902
rect 4852 60900 4858 60902
rect 4550 60891 4858 60900
rect 4804 60784 4856 60790
rect 4908 60772 4936 62240
rect 4856 60744 4936 60772
rect 4804 60726 4856 60732
rect 4436 60716 4488 60722
rect 4436 60658 4488 60664
rect 5000 60602 5028 65164
rect 5080 65146 5132 65152
rect 5184 65006 5212 65350
rect 5172 65000 5224 65006
rect 5172 64942 5224 64948
rect 5368 64938 5396 65583
rect 5356 64932 5408 64938
rect 5356 64874 5408 64880
rect 5080 64864 5132 64870
rect 5080 64806 5132 64812
rect 5092 64530 5120 64806
rect 5210 64764 5518 64773
rect 5210 64762 5216 64764
rect 5272 64762 5296 64764
rect 5352 64762 5376 64764
rect 5432 64762 5456 64764
rect 5512 64762 5518 64764
rect 5272 64710 5274 64762
rect 5454 64710 5456 64762
rect 5210 64708 5216 64710
rect 5272 64708 5296 64710
rect 5352 64708 5376 64710
rect 5432 64708 5456 64710
rect 5512 64708 5518 64710
rect 5210 64699 5518 64708
rect 5172 64660 5224 64666
rect 5172 64602 5224 64608
rect 5080 64524 5132 64530
rect 5080 64466 5132 64472
rect 5080 64320 5132 64326
rect 5080 64262 5132 64268
rect 5092 61282 5120 64262
rect 5184 64122 5212 64602
rect 5172 64116 5224 64122
rect 5172 64058 5224 64064
rect 5552 63782 5580 65912
rect 5644 65754 5672 65980
rect 5816 65962 5868 65968
rect 5632 65748 5684 65754
rect 5632 65690 5684 65696
rect 5724 65612 5776 65618
rect 5724 65554 5776 65560
rect 5632 65476 5684 65482
rect 5632 65418 5684 65424
rect 5540 63776 5592 63782
rect 5540 63718 5592 63724
rect 5210 63676 5518 63685
rect 5210 63674 5216 63676
rect 5272 63674 5296 63676
rect 5352 63674 5376 63676
rect 5432 63674 5456 63676
rect 5512 63674 5518 63676
rect 5272 63622 5274 63674
rect 5454 63622 5456 63674
rect 5210 63620 5216 63622
rect 5272 63620 5296 63622
rect 5352 63620 5376 63622
rect 5432 63620 5456 63622
rect 5512 63620 5518 63622
rect 5210 63611 5518 63620
rect 5172 63504 5224 63510
rect 5172 63446 5224 63452
rect 5184 62830 5212 63446
rect 5448 63436 5500 63442
rect 5448 63378 5500 63384
rect 5460 62830 5488 63378
rect 5540 63232 5592 63238
rect 5540 63174 5592 63180
rect 5172 62824 5224 62830
rect 5172 62766 5224 62772
rect 5448 62824 5500 62830
rect 5448 62766 5500 62772
rect 5210 62588 5518 62597
rect 5210 62586 5216 62588
rect 5272 62586 5296 62588
rect 5352 62586 5376 62588
rect 5432 62586 5456 62588
rect 5512 62586 5518 62588
rect 5272 62534 5274 62586
rect 5454 62534 5456 62586
rect 5210 62532 5216 62534
rect 5272 62532 5296 62534
rect 5352 62532 5376 62534
rect 5432 62532 5456 62534
rect 5512 62532 5518 62534
rect 5210 62523 5518 62532
rect 5448 62212 5500 62218
rect 5448 62154 5500 62160
rect 5460 61946 5488 62154
rect 5448 61940 5500 61946
rect 5448 61882 5500 61888
rect 5210 61500 5518 61509
rect 5210 61498 5216 61500
rect 5272 61498 5296 61500
rect 5352 61498 5376 61500
rect 5432 61498 5456 61500
rect 5512 61498 5518 61500
rect 5272 61446 5274 61498
rect 5454 61446 5456 61498
rect 5210 61444 5216 61446
rect 5272 61444 5296 61446
rect 5352 61444 5376 61446
rect 5432 61444 5456 61446
rect 5512 61444 5518 61446
rect 5210 61435 5518 61444
rect 5092 61254 5396 61282
rect 5264 61192 5316 61198
rect 5264 61134 5316 61140
rect 5172 61124 5224 61130
rect 5172 61066 5224 61072
rect 5184 60602 5212 61066
rect 4816 60574 5028 60602
rect 5092 60574 5212 60602
rect 4436 60512 4488 60518
rect 4436 60454 4488 60460
rect 4344 59084 4396 59090
rect 4344 59026 4396 59032
rect 4252 59016 4304 59022
rect 4448 58970 4476 60454
rect 4816 60314 4844 60574
rect 4896 60512 4948 60518
rect 5092 60466 5120 60574
rect 5276 60518 5304 61134
rect 5368 60518 5396 61254
rect 4896 60454 4948 60460
rect 4804 60308 4856 60314
rect 4804 60250 4856 60256
rect 4550 59868 4858 59877
rect 4550 59866 4556 59868
rect 4612 59866 4636 59868
rect 4692 59866 4716 59868
rect 4772 59866 4796 59868
rect 4852 59866 4858 59868
rect 4612 59814 4614 59866
rect 4794 59814 4796 59866
rect 4550 59812 4556 59814
rect 4612 59812 4636 59814
rect 4692 59812 4716 59814
rect 4772 59812 4796 59814
rect 4852 59812 4858 59814
rect 4550 59803 4858 59812
rect 4908 59752 4936 60454
rect 4816 59724 4936 59752
rect 5000 60438 5120 60466
rect 5264 60512 5316 60518
rect 5264 60454 5316 60460
rect 5356 60512 5408 60518
rect 5356 60454 5408 60460
rect 4528 59424 4580 59430
rect 4528 59366 4580 59372
rect 4540 59022 4568 59366
rect 4252 58958 4304 58964
rect 4160 57588 4212 57594
rect 4160 57530 4212 57536
rect 4264 57338 4292 58958
rect 4172 57310 4292 57338
rect 4356 58942 4476 58970
rect 4528 59016 4580 59022
rect 4528 58958 4580 58964
rect 4356 57322 4384 58942
rect 4816 58868 4844 59724
rect 4896 59560 4948 59566
rect 4896 59502 4948 59508
rect 4908 59022 4936 59502
rect 4896 59016 4948 59022
rect 4896 58958 4948 58964
rect 4448 58840 4844 58868
rect 4448 57526 4476 58840
rect 4550 58780 4858 58789
rect 4550 58778 4556 58780
rect 4612 58778 4636 58780
rect 4692 58778 4716 58780
rect 4772 58778 4796 58780
rect 4852 58778 4858 58780
rect 4612 58726 4614 58778
rect 4794 58726 4796 58778
rect 4550 58724 4556 58726
rect 4612 58724 4636 58726
rect 4692 58724 4716 58726
rect 4772 58724 4796 58726
rect 4852 58724 4858 58726
rect 4550 58715 4858 58724
rect 4908 58546 4936 58958
rect 4896 58540 4948 58546
rect 4896 58482 4948 58488
rect 4896 58404 4948 58410
rect 4896 58346 4948 58352
rect 4908 58138 4936 58346
rect 4896 58132 4948 58138
rect 4896 58074 4948 58080
rect 4550 57692 4858 57701
rect 4550 57690 4556 57692
rect 4612 57690 4636 57692
rect 4692 57690 4716 57692
rect 4772 57690 4796 57692
rect 4852 57690 4858 57692
rect 4612 57638 4614 57690
rect 4794 57638 4796 57690
rect 4550 57636 4556 57638
rect 4612 57636 4636 57638
rect 4692 57636 4716 57638
rect 4772 57636 4796 57638
rect 4852 57636 4858 57638
rect 4550 57627 4858 57636
rect 4436 57520 4488 57526
rect 4436 57462 4488 57468
rect 4896 57520 4948 57526
rect 4896 57462 4948 57468
rect 4344 57316 4396 57322
rect 4172 54233 4200 57310
rect 4344 57258 4396 57264
rect 4436 57316 4488 57322
rect 4436 57258 4488 57264
rect 4252 57248 4304 57254
rect 4252 57190 4304 57196
rect 4158 54224 4214 54233
rect 4158 54159 4214 54168
rect 4172 53582 4200 54159
rect 4160 53576 4212 53582
rect 4160 53518 4212 53524
rect 4160 53100 4212 53106
rect 4160 53042 4212 53048
rect 4172 48890 4200 53042
rect 4264 52426 4292 57190
rect 4252 52420 4304 52426
rect 4252 52362 4304 52368
rect 4252 51264 4304 51270
rect 4252 51206 4304 51212
rect 4160 48884 4212 48890
rect 4160 48826 4212 48832
rect 4264 48634 4292 51206
rect 4356 50250 4384 57258
rect 4448 56370 4476 57258
rect 4550 56604 4858 56613
rect 4550 56602 4556 56604
rect 4612 56602 4636 56604
rect 4692 56602 4716 56604
rect 4772 56602 4796 56604
rect 4852 56602 4858 56604
rect 4612 56550 4614 56602
rect 4794 56550 4796 56602
rect 4550 56548 4556 56550
rect 4612 56548 4636 56550
rect 4692 56548 4716 56550
rect 4772 56548 4796 56550
rect 4852 56548 4858 56550
rect 4550 56539 4858 56548
rect 4436 56364 4488 56370
rect 4436 56306 4488 56312
rect 4436 55684 4488 55690
rect 4436 55626 4488 55632
rect 4448 53582 4476 55626
rect 4550 55516 4858 55525
rect 4550 55514 4556 55516
rect 4612 55514 4636 55516
rect 4692 55514 4716 55516
rect 4772 55514 4796 55516
rect 4852 55514 4858 55516
rect 4612 55462 4614 55514
rect 4794 55462 4796 55514
rect 4550 55460 4556 55462
rect 4612 55460 4636 55462
rect 4692 55460 4716 55462
rect 4772 55460 4796 55462
rect 4852 55460 4858 55462
rect 4550 55451 4858 55460
rect 4550 54428 4858 54437
rect 4550 54426 4556 54428
rect 4612 54426 4636 54428
rect 4692 54426 4716 54428
rect 4772 54426 4796 54428
rect 4852 54426 4858 54428
rect 4612 54374 4614 54426
rect 4794 54374 4796 54426
rect 4550 54372 4556 54374
rect 4612 54372 4636 54374
rect 4692 54372 4716 54374
rect 4772 54372 4796 54374
rect 4852 54372 4858 54374
rect 4550 54363 4858 54372
rect 4908 53786 4936 57462
rect 5000 56370 5028 60438
rect 5210 60412 5518 60421
rect 5210 60410 5216 60412
rect 5272 60410 5296 60412
rect 5352 60410 5376 60412
rect 5432 60410 5456 60412
rect 5512 60410 5518 60412
rect 5272 60358 5274 60410
rect 5454 60358 5456 60410
rect 5210 60356 5216 60358
rect 5272 60356 5296 60358
rect 5352 60356 5376 60358
rect 5432 60356 5456 60358
rect 5512 60356 5518 60358
rect 5210 60347 5518 60356
rect 5080 60308 5132 60314
rect 5080 60250 5132 60256
rect 5092 59208 5120 60250
rect 5210 59324 5518 59333
rect 5210 59322 5216 59324
rect 5272 59322 5296 59324
rect 5352 59322 5376 59324
rect 5432 59322 5456 59324
rect 5512 59322 5518 59324
rect 5272 59270 5274 59322
rect 5454 59270 5456 59322
rect 5210 59268 5216 59270
rect 5272 59268 5296 59270
rect 5352 59268 5376 59270
rect 5432 59268 5456 59270
rect 5512 59268 5518 59270
rect 5210 59259 5518 59268
rect 5092 59180 5212 59208
rect 5080 58880 5132 58886
rect 5080 58822 5132 58828
rect 5092 56370 5120 58822
rect 5184 58410 5212 59180
rect 5172 58404 5224 58410
rect 5172 58346 5224 58352
rect 5210 58236 5518 58245
rect 5210 58234 5216 58236
rect 5272 58234 5296 58236
rect 5352 58234 5376 58236
rect 5432 58234 5456 58236
rect 5512 58234 5518 58236
rect 5272 58182 5274 58234
rect 5454 58182 5456 58234
rect 5210 58180 5216 58182
rect 5272 58180 5296 58182
rect 5352 58180 5376 58182
rect 5432 58180 5456 58182
rect 5512 58180 5518 58182
rect 5210 58171 5518 58180
rect 5172 58132 5224 58138
rect 5172 58074 5224 58080
rect 5184 57594 5212 58074
rect 5552 57974 5580 63174
rect 5368 57946 5580 57974
rect 5172 57588 5224 57594
rect 5172 57530 5224 57536
rect 5368 57322 5396 57946
rect 5448 57792 5500 57798
rect 5448 57734 5500 57740
rect 5356 57316 5408 57322
rect 5356 57258 5408 57264
rect 5460 57236 5488 57734
rect 5644 57322 5672 65418
rect 5736 64530 5764 65554
rect 5724 64524 5776 64530
rect 5724 64466 5776 64472
rect 5736 63986 5764 64466
rect 5828 64462 5856 65962
rect 5816 64456 5868 64462
rect 5816 64398 5868 64404
rect 5816 64320 5868 64326
rect 5816 64262 5868 64268
rect 5828 64122 5856 64262
rect 5816 64116 5868 64122
rect 5816 64058 5868 64064
rect 5724 63980 5776 63986
rect 5724 63922 5776 63928
rect 5920 63866 5948 66574
rect 6012 66162 6040 67050
rect 6104 66502 6132 67118
rect 6196 66570 6224 67340
rect 6460 67322 6512 67328
rect 6552 67380 6604 67386
rect 6552 67322 6604 67328
rect 6472 66706 6500 67322
rect 6460 66700 6512 66706
rect 6460 66642 6512 66648
rect 6564 66570 6592 67322
rect 6184 66564 6236 66570
rect 6184 66506 6236 66512
rect 6552 66564 6604 66570
rect 6552 66506 6604 66512
rect 6092 66496 6144 66502
rect 6092 66438 6144 66444
rect 6150 66396 6458 66405
rect 6150 66394 6156 66396
rect 6212 66394 6236 66396
rect 6292 66394 6316 66396
rect 6372 66394 6396 66396
rect 6452 66394 6458 66396
rect 6212 66342 6214 66394
rect 6394 66342 6396 66394
rect 6150 66340 6156 66342
rect 6212 66340 6236 66342
rect 6292 66340 6316 66342
rect 6372 66340 6396 66342
rect 6452 66340 6458 66342
rect 6150 66331 6458 66340
rect 6000 66156 6052 66162
rect 6000 66098 6052 66104
rect 6276 66088 6328 66094
rect 6276 66030 6328 66036
rect 6000 65544 6052 65550
rect 6000 65486 6052 65492
rect 5736 63838 5948 63866
rect 5736 59702 5764 63838
rect 5816 63776 5868 63782
rect 5816 63718 5868 63724
rect 5828 61198 5856 63718
rect 6012 63594 6040 65486
rect 6288 65414 6316 66030
rect 6276 65408 6328 65414
rect 6276 65350 6328 65356
rect 6150 65308 6458 65317
rect 6150 65306 6156 65308
rect 6212 65306 6236 65308
rect 6292 65306 6316 65308
rect 6372 65306 6396 65308
rect 6452 65306 6458 65308
rect 6212 65254 6214 65306
rect 6394 65254 6396 65306
rect 6150 65252 6156 65254
rect 6212 65252 6236 65254
rect 6292 65252 6316 65254
rect 6372 65252 6396 65254
rect 6452 65252 6458 65254
rect 6150 65243 6458 65252
rect 6564 65074 6592 66506
rect 6552 65068 6604 65074
rect 6552 65010 6604 65016
rect 6092 64932 6144 64938
rect 6092 64874 6144 64880
rect 6104 64326 6132 64874
rect 6552 64864 6604 64870
rect 6552 64806 6604 64812
rect 6092 64320 6144 64326
rect 6092 64262 6144 64268
rect 6150 64220 6458 64229
rect 6150 64218 6156 64220
rect 6212 64218 6236 64220
rect 6292 64218 6316 64220
rect 6372 64218 6396 64220
rect 6452 64218 6458 64220
rect 6212 64166 6214 64218
rect 6394 64166 6396 64218
rect 6150 64164 6156 64166
rect 6212 64164 6236 64166
rect 6292 64164 6316 64166
rect 6372 64164 6396 64166
rect 6452 64164 6458 64166
rect 6150 64155 6458 64164
rect 6276 64116 6328 64122
rect 6276 64058 6328 64064
rect 6092 63980 6144 63986
rect 6092 63922 6144 63928
rect 5920 63566 6040 63594
rect 5816 61192 5868 61198
rect 5816 61134 5868 61140
rect 5816 61056 5868 61062
rect 5816 60998 5868 61004
rect 5724 59696 5776 59702
rect 5724 59638 5776 59644
rect 5724 58948 5776 58954
rect 5724 58890 5776 58896
rect 5736 58682 5764 58890
rect 5724 58676 5776 58682
rect 5724 58618 5776 58624
rect 5724 58404 5776 58410
rect 5724 58346 5776 58352
rect 5632 57316 5684 57322
rect 5632 57258 5684 57264
rect 5460 57208 5580 57236
rect 5552 57202 5580 57208
rect 5552 57174 5672 57202
rect 5210 57148 5518 57157
rect 5210 57146 5216 57148
rect 5272 57146 5296 57148
rect 5352 57146 5376 57148
rect 5432 57146 5456 57148
rect 5512 57146 5518 57148
rect 5272 57094 5274 57146
rect 5454 57094 5456 57146
rect 5210 57092 5216 57094
rect 5272 57092 5296 57094
rect 5352 57092 5376 57094
rect 5432 57092 5456 57094
rect 5512 57092 5518 57094
rect 5210 57083 5518 57092
rect 4988 56364 5040 56370
rect 4988 56306 5040 56312
rect 5080 56364 5132 56370
rect 5080 56306 5132 56312
rect 5080 56160 5132 56166
rect 5080 56102 5132 56108
rect 4896 53780 4948 53786
rect 4896 53722 4948 53728
rect 4804 53712 4856 53718
rect 4804 53654 4856 53660
rect 4436 53576 4488 53582
rect 4436 53518 4488 53524
rect 4816 53530 4844 53654
rect 4344 50244 4396 50250
rect 4344 50186 4396 50192
rect 4448 50130 4476 53518
rect 4816 53502 4936 53530
rect 4550 53340 4858 53349
rect 4550 53338 4556 53340
rect 4612 53338 4636 53340
rect 4692 53338 4716 53340
rect 4772 53338 4796 53340
rect 4852 53338 4858 53340
rect 4612 53286 4614 53338
rect 4794 53286 4796 53338
rect 4550 53284 4556 53286
rect 4612 53284 4636 53286
rect 4692 53284 4716 53286
rect 4772 53284 4796 53286
rect 4852 53284 4858 53286
rect 4550 53275 4858 53284
rect 4804 53100 4856 53106
rect 4804 53042 4856 53048
rect 4816 52902 4844 53042
rect 4804 52896 4856 52902
rect 4804 52838 4856 52844
rect 4550 52252 4858 52261
rect 4550 52250 4556 52252
rect 4612 52250 4636 52252
rect 4692 52250 4716 52252
rect 4772 52250 4796 52252
rect 4852 52250 4858 52252
rect 4612 52198 4614 52250
rect 4794 52198 4796 52250
rect 4550 52196 4556 52198
rect 4612 52196 4636 52198
rect 4692 52196 4716 52198
rect 4772 52196 4796 52198
rect 4852 52196 4858 52198
rect 4550 52187 4858 52196
rect 4804 52148 4856 52154
rect 4804 52090 4856 52096
rect 4816 51354 4844 52090
rect 4908 51474 4936 53502
rect 5092 53174 5120 56102
rect 5210 56060 5518 56069
rect 5210 56058 5216 56060
rect 5272 56058 5296 56060
rect 5352 56058 5376 56060
rect 5432 56058 5456 56060
rect 5512 56058 5518 56060
rect 5272 56006 5274 56058
rect 5454 56006 5456 56058
rect 5210 56004 5216 56006
rect 5272 56004 5296 56006
rect 5352 56004 5376 56006
rect 5432 56004 5456 56006
rect 5512 56004 5518 56006
rect 5210 55995 5518 56004
rect 5540 55616 5592 55622
rect 5540 55558 5592 55564
rect 5210 54972 5518 54981
rect 5210 54970 5216 54972
rect 5272 54970 5296 54972
rect 5352 54970 5376 54972
rect 5432 54970 5456 54972
rect 5512 54970 5518 54972
rect 5272 54918 5274 54970
rect 5454 54918 5456 54970
rect 5210 54916 5216 54918
rect 5272 54916 5296 54918
rect 5352 54916 5376 54918
rect 5432 54916 5456 54918
rect 5512 54916 5518 54918
rect 5210 54907 5518 54916
rect 5210 53884 5518 53893
rect 5210 53882 5216 53884
rect 5272 53882 5296 53884
rect 5352 53882 5376 53884
rect 5432 53882 5456 53884
rect 5512 53882 5518 53884
rect 5272 53830 5274 53882
rect 5454 53830 5456 53882
rect 5210 53828 5216 53830
rect 5272 53828 5296 53830
rect 5352 53828 5376 53830
rect 5432 53828 5456 53830
rect 5512 53828 5518 53830
rect 5210 53819 5518 53828
rect 5080 53168 5132 53174
rect 5000 53128 5080 53156
rect 4896 51468 4948 51474
rect 4896 51410 4948 51416
rect 4816 51326 4936 51354
rect 4550 51164 4858 51173
rect 4550 51162 4556 51164
rect 4612 51162 4636 51164
rect 4692 51162 4716 51164
rect 4772 51162 4796 51164
rect 4852 51162 4858 51164
rect 4612 51110 4614 51162
rect 4794 51110 4796 51162
rect 4550 51108 4556 51110
rect 4612 51108 4636 51110
rect 4692 51108 4716 51110
rect 4772 51108 4796 51110
rect 4852 51108 4858 51110
rect 4550 51099 4858 51108
rect 4356 50102 4476 50130
rect 4356 49774 4384 50102
rect 4550 50076 4858 50085
rect 4550 50074 4556 50076
rect 4612 50074 4636 50076
rect 4692 50074 4716 50076
rect 4772 50074 4796 50076
rect 4852 50074 4858 50076
rect 4612 50022 4614 50074
rect 4794 50022 4796 50074
rect 4550 50020 4556 50022
rect 4612 50020 4636 50022
rect 4692 50020 4716 50022
rect 4772 50020 4796 50022
rect 4852 50020 4858 50022
rect 4550 50011 4858 50020
rect 4436 49972 4488 49978
rect 4436 49914 4488 49920
rect 4344 49768 4396 49774
rect 4344 49710 4396 49716
rect 4344 49632 4396 49638
rect 4344 49574 4396 49580
rect 4172 48606 4292 48634
rect 4172 45830 4200 48606
rect 4252 48544 4304 48550
rect 4252 48486 4304 48492
rect 4264 46986 4292 48486
rect 4252 46980 4304 46986
rect 4252 46922 4304 46928
rect 4356 46458 4384 49574
rect 4448 47025 4476 49914
rect 4712 49904 4764 49910
rect 4712 49846 4764 49852
rect 4724 49434 4752 49846
rect 4908 49756 4936 51326
rect 5000 49858 5028 53128
rect 5080 53110 5132 53116
rect 5080 52896 5132 52902
rect 5080 52838 5132 52844
rect 5092 51490 5120 52838
rect 5210 52796 5518 52805
rect 5210 52794 5216 52796
rect 5272 52794 5296 52796
rect 5352 52794 5376 52796
rect 5432 52794 5456 52796
rect 5512 52794 5518 52796
rect 5272 52742 5274 52794
rect 5454 52742 5456 52794
rect 5210 52740 5216 52742
rect 5272 52740 5296 52742
rect 5352 52740 5376 52742
rect 5432 52740 5456 52742
rect 5512 52740 5518 52742
rect 5210 52731 5518 52740
rect 5210 51708 5518 51717
rect 5210 51706 5216 51708
rect 5272 51706 5296 51708
rect 5352 51706 5376 51708
rect 5432 51706 5456 51708
rect 5512 51706 5518 51708
rect 5272 51654 5274 51706
rect 5454 51654 5456 51706
rect 5210 51652 5216 51654
rect 5272 51652 5296 51654
rect 5352 51652 5376 51654
rect 5432 51652 5456 51654
rect 5512 51652 5518 51654
rect 5210 51643 5518 51652
rect 5092 51462 5212 51490
rect 5080 51400 5132 51406
rect 5080 51342 5132 51348
rect 5092 49978 5120 51342
rect 5184 51074 5212 51462
rect 5184 51046 5488 51074
rect 5460 50708 5488 51046
rect 5552 50776 5580 55558
rect 5644 53122 5672 57174
rect 5736 53242 5764 58346
rect 5828 54262 5856 60998
rect 5920 58954 5948 63566
rect 6000 63504 6052 63510
rect 6000 63446 6052 63452
rect 6012 63034 6040 63446
rect 6104 63442 6132 63922
rect 6092 63436 6144 63442
rect 6092 63378 6144 63384
rect 6288 63374 6316 64058
rect 6368 63776 6420 63782
rect 6368 63718 6420 63724
rect 6276 63368 6328 63374
rect 6276 63310 6328 63316
rect 6380 63220 6408 63718
rect 6564 63510 6592 64806
rect 6552 63504 6604 63510
rect 6552 63446 6604 63452
rect 6564 63345 6592 63446
rect 6550 63336 6606 63345
rect 6550 63271 6606 63280
rect 6380 63192 6592 63220
rect 6150 63132 6458 63141
rect 6150 63130 6156 63132
rect 6212 63130 6236 63132
rect 6292 63130 6316 63132
rect 6372 63130 6396 63132
rect 6452 63130 6458 63132
rect 6212 63078 6214 63130
rect 6394 63078 6396 63130
rect 6150 63076 6156 63078
rect 6212 63076 6236 63078
rect 6292 63076 6316 63078
rect 6372 63076 6396 63078
rect 6452 63076 6458 63078
rect 6150 63067 6458 63076
rect 6000 63028 6052 63034
rect 6564 63016 6592 63192
rect 6000 62970 6052 62976
rect 6472 62988 6592 63016
rect 6092 62892 6144 62898
rect 6092 62834 6144 62840
rect 6104 62218 6132 62834
rect 6472 62490 6500 62988
rect 6552 62892 6604 62898
rect 6552 62834 6604 62840
rect 6460 62484 6512 62490
rect 6460 62426 6512 62432
rect 6092 62212 6144 62218
rect 6092 62154 6144 62160
rect 6000 62144 6052 62150
rect 6000 62086 6052 62092
rect 5908 58948 5960 58954
rect 5908 58890 5960 58896
rect 5908 58336 5960 58342
rect 5908 58278 5960 58284
rect 5816 54256 5868 54262
rect 5816 54198 5868 54204
rect 5724 53236 5776 53242
rect 5724 53178 5776 53184
rect 5644 53094 5856 53122
rect 5632 53032 5684 53038
rect 5632 52974 5684 52980
rect 5644 50930 5672 52974
rect 5724 52692 5776 52698
rect 5724 52634 5776 52640
rect 5632 50924 5684 50930
rect 5632 50866 5684 50872
rect 5552 50748 5672 50776
rect 5460 50680 5580 50708
rect 5210 50620 5518 50629
rect 5210 50618 5216 50620
rect 5272 50618 5296 50620
rect 5352 50618 5376 50620
rect 5432 50618 5456 50620
rect 5512 50618 5518 50620
rect 5272 50566 5274 50618
rect 5454 50566 5456 50618
rect 5210 50564 5216 50566
rect 5272 50564 5296 50566
rect 5352 50564 5376 50566
rect 5432 50564 5456 50566
rect 5512 50564 5518 50566
rect 5210 50555 5518 50564
rect 5552 50402 5580 50680
rect 5460 50374 5580 50402
rect 5080 49972 5132 49978
rect 5080 49914 5132 49920
rect 5000 49830 5120 49858
rect 4908 49728 5028 49756
rect 4896 49632 4948 49638
rect 4896 49574 4948 49580
rect 4712 49428 4764 49434
rect 4712 49370 4764 49376
rect 4550 48988 4858 48997
rect 4550 48986 4556 48988
rect 4612 48986 4636 48988
rect 4692 48986 4716 48988
rect 4772 48986 4796 48988
rect 4852 48986 4858 48988
rect 4612 48934 4614 48986
rect 4794 48934 4796 48986
rect 4550 48932 4556 48934
rect 4612 48932 4636 48934
rect 4692 48932 4716 48934
rect 4772 48932 4796 48934
rect 4852 48932 4858 48934
rect 4550 48923 4858 48932
rect 4908 48890 4936 49574
rect 4804 48884 4856 48890
rect 4804 48826 4856 48832
rect 4896 48884 4948 48890
rect 4896 48826 4948 48832
rect 4712 48612 4764 48618
rect 4712 48554 4764 48560
rect 4724 48346 4752 48554
rect 4712 48340 4764 48346
rect 4712 48282 4764 48288
rect 4816 48314 4844 48826
rect 4816 48286 4936 48314
rect 4550 47900 4858 47909
rect 4550 47898 4556 47900
rect 4612 47898 4636 47900
rect 4692 47898 4716 47900
rect 4772 47898 4796 47900
rect 4852 47898 4858 47900
rect 4612 47846 4614 47898
rect 4794 47846 4796 47898
rect 4550 47844 4556 47846
rect 4612 47844 4636 47846
rect 4692 47844 4716 47846
rect 4772 47844 4796 47846
rect 4852 47844 4858 47846
rect 4550 47835 4858 47844
rect 4908 47682 4936 48286
rect 4816 47654 4936 47682
rect 4434 47016 4490 47025
rect 4434 46951 4490 46960
rect 4816 46900 4844 47654
rect 4896 47524 4948 47530
rect 4896 47466 4948 47472
rect 4448 46872 4844 46900
rect 4448 46696 4476 46872
rect 4550 46812 4858 46821
rect 4550 46810 4556 46812
rect 4612 46810 4636 46812
rect 4692 46810 4716 46812
rect 4772 46810 4796 46812
rect 4852 46810 4858 46812
rect 4612 46758 4614 46810
rect 4794 46758 4796 46810
rect 4550 46756 4556 46758
rect 4612 46756 4636 46758
rect 4692 46756 4716 46758
rect 4772 46756 4796 46758
rect 4852 46756 4858 46758
rect 4550 46747 4858 46756
rect 4448 46668 4568 46696
rect 4434 46608 4490 46617
rect 4434 46543 4490 46552
rect 4264 46430 4384 46458
rect 4160 45824 4212 45830
rect 4160 45766 4212 45772
rect 4066 45520 4122 45529
rect 4264 45490 4292 46430
rect 4344 46368 4396 46374
rect 4344 46310 4396 46316
rect 4066 45455 4122 45464
rect 4252 45484 4304 45490
rect 4252 45426 4304 45432
rect 4356 45370 4384 46310
rect 4080 45342 4384 45370
rect 3974 44976 4030 44985
rect 3974 44911 4030 44920
rect 3528 44798 4016 44826
rect 3516 44736 3568 44742
rect 3516 44678 3568 44684
rect 3528 22778 3556 44678
rect 3610 44092 3918 44101
rect 3610 44090 3616 44092
rect 3672 44090 3696 44092
rect 3752 44090 3776 44092
rect 3832 44090 3856 44092
rect 3912 44090 3918 44092
rect 3672 44038 3674 44090
rect 3854 44038 3856 44090
rect 3610 44036 3616 44038
rect 3672 44036 3696 44038
rect 3752 44036 3776 44038
rect 3832 44036 3856 44038
rect 3912 44036 3918 44038
rect 3610 44027 3918 44036
rect 3610 43004 3918 43013
rect 3610 43002 3616 43004
rect 3672 43002 3696 43004
rect 3752 43002 3776 43004
rect 3832 43002 3856 43004
rect 3912 43002 3918 43004
rect 3672 42950 3674 43002
rect 3854 42950 3856 43002
rect 3610 42948 3616 42950
rect 3672 42948 3696 42950
rect 3752 42948 3776 42950
rect 3832 42948 3856 42950
rect 3912 42948 3918 42950
rect 3610 42939 3918 42948
rect 3988 42838 4016 44798
rect 4080 43994 4108 45342
rect 4160 45280 4212 45286
rect 4160 45222 4212 45228
rect 4252 45280 4304 45286
rect 4252 45222 4304 45228
rect 4068 43988 4120 43994
rect 4068 43930 4120 43936
rect 3976 42832 4028 42838
rect 3976 42774 4028 42780
rect 3884 42560 3936 42566
rect 3884 42502 3936 42508
rect 4068 42560 4120 42566
rect 4068 42502 4120 42508
rect 3896 42090 3924 42502
rect 3976 42356 4028 42362
rect 3976 42298 4028 42304
rect 3884 42084 3936 42090
rect 3884 42026 3936 42032
rect 3610 41916 3918 41925
rect 3610 41914 3616 41916
rect 3672 41914 3696 41916
rect 3752 41914 3776 41916
rect 3832 41914 3856 41916
rect 3912 41914 3918 41916
rect 3672 41862 3674 41914
rect 3854 41862 3856 41914
rect 3610 41860 3616 41862
rect 3672 41860 3696 41862
rect 3752 41860 3776 41862
rect 3832 41860 3856 41862
rect 3912 41860 3918 41862
rect 3610 41851 3918 41860
rect 3610 40828 3918 40837
rect 3610 40826 3616 40828
rect 3672 40826 3696 40828
rect 3752 40826 3776 40828
rect 3832 40826 3856 40828
rect 3912 40826 3918 40828
rect 3672 40774 3674 40826
rect 3854 40774 3856 40826
rect 3610 40772 3616 40774
rect 3672 40772 3696 40774
rect 3752 40772 3776 40774
rect 3832 40772 3856 40774
rect 3912 40772 3918 40774
rect 3610 40763 3918 40772
rect 3610 39740 3918 39749
rect 3610 39738 3616 39740
rect 3672 39738 3696 39740
rect 3752 39738 3776 39740
rect 3832 39738 3856 39740
rect 3912 39738 3918 39740
rect 3672 39686 3674 39738
rect 3854 39686 3856 39738
rect 3610 39684 3616 39686
rect 3672 39684 3696 39686
rect 3752 39684 3776 39686
rect 3832 39684 3856 39686
rect 3912 39684 3918 39686
rect 3610 39675 3918 39684
rect 3610 38652 3918 38661
rect 3610 38650 3616 38652
rect 3672 38650 3696 38652
rect 3752 38650 3776 38652
rect 3832 38650 3856 38652
rect 3912 38650 3918 38652
rect 3672 38598 3674 38650
rect 3854 38598 3856 38650
rect 3610 38596 3616 38598
rect 3672 38596 3696 38598
rect 3752 38596 3776 38598
rect 3832 38596 3856 38598
rect 3912 38596 3918 38598
rect 3610 38587 3918 38596
rect 3610 37564 3918 37573
rect 3610 37562 3616 37564
rect 3672 37562 3696 37564
rect 3752 37562 3776 37564
rect 3832 37562 3856 37564
rect 3912 37562 3918 37564
rect 3672 37510 3674 37562
rect 3854 37510 3856 37562
rect 3610 37508 3616 37510
rect 3672 37508 3696 37510
rect 3752 37508 3776 37510
rect 3832 37508 3856 37510
rect 3912 37508 3918 37510
rect 3610 37499 3918 37508
rect 3610 36476 3918 36485
rect 3610 36474 3616 36476
rect 3672 36474 3696 36476
rect 3752 36474 3776 36476
rect 3832 36474 3856 36476
rect 3912 36474 3918 36476
rect 3672 36422 3674 36474
rect 3854 36422 3856 36474
rect 3610 36420 3616 36422
rect 3672 36420 3696 36422
rect 3752 36420 3776 36422
rect 3832 36420 3856 36422
rect 3912 36420 3918 36422
rect 3610 36411 3918 36420
rect 3610 35388 3918 35397
rect 3610 35386 3616 35388
rect 3672 35386 3696 35388
rect 3752 35386 3776 35388
rect 3832 35386 3856 35388
rect 3912 35386 3918 35388
rect 3672 35334 3674 35386
rect 3854 35334 3856 35386
rect 3610 35332 3616 35334
rect 3672 35332 3696 35334
rect 3752 35332 3776 35334
rect 3832 35332 3856 35334
rect 3912 35332 3918 35334
rect 3610 35323 3918 35332
rect 3610 34300 3918 34309
rect 3610 34298 3616 34300
rect 3672 34298 3696 34300
rect 3752 34298 3776 34300
rect 3832 34298 3856 34300
rect 3912 34298 3918 34300
rect 3672 34246 3674 34298
rect 3854 34246 3856 34298
rect 3610 34244 3616 34246
rect 3672 34244 3696 34246
rect 3752 34244 3776 34246
rect 3832 34244 3856 34246
rect 3912 34244 3918 34246
rect 3610 34235 3918 34244
rect 3884 34196 3936 34202
rect 3884 34138 3936 34144
rect 3896 33658 3924 34138
rect 3884 33652 3936 33658
rect 3884 33594 3936 33600
rect 3610 33212 3918 33221
rect 3610 33210 3616 33212
rect 3672 33210 3696 33212
rect 3752 33210 3776 33212
rect 3832 33210 3856 33212
rect 3912 33210 3918 33212
rect 3672 33158 3674 33210
rect 3854 33158 3856 33210
rect 3610 33156 3616 33158
rect 3672 33156 3696 33158
rect 3752 33156 3776 33158
rect 3832 33156 3856 33158
rect 3912 33156 3918 33158
rect 3610 33147 3918 33156
rect 3610 32124 3918 32133
rect 3610 32122 3616 32124
rect 3672 32122 3696 32124
rect 3752 32122 3776 32124
rect 3832 32122 3856 32124
rect 3912 32122 3918 32124
rect 3672 32070 3674 32122
rect 3854 32070 3856 32122
rect 3610 32068 3616 32070
rect 3672 32068 3696 32070
rect 3752 32068 3776 32070
rect 3832 32068 3856 32070
rect 3912 32068 3918 32070
rect 3610 32059 3918 32068
rect 3610 31036 3918 31045
rect 3610 31034 3616 31036
rect 3672 31034 3696 31036
rect 3752 31034 3776 31036
rect 3832 31034 3856 31036
rect 3912 31034 3918 31036
rect 3672 30982 3674 31034
rect 3854 30982 3856 31034
rect 3610 30980 3616 30982
rect 3672 30980 3696 30982
rect 3752 30980 3776 30982
rect 3832 30980 3856 30982
rect 3912 30980 3918 30982
rect 3610 30971 3918 30980
rect 3610 29948 3918 29957
rect 3610 29946 3616 29948
rect 3672 29946 3696 29948
rect 3752 29946 3776 29948
rect 3832 29946 3856 29948
rect 3912 29946 3918 29948
rect 3672 29894 3674 29946
rect 3854 29894 3856 29946
rect 3610 29892 3616 29894
rect 3672 29892 3696 29894
rect 3752 29892 3776 29894
rect 3832 29892 3856 29894
rect 3912 29892 3918 29894
rect 3610 29883 3918 29892
rect 3610 28860 3918 28869
rect 3610 28858 3616 28860
rect 3672 28858 3696 28860
rect 3752 28858 3776 28860
rect 3832 28858 3856 28860
rect 3912 28858 3918 28860
rect 3672 28806 3674 28858
rect 3854 28806 3856 28858
rect 3610 28804 3616 28806
rect 3672 28804 3696 28806
rect 3752 28804 3776 28806
rect 3832 28804 3856 28806
rect 3912 28804 3918 28806
rect 3610 28795 3918 28804
rect 3610 27772 3918 27781
rect 3610 27770 3616 27772
rect 3672 27770 3696 27772
rect 3752 27770 3776 27772
rect 3832 27770 3856 27772
rect 3912 27770 3918 27772
rect 3672 27718 3674 27770
rect 3854 27718 3856 27770
rect 3610 27716 3616 27718
rect 3672 27716 3696 27718
rect 3752 27716 3776 27718
rect 3832 27716 3856 27718
rect 3912 27716 3918 27718
rect 3610 27707 3918 27716
rect 3610 26684 3918 26693
rect 3610 26682 3616 26684
rect 3672 26682 3696 26684
rect 3752 26682 3776 26684
rect 3832 26682 3856 26684
rect 3912 26682 3918 26684
rect 3672 26630 3674 26682
rect 3854 26630 3856 26682
rect 3610 26628 3616 26630
rect 3672 26628 3696 26630
rect 3752 26628 3776 26630
rect 3832 26628 3856 26630
rect 3912 26628 3918 26630
rect 3610 26619 3918 26628
rect 3988 26382 4016 42298
rect 4080 42265 4108 42502
rect 4066 42256 4122 42265
rect 4066 42191 4122 42200
rect 4172 41818 4200 45222
rect 4160 41812 4212 41818
rect 4160 41754 4212 41760
rect 4068 40928 4120 40934
rect 4068 40870 4120 40876
rect 4080 39030 4108 40870
rect 4160 39296 4212 39302
rect 4160 39238 4212 39244
rect 4068 39024 4120 39030
rect 4068 38966 4120 38972
rect 4068 35692 4120 35698
rect 4068 35634 4120 35640
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 3610 25596 3918 25605
rect 3610 25594 3616 25596
rect 3672 25594 3696 25596
rect 3752 25594 3776 25596
rect 3832 25594 3856 25596
rect 3912 25594 3918 25596
rect 3672 25542 3674 25594
rect 3854 25542 3856 25594
rect 3610 25540 3616 25542
rect 3672 25540 3696 25542
rect 3752 25540 3776 25542
rect 3832 25540 3856 25542
rect 3912 25540 3918 25542
rect 3610 25531 3918 25540
rect 3610 24508 3918 24517
rect 3610 24506 3616 24508
rect 3672 24506 3696 24508
rect 3752 24506 3776 24508
rect 3832 24506 3856 24508
rect 3912 24506 3918 24508
rect 3672 24454 3674 24506
rect 3854 24454 3856 24506
rect 3610 24452 3616 24454
rect 3672 24452 3696 24454
rect 3752 24452 3776 24454
rect 3832 24452 3856 24454
rect 3912 24452 3918 24454
rect 3610 24443 3918 24452
rect 3610 23420 3918 23429
rect 3610 23418 3616 23420
rect 3672 23418 3696 23420
rect 3752 23418 3776 23420
rect 3832 23418 3856 23420
rect 3912 23418 3918 23420
rect 3672 23366 3674 23418
rect 3854 23366 3856 23418
rect 3610 23364 3616 23366
rect 3672 23364 3696 23366
rect 3752 23364 3776 23366
rect 3832 23364 3856 23366
rect 3912 23364 3918 23366
rect 3610 23355 3918 23364
rect 3608 23316 3660 23322
rect 3608 23258 3660 23264
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3620 22658 3648 23258
rect 3528 22630 3648 22658
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3528 15502 3556 22630
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3610 22332 3918 22341
rect 3610 22330 3616 22332
rect 3672 22330 3696 22332
rect 3752 22330 3776 22332
rect 3832 22330 3856 22332
rect 3912 22330 3918 22332
rect 3672 22278 3674 22330
rect 3854 22278 3856 22330
rect 3610 22276 3616 22278
rect 3672 22276 3696 22278
rect 3752 22276 3776 22278
rect 3832 22276 3856 22278
rect 3912 22276 3918 22278
rect 3610 22267 3918 22276
rect 3610 21244 3918 21253
rect 3610 21242 3616 21244
rect 3672 21242 3696 21244
rect 3752 21242 3776 21244
rect 3832 21242 3856 21244
rect 3912 21242 3918 21244
rect 3672 21190 3674 21242
rect 3854 21190 3856 21242
rect 3610 21188 3616 21190
rect 3672 21188 3696 21190
rect 3752 21188 3776 21190
rect 3832 21188 3856 21190
rect 3912 21188 3918 21190
rect 3610 21179 3918 21188
rect 3610 20156 3918 20165
rect 3610 20154 3616 20156
rect 3672 20154 3696 20156
rect 3752 20154 3776 20156
rect 3832 20154 3856 20156
rect 3912 20154 3918 20156
rect 3672 20102 3674 20154
rect 3854 20102 3856 20154
rect 3610 20100 3616 20102
rect 3672 20100 3696 20102
rect 3752 20100 3776 20102
rect 3832 20100 3856 20102
rect 3912 20100 3918 20102
rect 3610 20091 3918 20100
rect 3610 19068 3918 19077
rect 3610 19066 3616 19068
rect 3672 19066 3696 19068
rect 3752 19066 3776 19068
rect 3832 19066 3856 19068
rect 3912 19066 3918 19068
rect 3672 19014 3674 19066
rect 3854 19014 3856 19066
rect 3610 19012 3616 19014
rect 3672 19012 3696 19014
rect 3752 19012 3776 19014
rect 3832 19012 3856 19014
rect 3912 19012 3918 19014
rect 3610 19003 3918 19012
rect 3610 17980 3918 17989
rect 3610 17978 3616 17980
rect 3672 17978 3696 17980
rect 3752 17978 3776 17980
rect 3832 17978 3856 17980
rect 3912 17978 3918 17980
rect 3672 17926 3674 17978
rect 3854 17926 3856 17978
rect 3610 17924 3616 17926
rect 3672 17924 3696 17926
rect 3752 17924 3776 17926
rect 3832 17924 3856 17926
rect 3912 17924 3918 17926
rect 3610 17915 3918 17924
rect 3610 16892 3918 16901
rect 3610 16890 3616 16892
rect 3672 16890 3696 16892
rect 3752 16890 3776 16892
rect 3832 16890 3856 16892
rect 3912 16890 3918 16892
rect 3672 16838 3674 16890
rect 3854 16838 3856 16890
rect 3610 16836 3616 16838
rect 3672 16836 3696 16838
rect 3752 16836 3776 16838
rect 3832 16836 3856 16838
rect 3912 16836 3918 16838
rect 3610 16827 3918 16836
rect 3610 15804 3918 15813
rect 3610 15802 3616 15804
rect 3672 15802 3696 15804
rect 3752 15802 3776 15804
rect 3832 15802 3856 15804
rect 3912 15802 3918 15804
rect 3672 15750 3674 15802
rect 3854 15750 3856 15802
rect 3610 15748 3616 15750
rect 3672 15748 3696 15750
rect 3752 15748 3776 15750
rect 3832 15748 3856 15750
rect 3912 15748 3918 15750
rect 3610 15739 3918 15748
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3610 14716 3918 14725
rect 3610 14714 3616 14716
rect 3672 14714 3696 14716
rect 3752 14714 3776 14716
rect 3832 14714 3856 14716
rect 3912 14714 3918 14716
rect 3672 14662 3674 14714
rect 3854 14662 3856 14714
rect 3610 14660 3616 14662
rect 3672 14660 3696 14662
rect 3752 14660 3776 14662
rect 3832 14660 3856 14662
rect 3912 14660 3918 14662
rect 3610 14651 3918 14660
rect 3610 13628 3918 13637
rect 3610 13626 3616 13628
rect 3672 13626 3696 13628
rect 3752 13626 3776 13628
rect 3832 13626 3856 13628
rect 3912 13626 3918 13628
rect 3672 13574 3674 13626
rect 3854 13574 3856 13626
rect 3610 13572 3616 13574
rect 3672 13572 3696 13574
rect 3752 13572 3776 13574
rect 3832 13572 3856 13574
rect 3912 13572 3918 13574
rect 3610 13563 3918 13572
rect 3610 12540 3918 12549
rect 3610 12538 3616 12540
rect 3672 12538 3696 12540
rect 3752 12538 3776 12540
rect 3832 12538 3856 12540
rect 3912 12538 3918 12540
rect 3672 12486 3674 12538
rect 3854 12486 3856 12538
rect 3610 12484 3616 12486
rect 3672 12484 3696 12486
rect 3752 12484 3776 12486
rect 3832 12484 3856 12486
rect 3912 12484 3918 12486
rect 3610 12475 3918 12484
rect 3610 11452 3918 11461
rect 3610 11450 3616 11452
rect 3672 11450 3696 11452
rect 3752 11450 3776 11452
rect 3832 11450 3856 11452
rect 3912 11450 3918 11452
rect 3672 11398 3674 11450
rect 3854 11398 3856 11450
rect 3610 11396 3616 11398
rect 3672 11396 3696 11398
rect 3752 11396 3776 11398
rect 3832 11396 3856 11398
rect 3912 11396 3918 11398
rect 3610 11387 3918 11396
rect 3610 10364 3918 10373
rect 3610 10362 3616 10364
rect 3672 10362 3696 10364
rect 3752 10362 3776 10364
rect 3832 10362 3856 10364
rect 3912 10362 3918 10364
rect 3672 10310 3674 10362
rect 3854 10310 3856 10362
rect 3610 10308 3616 10310
rect 3672 10308 3696 10310
rect 3752 10308 3776 10310
rect 3832 10308 3856 10310
rect 3912 10308 3918 10310
rect 3610 10299 3918 10308
rect 3610 9276 3918 9285
rect 3610 9274 3616 9276
rect 3672 9274 3696 9276
rect 3752 9274 3776 9276
rect 3832 9274 3856 9276
rect 3912 9274 3918 9276
rect 3672 9222 3674 9274
rect 3854 9222 3856 9274
rect 3610 9220 3616 9222
rect 3672 9220 3696 9222
rect 3752 9220 3776 9222
rect 3832 9220 3856 9222
rect 3912 9220 3918 9222
rect 3610 9211 3918 9220
rect 3610 8188 3918 8197
rect 3610 8186 3616 8188
rect 3672 8186 3696 8188
rect 3752 8186 3776 8188
rect 3832 8186 3856 8188
rect 3912 8186 3918 8188
rect 3672 8134 3674 8186
rect 3854 8134 3856 8186
rect 3610 8132 3616 8134
rect 3672 8132 3696 8134
rect 3752 8132 3776 8134
rect 3832 8132 3856 8134
rect 3912 8132 3918 8134
rect 3610 8123 3918 8132
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3610 7100 3918 7109
rect 3610 7098 3616 7100
rect 3672 7098 3696 7100
rect 3752 7098 3776 7100
rect 3832 7098 3856 7100
rect 3912 7098 3918 7100
rect 3672 7046 3674 7098
rect 3854 7046 3856 7098
rect 3610 7044 3616 7046
rect 3672 7044 3696 7046
rect 3752 7044 3776 7046
rect 3832 7044 3856 7046
rect 3912 7044 3918 7046
rect 3610 7035 3918 7044
rect 2950 6556 3258 6565
rect 2950 6554 2956 6556
rect 3012 6554 3036 6556
rect 3092 6554 3116 6556
rect 3172 6554 3196 6556
rect 3252 6554 3258 6556
rect 3012 6502 3014 6554
rect 3194 6502 3196 6554
rect 2950 6500 2956 6502
rect 3012 6500 3036 6502
rect 3092 6500 3116 6502
rect 3172 6500 3196 6502
rect 3252 6500 3258 6502
rect 2950 6491 3258 6500
rect 3610 6012 3918 6021
rect 3610 6010 3616 6012
rect 3672 6010 3696 6012
rect 3752 6010 3776 6012
rect 3832 6010 3856 6012
rect 3912 6010 3918 6012
rect 3672 5958 3674 6010
rect 3854 5958 3856 6010
rect 3610 5956 3616 5958
rect 3672 5956 3696 5958
rect 3752 5956 3776 5958
rect 3832 5956 3856 5958
rect 3912 5956 3918 5958
rect 3610 5947 3918 5956
rect 3988 5710 4016 22374
rect 4080 14414 4108 35634
rect 4172 30326 4200 39238
rect 4264 36530 4292 45222
rect 4344 45076 4396 45082
rect 4344 45018 4396 45024
rect 4356 44402 4384 45018
rect 4344 44396 4396 44402
rect 4344 44338 4396 44344
rect 4344 44192 4396 44198
rect 4344 44134 4396 44140
rect 4356 42786 4384 44134
rect 4448 42922 4476 46543
rect 4540 45966 4568 46668
rect 4528 45960 4580 45966
rect 4528 45902 4580 45908
rect 4550 45724 4858 45733
rect 4550 45722 4556 45724
rect 4612 45722 4636 45724
rect 4692 45722 4716 45724
rect 4772 45722 4796 45724
rect 4852 45722 4858 45724
rect 4612 45670 4614 45722
rect 4794 45670 4796 45722
rect 4550 45668 4556 45670
rect 4612 45668 4636 45670
rect 4692 45668 4716 45670
rect 4772 45668 4796 45670
rect 4852 45668 4858 45670
rect 4550 45659 4858 45668
rect 4908 45608 4936 47466
rect 4540 45580 4936 45608
rect 4540 44946 4568 45580
rect 5000 45490 5028 49728
rect 4620 45484 4672 45490
rect 4620 45426 4672 45432
rect 4988 45484 5040 45490
rect 4988 45426 5040 45432
rect 4632 45082 4660 45426
rect 4988 45348 5040 45354
rect 4988 45290 5040 45296
rect 4620 45076 4672 45082
rect 4620 45018 4672 45024
rect 4528 44940 4580 44946
rect 4528 44882 4580 44888
rect 4632 44878 4660 45018
rect 4620 44872 4672 44878
rect 4620 44814 4672 44820
rect 4550 44636 4858 44645
rect 4550 44634 4556 44636
rect 4612 44634 4636 44636
rect 4692 44634 4716 44636
rect 4772 44634 4796 44636
rect 4852 44634 4858 44636
rect 4612 44582 4614 44634
rect 4794 44582 4796 44634
rect 4550 44580 4556 44582
rect 4612 44580 4636 44582
rect 4692 44580 4716 44582
rect 4772 44580 4796 44582
rect 4852 44580 4858 44582
rect 4550 44571 4858 44580
rect 4712 44532 4764 44538
rect 4764 44492 4844 44520
rect 4712 44474 4764 44480
rect 4712 44396 4764 44402
rect 4712 44338 4764 44344
rect 4724 44266 4752 44338
rect 4712 44260 4764 44266
rect 4712 44202 4764 44208
rect 4816 44180 4844 44492
rect 4896 44328 4948 44334
rect 5000 44282 5028 45290
rect 5092 44402 5120 49830
rect 5460 49722 5488 50374
rect 5644 50266 5672 50748
rect 5552 50238 5672 50266
rect 5552 49910 5580 50238
rect 5632 50176 5684 50182
rect 5632 50118 5684 50124
rect 5540 49904 5592 49910
rect 5540 49846 5592 49852
rect 5460 49694 5580 49722
rect 5210 49532 5518 49541
rect 5210 49530 5216 49532
rect 5272 49530 5296 49532
rect 5352 49530 5376 49532
rect 5432 49530 5456 49532
rect 5512 49530 5518 49532
rect 5272 49478 5274 49530
rect 5454 49478 5456 49530
rect 5210 49476 5216 49478
rect 5272 49476 5296 49478
rect 5352 49476 5376 49478
rect 5432 49476 5456 49478
rect 5512 49476 5518 49478
rect 5210 49467 5518 49476
rect 5172 49428 5224 49434
rect 5172 49370 5224 49376
rect 5184 48618 5212 49370
rect 5552 49314 5580 49694
rect 5460 49286 5580 49314
rect 5460 48634 5488 49286
rect 5172 48612 5224 48618
rect 5460 48606 5580 48634
rect 5172 48554 5224 48560
rect 5210 48444 5518 48453
rect 5210 48442 5216 48444
rect 5272 48442 5296 48444
rect 5352 48442 5376 48444
rect 5432 48442 5456 48444
rect 5512 48442 5518 48444
rect 5272 48390 5274 48442
rect 5454 48390 5456 48442
rect 5210 48388 5216 48390
rect 5272 48388 5296 48390
rect 5352 48388 5376 48390
rect 5432 48388 5456 48390
rect 5512 48388 5518 48390
rect 5210 48379 5518 48388
rect 5172 48340 5224 48346
rect 5172 48282 5224 48288
rect 5184 47462 5212 48282
rect 5172 47456 5224 47462
rect 5172 47398 5224 47404
rect 5210 47356 5518 47365
rect 5210 47354 5216 47356
rect 5272 47354 5296 47356
rect 5352 47354 5376 47356
rect 5432 47354 5456 47356
rect 5512 47354 5518 47356
rect 5272 47302 5274 47354
rect 5454 47302 5456 47354
rect 5210 47300 5216 47302
rect 5272 47300 5296 47302
rect 5352 47300 5376 47302
rect 5432 47300 5456 47302
rect 5512 47300 5518 47302
rect 5210 47291 5518 47300
rect 5552 47104 5580 48606
rect 5460 47076 5580 47104
rect 5172 46912 5224 46918
rect 5172 46854 5224 46860
rect 5184 46374 5212 46854
rect 5172 46368 5224 46374
rect 5460 46356 5488 47076
rect 5540 46980 5592 46986
rect 5540 46922 5592 46928
rect 5552 46578 5580 46922
rect 5540 46572 5592 46578
rect 5540 46514 5592 46520
rect 5460 46328 5580 46356
rect 5172 46310 5224 46316
rect 5210 46268 5518 46277
rect 5210 46266 5216 46268
rect 5272 46266 5296 46268
rect 5352 46266 5376 46268
rect 5432 46266 5456 46268
rect 5512 46266 5518 46268
rect 5272 46214 5274 46266
rect 5454 46214 5456 46266
rect 5210 46212 5216 46214
rect 5272 46212 5296 46214
rect 5352 46212 5376 46214
rect 5432 46212 5456 46214
rect 5512 46212 5518 46214
rect 5210 46203 5518 46212
rect 5552 46016 5580 46328
rect 5460 45988 5580 46016
rect 5172 45960 5224 45966
rect 5172 45902 5224 45908
rect 5184 45393 5212 45902
rect 5460 45490 5488 45988
rect 5540 45892 5592 45898
rect 5540 45834 5592 45840
rect 5448 45484 5500 45490
rect 5448 45426 5500 45432
rect 5170 45384 5226 45393
rect 5170 45319 5226 45328
rect 5210 45180 5518 45189
rect 5210 45178 5216 45180
rect 5272 45178 5296 45180
rect 5352 45178 5376 45180
rect 5432 45178 5456 45180
rect 5512 45178 5518 45180
rect 5272 45126 5274 45178
rect 5454 45126 5456 45178
rect 5210 45124 5216 45126
rect 5272 45124 5296 45126
rect 5352 45124 5376 45126
rect 5432 45124 5456 45126
rect 5512 45124 5518 45126
rect 5210 45115 5518 45124
rect 5170 44976 5226 44985
rect 5170 44911 5226 44920
rect 5184 44402 5212 44911
rect 5264 44872 5316 44878
rect 5448 44872 5500 44878
rect 5264 44814 5316 44820
rect 5446 44840 5448 44849
rect 5500 44840 5502 44849
rect 5276 44538 5304 44814
rect 5446 44775 5502 44784
rect 5264 44532 5316 44538
rect 5264 44474 5316 44480
rect 5080 44396 5132 44402
rect 5080 44338 5132 44344
rect 5172 44396 5224 44402
rect 5172 44338 5224 44344
rect 4948 44276 5028 44282
rect 4896 44270 5028 44276
rect 4908 44254 5028 44270
rect 4816 44152 5028 44180
rect 4896 43648 4948 43654
rect 4896 43590 4948 43596
rect 4550 43548 4858 43557
rect 4550 43546 4556 43548
rect 4612 43546 4636 43548
rect 4692 43546 4716 43548
rect 4772 43546 4796 43548
rect 4852 43546 4858 43548
rect 4612 43494 4614 43546
rect 4794 43494 4796 43546
rect 4550 43492 4556 43494
rect 4612 43492 4636 43494
rect 4692 43492 4716 43494
rect 4772 43492 4796 43494
rect 4852 43492 4858 43494
rect 4550 43483 4858 43492
rect 4448 42894 4568 42922
rect 4356 42758 4476 42786
rect 4540 42770 4568 42894
rect 4344 42560 4396 42566
rect 4344 42502 4396 42508
rect 4356 40594 4384 42502
rect 4344 40588 4396 40594
rect 4344 40530 4396 40536
rect 4344 40452 4396 40458
rect 4344 40394 4396 40400
rect 4356 39642 4384 40394
rect 4344 39636 4396 39642
rect 4344 39578 4396 39584
rect 4344 37664 4396 37670
rect 4344 37606 4396 37612
rect 4356 36689 4384 37606
rect 4342 36680 4398 36689
rect 4342 36615 4398 36624
rect 4264 36502 4384 36530
rect 4250 36408 4306 36417
rect 4250 36343 4306 36352
rect 4160 30320 4212 30326
rect 4160 30262 4212 30268
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4172 27674 4200 30126
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 4160 26240 4212 26246
rect 4160 26182 4212 26188
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4172 9654 4200 26182
rect 4264 22778 4292 36343
rect 4356 22953 4384 36502
rect 4342 22944 4398 22953
rect 4342 22879 4398 22888
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 4250 22672 4306 22681
rect 4250 22607 4306 22616
rect 4264 22522 4292 22607
rect 4264 22494 4384 22522
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 2950 5468 3258 5477
rect 2950 5466 2956 5468
rect 3012 5466 3036 5468
rect 3092 5466 3116 5468
rect 3172 5466 3196 5468
rect 3252 5466 3258 5468
rect 3012 5414 3014 5466
rect 3194 5414 3196 5466
rect 2950 5412 2956 5414
rect 3012 5412 3036 5414
rect 3092 5412 3116 5414
rect 3172 5412 3196 5414
rect 3252 5412 3258 5414
rect 2950 5403 3258 5412
rect 3610 4924 3918 4933
rect 3610 4922 3616 4924
rect 3672 4922 3696 4924
rect 3752 4922 3776 4924
rect 3832 4922 3856 4924
rect 3912 4922 3918 4924
rect 3672 4870 3674 4922
rect 3854 4870 3856 4922
rect 3610 4868 3616 4870
rect 3672 4868 3696 4870
rect 3752 4868 3776 4870
rect 3832 4868 3856 4870
rect 3912 4868 3918 4870
rect 3610 4859 3918 4868
rect 4264 4622 4292 22102
rect 4356 16182 4384 22494
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4448 15094 4476 42758
rect 4528 42764 4580 42770
rect 4528 42706 4580 42712
rect 4550 42460 4858 42469
rect 4550 42458 4556 42460
rect 4612 42458 4636 42460
rect 4692 42458 4716 42460
rect 4772 42458 4796 42460
rect 4852 42458 4858 42460
rect 4612 42406 4614 42458
rect 4794 42406 4796 42458
rect 4550 42404 4556 42406
rect 4612 42404 4636 42406
rect 4692 42404 4716 42406
rect 4772 42404 4796 42406
rect 4852 42404 4858 42406
rect 4550 42395 4858 42404
rect 4618 42256 4674 42265
rect 4618 42191 4674 42200
rect 4528 41608 4580 41614
rect 4632 41596 4660 42191
rect 4908 41614 4936 43590
rect 4580 41568 4660 41596
rect 4896 41608 4948 41614
rect 4528 41550 4580 41556
rect 4896 41550 4948 41556
rect 4550 41372 4858 41381
rect 4550 41370 4556 41372
rect 4612 41370 4636 41372
rect 4692 41370 4716 41372
rect 4772 41370 4796 41372
rect 4852 41370 4858 41372
rect 4612 41318 4614 41370
rect 4794 41318 4796 41370
rect 4550 41316 4556 41318
rect 4612 41316 4636 41318
rect 4692 41316 4716 41318
rect 4772 41316 4796 41318
rect 4852 41316 4858 41318
rect 4550 41307 4858 41316
rect 4804 40588 4856 40594
rect 5000 40576 5028 44152
rect 5210 44092 5518 44101
rect 5210 44090 5216 44092
rect 5272 44090 5296 44092
rect 5352 44090 5376 44092
rect 5432 44090 5456 44092
rect 5512 44090 5518 44092
rect 5272 44038 5274 44090
rect 5454 44038 5456 44090
rect 5210 44036 5216 44038
rect 5272 44036 5296 44038
rect 5352 44036 5376 44038
rect 5432 44036 5456 44038
rect 5512 44036 5518 44038
rect 5210 44027 5518 44036
rect 5210 43004 5518 43013
rect 5210 43002 5216 43004
rect 5272 43002 5296 43004
rect 5352 43002 5376 43004
rect 5432 43002 5456 43004
rect 5512 43002 5518 43004
rect 5272 42950 5274 43002
rect 5454 42950 5456 43002
rect 5210 42948 5216 42950
rect 5272 42948 5296 42950
rect 5352 42948 5376 42950
rect 5432 42948 5456 42950
rect 5512 42948 5518 42950
rect 5210 42939 5518 42948
rect 5264 42696 5316 42702
rect 5262 42664 5264 42673
rect 5448 42696 5500 42702
rect 5316 42664 5318 42673
rect 5448 42638 5500 42644
rect 5262 42599 5318 42608
rect 5080 42560 5132 42566
rect 5080 42502 5132 42508
rect 5172 42560 5224 42566
rect 5172 42502 5224 42508
rect 5264 42560 5316 42566
rect 5264 42502 5316 42508
rect 5092 40712 5120 42502
rect 5184 42022 5212 42502
rect 5276 42362 5304 42502
rect 5264 42356 5316 42362
rect 5264 42298 5316 42304
rect 5460 42294 5488 42638
rect 5552 42634 5580 45834
rect 5644 45014 5672 50118
rect 5736 46918 5764 52634
rect 5724 46912 5776 46918
rect 5724 46854 5776 46860
rect 5724 46708 5776 46714
rect 5724 46650 5776 46656
rect 5632 45008 5684 45014
rect 5632 44950 5684 44956
rect 5630 44840 5686 44849
rect 5630 44775 5686 44784
rect 5540 42628 5592 42634
rect 5540 42570 5592 42576
rect 5448 42288 5500 42294
rect 5448 42230 5500 42236
rect 5172 42016 5224 42022
rect 5172 41958 5224 41964
rect 5540 42016 5592 42022
rect 5540 41958 5592 41964
rect 5210 41916 5518 41925
rect 5210 41914 5216 41916
rect 5272 41914 5296 41916
rect 5352 41914 5376 41916
rect 5432 41914 5456 41916
rect 5512 41914 5518 41916
rect 5272 41862 5274 41914
rect 5454 41862 5456 41914
rect 5210 41860 5216 41862
rect 5272 41860 5296 41862
rect 5352 41860 5376 41862
rect 5432 41860 5456 41862
rect 5512 41860 5518 41862
rect 5210 41851 5518 41860
rect 5210 40828 5518 40837
rect 5210 40826 5216 40828
rect 5272 40826 5296 40828
rect 5352 40826 5376 40828
rect 5432 40826 5456 40828
rect 5512 40826 5518 40828
rect 5272 40774 5274 40826
rect 5454 40774 5456 40826
rect 5210 40772 5216 40774
rect 5272 40772 5296 40774
rect 5352 40772 5376 40774
rect 5432 40772 5456 40774
rect 5512 40772 5518 40774
rect 5210 40763 5518 40772
rect 5092 40684 5304 40712
rect 5000 40548 5212 40576
rect 4804 40530 4856 40536
rect 4816 40390 4844 40530
rect 4804 40384 4856 40390
rect 4804 40326 4856 40332
rect 4988 40384 5040 40390
rect 4988 40326 5040 40332
rect 4550 40284 4858 40293
rect 4550 40282 4556 40284
rect 4612 40282 4636 40284
rect 4692 40282 4716 40284
rect 4772 40282 4796 40284
rect 4852 40282 4858 40284
rect 4612 40230 4614 40282
rect 4794 40230 4796 40282
rect 4550 40228 4556 40230
rect 4612 40228 4636 40230
rect 4692 40228 4716 40230
rect 4772 40228 4796 40230
rect 4852 40228 4858 40230
rect 4550 40219 4858 40228
rect 4804 40180 4856 40186
rect 4804 40122 4856 40128
rect 4816 39386 4844 40122
rect 4816 39358 4936 39386
rect 4550 39196 4858 39205
rect 4550 39194 4556 39196
rect 4612 39194 4636 39196
rect 4692 39194 4716 39196
rect 4772 39194 4796 39196
rect 4852 39194 4858 39196
rect 4612 39142 4614 39194
rect 4794 39142 4796 39194
rect 4550 39140 4556 39142
rect 4612 39140 4636 39142
rect 4692 39140 4716 39142
rect 4772 39140 4796 39142
rect 4852 39140 4858 39142
rect 4550 39131 4858 39140
rect 4550 38108 4858 38117
rect 4550 38106 4556 38108
rect 4612 38106 4636 38108
rect 4692 38106 4716 38108
rect 4772 38106 4796 38108
rect 4852 38106 4858 38108
rect 4612 38054 4614 38106
rect 4794 38054 4796 38106
rect 4550 38052 4556 38054
rect 4612 38052 4636 38054
rect 4692 38052 4716 38054
rect 4772 38052 4796 38054
rect 4852 38052 4858 38054
rect 4550 38043 4858 38052
rect 4550 37020 4858 37029
rect 4550 37018 4556 37020
rect 4612 37018 4636 37020
rect 4692 37018 4716 37020
rect 4772 37018 4796 37020
rect 4852 37018 4858 37020
rect 4612 36966 4614 37018
rect 4794 36966 4796 37018
rect 4550 36964 4556 36966
rect 4612 36964 4636 36966
rect 4692 36964 4716 36966
rect 4772 36964 4796 36966
rect 4852 36964 4858 36966
rect 4550 36955 4858 36964
rect 4550 35932 4858 35941
rect 4550 35930 4556 35932
rect 4612 35930 4636 35932
rect 4692 35930 4716 35932
rect 4772 35930 4796 35932
rect 4852 35930 4858 35932
rect 4612 35878 4614 35930
rect 4794 35878 4796 35930
rect 4550 35876 4556 35878
rect 4612 35876 4636 35878
rect 4692 35876 4716 35878
rect 4772 35876 4796 35878
rect 4852 35876 4858 35878
rect 4550 35867 4858 35876
rect 4908 35698 4936 39358
rect 5000 37262 5028 40326
rect 5184 40186 5212 40548
rect 5172 40180 5224 40186
rect 5172 40122 5224 40128
rect 5276 40066 5304 40684
rect 5092 40038 5304 40066
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 4988 36644 5040 36650
rect 4988 36586 5040 36592
rect 4896 35692 4948 35698
rect 4896 35634 4948 35640
rect 4550 34844 4858 34853
rect 4550 34842 4556 34844
rect 4612 34842 4636 34844
rect 4692 34842 4716 34844
rect 4772 34842 4796 34844
rect 4852 34842 4858 34844
rect 4612 34790 4614 34842
rect 4794 34790 4796 34842
rect 4550 34788 4556 34790
rect 4612 34788 4636 34790
rect 4692 34788 4716 34790
rect 4772 34788 4796 34790
rect 4852 34788 4858 34790
rect 4550 34779 4858 34788
rect 4550 33756 4858 33765
rect 4550 33754 4556 33756
rect 4612 33754 4636 33756
rect 4692 33754 4716 33756
rect 4772 33754 4796 33756
rect 4852 33754 4858 33756
rect 4612 33702 4614 33754
rect 4794 33702 4796 33754
rect 4550 33700 4556 33702
rect 4612 33700 4636 33702
rect 4692 33700 4716 33702
rect 4772 33700 4796 33702
rect 4852 33700 4858 33702
rect 4550 33691 4858 33700
rect 4550 32668 4858 32677
rect 4550 32666 4556 32668
rect 4612 32666 4636 32668
rect 4692 32666 4716 32668
rect 4772 32666 4796 32668
rect 4852 32666 4858 32668
rect 4612 32614 4614 32666
rect 4794 32614 4796 32666
rect 4550 32612 4556 32614
rect 4612 32612 4636 32614
rect 4692 32612 4716 32614
rect 4772 32612 4796 32614
rect 4852 32612 4858 32614
rect 4550 32603 4858 32612
rect 4896 32224 4948 32230
rect 4896 32166 4948 32172
rect 4550 31580 4858 31589
rect 4550 31578 4556 31580
rect 4612 31578 4636 31580
rect 4692 31578 4716 31580
rect 4772 31578 4796 31580
rect 4852 31578 4858 31580
rect 4612 31526 4614 31578
rect 4794 31526 4796 31578
rect 4550 31524 4556 31526
rect 4612 31524 4636 31526
rect 4692 31524 4716 31526
rect 4772 31524 4796 31526
rect 4852 31524 4858 31526
rect 4550 31515 4858 31524
rect 4550 30492 4858 30501
rect 4550 30490 4556 30492
rect 4612 30490 4636 30492
rect 4692 30490 4716 30492
rect 4772 30490 4796 30492
rect 4852 30490 4858 30492
rect 4612 30438 4614 30490
rect 4794 30438 4796 30490
rect 4550 30436 4556 30438
rect 4612 30436 4636 30438
rect 4692 30436 4716 30438
rect 4772 30436 4796 30438
rect 4852 30436 4858 30438
rect 4550 30427 4858 30436
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 4816 29578 4844 30262
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4550 29404 4858 29413
rect 4550 29402 4556 29404
rect 4612 29402 4636 29404
rect 4692 29402 4716 29404
rect 4772 29402 4796 29404
rect 4852 29402 4858 29404
rect 4612 29350 4614 29402
rect 4794 29350 4796 29402
rect 4550 29348 4556 29350
rect 4612 29348 4636 29350
rect 4692 29348 4716 29350
rect 4772 29348 4796 29350
rect 4852 29348 4858 29350
rect 4550 29339 4858 29348
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4816 28422 4844 28902
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 4550 28316 4858 28325
rect 4550 28314 4556 28316
rect 4612 28314 4636 28316
rect 4692 28314 4716 28316
rect 4772 28314 4796 28316
rect 4852 28314 4858 28316
rect 4612 28262 4614 28314
rect 4794 28262 4796 28314
rect 4550 28260 4556 28262
rect 4612 28260 4636 28262
rect 4692 28260 4716 28262
rect 4772 28260 4796 28262
rect 4852 28260 4858 28262
rect 4550 28251 4858 28260
rect 4550 27228 4858 27237
rect 4550 27226 4556 27228
rect 4612 27226 4636 27228
rect 4692 27226 4716 27228
rect 4772 27226 4796 27228
rect 4852 27226 4858 27228
rect 4612 27174 4614 27226
rect 4794 27174 4796 27226
rect 4550 27172 4556 27174
rect 4612 27172 4636 27174
rect 4692 27172 4716 27174
rect 4772 27172 4796 27174
rect 4852 27172 4858 27174
rect 4550 27163 4858 27172
rect 4550 26140 4858 26149
rect 4550 26138 4556 26140
rect 4612 26138 4636 26140
rect 4692 26138 4716 26140
rect 4772 26138 4796 26140
rect 4852 26138 4858 26140
rect 4612 26086 4614 26138
rect 4794 26086 4796 26138
rect 4550 26084 4556 26086
rect 4612 26084 4636 26086
rect 4692 26084 4716 26086
rect 4772 26084 4796 26086
rect 4852 26084 4858 26086
rect 4550 26075 4858 26084
rect 4550 25052 4858 25061
rect 4550 25050 4556 25052
rect 4612 25050 4636 25052
rect 4692 25050 4716 25052
rect 4772 25050 4796 25052
rect 4852 25050 4858 25052
rect 4612 24998 4614 25050
rect 4794 24998 4796 25050
rect 4550 24996 4556 24998
rect 4612 24996 4636 24998
rect 4692 24996 4716 24998
rect 4772 24996 4796 24998
rect 4852 24996 4858 24998
rect 4550 24987 4858 24996
rect 4550 23964 4858 23973
rect 4550 23962 4556 23964
rect 4612 23962 4636 23964
rect 4692 23962 4716 23964
rect 4772 23962 4796 23964
rect 4852 23962 4858 23964
rect 4612 23910 4614 23962
rect 4794 23910 4796 23962
rect 4550 23908 4556 23910
rect 4612 23908 4636 23910
rect 4692 23908 4716 23910
rect 4772 23908 4796 23910
rect 4852 23908 4858 23910
rect 4550 23899 4858 23908
rect 4550 22876 4858 22885
rect 4550 22874 4556 22876
rect 4612 22874 4636 22876
rect 4692 22874 4716 22876
rect 4772 22874 4796 22876
rect 4852 22874 4858 22876
rect 4612 22822 4614 22874
rect 4794 22822 4796 22874
rect 4550 22820 4556 22822
rect 4612 22820 4636 22822
rect 4692 22820 4716 22822
rect 4772 22820 4796 22822
rect 4852 22820 4858 22822
rect 4550 22811 4858 22820
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4540 22030 4568 22714
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4632 22166 4660 22374
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4550 21788 4858 21797
rect 4550 21786 4556 21788
rect 4612 21786 4636 21788
rect 4692 21786 4716 21788
rect 4772 21786 4796 21788
rect 4852 21786 4858 21788
rect 4612 21734 4614 21786
rect 4794 21734 4796 21786
rect 4550 21732 4556 21734
rect 4612 21732 4636 21734
rect 4692 21732 4716 21734
rect 4772 21732 4796 21734
rect 4852 21732 4858 21734
rect 4550 21723 4858 21732
rect 4550 20700 4858 20709
rect 4550 20698 4556 20700
rect 4612 20698 4636 20700
rect 4692 20698 4716 20700
rect 4772 20698 4796 20700
rect 4852 20698 4858 20700
rect 4612 20646 4614 20698
rect 4794 20646 4796 20698
rect 4550 20644 4556 20646
rect 4612 20644 4636 20646
rect 4692 20644 4716 20646
rect 4772 20644 4796 20646
rect 4852 20644 4858 20646
rect 4550 20635 4858 20644
rect 4550 19612 4858 19621
rect 4550 19610 4556 19612
rect 4612 19610 4636 19612
rect 4692 19610 4716 19612
rect 4772 19610 4796 19612
rect 4852 19610 4858 19612
rect 4612 19558 4614 19610
rect 4794 19558 4796 19610
rect 4550 19556 4556 19558
rect 4612 19556 4636 19558
rect 4692 19556 4716 19558
rect 4772 19556 4796 19558
rect 4852 19556 4858 19558
rect 4550 19547 4858 19556
rect 4908 18766 4936 32166
rect 5000 30190 5028 36586
rect 4988 30184 5040 30190
rect 4988 30126 5040 30132
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 5000 26382 5028 29990
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 5092 26296 5120 40038
rect 5210 39740 5518 39749
rect 5210 39738 5216 39740
rect 5272 39738 5296 39740
rect 5352 39738 5376 39740
rect 5432 39738 5456 39740
rect 5512 39738 5518 39740
rect 5272 39686 5274 39738
rect 5454 39686 5456 39738
rect 5210 39684 5216 39686
rect 5272 39684 5296 39686
rect 5352 39684 5376 39686
rect 5432 39684 5456 39686
rect 5512 39684 5518 39686
rect 5210 39675 5518 39684
rect 5552 39642 5580 41958
rect 5644 40730 5672 44775
rect 5736 42770 5764 46650
rect 5724 42764 5776 42770
rect 5724 42706 5776 42712
rect 5828 41414 5856 53094
rect 5920 52698 5948 58278
rect 6012 54194 6040 62086
rect 6150 62044 6458 62053
rect 6150 62042 6156 62044
rect 6212 62042 6236 62044
rect 6292 62042 6316 62044
rect 6372 62042 6396 62044
rect 6452 62042 6458 62044
rect 6212 61990 6214 62042
rect 6394 61990 6396 62042
rect 6150 61988 6156 61990
rect 6212 61988 6236 61990
rect 6292 61988 6316 61990
rect 6372 61988 6396 61990
rect 6452 61988 6458 61990
rect 6150 61979 6458 61988
rect 6564 61810 6592 62834
rect 6552 61804 6604 61810
rect 6552 61746 6604 61752
rect 6150 60956 6458 60965
rect 6150 60954 6156 60956
rect 6212 60954 6236 60956
rect 6292 60954 6316 60956
rect 6372 60954 6396 60956
rect 6452 60954 6458 60956
rect 6212 60902 6214 60954
rect 6394 60902 6396 60954
rect 6150 60900 6156 60902
rect 6212 60900 6236 60902
rect 6292 60900 6316 60902
rect 6372 60900 6396 60902
rect 6452 60900 6458 60902
rect 6150 60891 6458 60900
rect 6564 60722 6592 61746
rect 6552 60716 6604 60722
rect 6552 60658 6604 60664
rect 6552 60512 6604 60518
rect 6552 60454 6604 60460
rect 6150 59868 6458 59877
rect 6150 59866 6156 59868
rect 6212 59866 6236 59868
rect 6292 59866 6316 59868
rect 6372 59866 6396 59868
rect 6452 59866 6458 59868
rect 6212 59814 6214 59866
rect 6394 59814 6396 59866
rect 6150 59812 6156 59814
rect 6212 59812 6236 59814
rect 6292 59812 6316 59814
rect 6372 59812 6396 59814
rect 6452 59812 6458 59814
rect 6150 59803 6458 59812
rect 6564 59158 6592 60454
rect 6552 59152 6604 59158
rect 6552 59094 6604 59100
rect 6552 59016 6604 59022
rect 6552 58958 6604 58964
rect 6150 58780 6458 58789
rect 6150 58778 6156 58780
rect 6212 58778 6236 58780
rect 6292 58778 6316 58780
rect 6372 58778 6396 58780
rect 6452 58778 6458 58780
rect 6212 58726 6214 58778
rect 6394 58726 6396 58778
rect 6150 58724 6156 58726
rect 6212 58724 6236 58726
rect 6292 58724 6316 58726
rect 6372 58724 6396 58726
rect 6452 58724 6458 58726
rect 6150 58715 6458 58724
rect 6092 58676 6144 58682
rect 6092 58618 6144 58624
rect 6368 58676 6420 58682
rect 6368 58618 6420 58624
rect 6104 57798 6132 58618
rect 6380 57934 6408 58618
rect 6460 58336 6512 58342
rect 6460 58278 6512 58284
rect 6368 57928 6420 57934
rect 6472 57905 6500 58278
rect 6368 57870 6420 57876
rect 6458 57896 6514 57905
rect 6458 57831 6514 57840
rect 6092 57792 6144 57798
rect 6092 57734 6144 57740
rect 6150 57692 6458 57701
rect 6150 57690 6156 57692
rect 6212 57690 6236 57692
rect 6292 57690 6316 57692
rect 6372 57690 6396 57692
rect 6452 57690 6458 57692
rect 6212 57638 6214 57690
rect 6394 57638 6396 57690
rect 6150 57636 6156 57638
rect 6212 57636 6236 57638
rect 6292 57636 6316 57638
rect 6372 57636 6396 57638
rect 6452 57636 6458 57638
rect 6150 57627 6458 57636
rect 6564 57594 6592 58958
rect 6276 57588 6328 57594
rect 6276 57530 6328 57536
rect 6368 57588 6420 57594
rect 6368 57530 6420 57536
rect 6552 57588 6604 57594
rect 6552 57530 6604 57536
rect 6288 56914 6316 57530
rect 6380 57458 6408 57530
rect 6550 57488 6606 57497
rect 6368 57452 6420 57458
rect 6550 57423 6606 57432
rect 6368 57394 6420 57400
rect 6368 57316 6420 57322
rect 6368 57258 6420 57264
rect 6276 56908 6328 56914
rect 6276 56850 6328 56856
rect 6380 56710 6408 57258
rect 6368 56704 6420 56710
rect 6368 56646 6420 56652
rect 6150 56604 6458 56613
rect 6150 56602 6156 56604
rect 6212 56602 6236 56604
rect 6292 56602 6316 56604
rect 6372 56602 6396 56604
rect 6452 56602 6458 56604
rect 6212 56550 6214 56602
rect 6394 56550 6396 56602
rect 6150 56548 6156 56550
rect 6212 56548 6236 56550
rect 6292 56548 6316 56550
rect 6372 56548 6396 56550
rect 6452 56548 6458 56550
rect 6150 56539 6458 56548
rect 6150 55516 6458 55525
rect 6150 55514 6156 55516
rect 6212 55514 6236 55516
rect 6292 55514 6316 55516
rect 6372 55514 6396 55516
rect 6452 55514 6458 55516
rect 6212 55462 6214 55514
rect 6394 55462 6396 55514
rect 6150 55460 6156 55462
rect 6212 55460 6236 55462
rect 6292 55460 6316 55462
rect 6372 55460 6396 55462
rect 6452 55460 6458 55462
rect 6150 55451 6458 55460
rect 6150 54428 6458 54437
rect 6150 54426 6156 54428
rect 6212 54426 6236 54428
rect 6292 54426 6316 54428
rect 6372 54426 6396 54428
rect 6452 54426 6458 54428
rect 6212 54374 6214 54426
rect 6394 54374 6396 54426
rect 6150 54372 6156 54374
rect 6212 54372 6236 54374
rect 6292 54372 6316 54374
rect 6372 54372 6396 54374
rect 6452 54372 6458 54374
rect 6150 54363 6458 54372
rect 6000 54188 6052 54194
rect 6000 54130 6052 54136
rect 5998 53544 6054 53553
rect 5998 53479 6054 53488
rect 5908 52692 5960 52698
rect 5908 52634 5960 52640
rect 5908 52352 5960 52358
rect 5908 52294 5960 52300
rect 5920 52154 5948 52294
rect 5908 52148 5960 52154
rect 5908 52090 5960 52096
rect 5908 51400 5960 51406
rect 5908 51342 5960 51348
rect 6012 51354 6040 53479
rect 6150 53340 6458 53349
rect 6150 53338 6156 53340
rect 6212 53338 6236 53340
rect 6292 53338 6316 53340
rect 6372 53338 6396 53340
rect 6452 53338 6458 53340
rect 6212 53286 6214 53338
rect 6394 53286 6396 53338
rect 6150 53284 6156 53286
rect 6212 53284 6236 53286
rect 6292 53284 6316 53286
rect 6372 53284 6396 53286
rect 6452 53284 6458 53286
rect 6150 53275 6458 53284
rect 6460 53100 6512 53106
rect 6460 53042 6512 53048
rect 6184 52896 6236 52902
rect 6184 52838 6236 52844
rect 6196 52494 6224 52838
rect 6184 52488 6236 52494
rect 6184 52430 6236 52436
rect 6472 52358 6500 53042
rect 6460 52352 6512 52358
rect 6460 52294 6512 52300
rect 6150 52252 6458 52261
rect 6150 52250 6156 52252
rect 6212 52250 6236 52252
rect 6292 52250 6316 52252
rect 6372 52250 6396 52252
rect 6452 52250 6458 52252
rect 6212 52198 6214 52250
rect 6394 52198 6396 52250
rect 6150 52196 6156 52198
rect 6212 52196 6236 52198
rect 6292 52196 6316 52198
rect 6372 52196 6396 52198
rect 6452 52196 6458 52198
rect 6150 52187 6458 52196
rect 6564 52136 6592 57423
rect 6656 56778 6684 67544
rect 6748 67182 6776 67606
rect 6920 67594 6972 67600
rect 7012 67652 7064 67658
rect 7012 67594 7064 67600
rect 7104 67652 7156 67658
rect 7104 67594 7156 67600
rect 6932 67289 6960 67594
rect 7024 67386 7052 67594
rect 7012 67380 7064 67386
rect 7012 67322 7064 67328
rect 6918 67280 6974 67289
rect 6918 67215 6974 67224
rect 6736 67176 6788 67182
rect 6736 67118 6788 67124
rect 7116 67130 7144 67594
rect 7208 67250 7236 69838
rect 7300 67402 7328 69838
rect 7392 69426 7420 69838
rect 7380 69420 7432 69426
rect 7380 69362 7432 69368
rect 7392 68785 7420 69362
rect 7378 68776 7434 68785
rect 7378 68711 7434 68720
rect 7380 68332 7432 68338
rect 7380 68274 7432 68280
rect 7392 67726 7420 68274
rect 7484 67794 7512 72422
rect 7576 71126 7604 72791
rect 7656 72684 7708 72690
rect 7656 72626 7708 72632
rect 7932 72684 7984 72690
rect 7932 72626 7984 72632
rect 7668 72282 7696 72626
rect 7748 72480 7800 72486
rect 7748 72422 7800 72428
rect 7656 72276 7708 72282
rect 7656 72218 7708 72224
rect 7760 71924 7788 72422
rect 7944 72214 7972 72626
rect 8024 72616 8076 72622
rect 8024 72558 8076 72564
rect 7932 72208 7984 72214
rect 7930 72176 7932 72185
rect 7984 72176 7986 72185
rect 7930 72111 7986 72120
rect 8036 72078 8064 72558
rect 8024 72072 8076 72078
rect 8024 72014 8076 72020
rect 7668 71896 7788 71924
rect 7564 71120 7616 71126
rect 7564 71062 7616 71068
rect 7668 70904 7696 71896
rect 7750 71836 8058 71845
rect 7750 71834 7756 71836
rect 7812 71834 7836 71836
rect 7892 71834 7916 71836
rect 7972 71834 7996 71836
rect 8052 71834 8058 71836
rect 7812 71782 7814 71834
rect 7994 71782 7996 71834
rect 7750 71780 7756 71782
rect 7812 71780 7836 71782
rect 7892 71780 7916 71782
rect 7972 71780 7996 71782
rect 8052 71780 8058 71782
rect 7750 71771 8058 71780
rect 7838 71632 7894 71641
rect 7748 71596 7800 71602
rect 7838 71567 7894 71576
rect 7748 71538 7800 71544
rect 7576 70876 7696 70904
rect 7576 69018 7604 70876
rect 7760 70836 7788 71538
rect 7852 71194 7880 71567
rect 7932 71392 7984 71398
rect 7932 71334 7984 71340
rect 7840 71188 7892 71194
rect 7840 71130 7892 71136
rect 7944 71058 7972 71334
rect 7932 71052 7984 71058
rect 7932 70994 7984 71000
rect 7668 70808 7788 70836
rect 7668 70514 7696 70808
rect 7750 70748 8058 70757
rect 7750 70746 7756 70748
rect 7812 70746 7836 70748
rect 7892 70746 7916 70748
rect 7972 70746 7996 70748
rect 8052 70746 8058 70748
rect 7812 70694 7814 70746
rect 7994 70694 7996 70746
rect 7750 70692 7756 70694
rect 7812 70692 7836 70694
rect 7892 70692 7916 70694
rect 7972 70692 7996 70694
rect 8052 70692 8058 70694
rect 7750 70683 8058 70692
rect 7748 70644 7800 70650
rect 7748 70586 7800 70592
rect 7760 70553 7788 70586
rect 7746 70544 7802 70553
rect 7656 70508 7708 70514
rect 8022 70544 8078 70553
rect 7746 70479 7802 70488
rect 7944 70502 8022 70530
rect 7656 70450 7708 70456
rect 7656 70304 7708 70310
rect 7656 70246 7708 70252
rect 7564 69012 7616 69018
rect 7564 68954 7616 68960
rect 7668 68728 7696 70246
rect 7944 69970 7972 70502
rect 8022 70479 8078 70488
rect 8024 70372 8076 70378
rect 8024 70314 8076 70320
rect 7932 69964 7984 69970
rect 7932 69906 7984 69912
rect 7748 69760 7800 69766
rect 8036 69748 8064 70314
rect 7800 69720 8064 69748
rect 7748 69702 7800 69708
rect 7750 69660 8058 69669
rect 7750 69658 7756 69660
rect 7812 69658 7836 69660
rect 7892 69658 7916 69660
rect 7972 69658 7996 69660
rect 8052 69658 8058 69660
rect 7812 69606 7814 69658
rect 7994 69606 7996 69658
rect 7750 69604 7756 69606
rect 7812 69604 7836 69606
rect 7892 69604 7916 69606
rect 7972 69604 7996 69606
rect 8052 69604 8058 69606
rect 7750 69595 8058 69604
rect 7748 69556 7800 69562
rect 7748 69498 7800 69504
rect 7576 68700 7696 68728
rect 7576 67946 7604 68700
rect 7760 68660 7788 69498
rect 8024 69488 8076 69494
rect 8024 69430 8076 69436
rect 7932 69352 7984 69358
rect 7932 69294 7984 69300
rect 7944 68746 7972 69294
rect 7932 68740 7984 68746
rect 7932 68682 7984 68688
rect 8036 68678 8064 69430
rect 7668 68632 7788 68660
rect 8024 68672 8076 68678
rect 7668 68218 7696 68632
rect 8024 68614 8076 68620
rect 7750 68572 8058 68581
rect 7750 68570 7756 68572
rect 7812 68570 7836 68572
rect 7892 68570 7916 68572
rect 7972 68570 7996 68572
rect 8052 68570 8058 68572
rect 7812 68518 7814 68570
rect 7994 68518 7996 68570
rect 7750 68516 7756 68518
rect 7812 68516 7836 68518
rect 7892 68516 7916 68518
rect 7972 68516 7996 68518
rect 8052 68516 8058 68518
rect 7750 68507 8058 68516
rect 7932 68468 7984 68474
rect 7932 68410 7984 68416
rect 7944 68338 7972 68410
rect 8128 68354 8156 73086
rect 8220 72554 8248 73238
rect 8208 72548 8260 72554
rect 8208 72490 8260 72496
rect 8208 71596 8260 71602
rect 8208 71538 8260 71544
rect 8220 70961 8248 71538
rect 8206 70952 8262 70961
rect 8206 70887 8262 70896
rect 8220 70514 8248 70887
rect 8208 70508 8260 70514
rect 8208 70450 8260 70456
rect 8208 70032 8260 70038
rect 8208 69974 8260 69980
rect 8220 69494 8248 69974
rect 8208 69488 8260 69494
rect 8208 69430 8260 69436
rect 8208 69216 8260 69222
rect 8208 69158 8260 69164
rect 8036 68338 8156 68354
rect 7932 68332 7984 68338
rect 7932 68274 7984 68280
rect 8024 68332 8156 68338
rect 8076 68326 8156 68332
rect 8024 68274 8076 68280
rect 7930 68232 7986 68241
rect 7668 68190 7880 68218
rect 7576 67918 7696 67946
rect 7472 67788 7524 67794
rect 7472 67730 7524 67736
rect 7380 67720 7432 67726
rect 7380 67662 7432 67668
rect 7668 67634 7696 67918
rect 7852 67912 7880 68190
rect 7930 68167 7986 68176
rect 7944 67930 7972 68167
rect 8024 68128 8076 68134
rect 8024 68070 8076 68076
rect 7576 67606 7696 67634
rect 7760 67884 7880 67912
rect 7932 67924 7984 67930
rect 7300 67374 7512 67402
rect 7380 67312 7432 67318
rect 7380 67254 7432 67260
rect 7196 67244 7248 67250
rect 7196 67186 7248 67192
rect 7116 67102 7236 67130
rect 6736 67040 6788 67046
rect 6736 66982 6788 66988
rect 6748 63442 6776 66982
rect 6810 66940 7118 66949
rect 6810 66938 6816 66940
rect 6872 66938 6896 66940
rect 6952 66938 6976 66940
rect 7032 66938 7056 66940
rect 7112 66938 7118 66940
rect 6872 66886 6874 66938
rect 7054 66886 7056 66938
rect 6810 66884 6816 66886
rect 6872 66884 6896 66886
rect 6952 66884 6976 66886
rect 7032 66884 7056 66886
rect 7112 66884 7118 66886
rect 6810 66875 7118 66884
rect 7208 66774 7236 67102
rect 7196 66768 7248 66774
rect 7392 66756 7420 67254
rect 7356 66728 7420 66756
rect 7356 66722 7384 66728
rect 7196 66710 7248 66716
rect 7305 66694 7384 66722
rect 7305 66688 7333 66694
rect 7300 66660 7333 66688
rect 7012 66632 7064 66638
rect 7012 66574 7064 66580
rect 7024 65958 7052 66574
rect 7196 66496 7248 66502
rect 7196 66438 7248 66444
rect 7012 65952 7064 65958
rect 7012 65894 7064 65900
rect 6810 65852 7118 65861
rect 6810 65850 6816 65852
rect 6872 65850 6896 65852
rect 6952 65850 6976 65852
rect 7032 65850 7056 65852
rect 7112 65850 7118 65852
rect 6872 65798 6874 65850
rect 7054 65798 7056 65850
rect 6810 65796 6816 65798
rect 6872 65796 6896 65798
rect 6952 65796 6976 65798
rect 7032 65796 7056 65798
rect 7112 65796 7118 65798
rect 6810 65787 7118 65796
rect 7104 65748 7156 65754
rect 7104 65690 7156 65696
rect 7012 65476 7064 65482
rect 7012 65418 7064 65424
rect 6828 65408 6880 65414
rect 6828 65350 6880 65356
rect 6840 64870 6868 65350
rect 7024 64977 7052 65418
rect 7010 64968 7066 64977
rect 7116 64938 7144 65690
rect 7010 64903 7066 64912
rect 7104 64932 7156 64938
rect 7104 64874 7156 64880
rect 6828 64864 6880 64870
rect 6828 64806 6880 64812
rect 6810 64764 7118 64773
rect 6810 64762 6816 64764
rect 6872 64762 6896 64764
rect 6952 64762 6976 64764
rect 7032 64762 7056 64764
rect 7112 64762 7118 64764
rect 6872 64710 6874 64762
rect 7054 64710 7056 64762
rect 6810 64708 6816 64710
rect 6872 64708 6896 64710
rect 6952 64708 6976 64710
rect 7032 64708 7056 64710
rect 7112 64708 7118 64710
rect 6810 64699 7118 64708
rect 6826 64560 6882 64569
rect 6826 64495 6882 64504
rect 6840 63782 6868 64495
rect 7104 64456 7156 64462
rect 7104 64398 7156 64404
rect 6828 63776 6880 63782
rect 7116 63764 7144 64398
rect 7208 63986 7236 66438
rect 7300 66254 7328 66660
rect 7380 66632 7432 66638
rect 7484 66586 7512 67374
rect 7432 66580 7512 66586
rect 7380 66574 7512 66580
rect 7392 66558 7512 66574
rect 7576 66314 7604 67606
rect 7760 67572 7788 67884
rect 7932 67866 7984 67872
rect 7668 67544 7788 67572
rect 8036 67572 8064 68070
rect 8220 67708 8248 69158
rect 8312 67794 8340 73510
rect 8410 73468 8718 73477
rect 8410 73466 8416 73468
rect 8472 73466 8496 73468
rect 8552 73466 8576 73468
rect 8632 73466 8656 73468
rect 8712 73466 8718 73468
rect 8472 73414 8474 73466
rect 8654 73414 8656 73466
rect 8410 73412 8416 73414
rect 8472 73412 8496 73414
rect 8552 73412 8576 73414
rect 8632 73412 8656 73414
rect 8712 73412 8718 73414
rect 8410 73403 8718 73412
rect 8484 73364 8536 73370
rect 8484 73306 8536 73312
rect 8392 73296 8444 73302
rect 8392 73238 8444 73244
rect 8404 73166 8432 73238
rect 8392 73160 8444 73166
rect 8496 73137 8524 73306
rect 8666 73264 8722 73273
rect 8666 73199 8722 73208
rect 8392 73102 8444 73108
rect 8482 73128 8538 73137
rect 8404 72729 8432 73102
rect 8482 73063 8538 73072
rect 8484 73024 8536 73030
rect 8484 72966 8536 72972
rect 8496 72826 8524 72966
rect 8484 72820 8536 72826
rect 8484 72762 8536 72768
rect 8390 72720 8446 72729
rect 8496 72690 8524 72762
rect 8390 72655 8392 72664
rect 8444 72655 8446 72664
rect 8484 72684 8536 72690
rect 8392 72626 8444 72632
rect 8484 72626 8536 72632
rect 8680 72536 8708 73199
rect 8772 72978 8800 74666
rect 8864 73166 8892 76298
rect 8956 74390 8984 76434
rect 8944 74384 8996 74390
rect 8944 74326 8996 74332
rect 9048 74254 9076 77114
rect 9140 74780 9168 85546
rect 9232 75342 9260 85750
rect 10324 85468 10376 85474
rect 10324 85410 10376 85416
rect 10140 85332 10192 85338
rect 10140 85274 10192 85280
rect 9350 84892 9658 84901
rect 9350 84890 9356 84892
rect 9412 84890 9436 84892
rect 9492 84890 9516 84892
rect 9572 84890 9596 84892
rect 9652 84890 9658 84892
rect 9412 84838 9414 84890
rect 9594 84838 9596 84890
rect 9350 84836 9356 84838
rect 9412 84836 9436 84838
rect 9492 84836 9516 84838
rect 9572 84836 9596 84838
rect 9652 84836 9658 84838
rect 9350 84827 9658 84836
rect 9350 83804 9658 83813
rect 9350 83802 9356 83804
rect 9412 83802 9436 83804
rect 9492 83802 9516 83804
rect 9572 83802 9596 83804
rect 9652 83802 9658 83804
rect 9412 83750 9414 83802
rect 9594 83750 9596 83802
rect 9350 83748 9356 83750
rect 9412 83748 9436 83750
rect 9492 83748 9516 83750
rect 9572 83748 9596 83750
rect 9652 83748 9658 83750
rect 9350 83739 9658 83748
rect 9350 82716 9658 82725
rect 9350 82714 9356 82716
rect 9412 82714 9436 82716
rect 9492 82714 9516 82716
rect 9572 82714 9596 82716
rect 9652 82714 9658 82716
rect 9412 82662 9414 82714
rect 9594 82662 9596 82714
rect 9350 82660 9356 82662
rect 9412 82660 9436 82662
rect 9492 82660 9516 82662
rect 9572 82660 9596 82662
rect 9652 82660 9658 82662
rect 9350 82651 9658 82660
rect 9350 81628 9658 81637
rect 9350 81626 9356 81628
rect 9412 81626 9436 81628
rect 9492 81626 9516 81628
rect 9572 81626 9596 81628
rect 9652 81626 9658 81628
rect 9412 81574 9414 81626
rect 9594 81574 9596 81626
rect 9350 81572 9356 81574
rect 9412 81572 9436 81574
rect 9492 81572 9516 81574
rect 9572 81572 9596 81574
rect 9652 81572 9658 81574
rect 9350 81563 9658 81572
rect 9350 80540 9658 80549
rect 9350 80538 9356 80540
rect 9412 80538 9436 80540
rect 9492 80538 9516 80540
rect 9572 80538 9596 80540
rect 9652 80538 9658 80540
rect 9412 80486 9414 80538
rect 9594 80486 9596 80538
rect 9350 80484 9356 80486
rect 9412 80484 9436 80486
rect 9492 80484 9516 80486
rect 9572 80484 9596 80486
rect 9652 80484 9658 80486
rect 9350 80475 9658 80484
rect 9350 79452 9658 79461
rect 9350 79450 9356 79452
rect 9412 79450 9436 79452
rect 9492 79450 9516 79452
rect 9572 79450 9596 79452
rect 9652 79450 9658 79452
rect 9412 79398 9414 79450
rect 9594 79398 9596 79450
rect 9350 79396 9356 79398
rect 9412 79396 9436 79398
rect 9492 79396 9516 79398
rect 9572 79396 9596 79398
rect 9652 79396 9658 79398
rect 9350 79387 9658 79396
rect 9350 78364 9658 78373
rect 9350 78362 9356 78364
rect 9412 78362 9436 78364
rect 9492 78362 9516 78364
rect 9572 78362 9596 78364
rect 9652 78362 9658 78364
rect 9412 78310 9414 78362
rect 9594 78310 9596 78362
rect 9350 78308 9356 78310
rect 9412 78308 9436 78310
rect 9492 78308 9516 78310
rect 9572 78308 9596 78310
rect 9652 78308 9658 78310
rect 9350 78299 9658 78308
rect 9350 77276 9658 77285
rect 9350 77274 9356 77276
rect 9412 77274 9436 77276
rect 9492 77274 9516 77276
rect 9572 77274 9596 77276
rect 9652 77274 9658 77276
rect 9412 77222 9414 77274
rect 9594 77222 9596 77274
rect 9350 77220 9356 77222
rect 9412 77220 9436 77222
rect 9492 77220 9516 77222
rect 9572 77220 9596 77222
rect 9652 77220 9658 77222
rect 9350 77211 9658 77220
rect 10152 77042 10180 85274
rect 10232 83496 10284 83502
rect 10232 83438 10284 83444
rect 10140 77036 10192 77042
rect 10140 76978 10192 76984
rect 9350 76188 9658 76197
rect 9350 76186 9356 76188
rect 9412 76186 9436 76188
rect 9492 76186 9516 76188
rect 9572 76186 9596 76188
rect 9652 76186 9658 76188
rect 9412 76134 9414 76186
rect 9594 76134 9596 76186
rect 9350 76132 9356 76134
rect 9412 76132 9436 76134
rect 9492 76132 9516 76134
rect 9572 76132 9596 76134
rect 9652 76132 9658 76134
rect 9350 76123 9658 76132
rect 9220 75336 9272 75342
rect 9220 75278 9272 75284
rect 9496 75336 9548 75342
rect 9548 75296 9674 75324
rect 9496 75278 9548 75284
rect 9646 75256 9674 75296
rect 9646 75228 9720 75256
rect 9350 75100 9658 75109
rect 9350 75098 9356 75100
rect 9412 75098 9436 75100
rect 9492 75098 9516 75100
rect 9572 75098 9596 75100
rect 9652 75098 9658 75100
rect 9412 75046 9414 75098
rect 9594 75046 9596 75098
rect 9350 75044 9356 75046
rect 9412 75044 9436 75046
rect 9492 75044 9516 75046
rect 9572 75044 9596 75046
rect 9652 75044 9658 75046
rect 9350 75035 9658 75044
rect 9588 74928 9640 74934
rect 9692 74882 9720 75228
rect 9640 74876 9720 74882
rect 9588 74870 9720 74876
rect 9600 74854 9720 74870
rect 9312 74792 9364 74798
rect 9140 74752 9312 74780
rect 9312 74734 9364 74740
rect 9404 74792 9456 74798
rect 9404 74734 9456 74740
rect 9324 74458 9352 74734
rect 9312 74452 9364 74458
rect 9312 74394 9364 74400
rect 9220 74384 9272 74390
rect 9220 74326 9272 74332
rect 9036 74248 9088 74254
rect 9036 74190 9088 74196
rect 9128 74180 9180 74186
rect 9128 74122 9180 74128
rect 8944 74112 8996 74118
rect 8944 74054 8996 74060
rect 9036 74112 9088 74118
rect 9036 74054 9088 74060
rect 8852 73160 8904 73166
rect 8852 73102 8904 73108
rect 8772 72950 8892 72978
rect 8864 72690 8892 72950
rect 8852 72684 8904 72690
rect 8852 72626 8904 72632
rect 8680 72508 8892 72536
rect 8576 72480 8628 72486
rect 8628 72440 8800 72468
rect 8576 72422 8628 72428
rect 8410 72380 8718 72389
rect 8410 72378 8416 72380
rect 8472 72378 8496 72380
rect 8552 72378 8576 72380
rect 8632 72378 8656 72380
rect 8712 72378 8718 72380
rect 8472 72326 8474 72378
rect 8654 72326 8656 72378
rect 8410 72324 8416 72326
rect 8472 72324 8496 72326
rect 8552 72324 8576 72326
rect 8632 72324 8656 72326
rect 8712 72324 8718 72326
rect 8410 72315 8718 72324
rect 8576 72140 8628 72146
rect 8576 72082 8628 72088
rect 8392 71936 8444 71942
rect 8392 71878 8444 71884
rect 8404 71505 8432 71878
rect 8588 71534 8616 72082
rect 8576 71528 8628 71534
rect 8390 71496 8446 71505
rect 8576 71470 8628 71476
rect 8390 71431 8446 71440
rect 8410 71292 8718 71301
rect 8410 71290 8416 71292
rect 8472 71290 8496 71292
rect 8552 71290 8576 71292
rect 8632 71290 8656 71292
rect 8712 71290 8718 71292
rect 8472 71238 8474 71290
rect 8654 71238 8656 71290
rect 8410 71236 8416 71238
rect 8472 71236 8496 71238
rect 8552 71236 8576 71238
rect 8632 71236 8656 71238
rect 8712 71236 8718 71238
rect 8410 71227 8718 71236
rect 8482 71088 8538 71097
rect 8392 71052 8444 71058
rect 8772 71040 8800 72440
rect 8482 71023 8484 71032
rect 8392 70994 8444 71000
rect 8536 71023 8538 71032
rect 8484 70994 8536 71000
rect 8680 71012 8800 71040
rect 8404 70514 8432 70994
rect 8576 70916 8628 70922
rect 8576 70858 8628 70864
rect 8484 70848 8536 70854
rect 8484 70790 8536 70796
rect 8496 70553 8524 70790
rect 8588 70650 8616 70858
rect 8576 70644 8628 70650
rect 8576 70586 8628 70592
rect 8482 70544 8538 70553
rect 8392 70508 8444 70514
rect 8482 70479 8538 70488
rect 8576 70508 8628 70514
rect 8392 70450 8444 70456
rect 8576 70450 8628 70456
rect 8588 70417 8616 70450
rect 8574 70408 8630 70417
rect 8574 70343 8630 70352
rect 8680 70292 8708 71012
rect 8864 70854 8892 72508
rect 8852 70848 8904 70854
rect 8852 70790 8904 70796
rect 8680 70264 8800 70292
rect 8410 70204 8718 70213
rect 8410 70202 8416 70204
rect 8472 70202 8496 70204
rect 8552 70202 8576 70204
rect 8632 70202 8656 70204
rect 8712 70202 8718 70204
rect 8472 70150 8474 70202
rect 8654 70150 8656 70202
rect 8410 70148 8416 70150
rect 8472 70148 8496 70150
rect 8552 70148 8576 70150
rect 8632 70148 8656 70150
rect 8712 70148 8718 70150
rect 8410 70139 8718 70148
rect 8392 70032 8444 70038
rect 8772 70020 8800 70264
rect 8772 69992 8892 70020
rect 8392 69974 8444 69980
rect 8404 69358 8432 69974
rect 8668 69964 8720 69970
rect 8588 69924 8668 69952
rect 8484 69896 8536 69902
rect 8484 69838 8536 69844
rect 8496 69766 8524 69838
rect 8484 69760 8536 69766
rect 8484 69702 8536 69708
rect 8588 69494 8616 69924
rect 8668 69906 8720 69912
rect 8760 69556 8812 69562
rect 8760 69498 8812 69504
rect 8576 69488 8628 69494
rect 8576 69430 8628 69436
rect 8392 69352 8444 69358
rect 8392 69294 8444 69300
rect 8410 69116 8718 69125
rect 8410 69114 8416 69116
rect 8472 69114 8496 69116
rect 8552 69114 8576 69116
rect 8632 69114 8656 69116
rect 8712 69114 8718 69116
rect 8472 69062 8474 69114
rect 8654 69062 8656 69114
rect 8410 69060 8416 69062
rect 8472 69060 8496 69062
rect 8552 69060 8576 69062
rect 8632 69060 8656 69062
rect 8712 69060 8718 69062
rect 8410 69051 8718 69060
rect 8484 69012 8536 69018
rect 8484 68954 8536 68960
rect 8390 68912 8446 68921
rect 8390 68847 8446 68856
rect 8404 68814 8432 68847
rect 8392 68808 8444 68814
rect 8392 68750 8444 68756
rect 8392 68672 8444 68678
rect 8392 68614 8444 68620
rect 8404 68134 8432 68614
rect 8496 68241 8524 68954
rect 8576 68944 8628 68950
rect 8574 68912 8576 68921
rect 8628 68912 8630 68921
rect 8574 68847 8630 68856
rect 8482 68232 8538 68241
rect 8482 68167 8538 68176
rect 8392 68128 8444 68134
rect 8392 68070 8444 68076
rect 8410 68028 8718 68037
rect 8410 68026 8416 68028
rect 8472 68026 8496 68028
rect 8552 68026 8576 68028
rect 8632 68026 8656 68028
rect 8712 68026 8718 68028
rect 8472 67974 8474 68026
rect 8654 67974 8656 68026
rect 8410 67972 8416 67974
rect 8472 67972 8496 67974
rect 8552 67972 8576 67974
rect 8632 67972 8656 67974
rect 8712 67972 8718 67974
rect 8410 67963 8718 67972
rect 8300 67788 8352 67794
rect 8300 67730 8352 67736
rect 8392 67788 8444 67794
rect 8392 67730 8444 67736
rect 8128 67680 8248 67708
rect 8128 67640 8156 67680
rect 8128 67612 8294 67640
rect 8036 67544 8156 67572
rect 7668 67368 7696 67544
rect 7750 67484 8058 67493
rect 7750 67482 7756 67484
rect 7812 67482 7836 67484
rect 7892 67482 7916 67484
rect 7972 67482 7996 67484
rect 8052 67482 8058 67484
rect 7812 67430 7814 67482
rect 7994 67430 7996 67482
rect 7750 67428 7756 67430
rect 7812 67428 7836 67430
rect 7892 67428 7916 67430
rect 7972 67428 7996 67430
rect 8052 67428 8058 67430
rect 7750 67419 8058 67428
rect 7668 67340 7788 67368
rect 7760 67250 7788 67340
rect 7656 67244 7708 67250
rect 7656 67186 7708 67192
rect 7748 67244 7800 67250
rect 7748 67186 7800 67192
rect 7668 67114 7696 67186
rect 7656 67108 7708 67114
rect 7656 67050 7708 67056
rect 7567 66286 7604 66314
rect 7668 66298 7696 67050
rect 7760 66502 7788 67186
rect 7932 67176 7984 67182
rect 7932 67118 7984 67124
rect 7840 67108 7892 67114
rect 7840 67050 7892 67056
rect 7748 66496 7800 66502
rect 7852 66484 7880 67050
rect 7944 66774 7972 67118
rect 7932 66768 7984 66774
rect 7932 66710 7984 66716
rect 8128 66706 8156 67544
rect 8266 67300 8294 67612
rect 8220 67272 8294 67300
rect 8116 66700 8168 66706
rect 8116 66642 8168 66648
rect 7852 66456 8156 66484
rect 7748 66438 7800 66444
rect 7750 66396 8058 66405
rect 7750 66394 7756 66396
rect 7812 66394 7836 66396
rect 7892 66394 7916 66396
rect 7972 66394 7996 66396
rect 8052 66394 8058 66396
rect 7812 66342 7814 66394
rect 7994 66342 7996 66394
rect 7750 66340 7756 66342
rect 7812 66340 7836 66342
rect 7892 66340 7916 66342
rect 7972 66340 7996 66342
rect 8052 66340 8058 66342
rect 7750 66331 8058 66340
rect 7656 66292 7708 66298
rect 7300 66226 7512 66254
rect 7288 66156 7340 66162
rect 7288 66098 7340 66104
rect 7300 65618 7328 66098
rect 7378 66056 7434 66065
rect 7378 65991 7434 66000
rect 7288 65612 7340 65618
rect 7288 65554 7340 65560
rect 7288 65408 7340 65414
rect 7288 65350 7340 65356
rect 7196 63980 7248 63986
rect 7196 63922 7248 63928
rect 7116 63736 7236 63764
rect 6828 63718 6880 63724
rect 6810 63676 7118 63685
rect 6810 63674 6816 63676
rect 6872 63674 6896 63676
rect 6952 63674 6976 63676
rect 7032 63674 7056 63676
rect 7112 63674 7118 63676
rect 6872 63622 6874 63674
rect 7054 63622 7056 63674
rect 6810 63620 6816 63622
rect 6872 63620 6896 63622
rect 6952 63620 6976 63622
rect 7032 63620 7056 63622
rect 7112 63620 7118 63622
rect 6810 63611 7118 63620
rect 7208 63492 7236 63736
rect 7116 63464 7236 63492
rect 6736 63436 6788 63442
rect 6736 63378 6788 63384
rect 6828 63232 6880 63238
rect 6828 63174 6880 63180
rect 6736 63028 6788 63034
rect 6736 62970 6788 62976
rect 6748 56846 6776 62970
rect 6840 62898 6868 63174
rect 7116 62898 7144 63464
rect 7196 63368 7248 63374
rect 7196 63310 7248 63316
rect 6828 62892 6880 62898
rect 6828 62834 6880 62840
rect 7104 62892 7156 62898
rect 7104 62834 7156 62840
rect 6840 62801 6868 62834
rect 6826 62792 6882 62801
rect 6826 62727 6882 62736
rect 6810 62588 7118 62597
rect 6810 62586 6816 62588
rect 6872 62586 6896 62588
rect 6952 62586 6976 62588
rect 7032 62586 7056 62588
rect 7112 62586 7118 62588
rect 6872 62534 6874 62586
rect 7054 62534 7056 62586
rect 6810 62532 6816 62534
rect 6872 62532 6896 62534
rect 6952 62532 6976 62534
rect 7032 62532 7056 62534
rect 7112 62532 7118 62534
rect 6810 62523 7118 62532
rect 7208 62354 7236 63310
rect 7300 62354 7328 65350
rect 7196 62348 7248 62354
rect 7196 62290 7248 62296
rect 7288 62348 7340 62354
rect 7288 62290 7340 62296
rect 6810 61500 7118 61509
rect 6810 61498 6816 61500
rect 6872 61498 6896 61500
rect 6952 61498 6976 61500
rect 7032 61498 7056 61500
rect 7112 61498 7118 61500
rect 6872 61446 6874 61498
rect 7054 61446 7056 61498
rect 6810 61444 6816 61446
rect 6872 61444 6896 61446
rect 6952 61444 6976 61446
rect 7032 61444 7056 61446
rect 7112 61444 7118 61446
rect 6810 61435 7118 61444
rect 7208 61402 7236 62290
rect 7286 62248 7342 62257
rect 7286 62183 7342 62192
rect 7196 61396 7248 61402
rect 7196 61338 7248 61344
rect 7300 61198 7328 62183
rect 7288 61192 7340 61198
rect 7288 61134 7340 61140
rect 7392 61044 7420 65991
rect 7484 65754 7512 66226
rect 7567 66212 7595 66286
rect 7656 66234 7708 66240
rect 7840 66292 7892 66298
rect 7840 66234 7892 66240
rect 8024 66292 8076 66298
rect 8024 66234 8076 66240
rect 7567 66184 7604 66212
rect 7576 66178 7604 66184
rect 7576 66150 7696 66178
rect 7852 66162 7880 66234
rect 7932 66224 7984 66230
rect 7932 66166 7984 66172
rect 7564 66088 7616 66094
rect 7564 66030 7616 66036
rect 7576 65754 7604 66030
rect 7472 65748 7524 65754
rect 7472 65690 7524 65696
rect 7564 65748 7616 65754
rect 7564 65690 7616 65696
rect 7472 65612 7524 65618
rect 7472 65554 7524 65560
rect 7484 65074 7512 65554
rect 7564 65408 7616 65414
rect 7564 65350 7616 65356
rect 7472 65068 7524 65074
rect 7472 65010 7524 65016
rect 7472 64864 7524 64870
rect 7472 64806 7524 64812
rect 7484 64530 7512 64806
rect 7472 64524 7524 64530
rect 7472 64466 7524 64472
rect 7576 64410 7604 65350
rect 7668 65074 7696 66150
rect 7840 66156 7892 66162
rect 7840 66098 7892 66104
rect 7944 65754 7972 66166
rect 7932 65748 7984 65754
rect 7932 65690 7984 65696
rect 8036 65414 8064 66234
rect 8024 65408 8076 65414
rect 8024 65350 8076 65356
rect 7750 65308 8058 65317
rect 7750 65306 7756 65308
rect 7812 65306 7836 65308
rect 7892 65306 7916 65308
rect 7972 65306 7996 65308
rect 8052 65306 8058 65308
rect 7812 65254 7814 65306
rect 7994 65254 7996 65306
rect 7750 65252 7756 65254
rect 7812 65252 7836 65254
rect 7892 65252 7916 65254
rect 7972 65252 7996 65254
rect 8052 65252 8058 65254
rect 7750 65243 8058 65252
rect 7656 65068 7708 65074
rect 7656 65010 7708 65016
rect 8024 65068 8076 65074
rect 8024 65010 8076 65016
rect 7656 64932 7708 64938
rect 7656 64874 7708 64880
rect 7484 64382 7604 64410
rect 7484 62234 7512 64382
rect 7564 64320 7616 64326
rect 7564 64262 7616 64268
rect 7576 62354 7604 64262
rect 7668 63510 7696 64874
rect 8036 64462 8064 65010
rect 8024 64456 8076 64462
rect 8024 64398 8076 64404
rect 8128 64376 8156 66456
rect 8220 65074 8248 67272
rect 8404 67130 8432 67730
rect 8772 67726 8800 69498
rect 8760 67720 8812 67726
rect 8760 67662 8812 67668
rect 8576 67584 8628 67590
rect 8576 67526 8628 67532
rect 8482 67416 8538 67425
rect 8482 67351 8538 67360
rect 8496 67182 8524 67351
rect 8588 67289 8616 67526
rect 8574 67280 8630 67289
rect 8574 67215 8630 67224
rect 8760 67244 8812 67250
rect 8760 67186 8812 67192
rect 8312 67102 8432 67130
rect 8484 67176 8536 67182
rect 8484 67118 8536 67124
rect 8312 66178 8340 67102
rect 8410 66940 8718 66949
rect 8410 66938 8416 66940
rect 8472 66938 8496 66940
rect 8552 66938 8576 66940
rect 8632 66938 8656 66940
rect 8712 66938 8718 66940
rect 8472 66886 8474 66938
rect 8654 66886 8656 66938
rect 8410 66884 8416 66886
rect 8472 66884 8496 66886
rect 8552 66884 8576 66886
rect 8632 66884 8656 66886
rect 8712 66884 8718 66886
rect 8410 66875 8718 66884
rect 8484 66836 8536 66842
rect 8484 66778 8536 66784
rect 8392 66496 8444 66502
rect 8392 66438 8444 66444
rect 8404 66298 8432 66438
rect 8392 66292 8444 66298
rect 8392 66234 8444 66240
rect 8312 66150 8432 66178
rect 8300 66088 8352 66094
rect 8300 66030 8352 66036
rect 8208 65068 8260 65074
rect 8208 65010 8260 65016
rect 8312 65006 8340 66030
rect 8404 66026 8432 66150
rect 8496 66065 8524 66778
rect 8576 66700 8628 66706
rect 8628 66660 8708 66688
rect 8576 66642 8628 66648
rect 8680 66298 8708 66660
rect 8772 66502 8800 67186
rect 8760 66496 8812 66502
rect 8760 66438 8812 66444
rect 8668 66292 8720 66298
rect 8668 66234 8720 66240
rect 8482 66056 8538 66065
rect 8392 66020 8444 66026
rect 8482 65991 8538 66000
rect 8392 65962 8444 65968
rect 8410 65852 8718 65861
rect 8410 65850 8416 65852
rect 8472 65850 8496 65852
rect 8552 65850 8576 65852
rect 8632 65850 8656 65852
rect 8712 65850 8718 65852
rect 8472 65798 8474 65850
rect 8654 65798 8656 65850
rect 8410 65796 8416 65798
rect 8472 65796 8496 65798
rect 8552 65796 8576 65798
rect 8632 65796 8656 65798
rect 8712 65796 8718 65798
rect 8410 65787 8718 65796
rect 8484 65408 8536 65414
rect 8484 65350 8536 65356
rect 8496 65074 8524 65350
rect 8772 65090 8800 66438
rect 8864 66162 8892 69992
rect 8956 68474 8984 74054
rect 9048 71602 9076 74054
rect 9140 73681 9168 74122
rect 9126 73672 9182 73681
rect 9126 73607 9182 73616
rect 9128 71664 9180 71670
rect 9128 71606 9180 71612
rect 9036 71596 9088 71602
rect 9036 71538 9088 71544
rect 9036 71460 9088 71466
rect 9036 71402 9088 71408
rect 9048 70360 9076 71402
rect 9140 70938 9168 71606
rect 9232 71058 9260 74326
rect 9416 74118 9444 74734
rect 9600 74254 9628 74854
rect 9680 74656 9732 74662
rect 9680 74598 9732 74604
rect 9588 74248 9640 74254
rect 9588 74190 9640 74196
rect 9404 74112 9456 74118
rect 9404 74054 9456 74060
rect 9350 74012 9658 74021
rect 9350 74010 9356 74012
rect 9412 74010 9436 74012
rect 9492 74010 9516 74012
rect 9572 74010 9596 74012
rect 9652 74010 9658 74012
rect 9412 73958 9414 74010
rect 9594 73958 9596 74010
rect 9350 73956 9356 73958
rect 9412 73956 9436 73958
rect 9492 73956 9516 73958
rect 9572 73956 9596 73958
rect 9652 73956 9658 73958
rect 9350 73947 9658 73956
rect 9312 73568 9364 73574
rect 9312 73510 9364 73516
rect 9324 73030 9352 73510
rect 9312 73024 9364 73030
rect 9312 72966 9364 72972
rect 9350 72924 9658 72933
rect 9350 72922 9356 72924
rect 9412 72922 9436 72924
rect 9492 72922 9516 72924
rect 9572 72922 9596 72924
rect 9652 72922 9658 72924
rect 9412 72870 9414 72922
rect 9594 72870 9596 72922
rect 9350 72868 9356 72870
rect 9412 72868 9436 72870
rect 9492 72868 9516 72870
rect 9572 72868 9596 72870
rect 9652 72868 9658 72870
rect 9350 72859 9658 72868
rect 9404 72616 9456 72622
rect 9402 72584 9404 72593
rect 9456 72584 9458 72593
rect 9402 72519 9458 72528
rect 9404 72480 9456 72486
rect 9404 72422 9456 72428
rect 9416 72049 9444 72422
rect 9402 72040 9458 72049
rect 9402 71975 9458 71984
rect 9350 71836 9658 71845
rect 9350 71834 9356 71836
rect 9412 71834 9436 71836
rect 9492 71834 9516 71836
rect 9572 71834 9596 71836
rect 9652 71834 9658 71836
rect 9412 71782 9414 71834
rect 9594 71782 9596 71834
rect 9350 71780 9356 71782
rect 9412 71780 9436 71782
rect 9492 71780 9516 71782
rect 9572 71780 9596 71782
rect 9652 71780 9658 71782
rect 9350 71771 9658 71780
rect 9220 71052 9272 71058
rect 9272 71012 9352 71040
rect 9220 70994 9272 71000
rect 9218 70952 9274 70961
rect 9140 70910 9218 70938
rect 9218 70887 9274 70896
rect 9128 70848 9180 70854
rect 9324 70836 9352 71012
rect 9128 70790 9180 70796
rect 9232 70808 9352 70836
rect 9140 70650 9168 70790
rect 9128 70644 9180 70650
rect 9128 70586 9180 70592
rect 9232 70514 9260 70808
rect 9350 70748 9658 70757
rect 9350 70746 9356 70748
rect 9412 70746 9436 70748
rect 9492 70746 9516 70748
rect 9572 70746 9596 70748
rect 9652 70746 9658 70748
rect 9412 70694 9414 70746
rect 9594 70694 9596 70746
rect 9350 70692 9356 70694
rect 9412 70692 9436 70694
rect 9492 70692 9516 70694
rect 9572 70692 9596 70694
rect 9652 70692 9658 70694
rect 9350 70683 9658 70692
rect 9404 70576 9456 70582
rect 9324 70536 9404 70564
rect 9220 70508 9272 70514
rect 9220 70450 9272 70456
rect 9048 70332 9260 70360
rect 9126 70272 9182 70281
rect 9126 70207 9182 70216
rect 9036 70100 9088 70106
rect 9036 70042 9088 70048
rect 9048 69306 9076 70042
rect 9140 69426 9168 70207
rect 9232 69970 9260 70332
rect 9324 70145 9352 70536
rect 9404 70518 9456 70524
rect 9588 70372 9640 70378
rect 9588 70314 9640 70320
rect 9310 70136 9366 70145
rect 9600 70106 9628 70314
rect 9310 70071 9312 70080
rect 9364 70071 9366 70080
rect 9588 70100 9640 70106
rect 9312 70042 9364 70048
rect 9588 70042 9640 70048
rect 9586 70000 9642 70009
rect 9220 69964 9272 69970
rect 9692 69970 9720 74598
rect 9954 74352 10010 74361
rect 9954 74287 10010 74296
rect 9772 74112 9824 74118
rect 9772 74054 9824 74060
rect 9784 72214 9812 74054
rect 9968 73642 9996 74287
rect 9956 73636 10008 73642
rect 9956 73578 10008 73584
rect 9772 72208 9824 72214
rect 9772 72150 9824 72156
rect 9772 71120 9824 71126
rect 9772 71062 9824 71068
rect 9586 69935 9642 69944
rect 9680 69964 9732 69970
rect 9220 69906 9272 69912
rect 9600 69766 9628 69935
rect 9680 69906 9732 69912
rect 9680 69828 9732 69834
rect 9680 69770 9732 69776
rect 9220 69760 9272 69766
rect 9220 69702 9272 69708
rect 9588 69760 9640 69766
rect 9588 69702 9640 69708
rect 9232 69544 9260 69702
rect 9350 69660 9658 69669
rect 9350 69658 9356 69660
rect 9412 69658 9436 69660
rect 9492 69658 9516 69660
rect 9572 69658 9596 69660
rect 9652 69658 9658 69660
rect 9412 69606 9414 69658
rect 9594 69606 9596 69658
rect 9350 69604 9356 69606
rect 9412 69604 9436 69606
rect 9492 69604 9516 69606
rect 9572 69604 9596 69606
rect 9652 69604 9658 69606
rect 9350 69595 9658 69604
rect 9232 69516 9444 69544
rect 9416 69426 9444 69516
rect 9128 69420 9180 69426
rect 9128 69362 9180 69368
rect 9312 69420 9364 69426
rect 9312 69362 9364 69368
rect 9404 69420 9456 69426
rect 9404 69362 9456 69368
rect 9048 69278 9260 69306
rect 9036 69216 9088 69222
rect 9036 69158 9088 69164
rect 9048 68882 9076 69158
rect 9036 68876 9088 68882
rect 9036 68818 9088 68824
rect 8944 68468 8996 68474
rect 8944 68410 8996 68416
rect 8944 68332 8996 68338
rect 8944 68274 8996 68280
rect 8956 66638 8984 68274
rect 9048 67930 9076 68818
rect 9128 68672 9180 68678
rect 9128 68614 9180 68620
rect 9140 68377 9168 68614
rect 9126 68368 9182 68377
rect 9126 68303 9182 68312
rect 9128 68264 9180 68270
rect 9128 68206 9180 68212
rect 9036 67924 9088 67930
rect 9036 67866 9088 67872
rect 9048 67182 9076 67866
rect 9140 67386 9168 68206
rect 9232 67794 9260 69278
rect 9324 68746 9352 69362
rect 9416 69018 9444 69362
rect 9404 69012 9456 69018
rect 9404 68954 9456 68960
rect 9312 68740 9364 68746
rect 9312 68682 9364 68688
rect 9350 68572 9658 68581
rect 9350 68570 9356 68572
rect 9412 68570 9436 68572
rect 9492 68570 9516 68572
rect 9572 68570 9596 68572
rect 9652 68570 9658 68572
rect 9412 68518 9414 68570
rect 9594 68518 9596 68570
rect 9350 68516 9356 68518
rect 9412 68516 9436 68518
rect 9492 68516 9516 68518
rect 9572 68516 9596 68518
rect 9652 68516 9658 68518
rect 9350 68507 9658 68516
rect 9220 67788 9272 67794
rect 9220 67730 9272 67736
rect 9310 67688 9366 67697
rect 9310 67623 9366 67632
rect 9324 67572 9352 67623
rect 9232 67544 9352 67572
rect 9128 67380 9180 67386
rect 9232 67368 9260 67544
rect 9350 67484 9658 67493
rect 9350 67482 9356 67484
rect 9412 67482 9436 67484
rect 9492 67482 9516 67484
rect 9572 67482 9596 67484
rect 9652 67482 9658 67484
rect 9412 67430 9414 67482
rect 9594 67430 9596 67482
rect 9350 67428 9356 67430
rect 9412 67428 9436 67430
rect 9492 67428 9516 67430
rect 9572 67428 9596 67430
rect 9652 67428 9658 67430
rect 9350 67419 9658 67428
rect 9232 67340 9628 67368
rect 9128 67322 9180 67328
rect 9310 67280 9366 67289
rect 9310 67215 9366 67224
rect 9036 67176 9088 67182
rect 9128 67176 9180 67182
rect 9036 67118 9088 67124
rect 9126 67144 9128 67153
rect 9180 67144 9182 67153
rect 9048 66706 9076 67118
rect 9126 67079 9182 67088
rect 9220 66836 9272 66842
rect 9220 66778 9272 66784
rect 9036 66700 9088 66706
rect 9036 66642 9088 66648
rect 8944 66632 8996 66638
rect 8944 66574 8996 66580
rect 8944 66496 8996 66502
rect 8944 66438 8996 66444
rect 8852 66156 8904 66162
rect 8852 66098 8904 66104
rect 8852 66020 8904 66026
rect 8852 65962 8904 65968
rect 8484 65068 8536 65074
rect 8484 65010 8536 65016
rect 8588 65062 8800 65090
rect 8300 65000 8352 65006
rect 8300 64942 8352 64948
rect 8588 64852 8616 65062
rect 8760 65000 8812 65006
rect 8760 64942 8812 64948
rect 8312 64824 8616 64852
rect 8128 64348 8248 64376
rect 8024 64320 8076 64326
rect 8076 64280 8156 64308
rect 8024 64262 8076 64268
rect 7750 64220 8058 64229
rect 7750 64218 7756 64220
rect 7812 64218 7836 64220
rect 7892 64218 7916 64220
rect 7972 64218 7996 64220
rect 8052 64218 8058 64220
rect 7812 64166 7814 64218
rect 7994 64166 7996 64218
rect 7750 64164 7756 64166
rect 7812 64164 7836 64166
rect 7892 64164 7916 64166
rect 7972 64164 7996 64166
rect 8052 64164 8058 64166
rect 7750 64155 8058 64164
rect 8128 64104 8156 64280
rect 7852 64076 8156 64104
rect 7748 63980 7800 63986
rect 7748 63922 7800 63928
rect 7656 63504 7708 63510
rect 7656 63446 7708 63452
rect 7760 63356 7788 63922
rect 7668 63328 7788 63356
rect 7668 62898 7696 63328
rect 7852 63220 7880 64076
rect 7932 63980 7984 63986
rect 7932 63922 7984 63928
rect 7944 63374 7972 63922
rect 8116 63776 8168 63782
rect 8116 63718 8168 63724
rect 7932 63368 7984 63374
rect 7932 63310 7984 63316
rect 8128 63288 8156 63718
rect 8220 63481 8248 64348
rect 8312 63986 8340 64824
rect 8410 64764 8718 64773
rect 8410 64762 8416 64764
rect 8472 64762 8496 64764
rect 8552 64762 8576 64764
rect 8632 64762 8656 64764
rect 8712 64762 8718 64764
rect 8472 64710 8474 64762
rect 8654 64710 8656 64762
rect 8410 64708 8416 64710
rect 8472 64708 8496 64710
rect 8552 64708 8576 64710
rect 8632 64708 8656 64710
rect 8712 64708 8718 64710
rect 8410 64699 8718 64708
rect 8576 64524 8628 64530
rect 8576 64466 8628 64472
rect 8668 64524 8720 64530
rect 8668 64466 8720 64472
rect 8300 63980 8352 63986
rect 8300 63922 8352 63928
rect 8588 63918 8616 64466
rect 8680 63918 8708 64466
rect 8576 63912 8628 63918
rect 8576 63854 8628 63860
rect 8668 63912 8720 63918
rect 8668 63854 8720 63860
rect 8300 63844 8352 63850
rect 8300 63786 8352 63792
rect 8206 63472 8262 63481
rect 8206 63407 8262 63416
rect 8128 63260 8248 63288
rect 7852 63192 8156 63220
rect 7750 63132 8058 63141
rect 7750 63130 7756 63132
rect 7812 63130 7836 63132
rect 7892 63130 7916 63132
rect 7972 63130 7996 63132
rect 8052 63130 8058 63132
rect 7812 63078 7814 63130
rect 7994 63078 7996 63130
rect 7750 63076 7756 63078
rect 7812 63076 7836 63078
rect 7892 63076 7916 63078
rect 7972 63076 7996 63078
rect 8052 63076 8058 63078
rect 7750 63067 8058 63076
rect 7656 62892 7708 62898
rect 7656 62834 7708 62840
rect 7840 62824 7892 62830
rect 7840 62766 7892 62772
rect 7656 62688 7708 62694
rect 7656 62630 7708 62636
rect 7564 62348 7616 62354
rect 7564 62290 7616 62296
rect 7484 62206 7604 62234
rect 7472 61396 7524 61402
rect 7472 61338 7524 61344
rect 7208 61016 7420 61044
rect 6810 60412 7118 60421
rect 6810 60410 6816 60412
rect 6872 60410 6896 60412
rect 6952 60410 6976 60412
rect 7032 60410 7056 60412
rect 7112 60410 7118 60412
rect 6872 60358 6874 60410
rect 7054 60358 7056 60410
rect 6810 60356 6816 60358
rect 6872 60356 6896 60358
rect 6952 60356 6976 60358
rect 7032 60356 7056 60358
rect 7112 60356 7118 60358
rect 6810 60347 7118 60356
rect 6810 59324 7118 59333
rect 6810 59322 6816 59324
rect 6872 59322 6896 59324
rect 6952 59322 6976 59324
rect 7032 59322 7056 59324
rect 7112 59322 7118 59324
rect 6872 59270 6874 59322
rect 7054 59270 7056 59322
rect 6810 59268 6816 59270
rect 6872 59268 6896 59270
rect 6952 59268 6976 59270
rect 7032 59268 7056 59270
rect 7112 59268 7118 59270
rect 6810 59259 7118 59268
rect 6828 59084 6880 59090
rect 6880 59044 6960 59072
rect 6828 59026 6880 59032
rect 6828 58948 6880 58954
rect 6828 58890 6880 58896
rect 6840 58546 6868 58890
rect 6932 58682 6960 59044
rect 6920 58676 6972 58682
rect 6920 58618 6972 58624
rect 7208 58546 7236 61016
rect 7288 60716 7340 60722
rect 7288 60658 7340 60664
rect 7300 60178 7328 60658
rect 7288 60172 7340 60178
rect 7340 60132 7420 60160
rect 7288 60114 7340 60120
rect 7392 59770 7420 60132
rect 7380 59764 7432 59770
rect 7380 59706 7432 59712
rect 7288 59560 7340 59566
rect 7288 59502 7340 59508
rect 6828 58540 6880 58546
rect 6828 58482 6880 58488
rect 7196 58540 7248 58546
rect 7196 58482 7248 58488
rect 7196 58404 7248 58410
rect 7196 58346 7248 58352
rect 6810 58236 7118 58245
rect 6810 58234 6816 58236
rect 6872 58234 6896 58236
rect 6952 58234 6976 58236
rect 7032 58234 7056 58236
rect 7112 58234 7118 58236
rect 6872 58182 6874 58234
rect 7054 58182 7056 58234
rect 6810 58180 6816 58182
rect 6872 58180 6896 58182
rect 6952 58180 6976 58182
rect 7032 58180 7056 58182
rect 7112 58180 7118 58182
rect 6810 58171 7118 58180
rect 7208 58138 7236 58346
rect 7300 58138 7328 59502
rect 7392 59226 7420 59706
rect 7380 59220 7432 59226
rect 7380 59162 7432 59168
rect 7380 58880 7432 58886
rect 7380 58822 7432 58828
rect 7196 58132 7248 58138
rect 7196 58074 7248 58080
rect 7288 58132 7340 58138
rect 7288 58074 7340 58080
rect 7392 58018 7420 58822
rect 7484 58478 7512 61338
rect 7472 58472 7524 58478
rect 7472 58414 7524 58420
rect 7472 58336 7524 58342
rect 7472 58278 7524 58284
rect 7116 57990 7420 58018
rect 7116 57526 7144 57990
rect 7196 57792 7248 57798
rect 7196 57734 7248 57740
rect 7288 57792 7340 57798
rect 7288 57734 7340 57740
rect 7104 57520 7156 57526
rect 7104 57462 7156 57468
rect 7208 57458 7236 57734
rect 7196 57452 7248 57458
rect 7196 57394 7248 57400
rect 6810 57148 7118 57157
rect 6810 57146 6816 57148
rect 6872 57146 6896 57148
rect 6952 57146 6976 57148
rect 7032 57146 7056 57148
rect 7112 57146 7118 57148
rect 6872 57094 6874 57146
rect 7054 57094 7056 57146
rect 6810 57092 6816 57094
rect 6872 57092 6896 57094
rect 6952 57092 6976 57094
rect 7032 57092 7056 57094
rect 7112 57092 7118 57094
rect 6810 57083 7118 57092
rect 6828 56908 6880 56914
rect 6828 56850 6880 56856
rect 6736 56840 6788 56846
rect 6736 56782 6788 56788
rect 6644 56772 6696 56778
rect 6644 56714 6696 56720
rect 6736 56704 6788 56710
rect 6736 56646 6788 56652
rect 6644 56296 6696 56302
rect 6644 56238 6696 56244
rect 6656 54670 6684 56238
rect 6644 54664 6696 54670
rect 6644 54606 6696 54612
rect 6644 54188 6696 54194
rect 6644 54130 6696 54136
rect 6656 53106 6684 54130
rect 6644 53100 6696 53106
rect 6644 53042 6696 53048
rect 6644 52692 6696 52698
rect 6644 52634 6696 52640
rect 6472 52108 6592 52136
rect 6472 52018 6500 52108
rect 6460 52012 6512 52018
rect 6460 51954 6512 51960
rect 6552 51944 6604 51950
rect 6552 51886 6604 51892
rect 6368 51808 6420 51814
rect 6368 51750 6420 51756
rect 6380 51406 6408 51750
rect 6368 51400 6420 51406
rect 6090 51368 6146 51377
rect 5920 46714 5948 51342
rect 6012 51326 6090 51354
rect 6368 51342 6420 51348
rect 6090 51303 6146 51312
rect 6150 51164 6458 51173
rect 6150 51162 6156 51164
rect 6212 51162 6236 51164
rect 6292 51162 6316 51164
rect 6372 51162 6396 51164
rect 6452 51162 6458 51164
rect 6212 51110 6214 51162
rect 6394 51110 6396 51162
rect 6150 51108 6156 51110
rect 6212 51108 6236 51110
rect 6292 51108 6316 51110
rect 6372 51108 6396 51110
rect 6452 51108 6458 51110
rect 6150 51099 6458 51108
rect 6000 50992 6052 50998
rect 6000 50934 6052 50940
rect 6090 50960 6146 50969
rect 5908 46708 5960 46714
rect 5908 46650 5960 46656
rect 6012 46510 6040 50934
rect 6090 50895 6146 50904
rect 6104 50182 6132 50895
rect 6092 50176 6144 50182
rect 6092 50118 6144 50124
rect 6150 50076 6458 50085
rect 6150 50074 6156 50076
rect 6212 50074 6236 50076
rect 6292 50074 6316 50076
rect 6372 50074 6396 50076
rect 6452 50074 6458 50076
rect 6212 50022 6214 50074
rect 6394 50022 6396 50074
rect 6150 50020 6156 50022
rect 6212 50020 6236 50022
rect 6292 50020 6316 50022
rect 6372 50020 6396 50022
rect 6452 50020 6458 50022
rect 6150 50011 6458 50020
rect 6150 48988 6458 48997
rect 6150 48986 6156 48988
rect 6212 48986 6236 48988
rect 6292 48986 6316 48988
rect 6372 48986 6396 48988
rect 6452 48986 6458 48988
rect 6212 48934 6214 48986
rect 6394 48934 6396 48986
rect 6150 48932 6156 48934
rect 6212 48932 6236 48934
rect 6292 48932 6316 48934
rect 6372 48932 6396 48934
rect 6452 48932 6458 48934
rect 6150 48923 6458 48932
rect 6092 48748 6144 48754
rect 6092 48690 6144 48696
rect 6104 48006 6132 48690
rect 6092 48000 6144 48006
rect 6092 47942 6144 47948
rect 6150 47900 6458 47909
rect 6150 47898 6156 47900
rect 6212 47898 6236 47900
rect 6292 47898 6316 47900
rect 6372 47898 6396 47900
rect 6452 47898 6458 47900
rect 6212 47846 6214 47898
rect 6394 47846 6396 47898
rect 6150 47844 6156 47846
rect 6212 47844 6236 47846
rect 6292 47844 6316 47846
rect 6372 47844 6396 47846
rect 6452 47844 6458 47846
rect 6150 47835 6458 47844
rect 6460 47660 6512 47666
rect 6460 47602 6512 47608
rect 6472 46986 6500 47602
rect 6460 46980 6512 46986
rect 6460 46922 6512 46928
rect 6150 46812 6458 46821
rect 6150 46810 6156 46812
rect 6212 46810 6236 46812
rect 6292 46810 6316 46812
rect 6372 46810 6396 46812
rect 6452 46810 6458 46812
rect 6212 46758 6214 46810
rect 6394 46758 6396 46810
rect 6150 46756 6156 46758
rect 6212 46756 6236 46758
rect 6292 46756 6316 46758
rect 6372 46756 6396 46758
rect 6452 46756 6458 46758
rect 6150 46747 6458 46756
rect 6460 46640 6512 46646
rect 6460 46582 6512 46588
rect 6000 46504 6052 46510
rect 6000 46446 6052 46452
rect 6368 46504 6420 46510
rect 6368 46446 6420 46452
rect 6092 46436 6144 46442
rect 6092 46378 6144 46384
rect 5908 46368 5960 46374
rect 5908 46310 5960 46316
rect 5920 44878 5948 46310
rect 5998 45928 6054 45937
rect 6104 45914 6132 46378
rect 6276 46368 6328 46374
rect 6276 46310 6328 46316
rect 6054 45886 6132 45914
rect 5998 45863 6054 45872
rect 6288 45812 6316 46310
rect 6380 46034 6408 46446
rect 6368 46028 6420 46034
rect 6368 45970 6420 45976
rect 6472 45966 6500 46582
rect 6460 45960 6512 45966
rect 6460 45902 6512 45908
rect 6012 45784 6316 45812
rect 5908 44872 5960 44878
rect 5908 44814 5960 44820
rect 5908 44736 5960 44742
rect 5908 44678 5960 44684
rect 5920 42906 5948 44678
rect 5908 42900 5960 42906
rect 5908 42842 5960 42848
rect 5736 41386 5856 41414
rect 5632 40724 5684 40730
rect 5632 40666 5684 40672
rect 5632 40384 5684 40390
rect 5632 40326 5684 40332
rect 5540 39636 5592 39642
rect 5540 39578 5592 39584
rect 5448 39568 5500 39574
rect 5448 39510 5500 39516
rect 5460 38842 5488 39510
rect 5540 39432 5592 39438
rect 5540 39374 5592 39380
rect 5552 38962 5580 39374
rect 5540 38956 5592 38962
rect 5540 38898 5592 38904
rect 5460 38814 5580 38842
rect 5210 38652 5518 38661
rect 5210 38650 5216 38652
rect 5272 38650 5296 38652
rect 5352 38650 5376 38652
rect 5432 38650 5456 38652
rect 5512 38650 5518 38652
rect 5272 38598 5274 38650
rect 5454 38598 5456 38650
rect 5210 38596 5216 38598
rect 5272 38596 5296 38598
rect 5352 38596 5376 38598
rect 5432 38596 5456 38598
rect 5512 38596 5518 38598
rect 5210 38587 5518 38596
rect 5552 38434 5580 38814
rect 5460 38406 5580 38434
rect 5460 37652 5488 38406
rect 5460 37624 5580 37652
rect 5210 37564 5518 37573
rect 5210 37562 5216 37564
rect 5272 37562 5296 37564
rect 5352 37562 5376 37564
rect 5432 37562 5456 37564
rect 5512 37562 5518 37564
rect 5272 37510 5274 37562
rect 5454 37510 5456 37562
rect 5210 37508 5216 37510
rect 5272 37508 5296 37510
rect 5352 37508 5376 37510
rect 5432 37508 5456 37510
rect 5512 37508 5518 37510
rect 5210 37499 5518 37508
rect 5552 37346 5580 37624
rect 5460 37318 5580 37346
rect 5460 36650 5488 37318
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 5448 36644 5500 36650
rect 5448 36586 5500 36592
rect 5210 36476 5518 36485
rect 5210 36474 5216 36476
rect 5272 36474 5296 36476
rect 5352 36474 5376 36476
rect 5432 36474 5456 36476
rect 5512 36474 5518 36476
rect 5272 36422 5274 36474
rect 5454 36422 5456 36474
rect 5210 36420 5216 36422
rect 5272 36420 5296 36422
rect 5352 36420 5376 36422
rect 5432 36420 5456 36422
rect 5512 36420 5518 36422
rect 5210 36411 5518 36420
rect 5210 35388 5518 35397
rect 5210 35386 5216 35388
rect 5272 35386 5296 35388
rect 5352 35386 5376 35388
rect 5432 35386 5456 35388
rect 5512 35386 5518 35388
rect 5272 35334 5274 35386
rect 5454 35334 5456 35386
rect 5210 35332 5216 35334
rect 5272 35332 5296 35334
rect 5352 35332 5376 35334
rect 5432 35332 5456 35334
rect 5512 35332 5518 35334
rect 5210 35323 5518 35332
rect 5210 34300 5518 34309
rect 5210 34298 5216 34300
rect 5272 34298 5296 34300
rect 5352 34298 5376 34300
rect 5432 34298 5456 34300
rect 5512 34298 5518 34300
rect 5272 34246 5274 34298
rect 5454 34246 5456 34298
rect 5210 34244 5216 34246
rect 5272 34244 5296 34246
rect 5352 34244 5376 34246
rect 5432 34244 5456 34246
rect 5512 34244 5518 34246
rect 5210 34235 5518 34244
rect 5210 33212 5518 33221
rect 5210 33210 5216 33212
rect 5272 33210 5296 33212
rect 5352 33210 5376 33212
rect 5432 33210 5456 33212
rect 5512 33210 5518 33212
rect 5272 33158 5274 33210
rect 5454 33158 5456 33210
rect 5210 33156 5216 33158
rect 5272 33156 5296 33158
rect 5352 33156 5376 33158
rect 5432 33156 5456 33158
rect 5512 33156 5518 33158
rect 5210 33147 5518 33156
rect 5210 32124 5518 32133
rect 5210 32122 5216 32124
rect 5272 32122 5296 32124
rect 5352 32122 5376 32124
rect 5432 32122 5456 32124
rect 5512 32122 5518 32124
rect 5272 32070 5274 32122
rect 5454 32070 5456 32122
rect 5210 32068 5216 32070
rect 5272 32068 5296 32070
rect 5352 32068 5376 32070
rect 5432 32068 5456 32070
rect 5512 32068 5518 32070
rect 5210 32059 5518 32068
rect 5448 31952 5500 31958
rect 5448 31894 5500 31900
rect 5460 31346 5488 31894
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5210 31036 5518 31045
rect 5210 31034 5216 31036
rect 5272 31034 5296 31036
rect 5352 31034 5376 31036
rect 5432 31034 5456 31036
rect 5512 31034 5518 31036
rect 5272 30982 5274 31034
rect 5454 30982 5456 31034
rect 5210 30980 5216 30982
rect 5272 30980 5296 30982
rect 5352 30980 5376 30982
rect 5432 30980 5456 30982
rect 5512 30980 5518 30982
rect 5210 30971 5518 30980
rect 5210 29948 5518 29957
rect 5210 29946 5216 29948
rect 5272 29946 5296 29948
rect 5352 29946 5376 29948
rect 5432 29946 5456 29948
rect 5512 29946 5518 29948
rect 5272 29894 5274 29946
rect 5454 29894 5456 29946
rect 5210 29892 5216 29894
rect 5272 29892 5296 29894
rect 5352 29892 5376 29894
rect 5432 29892 5456 29894
rect 5512 29892 5518 29894
rect 5210 29883 5518 29892
rect 5552 29594 5580 37198
rect 5644 29714 5672 40326
rect 5736 29714 5764 41386
rect 6012 40458 6040 45784
rect 6150 45724 6458 45733
rect 6150 45722 6156 45724
rect 6212 45722 6236 45724
rect 6292 45722 6316 45724
rect 6372 45722 6396 45724
rect 6452 45722 6458 45724
rect 6212 45670 6214 45722
rect 6394 45670 6396 45722
rect 6150 45668 6156 45670
rect 6212 45668 6236 45670
rect 6292 45668 6316 45670
rect 6372 45668 6396 45670
rect 6452 45668 6458 45670
rect 6150 45659 6458 45668
rect 6090 45520 6146 45529
rect 6090 45455 6146 45464
rect 6104 44742 6132 45455
rect 6092 44736 6144 44742
rect 6092 44678 6144 44684
rect 6150 44636 6458 44645
rect 6150 44634 6156 44636
rect 6212 44634 6236 44636
rect 6292 44634 6316 44636
rect 6372 44634 6396 44636
rect 6452 44634 6458 44636
rect 6212 44582 6214 44634
rect 6394 44582 6396 44634
rect 6150 44580 6156 44582
rect 6212 44580 6236 44582
rect 6292 44580 6316 44582
rect 6372 44580 6396 44582
rect 6452 44580 6458 44582
rect 6150 44571 6458 44580
rect 6150 43548 6458 43557
rect 6150 43546 6156 43548
rect 6212 43546 6236 43548
rect 6292 43546 6316 43548
rect 6372 43546 6396 43548
rect 6452 43546 6458 43548
rect 6212 43494 6214 43546
rect 6394 43494 6396 43546
rect 6150 43492 6156 43494
rect 6212 43492 6236 43494
rect 6292 43492 6316 43494
rect 6372 43492 6396 43494
rect 6452 43492 6458 43494
rect 6150 43483 6458 43492
rect 6150 42460 6458 42469
rect 6150 42458 6156 42460
rect 6212 42458 6236 42460
rect 6292 42458 6316 42460
rect 6372 42458 6396 42460
rect 6452 42458 6458 42460
rect 6212 42406 6214 42458
rect 6394 42406 6396 42458
rect 6150 42404 6156 42406
rect 6212 42404 6236 42406
rect 6292 42404 6316 42406
rect 6372 42404 6396 42406
rect 6452 42404 6458 42406
rect 6150 42395 6458 42404
rect 6150 41372 6458 41381
rect 6150 41370 6156 41372
rect 6212 41370 6236 41372
rect 6292 41370 6316 41372
rect 6372 41370 6396 41372
rect 6452 41370 6458 41372
rect 6212 41318 6214 41370
rect 6394 41318 6396 41370
rect 6150 41316 6156 41318
rect 6212 41316 6236 41318
rect 6292 41316 6316 41318
rect 6372 41316 6396 41318
rect 6452 41316 6458 41318
rect 6150 41307 6458 41316
rect 5908 40452 5960 40458
rect 5908 40394 5960 40400
rect 6000 40452 6052 40458
rect 6000 40394 6052 40400
rect 5816 40180 5868 40186
rect 5816 40122 5868 40128
rect 5632 29708 5684 29714
rect 5632 29650 5684 29656
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5172 29572 5224 29578
rect 5552 29566 5764 29594
rect 5172 29514 5224 29520
rect 5184 28966 5212 29514
rect 5540 29504 5592 29510
rect 5540 29446 5592 29452
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 5210 28860 5518 28869
rect 5210 28858 5216 28860
rect 5272 28858 5296 28860
rect 5352 28858 5376 28860
rect 5432 28858 5456 28860
rect 5512 28858 5518 28860
rect 5272 28806 5274 28858
rect 5454 28806 5456 28858
rect 5210 28804 5216 28806
rect 5272 28804 5296 28806
rect 5352 28804 5376 28806
rect 5432 28804 5456 28806
rect 5512 28804 5518 28806
rect 5210 28795 5518 28804
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 27985 5488 28358
rect 5446 27976 5502 27985
rect 5446 27911 5502 27920
rect 5210 27772 5518 27781
rect 5210 27770 5216 27772
rect 5272 27770 5296 27772
rect 5352 27770 5376 27772
rect 5432 27770 5456 27772
rect 5512 27770 5518 27772
rect 5272 27718 5274 27770
rect 5454 27718 5456 27770
rect 5210 27716 5216 27718
rect 5272 27716 5296 27718
rect 5352 27716 5376 27718
rect 5432 27716 5456 27718
rect 5512 27716 5518 27718
rect 5210 27707 5518 27716
rect 5446 27568 5502 27577
rect 5446 27503 5502 27512
rect 5460 27010 5488 27503
rect 5552 27130 5580 29446
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5460 26982 5580 27010
rect 5210 26684 5518 26693
rect 5210 26682 5216 26684
rect 5272 26682 5296 26684
rect 5352 26682 5376 26684
rect 5432 26682 5456 26684
rect 5512 26682 5518 26684
rect 5272 26630 5274 26682
rect 5454 26630 5456 26682
rect 5210 26628 5216 26630
rect 5272 26628 5296 26630
rect 5352 26628 5376 26630
rect 5432 26628 5456 26630
rect 5512 26628 5518 26630
rect 5210 26619 5518 26628
rect 5552 26568 5580 26982
rect 5460 26540 5580 26568
rect 5356 26512 5408 26518
rect 5356 26454 5408 26460
rect 5092 26268 5304 26296
rect 5276 26058 5304 26268
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 5092 26030 5304 26058
rect 5368 26042 5396 26454
rect 5356 26036 5408 26042
rect 5000 25242 5028 25978
rect 5092 25378 5120 26030
rect 5356 25978 5408 25984
rect 5460 25786 5488 26540
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5552 25906 5580 26318
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5460 25758 5580 25786
rect 5210 25596 5518 25605
rect 5210 25594 5216 25596
rect 5272 25594 5296 25596
rect 5352 25594 5376 25596
rect 5432 25594 5456 25596
rect 5512 25594 5518 25596
rect 5272 25542 5274 25594
rect 5454 25542 5456 25594
rect 5210 25540 5216 25542
rect 5272 25540 5296 25542
rect 5352 25540 5376 25542
rect 5432 25540 5456 25542
rect 5512 25540 5518 25542
rect 5210 25531 5518 25540
rect 5092 25350 5212 25378
rect 5000 25214 5120 25242
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 5000 24070 5028 25094
rect 4988 24064 5040 24070
rect 4988 24006 5040 24012
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4550 18524 4858 18533
rect 4550 18522 4556 18524
rect 4612 18522 4636 18524
rect 4692 18522 4716 18524
rect 4772 18522 4796 18524
rect 4852 18522 4858 18524
rect 4612 18470 4614 18522
rect 4794 18470 4796 18522
rect 4550 18468 4556 18470
rect 4612 18468 4636 18470
rect 4692 18468 4716 18470
rect 4772 18468 4796 18470
rect 4852 18468 4858 18470
rect 4550 18459 4858 18468
rect 4550 17436 4858 17445
rect 4550 17434 4556 17436
rect 4612 17434 4636 17436
rect 4692 17434 4716 17436
rect 4772 17434 4796 17436
rect 4852 17434 4858 17436
rect 4612 17382 4614 17434
rect 4794 17382 4796 17434
rect 4550 17380 4556 17382
rect 4612 17380 4636 17382
rect 4692 17380 4716 17382
rect 4772 17380 4796 17382
rect 4852 17380 4858 17382
rect 4550 17371 4858 17380
rect 4550 16348 4858 16357
rect 4550 16346 4556 16348
rect 4612 16346 4636 16348
rect 4692 16346 4716 16348
rect 4772 16346 4796 16348
rect 4852 16346 4858 16348
rect 4612 16294 4614 16346
rect 4794 16294 4796 16346
rect 4550 16292 4556 16294
rect 4612 16292 4636 16294
rect 4692 16292 4716 16294
rect 4772 16292 4796 16294
rect 4852 16292 4858 16294
rect 4550 16283 4858 16292
rect 4550 15260 4858 15269
rect 4550 15258 4556 15260
rect 4612 15258 4636 15260
rect 4692 15258 4716 15260
rect 4772 15258 4796 15260
rect 4852 15258 4858 15260
rect 4612 15206 4614 15258
rect 4794 15206 4796 15258
rect 4550 15204 4556 15206
rect 4612 15204 4636 15206
rect 4692 15204 4716 15206
rect 4772 15204 4796 15206
rect 4852 15204 4858 15206
rect 4550 15195 4858 15204
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4550 14172 4858 14181
rect 4550 14170 4556 14172
rect 4612 14170 4636 14172
rect 4692 14170 4716 14172
rect 4772 14170 4796 14172
rect 4852 14170 4858 14172
rect 4612 14118 4614 14170
rect 4794 14118 4796 14170
rect 4550 14116 4556 14118
rect 4612 14116 4636 14118
rect 4692 14116 4716 14118
rect 4772 14116 4796 14118
rect 4852 14116 4858 14118
rect 4550 14107 4858 14116
rect 4550 13084 4858 13093
rect 4550 13082 4556 13084
rect 4612 13082 4636 13084
rect 4692 13082 4716 13084
rect 4772 13082 4796 13084
rect 4852 13082 4858 13084
rect 4612 13030 4614 13082
rect 4794 13030 4796 13082
rect 4550 13028 4556 13030
rect 4612 13028 4636 13030
rect 4692 13028 4716 13030
rect 4772 13028 4796 13030
rect 4852 13028 4858 13030
rect 4550 13019 4858 13028
rect 4550 11996 4858 12005
rect 4550 11994 4556 11996
rect 4612 11994 4636 11996
rect 4692 11994 4716 11996
rect 4772 11994 4796 11996
rect 4852 11994 4858 11996
rect 4612 11942 4614 11994
rect 4794 11942 4796 11994
rect 4550 11940 4556 11942
rect 4612 11940 4636 11942
rect 4692 11940 4716 11942
rect 4772 11940 4796 11942
rect 4852 11940 4858 11942
rect 4550 11931 4858 11940
rect 4550 10908 4858 10917
rect 4550 10906 4556 10908
rect 4612 10906 4636 10908
rect 4692 10906 4716 10908
rect 4772 10906 4796 10908
rect 4852 10906 4858 10908
rect 4612 10854 4614 10906
rect 4794 10854 4796 10906
rect 4550 10852 4556 10854
rect 4612 10852 4636 10854
rect 4692 10852 4716 10854
rect 4772 10852 4796 10854
rect 4852 10852 4858 10854
rect 4550 10843 4858 10852
rect 4550 9820 4858 9829
rect 4550 9818 4556 9820
rect 4612 9818 4636 9820
rect 4692 9818 4716 9820
rect 4772 9818 4796 9820
rect 4852 9818 4858 9820
rect 4612 9766 4614 9818
rect 4794 9766 4796 9818
rect 4550 9764 4556 9766
rect 4612 9764 4636 9766
rect 4692 9764 4716 9766
rect 4772 9764 4796 9766
rect 4852 9764 4858 9766
rect 4550 9755 4858 9764
rect 4550 8732 4858 8741
rect 4550 8730 4556 8732
rect 4612 8730 4636 8732
rect 4692 8730 4716 8732
rect 4772 8730 4796 8732
rect 4852 8730 4858 8732
rect 4612 8678 4614 8730
rect 4794 8678 4796 8730
rect 4550 8676 4556 8678
rect 4612 8676 4636 8678
rect 4692 8676 4716 8678
rect 4772 8676 4796 8678
rect 4852 8676 4858 8678
rect 4550 8667 4858 8676
rect 4550 7644 4858 7653
rect 4550 7642 4556 7644
rect 4612 7642 4636 7644
rect 4692 7642 4716 7644
rect 4772 7642 4796 7644
rect 4852 7642 4858 7644
rect 4612 7590 4614 7642
rect 4794 7590 4796 7642
rect 4550 7588 4556 7590
rect 4612 7588 4636 7590
rect 4692 7588 4716 7590
rect 4772 7588 4796 7590
rect 4852 7588 4858 7590
rect 4550 7579 4858 7588
rect 4550 6556 4858 6565
rect 4550 6554 4556 6556
rect 4612 6554 4636 6556
rect 4692 6554 4716 6556
rect 4772 6554 4796 6556
rect 4852 6554 4858 6556
rect 4612 6502 4614 6554
rect 4794 6502 4796 6554
rect 4550 6500 4556 6502
rect 4612 6500 4636 6502
rect 4692 6500 4716 6502
rect 4772 6500 4796 6502
rect 4852 6500 4858 6502
rect 4550 6491 4858 6500
rect 4550 5468 4858 5477
rect 4550 5466 4556 5468
rect 4612 5466 4636 5468
rect 4692 5466 4716 5468
rect 4772 5466 4796 5468
rect 4852 5466 4858 5468
rect 4612 5414 4614 5466
rect 4794 5414 4796 5466
rect 4550 5412 4556 5414
rect 4612 5412 4636 5414
rect 4692 5412 4716 5414
rect 4772 5412 4796 5414
rect 4852 5412 4858 5414
rect 4550 5403 4858 5412
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 2950 4380 3258 4389
rect 2950 4378 2956 4380
rect 3012 4378 3036 4380
rect 3092 4378 3116 4380
rect 3172 4378 3196 4380
rect 3252 4378 3258 4380
rect 3012 4326 3014 4378
rect 3194 4326 3196 4378
rect 2950 4324 2956 4326
rect 3012 4324 3036 4326
rect 3092 4324 3116 4326
rect 3172 4324 3196 4326
rect 3252 4324 3258 4326
rect 2950 4315 3258 4324
rect 4550 4380 4858 4389
rect 4550 4378 4556 4380
rect 4612 4378 4636 4380
rect 4692 4378 4716 4380
rect 4772 4378 4796 4380
rect 4852 4378 4858 4380
rect 4612 4326 4614 4378
rect 4794 4326 4796 4378
rect 4550 4324 4556 4326
rect 4612 4324 4636 4326
rect 4692 4324 4716 4326
rect 4772 4324 4796 4326
rect 4852 4324 4858 4326
rect 4550 4315 4858 4324
rect 3610 3836 3918 3845
rect 3610 3834 3616 3836
rect 3672 3834 3696 3836
rect 3752 3834 3776 3836
rect 3832 3834 3856 3836
rect 3912 3834 3918 3836
rect 3672 3782 3674 3834
rect 3854 3782 3856 3834
rect 3610 3780 3616 3782
rect 3672 3780 3696 3782
rect 3752 3780 3776 3782
rect 3832 3780 3856 3782
rect 3912 3780 3918 3782
rect 3610 3771 3918 3780
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2950 3292 3258 3301
rect 2950 3290 2956 3292
rect 3012 3290 3036 3292
rect 3092 3290 3116 3292
rect 3172 3290 3196 3292
rect 3252 3290 3258 3292
rect 3012 3238 3014 3290
rect 3194 3238 3196 3290
rect 2950 3236 2956 3238
rect 3012 3236 3036 3238
rect 3092 3236 3116 3238
rect 3172 3236 3196 3238
rect 3252 3236 3258 3238
rect 2950 3227 3258 3236
rect 4550 3292 4858 3301
rect 4550 3290 4556 3292
rect 4612 3290 4636 3292
rect 4692 3290 4716 3292
rect 4772 3290 4796 3292
rect 4852 3290 4858 3292
rect 4612 3238 4614 3290
rect 4794 3238 4796 3290
rect 4550 3236 4556 3238
rect 4612 3236 4636 3238
rect 4692 3236 4716 3238
rect 4772 3236 4796 3238
rect 4852 3236 4858 3238
rect 4550 3227 4858 3236
rect 3610 2748 3918 2757
rect 3610 2746 3616 2748
rect 3672 2746 3696 2748
rect 3752 2746 3776 2748
rect 3832 2746 3856 2748
rect 3912 2746 3918 2748
rect 3672 2694 3674 2746
rect 3854 2694 3856 2746
rect 3610 2692 3616 2694
rect 3672 2692 3696 2694
rect 3752 2692 3776 2694
rect 3832 2692 3856 2694
rect 3912 2692 3918 2694
rect 3610 2683 3918 2692
rect 2950 2204 3258 2213
rect 2950 2202 2956 2204
rect 3012 2202 3036 2204
rect 3092 2202 3116 2204
rect 3172 2202 3196 2204
rect 3252 2202 3258 2204
rect 3012 2150 3014 2202
rect 3194 2150 3196 2202
rect 2950 2148 2956 2150
rect 3012 2148 3036 2150
rect 3092 2148 3116 2150
rect 3172 2148 3196 2150
rect 3252 2148 3258 2150
rect 2950 2139 3258 2148
rect 4550 2204 4858 2213
rect 4550 2202 4556 2204
rect 4612 2202 4636 2204
rect 4692 2202 4716 2204
rect 4772 2202 4796 2204
rect 4852 2202 4858 2204
rect 4612 2150 4614 2202
rect 4794 2150 4796 2202
rect 4550 2148 4556 2150
rect 4612 2148 4636 2150
rect 4692 2148 4716 2150
rect 4772 2148 4796 2150
rect 4852 2148 4858 2150
rect 4550 2139 4858 2148
rect 1674 2000 1730 2009
rect 1674 1935 1730 1944
rect 3610 1660 3918 1669
rect 3610 1658 3616 1660
rect 3672 1658 3696 1660
rect 3752 1658 3776 1660
rect 3832 1658 3856 1660
rect 3912 1658 3918 1660
rect 3672 1606 3674 1658
rect 3854 1606 3856 1658
rect 3610 1604 3616 1606
rect 3672 1604 3696 1606
rect 3752 1604 3776 1606
rect 3832 1604 3856 1606
rect 3912 1604 3918 1606
rect 3610 1595 3918 1604
rect 2950 1116 3258 1125
rect 2950 1114 2956 1116
rect 3012 1114 3036 1116
rect 3092 1114 3116 1116
rect 3172 1114 3196 1116
rect 3252 1114 3258 1116
rect 3012 1062 3014 1114
rect 3194 1062 3196 1114
rect 2950 1060 2956 1062
rect 3012 1060 3036 1062
rect 3092 1060 3116 1062
rect 3172 1060 3196 1062
rect 3252 1060 3258 1062
rect 2950 1051 3258 1060
rect 4550 1116 4858 1125
rect 4550 1114 4556 1116
rect 4612 1114 4636 1116
rect 4692 1114 4716 1116
rect 4772 1114 4796 1116
rect 4852 1114 4858 1116
rect 4612 1062 4614 1114
rect 4794 1062 4796 1114
rect 4550 1060 4556 1062
rect 4612 1060 4636 1062
rect 4692 1060 4716 1062
rect 4772 1060 4796 1062
rect 4852 1060 4858 1062
rect 4550 1051 4858 1060
rect 5000 785 5028 23530
rect 5092 3602 5120 25214
rect 5184 24834 5212 25350
rect 5552 24954 5580 25758
rect 5540 24948 5592 24954
rect 5540 24890 5592 24896
rect 5184 24806 5580 24834
rect 5210 24508 5518 24517
rect 5210 24506 5216 24508
rect 5272 24506 5296 24508
rect 5352 24506 5376 24508
rect 5432 24506 5456 24508
rect 5512 24506 5518 24508
rect 5272 24454 5274 24506
rect 5454 24454 5456 24506
rect 5210 24452 5216 24454
rect 5272 24452 5296 24454
rect 5352 24452 5376 24454
rect 5432 24452 5456 24454
rect 5512 24452 5518 24454
rect 5210 24443 5518 24452
rect 5210 23420 5518 23429
rect 5210 23418 5216 23420
rect 5272 23418 5296 23420
rect 5352 23418 5376 23420
rect 5432 23418 5456 23420
rect 5512 23418 5518 23420
rect 5272 23366 5274 23418
rect 5454 23366 5456 23418
rect 5210 23364 5216 23366
rect 5272 23364 5296 23366
rect 5352 23364 5376 23366
rect 5432 23364 5456 23366
rect 5512 23364 5518 23366
rect 5210 23355 5518 23364
rect 5210 22332 5518 22341
rect 5210 22330 5216 22332
rect 5272 22330 5296 22332
rect 5352 22330 5376 22332
rect 5432 22330 5456 22332
rect 5512 22330 5518 22332
rect 5272 22278 5274 22330
rect 5454 22278 5456 22330
rect 5210 22276 5216 22278
rect 5272 22276 5296 22278
rect 5352 22276 5376 22278
rect 5432 22276 5456 22278
rect 5512 22276 5518 22278
rect 5210 22267 5518 22276
rect 5210 21244 5518 21253
rect 5210 21242 5216 21244
rect 5272 21242 5296 21244
rect 5352 21242 5376 21244
rect 5432 21242 5456 21244
rect 5512 21242 5518 21244
rect 5272 21190 5274 21242
rect 5454 21190 5456 21242
rect 5210 21188 5216 21190
rect 5272 21188 5296 21190
rect 5352 21188 5376 21190
rect 5432 21188 5456 21190
rect 5512 21188 5518 21190
rect 5210 21179 5518 21188
rect 5210 20156 5518 20165
rect 5210 20154 5216 20156
rect 5272 20154 5296 20156
rect 5352 20154 5376 20156
rect 5432 20154 5456 20156
rect 5512 20154 5518 20156
rect 5272 20102 5274 20154
rect 5454 20102 5456 20154
rect 5210 20100 5216 20102
rect 5272 20100 5296 20102
rect 5352 20100 5376 20102
rect 5432 20100 5456 20102
rect 5512 20100 5518 20102
rect 5210 20091 5518 20100
rect 5210 19068 5518 19077
rect 5210 19066 5216 19068
rect 5272 19066 5296 19068
rect 5352 19066 5376 19068
rect 5432 19066 5456 19068
rect 5512 19066 5518 19068
rect 5272 19014 5274 19066
rect 5454 19014 5456 19066
rect 5210 19012 5216 19014
rect 5272 19012 5296 19014
rect 5352 19012 5376 19014
rect 5432 19012 5456 19014
rect 5512 19012 5518 19014
rect 5210 19003 5518 19012
rect 5210 17980 5518 17989
rect 5210 17978 5216 17980
rect 5272 17978 5296 17980
rect 5352 17978 5376 17980
rect 5432 17978 5456 17980
rect 5512 17978 5518 17980
rect 5272 17926 5274 17978
rect 5454 17926 5456 17978
rect 5210 17924 5216 17926
rect 5272 17924 5296 17926
rect 5352 17924 5376 17926
rect 5432 17924 5456 17926
rect 5512 17924 5518 17926
rect 5210 17915 5518 17924
rect 5210 16892 5518 16901
rect 5210 16890 5216 16892
rect 5272 16890 5296 16892
rect 5352 16890 5376 16892
rect 5432 16890 5456 16892
rect 5512 16890 5518 16892
rect 5272 16838 5274 16890
rect 5454 16838 5456 16890
rect 5210 16836 5216 16838
rect 5272 16836 5296 16838
rect 5352 16836 5376 16838
rect 5432 16836 5456 16838
rect 5512 16836 5518 16838
rect 5210 16827 5518 16836
rect 5210 15804 5518 15813
rect 5210 15802 5216 15804
rect 5272 15802 5296 15804
rect 5352 15802 5376 15804
rect 5432 15802 5456 15804
rect 5512 15802 5518 15804
rect 5272 15750 5274 15802
rect 5454 15750 5456 15802
rect 5210 15748 5216 15750
rect 5272 15748 5296 15750
rect 5352 15748 5376 15750
rect 5432 15748 5456 15750
rect 5512 15748 5518 15750
rect 5210 15739 5518 15748
rect 5210 14716 5518 14725
rect 5210 14714 5216 14716
rect 5272 14714 5296 14716
rect 5352 14714 5376 14716
rect 5432 14714 5456 14716
rect 5512 14714 5518 14716
rect 5272 14662 5274 14714
rect 5454 14662 5456 14714
rect 5210 14660 5216 14662
rect 5272 14660 5296 14662
rect 5352 14660 5376 14662
rect 5432 14660 5456 14662
rect 5512 14660 5518 14662
rect 5210 14651 5518 14660
rect 5210 13628 5518 13637
rect 5210 13626 5216 13628
rect 5272 13626 5296 13628
rect 5352 13626 5376 13628
rect 5432 13626 5456 13628
rect 5512 13626 5518 13628
rect 5272 13574 5274 13626
rect 5454 13574 5456 13626
rect 5210 13572 5216 13574
rect 5272 13572 5296 13574
rect 5352 13572 5376 13574
rect 5432 13572 5456 13574
rect 5512 13572 5518 13574
rect 5210 13563 5518 13572
rect 5210 12540 5518 12549
rect 5210 12538 5216 12540
rect 5272 12538 5296 12540
rect 5352 12538 5376 12540
rect 5432 12538 5456 12540
rect 5512 12538 5518 12540
rect 5272 12486 5274 12538
rect 5454 12486 5456 12538
rect 5210 12484 5216 12486
rect 5272 12484 5296 12486
rect 5352 12484 5376 12486
rect 5432 12484 5456 12486
rect 5512 12484 5518 12486
rect 5210 12475 5518 12484
rect 5210 11452 5518 11461
rect 5210 11450 5216 11452
rect 5272 11450 5296 11452
rect 5352 11450 5376 11452
rect 5432 11450 5456 11452
rect 5512 11450 5518 11452
rect 5272 11398 5274 11450
rect 5454 11398 5456 11450
rect 5210 11396 5216 11398
rect 5272 11396 5296 11398
rect 5352 11396 5376 11398
rect 5432 11396 5456 11398
rect 5512 11396 5518 11398
rect 5210 11387 5518 11396
rect 5552 11354 5580 24806
rect 5644 23730 5672 29446
rect 5736 24206 5764 29566
rect 5828 28422 5856 40122
rect 5920 31958 5948 40394
rect 6150 40284 6458 40293
rect 6150 40282 6156 40284
rect 6212 40282 6236 40284
rect 6292 40282 6316 40284
rect 6372 40282 6396 40284
rect 6452 40282 6458 40284
rect 6212 40230 6214 40282
rect 6394 40230 6396 40282
rect 6150 40228 6156 40230
rect 6212 40228 6236 40230
rect 6292 40228 6316 40230
rect 6372 40228 6396 40230
rect 6452 40228 6458 40230
rect 6150 40219 6458 40228
rect 6000 39296 6052 39302
rect 6000 39238 6052 39244
rect 5908 31952 5960 31958
rect 6012 31929 6040 39238
rect 6150 39196 6458 39205
rect 6150 39194 6156 39196
rect 6212 39194 6236 39196
rect 6292 39194 6316 39196
rect 6372 39194 6396 39196
rect 6452 39194 6458 39196
rect 6212 39142 6214 39194
rect 6394 39142 6396 39194
rect 6150 39140 6156 39142
rect 6212 39140 6236 39142
rect 6292 39140 6316 39142
rect 6372 39140 6396 39142
rect 6452 39140 6458 39142
rect 6150 39131 6458 39140
rect 6150 38108 6458 38117
rect 6150 38106 6156 38108
rect 6212 38106 6236 38108
rect 6292 38106 6316 38108
rect 6372 38106 6396 38108
rect 6452 38106 6458 38108
rect 6212 38054 6214 38106
rect 6394 38054 6396 38106
rect 6150 38052 6156 38054
rect 6212 38052 6236 38054
rect 6292 38052 6316 38054
rect 6372 38052 6396 38054
rect 6452 38052 6458 38054
rect 6150 38043 6458 38052
rect 6150 37020 6458 37029
rect 6150 37018 6156 37020
rect 6212 37018 6236 37020
rect 6292 37018 6316 37020
rect 6372 37018 6396 37020
rect 6452 37018 6458 37020
rect 6212 36966 6214 37018
rect 6394 36966 6396 37018
rect 6150 36964 6156 36966
rect 6212 36964 6236 36966
rect 6292 36964 6316 36966
rect 6372 36964 6396 36966
rect 6452 36964 6458 36966
rect 6150 36955 6458 36964
rect 6460 36644 6512 36650
rect 6460 36586 6512 36592
rect 6472 36122 6500 36586
rect 6564 36394 6592 51886
rect 6656 49434 6684 52634
rect 6748 52578 6776 56646
rect 6840 56166 6868 56850
rect 7196 56704 7248 56710
rect 7196 56646 7248 56652
rect 6828 56160 6880 56166
rect 6828 56102 6880 56108
rect 6810 56060 7118 56069
rect 6810 56058 6816 56060
rect 6872 56058 6896 56060
rect 6952 56058 6976 56060
rect 7032 56058 7056 56060
rect 7112 56058 7118 56060
rect 6872 56006 6874 56058
rect 7054 56006 7056 56058
rect 6810 56004 6816 56006
rect 6872 56004 6896 56006
rect 6952 56004 6976 56006
rect 7032 56004 7056 56006
rect 7112 56004 7118 56006
rect 6810 55995 7118 56004
rect 6810 54972 7118 54981
rect 6810 54970 6816 54972
rect 6872 54970 6896 54972
rect 6952 54970 6976 54972
rect 7032 54970 7056 54972
rect 7112 54970 7118 54972
rect 6872 54918 6874 54970
rect 7054 54918 7056 54970
rect 6810 54916 6816 54918
rect 6872 54916 6896 54918
rect 6952 54916 6976 54918
rect 7032 54916 7056 54918
rect 7112 54916 7118 54918
rect 6810 54907 7118 54916
rect 6810 53884 7118 53893
rect 6810 53882 6816 53884
rect 6872 53882 6896 53884
rect 6952 53882 6976 53884
rect 7032 53882 7056 53884
rect 7112 53882 7118 53884
rect 6872 53830 6874 53882
rect 7054 53830 7056 53882
rect 6810 53828 6816 53830
rect 6872 53828 6896 53830
rect 6952 53828 6976 53830
rect 7032 53828 7056 53830
rect 7112 53828 7118 53830
rect 6810 53819 7118 53828
rect 7012 53780 7064 53786
rect 7012 53722 7064 53728
rect 7024 53242 7052 53722
rect 7104 53576 7156 53582
rect 7102 53544 7104 53553
rect 7156 53544 7158 53553
rect 7102 53479 7158 53488
rect 7104 53440 7156 53446
rect 7104 53382 7156 53388
rect 7012 53236 7064 53242
rect 7012 53178 7064 53184
rect 7116 53174 7144 53382
rect 7208 53242 7236 56646
rect 7300 53582 7328 57734
rect 7380 57316 7432 57322
rect 7380 57258 7432 57264
rect 7392 53582 7420 57258
rect 7484 54262 7512 58278
rect 7576 57934 7604 62206
rect 7668 61266 7696 62630
rect 7852 62286 7880 62766
rect 7840 62280 7892 62286
rect 7840 62222 7892 62228
rect 7750 62044 8058 62053
rect 7750 62042 7756 62044
rect 7812 62042 7836 62044
rect 7892 62042 7916 62044
rect 7972 62042 7996 62044
rect 8052 62042 8058 62044
rect 7812 61990 7814 62042
rect 7994 61990 7996 62042
rect 7750 61988 7756 61990
rect 7812 61988 7836 61990
rect 7892 61988 7916 61990
rect 7972 61988 7996 61990
rect 8052 61988 8058 61990
rect 7750 61979 8058 61988
rect 7748 61804 7800 61810
rect 7748 61746 7800 61752
rect 7656 61260 7708 61266
rect 7656 61202 7708 61208
rect 7760 61044 7788 61746
rect 8128 61690 8156 63192
rect 8220 61826 8248 63260
rect 8312 63034 8340 63786
rect 8410 63676 8718 63685
rect 8410 63674 8416 63676
rect 8472 63674 8496 63676
rect 8552 63674 8576 63676
rect 8632 63674 8656 63676
rect 8712 63674 8718 63676
rect 8472 63622 8474 63674
rect 8654 63622 8656 63674
rect 8410 63620 8416 63622
rect 8472 63620 8496 63622
rect 8552 63620 8576 63622
rect 8632 63620 8656 63622
rect 8712 63620 8718 63622
rect 8410 63611 8718 63620
rect 8392 63436 8444 63442
rect 8772 63424 8800 64942
rect 8864 64394 8892 65962
rect 8852 64388 8904 64394
rect 8852 64330 8904 64336
rect 8852 64116 8904 64122
rect 8852 64058 8904 64064
rect 8444 63396 8800 63424
rect 8392 63378 8444 63384
rect 8864 63374 8892 64058
rect 8956 63442 8984 66438
rect 9048 66162 9076 66642
rect 9232 66638 9260 66778
rect 9324 66638 9352 67215
rect 9404 67176 9456 67182
rect 9402 67144 9404 67153
rect 9456 67144 9458 67153
rect 9402 67079 9458 67088
rect 9600 66638 9628 67340
rect 9220 66632 9272 66638
rect 9220 66574 9272 66580
rect 9312 66632 9364 66638
rect 9312 66574 9364 66580
rect 9588 66632 9640 66638
rect 9588 66574 9640 66580
rect 9128 66292 9180 66298
rect 9128 66234 9180 66240
rect 9036 66156 9088 66162
rect 9036 66098 9088 66104
rect 9036 66020 9088 66026
rect 9036 65962 9088 65968
rect 9048 65090 9076 65962
rect 9140 65210 9168 66234
rect 9128 65204 9180 65210
rect 9128 65146 9180 65152
rect 9048 65062 9168 65090
rect 9036 65000 9088 65006
rect 9036 64942 9088 64948
rect 9048 64530 9076 64942
rect 9036 64524 9088 64530
rect 9036 64466 9088 64472
rect 9036 64388 9088 64394
rect 9036 64330 9088 64336
rect 9048 63442 9076 64330
rect 9140 64326 9168 65062
rect 9232 64988 9260 66574
rect 9350 66396 9658 66405
rect 9350 66394 9356 66396
rect 9412 66394 9436 66396
rect 9492 66394 9516 66396
rect 9572 66394 9596 66396
rect 9652 66394 9658 66396
rect 9412 66342 9414 66394
rect 9594 66342 9596 66394
rect 9350 66340 9356 66342
rect 9412 66340 9436 66342
rect 9492 66340 9516 66342
rect 9572 66340 9596 66342
rect 9652 66340 9658 66342
rect 9350 66331 9658 66340
rect 9312 66292 9364 66298
rect 9312 66234 9364 66240
rect 9324 65414 9352 66234
rect 9312 65408 9364 65414
rect 9312 65350 9364 65356
rect 9350 65308 9658 65317
rect 9350 65306 9356 65308
rect 9412 65306 9436 65308
rect 9492 65306 9516 65308
rect 9572 65306 9596 65308
rect 9652 65306 9658 65308
rect 9412 65254 9414 65306
rect 9594 65254 9596 65306
rect 9350 65252 9356 65254
rect 9412 65252 9436 65254
rect 9492 65252 9516 65254
rect 9572 65252 9596 65254
rect 9652 65252 9658 65254
rect 9350 65243 9658 65252
rect 9312 65000 9364 65006
rect 9232 64960 9312 64988
rect 9128 64320 9180 64326
rect 9128 64262 9180 64268
rect 9232 64138 9260 64960
rect 9312 64942 9364 64948
rect 9496 65000 9548 65006
rect 9496 64942 9548 64948
rect 9508 64870 9536 64942
rect 9496 64864 9548 64870
rect 9496 64806 9548 64812
rect 9350 64220 9658 64229
rect 9350 64218 9356 64220
rect 9412 64218 9436 64220
rect 9492 64218 9516 64220
rect 9572 64218 9596 64220
rect 9652 64218 9658 64220
rect 9412 64166 9414 64218
rect 9594 64166 9596 64218
rect 9350 64164 9356 64166
rect 9412 64164 9436 64166
rect 9492 64164 9516 64166
rect 9572 64164 9596 64166
rect 9652 64164 9658 64166
rect 9350 64155 9658 64164
rect 9140 64110 9260 64138
rect 8944 63436 8996 63442
rect 8944 63378 8996 63384
rect 9036 63436 9088 63442
rect 9036 63378 9088 63384
rect 8852 63368 8904 63374
rect 8390 63336 8446 63345
rect 8852 63310 8904 63316
rect 8942 63336 8998 63345
rect 8390 63271 8446 63280
rect 8998 63294 9076 63322
rect 8942 63271 8998 63280
rect 8300 63028 8352 63034
rect 8300 62970 8352 62976
rect 8404 62812 8432 63271
rect 8760 63232 8812 63238
rect 8760 63174 8812 63180
rect 8944 63232 8996 63238
rect 8944 63174 8996 63180
rect 8772 63034 8800 63174
rect 8760 63028 8812 63034
rect 8760 62970 8812 62976
rect 8666 62928 8722 62937
rect 8666 62863 8668 62872
rect 8720 62863 8722 62872
rect 8668 62834 8720 62840
rect 8484 62824 8536 62830
rect 8312 62784 8484 62812
rect 8312 61946 8340 62784
rect 8484 62766 8536 62772
rect 8760 62824 8812 62830
rect 8760 62766 8812 62772
rect 8410 62588 8718 62597
rect 8410 62586 8416 62588
rect 8472 62586 8496 62588
rect 8552 62586 8576 62588
rect 8632 62586 8656 62588
rect 8712 62586 8718 62588
rect 8472 62534 8474 62586
rect 8654 62534 8656 62586
rect 8410 62532 8416 62534
rect 8472 62532 8496 62534
rect 8552 62532 8576 62534
rect 8632 62532 8656 62534
rect 8712 62532 8718 62534
rect 8410 62523 8718 62532
rect 8772 62286 8800 62766
rect 8852 62484 8904 62490
rect 8852 62426 8904 62432
rect 8760 62280 8812 62286
rect 8760 62222 8812 62228
rect 8300 61940 8352 61946
rect 8300 61882 8352 61888
rect 8772 61878 8800 62222
rect 8392 61872 8444 61878
rect 8220 61820 8392 61826
rect 8220 61814 8444 61820
rect 8760 61872 8812 61878
rect 8760 61814 8812 61820
rect 8220 61810 8432 61814
rect 8208 61804 8432 61810
rect 8260 61798 8432 61804
rect 8208 61746 8260 61752
rect 7944 61662 8156 61690
rect 8300 61736 8352 61742
rect 8300 61678 8352 61684
rect 8760 61736 8812 61742
rect 8760 61678 8812 61684
rect 7944 61146 7972 61662
rect 8024 61600 8076 61606
rect 8024 61542 8076 61548
rect 8116 61600 8168 61606
rect 8116 61542 8168 61548
rect 8036 61402 8064 61542
rect 8024 61396 8076 61402
rect 8024 61338 8076 61344
rect 8128 61282 8156 61542
rect 8128 61254 8248 61282
rect 7944 61118 8156 61146
rect 7668 61016 7788 61044
rect 7668 60790 7696 61016
rect 7750 60956 8058 60965
rect 7750 60954 7756 60956
rect 7812 60954 7836 60956
rect 7892 60954 7916 60956
rect 7972 60954 7996 60956
rect 8052 60954 8058 60956
rect 7812 60902 7814 60954
rect 7994 60902 7996 60954
rect 7750 60900 7756 60902
rect 7812 60900 7836 60902
rect 7892 60900 7916 60902
rect 7972 60900 7996 60902
rect 8052 60900 8058 60902
rect 7750 60891 8058 60900
rect 7656 60784 7708 60790
rect 7656 60726 7708 60732
rect 7656 60308 7708 60314
rect 7656 60250 7708 60256
rect 7668 59650 7696 60250
rect 7750 59868 8058 59877
rect 7750 59866 7756 59868
rect 7812 59866 7836 59868
rect 7892 59866 7916 59868
rect 7972 59866 7996 59868
rect 8052 59866 8058 59868
rect 7812 59814 7814 59866
rect 7994 59814 7996 59866
rect 7750 59812 7756 59814
rect 7812 59812 7836 59814
rect 7892 59812 7916 59814
rect 7972 59812 7996 59814
rect 8052 59812 8058 59814
rect 7750 59803 8058 59812
rect 7668 59622 7788 59650
rect 7656 59016 7708 59022
rect 7656 58958 7708 58964
rect 7668 58664 7696 58958
rect 7760 58886 7788 59622
rect 7748 58880 7800 58886
rect 7748 58822 7800 58828
rect 7750 58780 8058 58789
rect 7750 58778 7756 58780
rect 7812 58778 7836 58780
rect 7892 58778 7916 58780
rect 7972 58778 7996 58780
rect 8052 58778 8058 58780
rect 7812 58726 7814 58778
rect 7994 58726 7996 58778
rect 7750 58724 7756 58726
rect 7812 58724 7836 58726
rect 7892 58724 7916 58726
rect 7972 58724 7996 58726
rect 8052 58724 8058 58726
rect 7750 58715 8058 58724
rect 7668 58636 7788 58664
rect 7656 58472 7708 58478
rect 7656 58414 7708 58420
rect 7564 57928 7616 57934
rect 7564 57870 7616 57876
rect 7564 57384 7616 57390
rect 7564 57326 7616 57332
rect 7576 55758 7604 57326
rect 7668 56506 7696 58414
rect 7760 57934 7788 58636
rect 7748 57928 7800 57934
rect 7748 57870 7800 57876
rect 7750 57692 8058 57701
rect 7750 57690 7756 57692
rect 7812 57690 7836 57692
rect 7892 57690 7916 57692
rect 7972 57690 7996 57692
rect 8052 57690 8058 57692
rect 7812 57638 7814 57690
rect 7994 57638 7996 57690
rect 7750 57636 7756 57638
rect 7812 57636 7836 57638
rect 7892 57636 7916 57638
rect 7972 57636 7996 57638
rect 8052 57636 8058 57638
rect 7750 57627 8058 57636
rect 7750 56604 8058 56613
rect 7750 56602 7756 56604
rect 7812 56602 7836 56604
rect 7892 56602 7916 56604
rect 7972 56602 7996 56604
rect 8052 56602 8058 56604
rect 7812 56550 7814 56602
rect 7994 56550 7996 56602
rect 7750 56548 7756 56550
rect 7812 56548 7836 56550
rect 7892 56548 7916 56550
rect 7972 56548 7996 56550
rect 8052 56548 8058 56550
rect 7750 56539 8058 56548
rect 7656 56500 7708 56506
rect 7656 56442 7708 56448
rect 7656 56160 7708 56166
rect 7656 56102 7708 56108
rect 7564 55752 7616 55758
rect 7564 55694 7616 55700
rect 7576 55418 7604 55694
rect 7564 55412 7616 55418
rect 7564 55354 7616 55360
rect 7668 54312 7696 56102
rect 8128 55758 8156 61118
rect 8220 60314 8248 61254
rect 8312 60586 8340 61678
rect 8410 61500 8718 61509
rect 8410 61498 8416 61500
rect 8472 61498 8496 61500
rect 8552 61498 8576 61500
rect 8632 61498 8656 61500
rect 8712 61498 8718 61500
rect 8472 61446 8474 61498
rect 8654 61446 8656 61498
rect 8410 61444 8416 61446
rect 8472 61444 8496 61446
rect 8552 61444 8576 61446
rect 8632 61444 8656 61446
rect 8712 61444 8718 61446
rect 8410 61435 8718 61444
rect 8772 61266 8800 61678
rect 8760 61260 8812 61266
rect 8760 61202 8812 61208
rect 8760 61124 8812 61130
rect 8760 61066 8812 61072
rect 8300 60580 8352 60586
rect 8300 60522 8352 60528
rect 8410 60412 8718 60421
rect 8410 60410 8416 60412
rect 8472 60410 8496 60412
rect 8552 60410 8576 60412
rect 8632 60410 8656 60412
rect 8712 60410 8718 60412
rect 8472 60358 8474 60410
rect 8654 60358 8656 60410
rect 8410 60356 8416 60358
rect 8472 60356 8496 60358
rect 8552 60356 8576 60358
rect 8632 60356 8656 60358
rect 8712 60356 8718 60358
rect 8410 60347 8718 60356
rect 8208 60308 8260 60314
rect 8208 60250 8260 60256
rect 8208 60036 8260 60042
rect 8208 59978 8260 59984
rect 8220 58546 8248 59978
rect 8300 59968 8352 59974
rect 8300 59910 8352 59916
rect 8312 58682 8340 59910
rect 8410 59324 8718 59333
rect 8410 59322 8416 59324
rect 8472 59322 8496 59324
rect 8552 59322 8576 59324
rect 8632 59322 8656 59324
rect 8712 59322 8718 59324
rect 8472 59270 8474 59322
rect 8654 59270 8656 59322
rect 8410 59268 8416 59270
rect 8472 59268 8496 59270
rect 8552 59268 8576 59270
rect 8632 59268 8656 59270
rect 8712 59268 8718 59270
rect 8410 59259 8718 59268
rect 8392 58880 8444 58886
rect 8392 58822 8444 58828
rect 8300 58676 8352 58682
rect 8300 58618 8352 58624
rect 8208 58540 8260 58546
rect 8208 58482 8260 58488
rect 8404 58426 8432 58822
rect 8772 58478 8800 61066
rect 8864 60330 8892 62426
rect 8956 61674 8984 63174
rect 8944 61668 8996 61674
rect 8944 61610 8996 61616
rect 8956 61402 8984 61610
rect 8944 61396 8996 61402
rect 8944 61338 8996 61344
rect 8944 61192 8996 61198
rect 8944 61134 8996 61140
rect 8956 60858 8984 61134
rect 8944 60852 8996 60858
rect 8944 60794 8996 60800
rect 9048 60489 9076 63294
rect 9140 61266 9168 64110
rect 9220 63776 9272 63782
rect 9220 63718 9272 63724
rect 9128 61260 9180 61266
rect 9128 61202 9180 61208
rect 9128 61056 9180 61062
rect 9128 60998 9180 61004
rect 9034 60480 9090 60489
rect 9034 60415 9090 60424
rect 8864 60302 9076 60330
rect 8852 60240 8904 60246
rect 8852 60182 8904 60188
rect 8942 60208 8998 60217
rect 8208 58404 8260 58410
rect 8208 58346 8260 58352
rect 8312 58398 8432 58426
rect 8760 58472 8812 58478
rect 8760 58414 8812 58420
rect 8220 57866 8248 58346
rect 8312 58002 8340 58398
rect 8760 58336 8812 58342
rect 8760 58278 8812 58284
rect 8410 58236 8718 58245
rect 8410 58234 8416 58236
rect 8472 58234 8496 58236
rect 8552 58234 8576 58236
rect 8632 58234 8656 58236
rect 8712 58234 8718 58236
rect 8472 58182 8474 58234
rect 8654 58182 8656 58234
rect 8410 58180 8416 58182
rect 8472 58180 8496 58182
rect 8552 58180 8576 58182
rect 8632 58180 8656 58182
rect 8712 58180 8718 58182
rect 8410 58171 8718 58180
rect 8300 57996 8352 58002
rect 8772 57974 8800 58278
rect 8300 57938 8352 57944
rect 8680 57946 8800 57974
rect 8298 57896 8354 57905
rect 8208 57860 8260 57866
rect 8298 57831 8354 57840
rect 8208 57802 8260 57808
rect 8206 57760 8262 57769
rect 8206 57695 8262 57704
rect 8220 56302 8248 57695
rect 8208 56296 8260 56302
rect 8208 56238 8260 56244
rect 8208 55820 8260 55826
rect 8312 55808 8340 57831
rect 8576 57792 8628 57798
rect 8576 57734 8628 57740
rect 8680 57746 8708 57946
rect 8864 57905 8892 60182
rect 8942 60143 8998 60152
rect 8850 57896 8906 57905
rect 8850 57831 8906 57840
rect 8852 57792 8904 57798
rect 8588 57322 8616 57734
rect 8680 57718 8800 57746
rect 8852 57734 8904 57740
rect 8576 57316 8628 57322
rect 8576 57258 8628 57264
rect 8410 57148 8718 57157
rect 8410 57146 8416 57148
rect 8472 57146 8496 57148
rect 8552 57146 8576 57148
rect 8632 57146 8656 57148
rect 8712 57146 8718 57148
rect 8472 57094 8474 57146
rect 8654 57094 8656 57146
rect 8410 57092 8416 57094
rect 8472 57092 8496 57094
rect 8552 57092 8576 57094
rect 8632 57092 8656 57094
rect 8712 57092 8718 57094
rect 8410 57083 8718 57092
rect 8410 56060 8718 56069
rect 8410 56058 8416 56060
rect 8472 56058 8496 56060
rect 8552 56058 8576 56060
rect 8632 56058 8656 56060
rect 8712 56058 8718 56060
rect 8472 56006 8474 56058
rect 8654 56006 8656 56058
rect 8410 56004 8416 56006
rect 8472 56004 8496 56006
rect 8552 56004 8576 56006
rect 8632 56004 8656 56006
rect 8712 56004 8718 56006
rect 8410 55995 8718 56004
rect 8260 55780 8340 55808
rect 8208 55762 8260 55768
rect 8116 55752 8168 55758
rect 8116 55694 8168 55700
rect 8208 55616 8260 55622
rect 8208 55558 8260 55564
rect 7750 55516 8058 55525
rect 7750 55514 7756 55516
rect 7812 55514 7836 55516
rect 7892 55514 7916 55516
rect 7972 55514 7996 55516
rect 8052 55514 8058 55516
rect 7812 55462 7814 55514
rect 7994 55462 7996 55514
rect 7750 55460 7756 55462
rect 7812 55460 7836 55462
rect 7892 55460 7916 55462
rect 7972 55460 7996 55462
rect 8052 55460 8058 55462
rect 7750 55451 8058 55460
rect 8116 55412 8168 55418
rect 8116 55354 8168 55360
rect 7750 54428 8058 54437
rect 7750 54426 7756 54428
rect 7812 54426 7836 54428
rect 7892 54426 7916 54428
rect 7972 54426 7996 54428
rect 8052 54426 8058 54428
rect 7812 54374 7814 54426
rect 7994 54374 7996 54426
rect 7750 54372 7756 54374
rect 7812 54372 7836 54374
rect 7892 54372 7916 54374
rect 7972 54372 7996 54374
rect 8052 54372 8058 54374
rect 7750 54363 8058 54372
rect 7668 54284 7788 54312
rect 7472 54256 7524 54262
rect 7472 54198 7524 54204
rect 7564 53984 7616 53990
rect 7564 53926 7616 53932
rect 7656 53984 7708 53990
rect 7656 53926 7708 53932
rect 7288 53576 7340 53582
rect 7288 53518 7340 53524
rect 7380 53576 7432 53582
rect 7380 53518 7432 53524
rect 7380 53440 7432 53446
rect 7380 53382 7432 53388
rect 7472 53440 7524 53446
rect 7472 53382 7524 53388
rect 7392 53242 7420 53382
rect 7196 53236 7248 53242
rect 7196 53178 7248 53184
rect 7380 53236 7432 53242
rect 7380 53178 7432 53184
rect 7104 53168 7156 53174
rect 7104 53110 7156 53116
rect 7484 53009 7512 53382
rect 7576 53242 7604 53926
rect 7564 53236 7616 53242
rect 7564 53178 7616 53184
rect 7668 53106 7696 53926
rect 7760 53582 7788 54284
rect 7838 54224 7894 54233
rect 7838 54159 7840 54168
rect 7892 54159 7894 54168
rect 7840 54130 7892 54136
rect 7748 53576 7800 53582
rect 7748 53518 7800 53524
rect 7750 53340 8058 53349
rect 7750 53338 7756 53340
rect 7812 53338 7836 53340
rect 7892 53338 7916 53340
rect 7972 53338 7996 53340
rect 8052 53338 8058 53340
rect 7812 53286 7814 53338
rect 7994 53286 7996 53338
rect 7750 53284 7756 53286
rect 7812 53284 7836 53286
rect 7892 53284 7916 53286
rect 7972 53284 7996 53286
rect 8052 53284 8058 53286
rect 7750 53275 8058 53284
rect 7656 53100 7708 53106
rect 7656 53042 7708 53048
rect 7194 53000 7250 53009
rect 7470 53000 7526 53009
rect 7194 52935 7250 52944
rect 7288 52964 7340 52970
rect 6810 52796 7118 52805
rect 6810 52794 6816 52796
rect 6872 52794 6896 52796
rect 6952 52794 6976 52796
rect 7032 52794 7056 52796
rect 7112 52794 7118 52796
rect 6872 52742 6874 52794
rect 7054 52742 7056 52794
rect 6810 52740 6816 52742
rect 6872 52740 6896 52742
rect 6952 52740 6976 52742
rect 7032 52740 7056 52742
rect 7112 52740 7118 52742
rect 6810 52731 7118 52740
rect 6748 52550 6868 52578
rect 6736 52488 6788 52494
rect 6736 52430 6788 52436
rect 6748 51950 6776 52430
rect 6840 52018 6868 52550
rect 6828 52012 6880 52018
rect 6828 51954 6880 51960
rect 6736 51944 6788 51950
rect 6736 51886 6788 51892
rect 6748 51406 6776 51886
rect 6810 51708 7118 51717
rect 6810 51706 6816 51708
rect 6872 51706 6896 51708
rect 6952 51706 6976 51708
rect 7032 51706 7056 51708
rect 7112 51706 7118 51708
rect 6872 51654 6874 51706
rect 7054 51654 7056 51706
rect 6810 51652 6816 51654
rect 6872 51652 6896 51654
rect 6952 51652 6976 51654
rect 7032 51652 7056 51654
rect 7112 51652 7118 51654
rect 6810 51643 7118 51652
rect 7012 51604 7064 51610
rect 7012 51546 7064 51552
rect 6736 51400 6788 51406
rect 6736 51342 6788 51348
rect 6748 50930 6776 51342
rect 7024 51066 7052 51546
rect 7012 51060 7064 51066
rect 7012 51002 7064 51008
rect 6736 50924 6788 50930
rect 6736 50866 6788 50872
rect 6748 49842 6776 50866
rect 7208 50844 7236 52935
rect 8128 52986 8156 55354
rect 7470 52935 7526 52944
rect 7564 52964 7616 52970
rect 7288 52906 7340 52912
rect 7564 52906 7616 52912
rect 7668 52958 8156 52986
rect 7300 52442 7328 52906
rect 7472 52896 7524 52902
rect 7472 52838 7524 52844
rect 7300 52414 7420 52442
rect 7288 52352 7340 52358
rect 7288 52294 7340 52300
rect 7300 51338 7328 52294
rect 7392 52193 7420 52414
rect 7378 52184 7434 52193
rect 7378 52119 7434 52128
rect 7484 52018 7512 52838
rect 7576 52086 7604 52906
rect 7564 52080 7616 52086
rect 7564 52022 7616 52028
rect 7472 52012 7524 52018
rect 7472 51954 7524 51960
rect 7562 51912 7618 51921
rect 7562 51847 7618 51856
rect 7288 51332 7340 51338
rect 7288 51274 7340 51280
rect 7472 51332 7524 51338
rect 7472 51274 7524 51280
rect 7484 50998 7512 51274
rect 7472 50992 7524 50998
rect 7472 50934 7524 50940
rect 7208 50816 7420 50844
rect 7012 50720 7064 50726
rect 7288 50720 7340 50726
rect 7064 50680 7236 50708
rect 7012 50662 7064 50668
rect 6810 50620 7118 50629
rect 6810 50618 6816 50620
rect 6872 50618 6896 50620
rect 6952 50618 6976 50620
rect 7032 50618 7056 50620
rect 7112 50618 7118 50620
rect 6872 50566 6874 50618
rect 7054 50566 7056 50618
rect 6810 50564 6816 50566
rect 6872 50564 6896 50566
rect 6952 50564 6976 50566
rect 7032 50564 7056 50566
rect 7112 50564 7118 50566
rect 6810 50555 7118 50564
rect 6736 49836 6788 49842
rect 6736 49778 6788 49784
rect 6644 49428 6696 49434
rect 6644 49370 6696 49376
rect 6748 49230 6776 49778
rect 6810 49532 7118 49541
rect 6810 49530 6816 49532
rect 6872 49530 6896 49532
rect 6952 49530 6976 49532
rect 7032 49530 7056 49532
rect 7112 49530 7118 49532
rect 6872 49478 6874 49530
rect 7054 49478 7056 49530
rect 6810 49476 6816 49478
rect 6872 49476 6896 49478
rect 6952 49476 6976 49478
rect 7032 49476 7056 49478
rect 7112 49476 7118 49478
rect 6810 49467 7118 49476
rect 6736 49224 6788 49230
rect 6736 49166 6788 49172
rect 6644 49088 6696 49094
rect 6644 49030 6696 49036
rect 6656 46356 6684 49030
rect 6748 48754 6776 49166
rect 6736 48748 6788 48754
rect 6736 48690 6788 48696
rect 6748 48142 6776 48690
rect 6810 48444 7118 48453
rect 6810 48442 6816 48444
rect 6872 48442 6896 48444
rect 6952 48442 6976 48444
rect 7032 48442 7056 48444
rect 7112 48442 7118 48444
rect 6872 48390 6874 48442
rect 7054 48390 7056 48442
rect 6810 48388 6816 48390
rect 6872 48388 6896 48390
rect 6952 48388 6976 48390
rect 7032 48388 7056 48390
rect 7112 48388 7118 48390
rect 6810 48379 7118 48388
rect 7208 48142 7236 50680
rect 7288 50662 7340 50668
rect 6736 48136 6788 48142
rect 6736 48078 6788 48084
rect 7196 48136 7248 48142
rect 7196 48078 7248 48084
rect 6748 47138 6776 48078
rect 6828 48000 6880 48006
rect 6828 47942 6880 47948
rect 7196 48000 7248 48006
rect 7196 47942 7248 47948
rect 6840 47666 6868 47942
rect 6828 47660 6880 47666
rect 6828 47602 6880 47608
rect 6810 47356 7118 47365
rect 6810 47354 6816 47356
rect 6872 47354 6896 47356
rect 6952 47354 6976 47356
rect 7032 47354 7056 47356
rect 7112 47354 7118 47356
rect 6872 47302 6874 47354
rect 7054 47302 7056 47354
rect 6810 47300 6816 47302
rect 6872 47300 6896 47302
rect 6952 47300 6976 47302
rect 7032 47300 7056 47302
rect 7112 47300 7118 47302
rect 6810 47291 7118 47300
rect 6748 47110 6868 47138
rect 6840 47054 6868 47110
rect 6828 47048 6880 47054
rect 6828 46990 6880 46996
rect 6736 46912 6788 46918
rect 6736 46854 6788 46860
rect 6748 46646 6776 46854
rect 6840 46714 6868 46990
rect 7104 46980 7156 46986
rect 7104 46922 7156 46928
rect 6828 46708 6880 46714
rect 6828 46650 6880 46656
rect 6736 46640 6788 46646
rect 6736 46582 6788 46588
rect 7116 46481 7144 46922
rect 7208 46730 7236 47942
rect 7300 47462 7328 50662
rect 7288 47456 7340 47462
rect 7288 47398 7340 47404
rect 7208 46702 7328 46730
rect 7196 46640 7248 46646
rect 7196 46582 7248 46588
rect 7102 46472 7158 46481
rect 7102 46407 7158 46416
rect 6656 46328 6776 46356
rect 6644 46028 6696 46034
rect 6644 45970 6696 45976
rect 6656 44402 6684 45970
rect 6644 44396 6696 44402
rect 6644 44338 6696 44344
rect 6656 43858 6684 44338
rect 6748 44266 6776 46328
rect 6810 46268 7118 46277
rect 6810 46266 6816 46268
rect 6872 46266 6896 46268
rect 6952 46266 6976 46268
rect 7032 46266 7056 46268
rect 7112 46266 7118 46268
rect 6872 46214 6874 46266
rect 7054 46214 7056 46266
rect 6810 46212 6816 46214
rect 6872 46212 6896 46214
rect 6952 46212 6976 46214
rect 7032 46212 7056 46214
rect 7112 46212 7118 46214
rect 6810 46203 7118 46212
rect 7012 46164 7064 46170
rect 7012 46106 7064 46112
rect 7024 45490 7052 46106
rect 7012 45484 7064 45490
rect 7012 45426 7064 45432
rect 6810 45180 7118 45189
rect 6810 45178 6816 45180
rect 6872 45178 6896 45180
rect 6952 45178 6976 45180
rect 7032 45178 7056 45180
rect 7112 45178 7118 45180
rect 6872 45126 6874 45178
rect 7054 45126 7056 45178
rect 6810 45124 6816 45126
rect 6872 45124 6896 45126
rect 6952 45124 6976 45126
rect 7032 45124 7056 45126
rect 7112 45124 7118 45126
rect 6810 45115 7118 45124
rect 6736 44260 6788 44266
rect 6736 44202 6788 44208
rect 6810 44092 7118 44101
rect 6810 44090 6816 44092
rect 6872 44090 6896 44092
rect 6952 44090 6976 44092
rect 7032 44090 7056 44092
rect 7112 44090 7118 44092
rect 6872 44038 6874 44090
rect 7054 44038 7056 44090
rect 6810 44036 6816 44038
rect 6872 44036 6896 44038
rect 6952 44036 6976 44038
rect 7032 44036 7056 44038
rect 7112 44036 7118 44038
rect 6810 44027 7118 44036
rect 7208 43897 7236 46582
rect 7300 46170 7328 46702
rect 7288 46164 7340 46170
rect 7288 46106 7340 46112
rect 7392 45914 7420 50816
rect 7472 49224 7524 49230
rect 7472 49166 7524 49172
rect 7484 48142 7512 49166
rect 7472 48136 7524 48142
rect 7472 48078 7524 48084
rect 7472 48000 7524 48006
rect 7472 47942 7524 47948
rect 7300 45886 7420 45914
rect 6734 43888 6790 43897
rect 6644 43852 6696 43858
rect 6734 43823 6790 43832
rect 7194 43888 7250 43897
rect 7194 43823 7250 43832
rect 6644 43794 6696 43800
rect 6656 43314 6684 43794
rect 6644 43308 6696 43314
rect 6644 43250 6696 43256
rect 6656 42226 6684 43250
rect 6644 42220 6696 42226
rect 6644 42162 6696 42168
rect 6656 38842 6684 42162
rect 6748 39030 6776 43823
rect 7196 43648 7248 43654
rect 7196 43590 7248 43596
rect 6810 43004 7118 43013
rect 6810 43002 6816 43004
rect 6872 43002 6896 43004
rect 6952 43002 6976 43004
rect 7032 43002 7056 43004
rect 7112 43002 7118 43004
rect 6872 42950 6874 43002
rect 7054 42950 7056 43002
rect 6810 42948 6816 42950
rect 6872 42948 6896 42950
rect 6952 42948 6976 42950
rect 7032 42948 7056 42950
rect 7112 42948 7118 42950
rect 6810 42939 7118 42948
rect 7208 42838 7236 43590
rect 7196 42832 7248 42838
rect 7196 42774 7248 42780
rect 7300 42294 7328 45886
rect 7380 45824 7432 45830
rect 7380 45766 7432 45772
rect 7392 42566 7420 45766
rect 7484 45286 7512 47942
rect 7472 45280 7524 45286
rect 7472 45222 7524 45228
rect 7576 44402 7604 51847
rect 7668 49978 7696 52958
rect 7748 52896 7800 52902
rect 7748 52838 7800 52844
rect 7760 52358 7788 52838
rect 7748 52352 7800 52358
rect 7748 52294 7800 52300
rect 7750 52252 8058 52261
rect 7750 52250 7756 52252
rect 7812 52250 7836 52252
rect 7892 52250 7916 52252
rect 7972 52250 7996 52252
rect 8052 52250 8058 52252
rect 7812 52198 7814 52250
rect 7994 52198 7996 52250
rect 7750 52196 7756 52198
rect 7812 52196 7836 52198
rect 7892 52196 7916 52198
rect 7972 52196 7996 52198
rect 8052 52196 8058 52198
rect 7750 52187 8058 52196
rect 7748 52012 7800 52018
rect 7748 51954 7800 51960
rect 7760 51338 7788 51954
rect 8116 51808 8168 51814
rect 8116 51750 8168 51756
rect 7748 51332 7800 51338
rect 7748 51274 7800 51280
rect 7750 51164 8058 51173
rect 7750 51162 7756 51164
rect 7812 51162 7836 51164
rect 7892 51162 7916 51164
rect 7972 51162 7996 51164
rect 8052 51162 8058 51164
rect 7812 51110 7814 51162
rect 7994 51110 7996 51162
rect 7750 51108 7756 51110
rect 7812 51108 7836 51110
rect 7892 51108 7916 51110
rect 7972 51108 7996 51110
rect 8052 51108 8058 51110
rect 7750 51099 8058 51108
rect 7750 50076 8058 50085
rect 7750 50074 7756 50076
rect 7812 50074 7836 50076
rect 7892 50074 7916 50076
rect 7972 50074 7996 50076
rect 8052 50074 8058 50076
rect 7812 50022 7814 50074
rect 7994 50022 7996 50074
rect 7750 50020 7756 50022
rect 7812 50020 7836 50022
rect 7892 50020 7916 50022
rect 7972 50020 7996 50022
rect 8052 50020 8058 50022
rect 7750 50011 8058 50020
rect 7656 49972 7708 49978
rect 7656 49914 7708 49920
rect 8128 49434 8156 51750
rect 8220 51406 8248 55558
rect 8410 54972 8718 54981
rect 8410 54970 8416 54972
rect 8472 54970 8496 54972
rect 8552 54970 8576 54972
rect 8632 54970 8656 54972
rect 8712 54970 8718 54972
rect 8472 54918 8474 54970
rect 8654 54918 8656 54970
rect 8410 54916 8416 54918
rect 8472 54916 8496 54918
rect 8552 54916 8576 54918
rect 8632 54916 8656 54918
rect 8712 54916 8718 54918
rect 8410 54907 8718 54916
rect 8410 53884 8718 53893
rect 8410 53882 8416 53884
rect 8472 53882 8496 53884
rect 8552 53882 8576 53884
rect 8632 53882 8656 53884
rect 8712 53882 8718 53884
rect 8472 53830 8474 53882
rect 8654 53830 8656 53882
rect 8410 53828 8416 53830
rect 8472 53828 8496 53830
rect 8552 53828 8576 53830
rect 8632 53828 8656 53830
rect 8712 53828 8718 53830
rect 8410 53819 8718 53828
rect 8300 53032 8352 53038
rect 8300 52974 8352 52980
rect 8312 51406 8340 52974
rect 8410 52796 8718 52805
rect 8410 52794 8416 52796
rect 8472 52794 8496 52796
rect 8552 52794 8576 52796
rect 8632 52794 8656 52796
rect 8712 52794 8718 52796
rect 8472 52742 8474 52794
rect 8654 52742 8656 52794
rect 8410 52740 8416 52742
rect 8472 52740 8496 52742
rect 8552 52740 8576 52742
rect 8632 52740 8656 52742
rect 8712 52740 8718 52742
rect 8410 52731 8718 52740
rect 8410 51708 8718 51717
rect 8410 51706 8416 51708
rect 8472 51706 8496 51708
rect 8552 51706 8576 51708
rect 8632 51706 8656 51708
rect 8712 51706 8718 51708
rect 8472 51654 8474 51706
rect 8654 51654 8656 51706
rect 8410 51652 8416 51654
rect 8472 51652 8496 51654
rect 8552 51652 8576 51654
rect 8632 51652 8656 51654
rect 8712 51652 8718 51654
rect 8410 51643 8718 51652
rect 8668 51604 8720 51610
rect 8668 51546 8720 51552
rect 8208 51400 8260 51406
rect 8208 51342 8260 51348
rect 8300 51400 8352 51406
rect 8300 51342 8352 51348
rect 8576 51332 8628 51338
rect 8576 51274 8628 51280
rect 8208 51264 8260 51270
rect 8208 51206 8260 51212
rect 8300 51264 8352 51270
rect 8300 51206 8352 51212
rect 8116 49428 8168 49434
rect 8116 49370 8168 49376
rect 7656 49156 7708 49162
rect 7656 49098 7708 49104
rect 7668 45370 7696 49098
rect 8116 49088 8168 49094
rect 8116 49030 8168 49036
rect 7750 48988 8058 48997
rect 7750 48986 7756 48988
rect 7812 48986 7836 48988
rect 7892 48986 7916 48988
rect 7972 48986 7996 48988
rect 8052 48986 8058 48988
rect 7812 48934 7814 48986
rect 7994 48934 7996 48986
rect 7750 48932 7756 48934
rect 7812 48932 7836 48934
rect 7892 48932 7916 48934
rect 7972 48932 7996 48934
rect 8052 48932 8058 48934
rect 7750 48923 8058 48932
rect 7750 47900 8058 47909
rect 7750 47898 7756 47900
rect 7812 47898 7836 47900
rect 7892 47898 7916 47900
rect 7972 47898 7996 47900
rect 8052 47898 8058 47900
rect 7812 47846 7814 47898
rect 7994 47846 7996 47898
rect 7750 47844 7756 47846
rect 7812 47844 7836 47846
rect 7892 47844 7916 47846
rect 7972 47844 7996 47846
rect 8052 47844 8058 47846
rect 7750 47835 8058 47844
rect 7750 46812 8058 46821
rect 7750 46810 7756 46812
rect 7812 46810 7836 46812
rect 7892 46810 7916 46812
rect 7972 46810 7996 46812
rect 8052 46810 8058 46812
rect 7812 46758 7814 46810
rect 7994 46758 7996 46810
rect 7750 46756 7756 46758
rect 7812 46756 7836 46758
rect 7892 46756 7916 46758
rect 7972 46756 7996 46758
rect 8052 46756 8058 46758
rect 7750 46747 8058 46756
rect 8128 45880 8156 49030
rect 8220 48822 8248 51206
rect 8312 49842 8340 51206
rect 8588 50708 8616 51274
rect 8680 50862 8708 51546
rect 8772 51252 8800 57718
rect 8864 56370 8892 57734
rect 8956 57458 8984 60143
rect 9048 58682 9076 60302
rect 9036 58676 9088 58682
rect 9036 58618 9088 58624
rect 9140 57882 9168 60998
rect 9232 60246 9260 63718
rect 9692 63510 9720 69770
rect 9680 63504 9732 63510
rect 9680 63446 9732 63452
rect 9350 63132 9658 63141
rect 9350 63130 9356 63132
rect 9412 63130 9436 63132
rect 9492 63130 9516 63132
rect 9572 63130 9596 63132
rect 9652 63130 9658 63132
rect 9412 63078 9414 63130
rect 9594 63078 9596 63130
rect 9350 63076 9356 63078
rect 9412 63076 9436 63078
rect 9492 63076 9516 63078
rect 9572 63076 9596 63078
rect 9652 63076 9658 63078
rect 9350 63067 9658 63076
rect 9784 62234 9812 71062
rect 9968 70394 9996 73578
rect 10140 73160 10192 73166
rect 10140 73102 10192 73108
rect 10152 72622 10180 73102
rect 10140 72616 10192 72622
rect 10140 72558 10192 72564
rect 10048 70644 10100 70650
rect 10048 70586 10100 70592
rect 9876 70366 9996 70394
rect 9876 67182 9904 70366
rect 9956 69420 10008 69426
rect 9956 69362 10008 69368
rect 9864 67176 9916 67182
rect 9864 67118 9916 67124
rect 9864 67040 9916 67046
rect 9864 66982 9916 66988
rect 9876 66298 9904 66982
rect 9864 66292 9916 66298
rect 9864 66234 9916 66240
rect 9864 65952 9916 65958
rect 9864 65894 9916 65900
rect 9876 65074 9904 65894
rect 9968 65482 9996 69362
rect 9956 65476 10008 65482
rect 9956 65418 10008 65424
rect 10060 65346 10088 70586
rect 10152 67250 10180 72558
rect 10244 71097 10272 83438
rect 10230 71088 10286 71097
rect 10230 71023 10286 71032
rect 10232 70984 10284 70990
rect 10232 70926 10284 70932
rect 10140 67244 10192 67250
rect 10140 67186 10192 67192
rect 10244 65770 10272 70926
rect 10336 67386 10364 85410
rect 10324 67380 10376 67386
rect 10324 67322 10376 67328
rect 10152 65742 10272 65770
rect 10048 65340 10100 65346
rect 10048 65282 10100 65288
rect 9864 65068 9916 65074
rect 10152 65056 10180 65742
rect 10324 65340 10376 65346
rect 10324 65282 10376 65288
rect 9864 65010 9916 65016
rect 10060 65028 10180 65056
rect 10232 65068 10284 65074
rect 9864 64320 9916 64326
rect 9864 64262 9916 64268
rect 9692 62206 9812 62234
rect 9350 62044 9658 62053
rect 9350 62042 9356 62044
rect 9412 62042 9436 62044
rect 9492 62042 9516 62044
rect 9572 62042 9596 62044
rect 9652 62042 9658 62044
rect 9412 61990 9414 62042
rect 9594 61990 9596 62042
rect 9350 61988 9356 61990
rect 9412 61988 9436 61990
rect 9492 61988 9516 61990
rect 9572 61988 9596 61990
rect 9652 61988 9658 61990
rect 9350 61979 9658 61988
rect 9692 61826 9720 62206
rect 9312 61804 9364 61810
rect 9312 61746 9364 61752
rect 9600 61798 9720 61826
rect 9324 61130 9352 61746
rect 9600 61146 9628 61798
rect 9772 61260 9824 61266
rect 9772 61202 9824 61208
rect 9312 61124 9364 61130
rect 9600 61118 9720 61146
rect 9312 61066 9364 61072
rect 9350 60956 9658 60965
rect 9350 60954 9356 60956
rect 9412 60954 9436 60956
rect 9492 60954 9516 60956
rect 9572 60954 9596 60956
rect 9652 60954 9658 60956
rect 9412 60902 9414 60954
rect 9594 60902 9596 60954
rect 9350 60900 9356 60902
rect 9412 60900 9436 60902
rect 9492 60900 9516 60902
rect 9572 60900 9596 60902
rect 9652 60900 9658 60902
rect 9350 60891 9658 60900
rect 9404 60852 9456 60858
rect 9404 60794 9456 60800
rect 9220 60240 9272 60246
rect 9220 60182 9272 60188
rect 9416 60178 9444 60794
rect 9692 60738 9720 61118
rect 9600 60710 9720 60738
rect 9784 60734 9812 61202
rect 9876 60858 9904 64262
rect 10060 62830 10088 65028
rect 10232 65010 10284 65016
rect 10140 64932 10192 64938
rect 10140 64874 10192 64880
rect 10048 62824 10100 62830
rect 10048 62766 10100 62772
rect 9956 62688 10008 62694
rect 9956 62630 10008 62636
rect 10048 62688 10100 62694
rect 10048 62630 10100 62636
rect 9864 60852 9916 60858
rect 9864 60794 9916 60800
rect 9404 60172 9456 60178
rect 9404 60114 9456 60120
rect 9600 60058 9628 60710
rect 9784 60706 9904 60734
rect 9048 57854 9168 57882
rect 9232 60030 9628 60058
rect 8944 57452 8996 57458
rect 8944 57394 8996 57400
rect 8944 57316 8996 57322
rect 8944 57258 8996 57264
rect 8852 56364 8904 56370
rect 8852 56306 8904 56312
rect 8864 51406 8892 56306
rect 8956 54670 8984 57258
rect 8944 54664 8996 54670
rect 8944 54606 8996 54612
rect 8944 54188 8996 54194
rect 8944 54130 8996 54136
rect 8852 51400 8904 51406
rect 8852 51342 8904 51348
rect 8772 51224 8892 51252
rect 8668 50856 8720 50862
rect 8668 50798 8720 50804
rect 8588 50680 8800 50708
rect 8410 50620 8718 50629
rect 8410 50618 8416 50620
rect 8472 50618 8496 50620
rect 8552 50618 8576 50620
rect 8632 50618 8656 50620
rect 8712 50618 8718 50620
rect 8472 50566 8474 50618
rect 8654 50566 8656 50618
rect 8410 50564 8416 50566
rect 8472 50564 8496 50566
rect 8552 50564 8576 50566
rect 8632 50564 8656 50566
rect 8712 50564 8718 50566
rect 8410 50555 8718 50564
rect 8300 49836 8352 49842
rect 8300 49778 8352 49784
rect 8300 49632 8352 49638
rect 8300 49574 8352 49580
rect 8208 48816 8260 48822
rect 8208 48758 8260 48764
rect 8208 48544 8260 48550
rect 8208 48486 8260 48492
rect 8220 46170 8248 48486
rect 8312 46170 8340 49574
rect 8410 49532 8718 49541
rect 8410 49530 8416 49532
rect 8472 49530 8496 49532
rect 8552 49530 8576 49532
rect 8632 49530 8656 49532
rect 8712 49530 8718 49532
rect 8472 49478 8474 49530
rect 8654 49478 8656 49530
rect 8410 49476 8416 49478
rect 8472 49476 8496 49478
rect 8552 49476 8576 49478
rect 8632 49476 8656 49478
rect 8712 49476 8718 49478
rect 8410 49467 8718 49476
rect 8576 49292 8628 49298
rect 8576 49234 8628 49240
rect 8588 48550 8616 49234
rect 8772 49178 8800 50680
rect 8680 49150 8800 49178
rect 8680 48754 8708 49150
rect 8760 49088 8812 49094
rect 8760 49030 8812 49036
rect 8668 48748 8720 48754
rect 8668 48690 8720 48696
rect 8576 48544 8628 48550
rect 8576 48486 8628 48492
rect 8410 48444 8718 48453
rect 8410 48442 8416 48444
rect 8472 48442 8496 48444
rect 8552 48442 8576 48444
rect 8632 48442 8656 48444
rect 8712 48442 8718 48444
rect 8472 48390 8474 48442
rect 8654 48390 8656 48442
rect 8410 48388 8416 48390
rect 8472 48388 8496 48390
rect 8552 48388 8576 48390
rect 8632 48388 8656 48390
rect 8712 48388 8718 48390
rect 8410 48379 8718 48388
rect 8410 47356 8718 47365
rect 8410 47354 8416 47356
rect 8472 47354 8496 47356
rect 8552 47354 8576 47356
rect 8632 47354 8656 47356
rect 8712 47354 8718 47356
rect 8472 47302 8474 47354
rect 8654 47302 8656 47354
rect 8410 47300 8416 47302
rect 8472 47300 8496 47302
rect 8552 47300 8576 47302
rect 8632 47300 8656 47302
rect 8712 47300 8718 47302
rect 8410 47291 8718 47300
rect 8410 46268 8718 46277
rect 8410 46266 8416 46268
rect 8472 46266 8496 46268
rect 8552 46266 8576 46268
rect 8632 46266 8656 46268
rect 8712 46266 8718 46268
rect 8472 46214 8474 46266
rect 8654 46214 8656 46266
rect 8410 46212 8416 46214
rect 8472 46212 8496 46214
rect 8552 46212 8576 46214
rect 8632 46212 8656 46214
rect 8712 46212 8718 46214
rect 8410 46203 8718 46212
rect 8208 46164 8260 46170
rect 8208 46106 8260 46112
rect 8300 46164 8352 46170
rect 8300 46106 8352 46112
rect 8668 46164 8720 46170
rect 8668 46106 8720 46112
rect 8392 45892 8444 45898
rect 8128 45852 8248 45880
rect 8220 45778 8248 45852
rect 8392 45834 8444 45840
rect 8128 45750 8248 45778
rect 8300 45824 8352 45830
rect 8300 45766 8352 45772
rect 7750 45724 8058 45733
rect 7750 45722 7756 45724
rect 7812 45722 7836 45724
rect 7892 45722 7916 45724
rect 7972 45722 7996 45724
rect 8052 45722 8058 45724
rect 7812 45670 7814 45722
rect 7994 45670 7996 45722
rect 7750 45668 7756 45670
rect 7812 45668 7836 45670
rect 7892 45668 7916 45670
rect 7972 45668 7996 45670
rect 8052 45668 8058 45670
rect 7750 45659 8058 45668
rect 7840 45620 7892 45626
rect 7840 45562 7892 45568
rect 7668 45342 7788 45370
rect 7656 45280 7708 45286
rect 7656 45222 7708 45228
rect 7668 44538 7696 45222
rect 7760 44810 7788 45342
rect 7852 44946 7880 45562
rect 8128 44946 8156 45750
rect 8206 45656 8262 45665
rect 8206 45591 8262 45600
rect 7840 44940 7892 44946
rect 7840 44882 7892 44888
rect 8116 44940 8168 44946
rect 8116 44882 8168 44888
rect 7748 44804 7800 44810
rect 7748 44746 7800 44752
rect 7852 44724 7880 44882
rect 7852 44696 8156 44724
rect 7750 44636 8058 44645
rect 7750 44634 7756 44636
rect 7812 44634 7836 44636
rect 7892 44634 7916 44636
rect 7972 44634 7996 44636
rect 8052 44634 8058 44636
rect 7812 44582 7814 44634
rect 7994 44582 7996 44634
rect 7750 44580 7756 44582
rect 7812 44580 7836 44582
rect 7892 44580 7916 44582
rect 7972 44580 7996 44582
rect 8052 44580 8058 44582
rect 7750 44571 8058 44580
rect 7656 44532 7708 44538
rect 7656 44474 7708 44480
rect 7748 44532 7800 44538
rect 7748 44474 7800 44480
rect 7564 44396 7616 44402
rect 7564 44338 7616 44344
rect 7576 44282 7604 44338
rect 7484 44254 7604 44282
rect 7380 42560 7432 42566
rect 7380 42502 7432 42508
rect 7288 42288 7340 42294
rect 7208 42236 7288 42242
rect 7208 42230 7340 42236
rect 7208 42214 7328 42230
rect 6810 41916 7118 41925
rect 6810 41914 6816 41916
rect 6872 41914 6896 41916
rect 6952 41914 6976 41916
rect 7032 41914 7056 41916
rect 7112 41914 7118 41916
rect 6872 41862 6874 41914
rect 7054 41862 7056 41914
rect 6810 41860 6816 41862
rect 6872 41860 6896 41862
rect 6952 41860 6976 41862
rect 7032 41860 7056 41862
rect 7112 41860 7118 41862
rect 6810 41851 7118 41860
rect 6810 40828 7118 40837
rect 6810 40826 6816 40828
rect 6872 40826 6896 40828
rect 6952 40826 6976 40828
rect 7032 40826 7056 40828
rect 7112 40826 7118 40828
rect 6872 40774 6874 40826
rect 7054 40774 7056 40826
rect 6810 40772 6816 40774
rect 6872 40772 6896 40774
rect 6952 40772 6976 40774
rect 7032 40772 7056 40774
rect 7112 40772 7118 40774
rect 6810 40763 7118 40772
rect 6828 40724 6880 40730
rect 6828 40666 6880 40672
rect 6840 39914 6868 40666
rect 7104 40452 7156 40458
rect 7104 40394 7156 40400
rect 7116 40186 7144 40394
rect 7104 40180 7156 40186
rect 7104 40122 7156 40128
rect 6828 39908 6880 39914
rect 6828 39850 6880 39856
rect 6810 39740 7118 39749
rect 6810 39738 6816 39740
rect 6872 39738 6896 39740
rect 6952 39738 6976 39740
rect 7032 39738 7056 39740
rect 7112 39738 7118 39740
rect 6872 39686 6874 39738
rect 7054 39686 7056 39738
rect 6810 39684 6816 39686
rect 6872 39684 6896 39686
rect 6952 39684 6976 39686
rect 7032 39684 7056 39686
rect 7112 39684 7118 39686
rect 6810 39675 7118 39684
rect 6920 39636 6972 39642
rect 6920 39578 6972 39584
rect 6932 39302 6960 39578
rect 6920 39296 6972 39302
rect 6920 39238 6972 39244
rect 6736 39024 6788 39030
rect 6736 38966 6788 38972
rect 6656 38826 6868 38842
rect 6656 38820 6880 38826
rect 6656 38814 6828 38820
rect 6828 38762 6880 38768
rect 6644 38752 6696 38758
rect 6644 38694 6696 38700
rect 6656 36650 6684 38694
rect 6810 38652 7118 38661
rect 6810 38650 6816 38652
rect 6872 38650 6896 38652
rect 6952 38650 6976 38652
rect 7032 38650 7056 38652
rect 7112 38650 7118 38652
rect 6872 38598 6874 38650
rect 7054 38598 7056 38650
rect 6810 38596 6816 38598
rect 6872 38596 6896 38598
rect 6952 38596 6976 38598
rect 7032 38596 7056 38598
rect 7112 38596 7118 38598
rect 6810 38587 7118 38596
rect 7104 38276 7156 38282
rect 7104 38218 7156 38224
rect 7116 37890 7144 38218
rect 7208 38010 7236 42214
rect 7380 42016 7432 42022
rect 7380 41958 7432 41964
rect 7288 41608 7340 41614
rect 7288 41550 7340 41556
rect 7300 39438 7328 41550
rect 7288 39432 7340 39438
rect 7288 39374 7340 39380
rect 7288 38956 7340 38962
rect 7288 38898 7340 38904
rect 7196 38004 7248 38010
rect 7196 37946 7248 37952
rect 7116 37862 7236 37890
rect 6810 37564 7118 37573
rect 6810 37562 6816 37564
rect 6872 37562 6896 37564
rect 6952 37562 6976 37564
rect 7032 37562 7056 37564
rect 7112 37562 7118 37564
rect 6872 37510 6874 37562
rect 7054 37510 7056 37562
rect 6810 37508 6816 37510
rect 6872 37508 6896 37510
rect 6952 37508 6976 37510
rect 7032 37508 7056 37510
rect 7112 37508 7118 37510
rect 6810 37499 7118 37508
rect 6918 37360 6974 37369
rect 6918 37295 6920 37304
rect 6972 37295 6974 37304
rect 6920 37266 6972 37272
rect 7104 37120 7156 37126
rect 7104 37062 7156 37068
rect 7116 36854 7144 37062
rect 7104 36848 7156 36854
rect 7104 36790 7156 36796
rect 6644 36644 6696 36650
rect 6644 36586 6696 36592
rect 6810 36476 7118 36485
rect 6810 36474 6816 36476
rect 6872 36474 6896 36476
rect 6952 36474 6976 36476
rect 7032 36474 7056 36476
rect 7112 36474 7118 36476
rect 6872 36422 6874 36474
rect 7054 36422 7056 36474
rect 6810 36420 6816 36422
rect 6872 36420 6896 36422
rect 6952 36420 6976 36422
rect 7032 36420 7056 36422
rect 7112 36420 7118 36422
rect 6810 36411 7118 36420
rect 6564 36366 6776 36394
rect 6472 36094 6684 36122
rect 6552 36032 6604 36038
rect 6552 35974 6604 35980
rect 6150 35932 6458 35941
rect 6150 35930 6156 35932
rect 6212 35930 6236 35932
rect 6292 35930 6316 35932
rect 6372 35930 6396 35932
rect 6452 35930 6458 35932
rect 6212 35878 6214 35930
rect 6394 35878 6396 35930
rect 6150 35876 6156 35878
rect 6212 35876 6236 35878
rect 6292 35876 6316 35878
rect 6372 35876 6396 35878
rect 6452 35876 6458 35878
rect 6150 35867 6458 35876
rect 6150 34844 6458 34853
rect 6150 34842 6156 34844
rect 6212 34842 6236 34844
rect 6292 34842 6316 34844
rect 6372 34842 6396 34844
rect 6452 34842 6458 34844
rect 6212 34790 6214 34842
rect 6394 34790 6396 34842
rect 6150 34788 6156 34790
rect 6212 34788 6236 34790
rect 6292 34788 6316 34790
rect 6372 34788 6396 34790
rect 6452 34788 6458 34790
rect 6150 34779 6458 34788
rect 6150 33756 6458 33765
rect 6150 33754 6156 33756
rect 6212 33754 6236 33756
rect 6292 33754 6316 33756
rect 6372 33754 6396 33756
rect 6452 33754 6458 33756
rect 6212 33702 6214 33754
rect 6394 33702 6396 33754
rect 6150 33700 6156 33702
rect 6212 33700 6236 33702
rect 6292 33700 6316 33702
rect 6372 33700 6396 33702
rect 6452 33700 6458 33702
rect 6150 33691 6458 33700
rect 6564 33114 6592 35974
rect 6552 33108 6604 33114
rect 6552 33050 6604 33056
rect 6656 32994 6684 36094
rect 6564 32966 6684 32994
rect 6150 32668 6458 32677
rect 6150 32666 6156 32668
rect 6212 32666 6236 32668
rect 6292 32666 6316 32668
rect 6372 32666 6396 32668
rect 6452 32666 6458 32668
rect 6212 32614 6214 32666
rect 6394 32614 6396 32666
rect 6150 32612 6156 32614
rect 6212 32612 6236 32614
rect 6292 32612 6316 32614
rect 6372 32612 6396 32614
rect 6452 32612 6458 32614
rect 6150 32603 6458 32612
rect 6564 32502 6592 32966
rect 6644 32836 6696 32842
rect 6644 32778 6696 32784
rect 6552 32496 6604 32502
rect 6552 32438 6604 32444
rect 5908 31894 5960 31900
rect 5998 31920 6054 31929
rect 5998 31855 6054 31864
rect 6150 31580 6458 31589
rect 6150 31578 6156 31580
rect 6212 31578 6236 31580
rect 6292 31578 6316 31580
rect 6372 31578 6396 31580
rect 6452 31578 6458 31580
rect 6212 31526 6214 31578
rect 6394 31526 6396 31578
rect 6150 31524 6156 31526
rect 6212 31524 6236 31526
rect 6292 31524 6316 31526
rect 6372 31524 6396 31526
rect 6452 31524 6458 31526
rect 6150 31515 6458 31524
rect 5908 31408 5960 31414
rect 5908 31350 5960 31356
rect 5998 31376 6054 31385
rect 5920 28529 5948 31350
rect 5998 31311 6054 31320
rect 6092 31340 6144 31346
rect 6012 28642 6040 31311
rect 6092 31282 6144 31288
rect 6104 30705 6132 31282
rect 6090 30696 6146 30705
rect 6090 30631 6146 30640
rect 6150 30492 6458 30501
rect 6150 30490 6156 30492
rect 6212 30490 6236 30492
rect 6292 30490 6316 30492
rect 6372 30490 6396 30492
rect 6452 30490 6458 30492
rect 6212 30438 6214 30490
rect 6394 30438 6396 30490
rect 6150 30436 6156 30438
rect 6212 30436 6236 30438
rect 6292 30436 6316 30438
rect 6372 30436 6396 30438
rect 6452 30436 6458 30438
rect 6150 30427 6458 30436
rect 6150 29404 6458 29413
rect 6150 29402 6156 29404
rect 6212 29402 6236 29404
rect 6292 29402 6316 29404
rect 6372 29402 6396 29404
rect 6452 29402 6458 29404
rect 6212 29350 6214 29402
rect 6394 29350 6396 29402
rect 6150 29348 6156 29350
rect 6212 29348 6236 29350
rect 6292 29348 6316 29350
rect 6372 29348 6396 29350
rect 6452 29348 6458 29350
rect 6150 29339 6458 29348
rect 6090 29200 6146 29209
rect 6090 29135 6146 29144
rect 6104 28762 6132 29135
rect 6092 28756 6144 28762
rect 6092 28698 6144 28704
rect 6012 28614 6132 28642
rect 6104 28558 6132 28614
rect 6092 28552 6144 28558
rect 5906 28520 5962 28529
rect 6092 28494 6144 28500
rect 5906 28455 5962 28464
rect 5816 28416 5868 28422
rect 5816 28358 5868 28364
rect 6000 28416 6052 28422
rect 6000 28358 6052 28364
rect 5906 28248 5962 28257
rect 5816 28212 5868 28218
rect 5906 28183 5962 28192
rect 5816 28154 5868 28160
rect 5828 26042 5856 28154
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 5920 25974 5948 28183
rect 6012 26024 6040 28358
rect 6150 28316 6458 28325
rect 6150 28314 6156 28316
rect 6212 28314 6236 28316
rect 6292 28314 6316 28316
rect 6372 28314 6396 28316
rect 6452 28314 6458 28316
rect 6212 28262 6214 28314
rect 6394 28262 6396 28314
rect 6150 28260 6156 28262
rect 6212 28260 6236 28262
rect 6292 28260 6316 28262
rect 6372 28260 6396 28262
rect 6452 28260 6458 28262
rect 6150 28251 6458 28260
rect 6150 27228 6458 27237
rect 6150 27226 6156 27228
rect 6212 27226 6236 27228
rect 6292 27226 6316 27228
rect 6372 27226 6396 27228
rect 6452 27226 6458 27228
rect 6212 27174 6214 27226
rect 6394 27174 6396 27226
rect 6150 27172 6156 27174
rect 6212 27172 6236 27174
rect 6292 27172 6316 27174
rect 6372 27172 6396 27174
rect 6452 27172 6458 27174
rect 6150 27163 6458 27172
rect 6460 26988 6512 26994
rect 6460 26930 6512 26936
rect 6092 26920 6144 26926
rect 6092 26862 6144 26868
rect 6104 26353 6132 26862
rect 6472 26518 6500 26930
rect 6460 26512 6512 26518
rect 6460 26454 6512 26460
rect 6564 26382 6592 32438
rect 6656 26874 6684 32778
rect 6748 29306 6776 36366
rect 7208 36038 7236 37862
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 6810 35388 7118 35397
rect 6810 35386 6816 35388
rect 6872 35386 6896 35388
rect 6952 35386 6976 35388
rect 7032 35386 7056 35388
rect 7112 35386 7118 35388
rect 6872 35334 6874 35386
rect 7054 35334 7056 35386
rect 6810 35332 6816 35334
rect 6872 35332 6896 35334
rect 6952 35332 6976 35334
rect 7032 35332 7056 35334
rect 7112 35332 7118 35334
rect 6810 35323 7118 35332
rect 6810 34300 7118 34309
rect 6810 34298 6816 34300
rect 6872 34298 6896 34300
rect 6952 34298 6976 34300
rect 7032 34298 7056 34300
rect 7112 34298 7118 34300
rect 6872 34246 6874 34298
rect 7054 34246 7056 34298
rect 6810 34244 6816 34246
rect 6872 34244 6896 34246
rect 6952 34244 6976 34246
rect 7032 34244 7056 34246
rect 7112 34244 7118 34246
rect 6810 34235 7118 34244
rect 7208 33930 7236 35770
rect 7196 33924 7248 33930
rect 7196 33866 7248 33872
rect 7300 33810 7328 38898
rect 7392 38010 7420 41958
rect 7484 40186 7512 44254
rect 7760 44180 7788 44474
rect 8128 44402 8156 44696
rect 8220 44538 8248 45591
rect 8208 44532 8260 44538
rect 8208 44474 8260 44480
rect 8116 44396 8168 44402
rect 8116 44338 8168 44344
rect 7576 44152 7788 44180
rect 8116 44192 8168 44198
rect 7576 40662 7604 44152
rect 8116 44134 8168 44140
rect 8208 44192 8260 44198
rect 8208 44134 8260 44140
rect 7750 43548 8058 43557
rect 7750 43546 7756 43548
rect 7812 43546 7836 43548
rect 7892 43546 7916 43548
rect 7972 43546 7996 43548
rect 8052 43546 8058 43548
rect 7812 43494 7814 43546
rect 7994 43494 7996 43546
rect 7750 43492 7756 43494
rect 7812 43492 7836 43494
rect 7892 43492 7916 43494
rect 7972 43492 7996 43494
rect 8052 43492 8058 43494
rect 7750 43483 8058 43492
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 7656 43376 7708 43382
rect 7656 43318 7708 43324
rect 7668 41614 7696 43318
rect 7760 42770 7788 43386
rect 8128 43194 8156 44134
rect 8220 43994 8248 44134
rect 8208 43988 8260 43994
rect 8208 43930 8260 43936
rect 8220 43450 8248 43930
rect 8208 43444 8260 43450
rect 8208 43386 8260 43392
rect 8128 43166 8248 43194
rect 8116 43104 8168 43110
rect 8116 43046 8168 43052
rect 7748 42764 7800 42770
rect 7748 42706 7800 42712
rect 7760 42566 7788 42706
rect 7748 42560 7800 42566
rect 7748 42502 7800 42508
rect 7750 42460 8058 42469
rect 7750 42458 7756 42460
rect 7812 42458 7836 42460
rect 7892 42458 7916 42460
rect 7972 42458 7996 42460
rect 8052 42458 8058 42460
rect 7812 42406 7814 42458
rect 7994 42406 7996 42458
rect 7750 42404 7756 42406
rect 7812 42404 7836 42406
rect 7892 42404 7916 42406
rect 7972 42404 7996 42406
rect 8052 42404 8058 42406
rect 7750 42395 8058 42404
rect 7748 42356 7800 42362
rect 7748 42298 7800 42304
rect 7656 41608 7708 41614
rect 7656 41550 7708 41556
rect 7760 41460 7788 42298
rect 7668 41432 7788 41460
rect 7564 40656 7616 40662
rect 7564 40598 7616 40604
rect 7564 40520 7616 40526
rect 7564 40462 7616 40468
rect 7472 40180 7524 40186
rect 7472 40122 7524 40128
rect 7472 39976 7524 39982
rect 7472 39918 7524 39924
rect 7484 39574 7512 39918
rect 7472 39568 7524 39574
rect 7472 39510 7524 39516
rect 7380 38004 7432 38010
rect 7380 37946 7432 37952
rect 7484 37806 7512 39510
rect 7576 39506 7604 40462
rect 7668 40118 7696 41432
rect 7750 41372 8058 41381
rect 7750 41370 7756 41372
rect 7812 41370 7836 41372
rect 7892 41370 7916 41372
rect 7972 41370 7996 41372
rect 8052 41370 8058 41372
rect 7812 41318 7814 41370
rect 7994 41318 7996 41370
rect 7750 41316 7756 41318
rect 7812 41316 7836 41318
rect 7892 41316 7916 41318
rect 7972 41316 7996 41318
rect 8052 41316 8058 41318
rect 7750 41307 8058 41316
rect 8128 41256 8156 43046
rect 8036 41228 8156 41256
rect 8036 40662 8064 41228
rect 8220 41154 8248 43166
rect 8312 42702 8340 45766
rect 8404 45626 8432 45834
rect 8392 45620 8444 45626
rect 8392 45562 8444 45568
rect 8680 45268 8708 46106
rect 8772 45490 8800 49030
rect 8864 47122 8892 51224
rect 8956 48634 8984 54130
rect 9048 49042 9076 57854
rect 9128 57792 9180 57798
rect 9128 57734 9180 57740
rect 9140 49298 9168 57734
rect 9232 56846 9260 60030
rect 9350 59868 9658 59877
rect 9350 59866 9356 59868
rect 9412 59866 9436 59868
rect 9492 59866 9516 59868
rect 9572 59866 9596 59868
rect 9652 59866 9658 59868
rect 9412 59814 9414 59866
rect 9594 59814 9596 59866
rect 9350 59812 9356 59814
rect 9412 59812 9436 59814
rect 9492 59812 9516 59814
rect 9572 59812 9596 59814
rect 9652 59812 9658 59814
rect 9350 59803 9658 59812
rect 9876 59650 9904 60706
rect 9600 59622 9904 59650
rect 9600 59022 9628 59622
rect 9588 59016 9640 59022
rect 9588 58958 9640 58964
rect 9350 58780 9658 58789
rect 9350 58778 9356 58780
rect 9412 58778 9436 58780
rect 9492 58778 9516 58780
rect 9572 58778 9596 58780
rect 9652 58778 9658 58780
rect 9412 58726 9414 58778
rect 9594 58726 9596 58778
rect 9350 58724 9356 58726
rect 9412 58724 9436 58726
rect 9492 58724 9516 58726
rect 9572 58724 9596 58726
rect 9652 58724 9658 58726
rect 9350 58715 9658 58724
rect 9312 58676 9364 58682
rect 9312 58618 9364 58624
rect 9324 57905 9352 58618
rect 9968 57974 9996 62630
rect 9876 57946 9996 57974
rect 9310 57896 9366 57905
rect 9310 57831 9366 57840
rect 9350 57692 9658 57701
rect 9350 57690 9356 57692
rect 9412 57690 9436 57692
rect 9492 57690 9516 57692
rect 9572 57690 9596 57692
rect 9652 57690 9658 57692
rect 9412 57638 9414 57690
rect 9594 57638 9596 57690
rect 9350 57636 9356 57638
rect 9412 57636 9436 57638
rect 9492 57636 9516 57638
rect 9572 57636 9596 57638
rect 9652 57636 9658 57638
rect 9350 57627 9658 57636
rect 9220 56840 9272 56846
rect 9220 56782 9272 56788
rect 9350 56604 9658 56613
rect 9350 56602 9356 56604
rect 9412 56602 9436 56604
rect 9492 56602 9516 56604
rect 9572 56602 9596 56604
rect 9652 56602 9658 56604
rect 9412 56550 9414 56602
rect 9594 56550 9596 56602
rect 9350 56548 9356 56550
rect 9412 56548 9436 56550
rect 9492 56548 9516 56550
rect 9572 56548 9596 56550
rect 9652 56548 9658 56550
rect 9350 56539 9658 56548
rect 9680 55888 9732 55894
rect 9680 55830 9732 55836
rect 9350 55516 9658 55525
rect 9350 55514 9356 55516
rect 9412 55514 9436 55516
rect 9492 55514 9516 55516
rect 9572 55514 9596 55516
rect 9652 55514 9658 55516
rect 9412 55462 9414 55514
rect 9594 55462 9596 55514
rect 9350 55460 9356 55462
rect 9412 55460 9436 55462
rect 9492 55460 9516 55462
rect 9572 55460 9596 55462
rect 9652 55460 9658 55462
rect 9350 55451 9658 55460
rect 9692 55282 9720 55830
rect 9876 55434 9904 57946
rect 9876 55406 9996 55434
rect 9680 55276 9732 55282
rect 9680 55218 9732 55224
rect 9864 55276 9916 55282
rect 9864 55218 9916 55224
rect 9220 54596 9272 54602
rect 9220 54538 9272 54544
rect 9232 51388 9260 54538
rect 9350 54428 9658 54437
rect 9350 54426 9356 54428
rect 9412 54426 9436 54428
rect 9492 54426 9516 54428
rect 9572 54426 9596 54428
rect 9652 54426 9658 54428
rect 9412 54374 9414 54426
rect 9594 54374 9596 54426
rect 9350 54372 9356 54374
rect 9412 54372 9436 54374
rect 9492 54372 9516 54374
rect 9572 54372 9596 54374
rect 9652 54372 9658 54374
rect 9350 54363 9658 54372
rect 9680 54324 9732 54330
rect 9680 54266 9732 54272
rect 9350 53340 9658 53349
rect 9350 53338 9356 53340
rect 9412 53338 9436 53340
rect 9492 53338 9516 53340
rect 9572 53338 9596 53340
rect 9652 53338 9658 53340
rect 9412 53286 9414 53338
rect 9594 53286 9596 53338
rect 9350 53284 9356 53286
rect 9412 53284 9436 53286
rect 9492 53284 9516 53286
rect 9572 53284 9596 53286
rect 9652 53284 9658 53286
rect 9350 53275 9658 53284
rect 9692 53122 9720 54266
rect 9600 53094 9720 53122
rect 9772 53168 9824 53174
rect 9772 53110 9824 53116
rect 9600 52442 9628 53094
rect 9600 52414 9720 52442
rect 9350 52252 9658 52261
rect 9350 52250 9356 52252
rect 9412 52250 9436 52252
rect 9492 52250 9516 52252
rect 9572 52250 9596 52252
rect 9652 52250 9658 52252
rect 9412 52198 9414 52250
rect 9594 52198 9596 52250
rect 9350 52196 9356 52198
rect 9412 52196 9436 52198
rect 9492 52196 9516 52198
rect 9572 52196 9596 52198
rect 9652 52196 9658 52198
rect 9350 52187 9658 52196
rect 9692 52034 9720 52414
rect 9600 52006 9720 52034
rect 9600 51610 9628 52006
rect 9588 51604 9640 51610
rect 9588 51546 9640 51552
rect 9232 51360 9628 51388
rect 9600 51354 9628 51360
rect 9600 51326 9720 51354
rect 9220 51264 9272 51270
rect 9220 51206 9272 51212
rect 9232 49434 9260 51206
rect 9350 51164 9658 51173
rect 9350 51162 9356 51164
rect 9412 51162 9436 51164
rect 9492 51162 9516 51164
rect 9572 51162 9596 51164
rect 9652 51162 9658 51164
rect 9412 51110 9414 51162
rect 9594 51110 9596 51162
rect 9350 51108 9356 51110
rect 9412 51108 9436 51110
rect 9492 51108 9516 51110
rect 9572 51108 9596 51110
rect 9652 51108 9658 51110
rect 9350 51099 9658 51108
rect 9692 51048 9720 51326
rect 9508 51020 9720 51048
rect 9508 50289 9536 51020
rect 9588 50856 9640 50862
rect 9588 50798 9640 50804
rect 9494 50280 9550 50289
rect 9600 50266 9628 50798
rect 9600 50238 9720 50266
rect 9494 50215 9550 50224
rect 9350 50076 9658 50085
rect 9350 50074 9356 50076
rect 9412 50074 9436 50076
rect 9492 50074 9516 50076
rect 9572 50074 9596 50076
rect 9652 50074 9658 50076
rect 9412 50022 9414 50074
rect 9594 50022 9596 50074
rect 9350 50020 9356 50022
rect 9412 50020 9436 50022
rect 9492 50020 9516 50022
rect 9572 50020 9596 50022
rect 9652 50020 9658 50022
rect 9350 50011 9658 50020
rect 9692 49892 9720 50238
rect 9600 49864 9720 49892
rect 9220 49428 9272 49434
rect 9220 49370 9272 49376
rect 9128 49292 9180 49298
rect 9128 49234 9180 49240
rect 9600 49178 9628 49864
rect 9600 49150 9720 49178
rect 9048 49014 9260 49042
rect 9128 48748 9180 48754
rect 9128 48690 9180 48696
rect 8956 48606 9076 48634
rect 8944 48544 8996 48550
rect 8944 48486 8996 48492
rect 8852 47116 8904 47122
rect 8852 47058 8904 47064
rect 8852 46912 8904 46918
rect 8852 46854 8904 46860
rect 8760 45484 8812 45490
rect 8760 45426 8812 45432
rect 8680 45240 8800 45268
rect 8410 45180 8718 45189
rect 8410 45178 8416 45180
rect 8472 45178 8496 45180
rect 8552 45178 8576 45180
rect 8632 45178 8656 45180
rect 8712 45178 8718 45180
rect 8472 45126 8474 45178
rect 8654 45126 8656 45178
rect 8410 45124 8416 45126
rect 8472 45124 8496 45126
rect 8552 45124 8576 45126
rect 8632 45124 8656 45126
rect 8712 45124 8718 45126
rect 8410 45115 8718 45124
rect 8410 44092 8718 44101
rect 8410 44090 8416 44092
rect 8472 44090 8496 44092
rect 8552 44090 8576 44092
rect 8632 44090 8656 44092
rect 8712 44090 8718 44092
rect 8472 44038 8474 44090
rect 8654 44038 8656 44090
rect 8410 44036 8416 44038
rect 8472 44036 8496 44038
rect 8552 44036 8576 44038
rect 8632 44036 8656 44038
rect 8712 44036 8718 44038
rect 8410 44027 8718 44036
rect 8772 43874 8800 45240
rect 8680 43846 8800 43874
rect 8680 43382 8708 43846
rect 8760 43784 8812 43790
rect 8760 43726 8812 43732
rect 8668 43376 8720 43382
rect 8668 43318 8720 43324
rect 8410 43004 8718 43013
rect 8410 43002 8416 43004
rect 8472 43002 8496 43004
rect 8552 43002 8576 43004
rect 8632 43002 8656 43004
rect 8712 43002 8718 43004
rect 8472 42950 8474 43002
rect 8654 42950 8656 43002
rect 8410 42948 8416 42950
rect 8472 42948 8496 42950
rect 8552 42948 8576 42950
rect 8632 42948 8656 42950
rect 8712 42948 8718 42950
rect 8410 42939 8718 42948
rect 8668 42832 8720 42838
rect 8668 42774 8720 42780
rect 8300 42696 8352 42702
rect 8300 42638 8352 42644
rect 8576 42696 8628 42702
rect 8576 42638 8628 42644
rect 8300 42560 8352 42566
rect 8300 42502 8352 42508
rect 8128 41126 8248 41154
rect 8024 40656 8076 40662
rect 8024 40598 8076 40604
rect 7750 40284 8058 40293
rect 7750 40282 7756 40284
rect 7812 40282 7836 40284
rect 7892 40282 7916 40284
rect 7972 40282 7996 40284
rect 8052 40282 8058 40284
rect 7812 40230 7814 40282
rect 7994 40230 7996 40282
rect 7750 40228 7756 40230
rect 7812 40228 7836 40230
rect 7892 40228 7916 40230
rect 7972 40228 7996 40230
rect 8052 40228 8058 40230
rect 7750 40219 8058 40228
rect 7656 40112 7708 40118
rect 7656 40054 7708 40060
rect 8128 39982 8156 41126
rect 8312 40712 8340 42502
rect 8588 42022 8616 42638
rect 8680 42378 8708 42774
rect 8772 42548 8800 43726
rect 8864 42702 8892 46854
rect 8956 46170 8984 48486
rect 9048 47530 9076 48606
rect 9036 47524 9088 47530
rect 9036 47466 9088 47472
rect 9036 47116 9088 47122
rect 9036 47058 9088 47064
rect 8944 46164 8996 46170
rect 8944 46106 8996 46112
rect 8944 45824 8996 45830
rect 8944 45766 8996 45772
rect 8852 42696 8904 42702
rect 8956 42673 8984 45766
rect 9048 43790 9076 47058
rect 9140 45558 9168 48690
rect 9232 47122 9260 49014
rect 9350 48988 9658 48997
rect 9350 48986 9356 48988
rect 9412 48986 9436 48988
rect 9492 48986 9516 48988
rect 9572 48986 9596 48988
rect 9652 48986 9658 48988
rect 9412 48934 9414 48986
rect 9594 48934 9596 48986
rect 9350 48932 9356 48934
rect 9412 48932 9436 48934
rect 9492 48932 9516 48934
rect 9572 48932 9596 48934
rect 9652 48932 9658 48934
rect 9350 48923 9658 48932
rect 9310 48784 9366 48793
rect 9692 48770 9720 49150
rect 9310 48719 9366 48728
rect 9600 48742 9720 48770
rect 9324 48113 9352 48719
rect 9310 48104 9366 48113
rect 9600 48090 9628 48742
rect 9600 48062 9720 48090
rect 9310 48039 9366 48048
rect 9350 47900 9658 47909
rect 9350 47898 9356 47900
rect 9412 47898 9436 47900
rect 9492 47898 9516 47900
rect 9572 47898 9596 47900
rect 9652 47898 9658 47900
rect 9412 47846 9414 47898
rect 9594 47846 9596 47898
rect 9350 47844 9356 47846
rect 9412 47844 9436 47846
rect 9492 47844 9516 47846
rect 9572 47844 9596 47846
rect 9652 47844 9658 47846
rect 9350 47835 9658 47844
rect 9692 47716 9720 48062
rect 9600 47688 9720 47716
rect 9312 47524 9364 47530
rect 9312 47466 9364 47472
rect 9220 47116 9272 47122
rect 9220 47058 9272 47064
rect 9324 47002 9352 47466
rect 9232 46974 9352 47002
rect 9600 47002 9628 47688
rect 9600 46974 9720 47002
rect 9128 45552 9180 45558
rect 9128 45494 9180 45500
rect 9128 45348 9180 45354
rect 9128 45290 9180 45296
rect 9036 43784 9088 43790
rect 9036 43726 9088 43732
rect 9036 43648 9088 43654
rect 9036 43590 9088 43596
rect 8852 42638 8904 42644
rect 8942 42664 8998 42673
rect 8942 42599 8998 42608
rect 8772 42520 8984 42548
rect 8680 42350 8800 42378
rect 8576 42016 8628 42022
rect 8576 41958 8628 41964
rect 8410 41916 8718 41925
rect 8410 41914 8416 41916
rect 8472 41914 8496 41916
rect 8552 41914 8576 41916
rect 8632 41914 8656 41916
rect 8712 41914 8718 41916
rect 8472 41862 8474 41914
rect 8654 41862 8656 41914
rect 8410 41860 8416 41862
rect 8472 41860 8496 41862
rect 8552 41860 8576 41862
rect 8632 41860 8656 41862
rect 8712 41860 8718 41862
rect 8410 41851 8718 41860
rect 8410 40828 8718 40837
rect 8410 40826 8416 40828
rect 8472 40826 8496 40828
rect 8552 40826 8576 40828
rect 8632 40826 8656 40828
rect 8712 40826 8718 40828
rect 8472 40774 8474 40826
rect 8654 40774 8656 40826
rect 8410 40772 8416 40774
rect 8472 40772 8496 40774
rect 8552 40772 8576 40774
rect 8632 40772 8656 40774
rect 8712 40772 8718 40774
rect 8410 40763 8718 40772
rect 8220 40684 8340 40712
rect 8220 40066 8248 40684
rect 8392 40384 8444 40390
rect 8392 40326 8444 40332
rect 8220 40038 8340 40066
rect 8312 39982 8340 40038
rect 8024 39976 8076 39982
rect 7838 39944 7894 39953
rect 8024 39918 8076 39924
rect 8116 39976 8168 39982
rect 8116 39918 8168 39924
rect 8300 39976 8352 39982
rect 8300 39918 8352 39924
rect 7838 39879 7894 39888
rect 7852 39506 7880 39879
rect 8036 39828 8064 39918
rect 8404 39828 8432 40326
rect 8036 39800 8156 39828
rect 7564 39500 7616 39506
rect 7564 39442 7616 39448
rect 7656 39500 7708 39506
rect 7656 39442 7708 39448
rect 7840 39500 7892 39506
rect 7840 39442 7892 39448
rect 7564 39296 7616 39302
rect 7564 39238 7616 39244
rect 7472 37800 7524 37806
rect 7472 37742 7524 37748
rect 7472 37664 7524 37670
rect 7472 37606 7524 37612
rect 7380 37460 7432 37466
rect 7380 37402 7432 37408
rect 7392 37126 7420 37402
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 7208 33782 7328 33810
rect 6810 33212 7118 33221
rect 6810 33210 6816 33212
rect 6872 33210 6896 33212
rect 6952 33210 6976 33212
rect 7032 33210 7056 33212
rect 7112 33210 7118 33212
rect 6872 33158 6874 33210
rect 7054 33158 7056 33210
rect 6810 33156 6816 33158
rect 6872 33156 6896 33158
rect 6952 33156 6976 33158
rect 7032 33156 7056 33158
rect 7112 33156 7118 33158
rect 6810 33147 7118 33156
rect 7104 33108 7156 33114
rect 7104 33050 7156 33056
rect 7116 32314 7144 33050
rect 7208 32434 7236 33782
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7300 32337 7328 33390
rect 7286 32328 7342 32337
rect 7116 32286 7236 32314
rect 6810 32124 7118 32133
rect 6810 32122 6816 32124
rect 6872 32122 6896 32124
rect 6952 32122 6976 32124
rect 7032 32122 7056 32124
rect 7112 32122 7118 32124
rect 6872 32070 6874 32122
rect 7054 32070 7056 32122
rect 6810 32068 6816 32070
rect 6872 32068 6896 32070
rect 6952 32068 6976 32070
rect 7032 32068 7056 32070
rect 7112 32068 7118 32070
rect 6810 32059 7118 32068
rect 7010 31920 7066 31929
rect 7010 31855 7066 31864
rect 7024 31414 7052 31855
rect 7208 31822 7236 32286
rect 7286 32263 7342 32272
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 7300 31464 7328 32166
rect 7392 31482 7420 37062
rect 7484 33318 7512 37606
rect 7472 33312 7524 33318
rect 7472 33254 7524 33260
rect 7484 32434 7512 33254
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7472 31952 7524 31958
rect 7472 31894 7524 31900
rect 7116 31436 7328 31464
rect 7380 31476 7432 31482
rect 7012 31408 7064 31414
rect 7012 31350 7064 31356
rect 7116 31124 7144 31436
rect 7380 31418 7432 31424
rect 7484 31226 7512 31894
rect 7576 31754 7604 39238
rect 7668 38894 7696 39442
rect 7750 39196 8058 39205
rect 7750 39194 7756 39196
rect 7812 39194 7836 39196
rect 7892 39194 7916 39196
rect 7972 39194 7996 39196
rect 8052 39194 8058 39196
rect 7812 39142 7814 39194
rect 7994 39142 7996 39194
rect 7750 39140 7756 39142
rect 7812 39140 7836 39142
rect 7892 39140 7916 39142
rect 7972 39140 7996 39142
rect 8052 39140 8058 39142
rect 7750 39131 8058 39140
rect 7656 38888 7708 38894
rect 7656 38830 7708 38836
rect 7668 38282 7696 38830
rect 7656 38276 7708 38282
rect 7656 38218 7708 38224
rect 7668 37176 7696 38218
rect 8128 38214 8156 39800
rect 8312 39800 8432 39828
rect 8206 38448 8262 38457
rect 8206 38383 8262 38392
rect 8116 38208 8168 38214
rect 8116 38150 8168 38156
rect 7750 38108 8058 38117
rect 7750 38106 7756 38108
rect 7812 38106 7836 38108
rect 7892 38106 7916 38108
rect 7972 38106 7996 38108
rect 8052 38106 8058 38108
rect 7812 38054 7814 38106
rect 7994 38054 7996 38106
rect 7750 38052 7756 38054
rect 7812 38052 7836 38054
rect 7892 38052 7916 38054
rect 7972 38052 7996 38054
rect 8052 38052 8058 38054
rect 7750 38043 8058 38052
rect 8220 38010 8248 38383
rect 8208 38004 8260 38010
rect 8208 37946 8260 37952
rect 8116 37800 8168 37806
rect 8116 37742 8168 37748
rect 7748 37324 7800 37330
rect 7748 37266 7800 37272
rect 7760 37176 7788 37266
rect 7668 37148 7788 37176
rect 7668 36038 7696 37148
rect 7750 37020 8058 37029
rect 7750 37018 7756 37020
rect 7812 37018 7836 37020
rect 7892 37018 7916 37020
rect 7972 37018 7996 37020
rect 8052 37018 8058 37020
rect 7812 36966 7814 37018
rect 7994 36966 7996 37018
rect 7750 36964 7756 36966
rect 7812 36964 7836 36966
rect 7892 36964 7916 36966
rect 7972 36964 7996 36966
rect 8052 36964 8058 36966
rect 7750 36955 8058 36964
rect 7656 36032 7708 36038
rect 7656 35974 7708 35980
rect 7668 31958 7696 35974
rect 7750 35932 8058 35941
rect 7750 35930 7756 35932
rect 7812 35930 7836 35932
rect 7892 35930 7916 35932
rect 7972 35930 7996 35932
rect 8052 35930 8058 35932
rect 7812 35878 7814 35930
rect 7994 35878 7996 35930
rect 7750 35876 7756 35878
rect 7812 35876 7836 35878
rect 7892 35876 7916 35878
rect 7972 35876 7996 35878
rect 8052 35876 8058 35878
rect 7750 35867 8058 35876
rect 7750 34844 8058 34853
rect 7750 34842 7756 34844
rect 7812 34842 7836 34844
rect 7892 34842 7916 34844
rect 7972 34842 7996 34844
rect 8052 34842 8058 34844
rect 7812 34790 7814 34842
rect 7994 34790 7996 34842
rect 7750 34788 7756 34790
rect 7812 34788 7836 34790
rect 7892 34788 7916 34790
rect 7972 34788 7996 34790
rect 8052 34788 8058 34790
rect 7750 34779 8058 34788
rect 7750 33756 8058 33765
rect 7750 33754 7756 33756
rect 7812 33754 7836 33756
rect 7892 33754 7916 33756
rect 7972 33754 7996 33756
rect 8052 33754 8058 33756
rect 7812 33702 7814 33754
rect 7994 33702 7996 33754
rect 7750 33700 7756 33702
rect 7812 33700 7836 33702
rect 7892 33700 7916 33702
rect 7972 33700 7996 33702
rect 8052 33700 8058 33702
rect 7750 33691 8058 33700
rect 8128 33590 8156 37742
rect 8312 37210 8340 39800
rect 8410 39740 8718 39749
rect 8410 39738 8416 39740
rect 8472 39738 8496 39740
rect 8552 39738 8576 39740
rect 8632 39738 8656 39740
rect 8712 39738 8718 39740
rect 8472 39686 8474 39738
rect 8654 39686 8656 39738
rect 8410 39684 8416 39686
rect 8472 39684 8496 39686
rect 8552 39684 8576 39686
rect 8632 39684 8656 39686
rect 8712 39684 8718 39686
rect 8410 39675 8718 39684
rect 8410 38652 8718 38661
rect 8410 38650 8416 38652
rect 8472 38650 8496 38652
rect 8552 38650 8576 38652
rect 8632 38650 8656 38652
rect 8712 38650 8718 38652
rect 8472 38598 8474 38650
rect 8654 38598 8656 38650
rect 8410 38596 8416 38598
rect 8472 38596 8496 38598
rect 8552 38596 8576 38598
rect 8632 38596 8656 38598
rect 8712 38596 8718 38598
rect 8410 38587 8718 38596
rect 8410 37564 8718 37573
rect 8410 37562 8416 37564
rect 8472 37562 8496 37564
rect 8552 37562 8576 37564
rect 8632 37562 8656 37564
rect 8712 37562 8718 37564
rect 8472 37510 8474 37562
rect 8654 37510 8656 37562
rect 8410 37508 8416 37510
rect 8472 37508 8496 37510
rect 8552 37508 8576 37510
rect 8632 37508 8656 37510
rect 8712 37508 8718 37510
rect 8410 37499 8718 37508
rect 8312 37182 8432 37210
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8312 36825 8340 36858
rect 8298 36816 8354 36825
rect 8298 36751 8354 36760
rect 8404 36666 8432 37182
rect 8312 36638 8432 36666
rect 8312 35850 8340 36638
rect 8410 36476 8718 36485
rect 8410 36474 8416 36476
rect 8472 36474 8496 36476
rect 8552 36474 8576 36476
rect 8632 36474 8656 36476
rect 8712 36474 8718 36476
rect 8472 36422 8474 36474
rect 8654 36422 8656 36474
rect 8410 36420 8416 36422
rect 8472 36420 8496 36422
rect 8552 36420 8576 36422
rect 8632 36420 8656 36422
rect 8712 36420 8718 36422
rect 8410 36411 8718 36420
rect 8220 35822 8340 35850
rect 8220 35034 8248 35822
rect 8300 35760 8352 35766
rect 8300 35702 8352 35708
rect 8312 35193 8340 35702
rect 8410 35388 8718 35397
rect 8410 35386 8416 35388
rect 8472 35386 8496 35388
rect 8552 35386 8576 35388
rect 8632 35386 8656 35388
rect 8712 35386 8718 35388
rect 8472 35334 8474 35386
rect 8654 35334 8656 35386
rect 8410 35332 8416 35334
rect 8472 35332 8496 35334
rect 8552 35332 8576 35334
rect 8632 35332 8656 35334
rect 8712 35332 8718 35334
rect 8410 35323 8718 35332
rect 8298 35184 8354 35193
rect 8298 35119 8354 35128
rect 8220 35006 8340 35034
rect 8116 33584 8168 33590
rect 8312 33538 8340 35006
rect 8410 34300 8718 34309
rect 8410 34298 8416 34300
rect 8472 34298 8496 34300
rect 8552 34298 8576 34300
rect 8632 34298 8656 34300
rect 8712 34298 8718 34300
rect 8472 34246 8474 34298
rect 8654 34246 8656 34298
rect 8410 34244 8416 34246
rect 8472 34244 8496 34246
rect 8552 34244 8576 34246
rect 8632 34244 8656 34246
rect 8712 34244 8718 34246
rect 8410 34235 8718 34244
rect 8576 34060 8628 34066
rect 8576 34002 8628 34008
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8116 33526 8168 33532
rect 8220 33510 8340 33538
rect 8392 33516 8444 33522
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 7750 32668 8058 32677
rect 7750 32666 7756 32668
rect 7812 32666 7836 32668
rect 7892 32666 7916 32668
rect 7972 32666 7996 32668
rect 8052 32666 8058 32668
rect 7812 32614 7814 32666
rect 7994 32614 7996 32666
rect 7750 32612 7756 32614
rect 7812 32612 7836 32614
rect 7892 32612 7916 32614
rect 7972 32612 7996 32614
rect 8052 32612 8058 32614
rect 7750 32603 8058 32612
rect 8024 32496 8076 32502
rect 8024 32438 8076 32444
rect 7748 32360 7800 32366
rect 7748 32302 7800 32308
rect 7656 31952 7708 31958
rect 7656 31894 7708 31900
rect 7760 31890 7788 32302
rect 7840 32224 7892 32230
rect 7840 32166 7892 32172
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 7576 31726 7696 31754
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7576 31346 7604 31622
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7380 31204 7432 31210
rect 7484 31198 7604 31226
rect 7380 31146 7432 31152
rect 7116 31096 7236 31124
rect 6810 31036 7118 31045
rect 6810 31034 6816 31036
rect 6872 31034 6896 31036
rect 6952 31034 6976 31036
rect 7032 31034 7056 31036
rect 7112 31034 7118 31036
rect 6872 30982 6874 31034
rect 7054 30982 7056 31034
rect 6810 30980 6816 30982
rect 6872 30980 6896 30982
rect 6952 30980 6976 30982
rect 7032 30980 7056 30982
rect 7112 30980 7118 30982
rect 6810 30971 7118 30980
rect 6810 29948 7118 29957
rect 6810 29946 6816 29948
rect 6872 29946 6896 29948
rect 6952 29946 6976 29948
rect 7032 29946 7056 29948
rect 7112 29946 7118 29948
rect 6872 29894 6874 29946
rect 7054 29894 7056 29946
rect 6810 29892 6816 29894
rect 6872 29892 6896 29894
rect 6952 29892 6976 29894
rect 7032 29892 7056 29894
rect 7112 29892 7118 29894
rect 6810 29883 7118 29892
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6840 28966 6868 29650
rect 6828 28960 6880 28966
rect 6828 28902 6880 28908
rect 6810 28860 7118 28869
rect 6810 28858 6816 28860
rect 6872 28858 6896 28860
rect 6952 28858 6976 28860
rect 7032 28858 7056 28860
rect 7112 28858 7118 28860
rect 6872 28806 6874 28858
rect 7054 28806 7056 28858
rect 6810 28804 6816 28806
rect 6872 28804 6896 28806
rect 6952 28804 6976 28806
rect 7032 28804 7056 28806
rect 7112 28804 7118 28806
rect 6810 28795 7118 28804
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6840 28370 6868 28494
rect 6748 28342 6868 28370
rect 6748 27554 6776 28342
rect 7024 27985 7052 28698
rect 7208 28694 7236 31096
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7300 29170 7328 30194
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7196 28688 7248 28694
rect 7196 28630 7248 28636
rect 7196 28416 7248 28422
rect 7196 28358 7248 28364
rect 7010 27976 7066 27985
rect 7010 27911 7066 27920
rect 6810 27772 7118 27781
rect 6810 27770 6816 27772
rect 6872 27770 6896 27772
rect 6952 27770 6976 27772
rect 7032 27770 7056 27772
rect 7112 27770 7118 27772
rect 6872 27718 6874 27770
rect 7054 27718 7056 27770
rect 6810 27716 6816 27718
rect 6872 27716 6896 27718
rect 6952 27716 6976 27718
rect 7032 27716 7056 27718
rect 7112 27716 7118 27718
rect 6810 27707 7118 27716
rect 7208 27656 7236 28358
rect 7116 27628 7236 27656
rect 6748 27526 6868 27554
rect 6656 26846 6776 26874
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6552 26376 6604 26382
rect 6090 26344 6146 26353
rect 6552 26318 6604 26324
rect 6090 26279 6146 26288
rect 6656 26194 6684 26726
rect 6564 26166 6684 26194
rect 6150 26140 6458 26149
rect 6150 26138 6156 26140
rect 6212 26138 6236 26140
rect 6292 26138 6316 26140
rect 6372 26138 6396 26140
rect 6452 26138 6458 26140
rect 6212 26086 6214 26138
rect 6394 26086 6396 26138
rect 6150 26084 6156 26086
rect 6212 26084 6236 26086
rect 6292 26084 6316 26086
rect 6372 26084 6396 26086
rect 6452 26084 6458 26086
rect 6150 26075 6458 26084
rect 6012 25996 6132 26024
rect 5908 25968 5960 25974
rect 5814 25936 5870 25945
rect 5908 25910 5960 25916
rect 5814 25871 5816 25880
rect 5868 25871 5870 25880
rect 5816 25842 5868 25848
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5828 24138 5856 25842
rect 5908 25832 5960 25838
rect 6104 25820 6132 25996
rect 6184 25900 6236 25906
rect 6184 25842 6236 25848
rect 5908 25774 5960 25780
rect 6012 25792 6132 25820
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5724 24064 5776 24070
rect 5724 24006 5776 24012
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5736 21554 5764 24006
rect 5816 23248 5868 23254
rect 5816 23190 5868 23196
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5210 10364 5518 10373
rect 5210 10362 5216 10364
rect 5272 10362 5296 10364
rect 5352 10362 5376 10364
rect 5432 10362 5456 10364
rect 5512 10362 5518 10364
rect 5272 10310 5274 10362
rect 5454 10310 5456 10362
rect 5210 10308 5216 10310
rect 5272 10308 5296 10310
rect 5352 10308 5376 10310
rect 5432 10308 5456 10310
rect 5512 10308 5518 10310
rect 5210 10299 5518 10308
rect 5210 9276 5518 9285
rect 5210 9274 5216 9276
rect 5272 9274 5296 9276
rect 5352 9274 5376 9276
rect 5432 9274 5456 9276
rect 5512 9274 5518 9276
rect 5272 9222 5274 9274
rect 5454 9222 5456 9274
rect 5210 9220 5216 9222
rect 5272 9220 5296 9222
rect 5352 9220 5376 9222
rect 5432 9220 5456 9222
rect 5512 9220 5518 9222
rect 5210 9211 5518 9220
rect 5210 8188 5518 8197
rect 5210 8186 5216 8188
rect 5272 8186 5296 8188
rect 5352 8186 5376 8188
rect 5432 8186 5456 8188
rect 5512 8186 5518 8188
rect 5272 8134 5274 8186
rect 5454 8134 5456 8186
rect 5210 8132 5216 8134
rect 5272 8132 5296 8134
rect 5352 8132 5376 8134
rect 5432 8132 5456 8134
rect 5512 8132 5518 8134
rect 5210 8123 5518 8132
rect 5210 7100 5518 7109
rect 5210 7098 5216 7100
rect 5272 7098 5296 7100
rect 5352 7098 5376 7100
rect 5432 7098 5456 7100
rect 5512 7098 5518 7100
rect 5272 7046 5274 7098
rect 5454 7046 5456 7098
rect 5210 7044 5216 7046
rect 5272 7044 5296 7046
rect 5352 7044 5376 7046
rect 5432 7044 5456 7046
rect 5512 7044 5518 7046
rect 5210 7035 5518 7044
rect 5210 6012 5518 6021
rect 5210 6010 5216 6012
rect 5272 6010 5296 6012
rect 5352 6010 5376 6012
rect 5432 6010 5456 6012
rect 5512 6010 5518 6012
rect 5272 5958 5274 6010
rect 5454 5958 5456 6010
rect 5210 5956 5216 5958
rect 5272 5956 5296 5958
rect 5352 5956 5376 5958
rect 5432 5956 5456 5958
rect 5512 5956 5518 5958
rect 5210 5947 5518 5956
rect 5210 4924 5518 4933
rect 5210 4922 5216 4924
rect 5272 4922 5296 4924
rect 5352 4922 5376 4924
rect 5432 4922 5456 4924
rect 5512 4922 5518 4924
rect 5272 4870 5274 4922
rect 5454 4870 5456 4922
rect 5210 4868 5216 4870
rect 5272 4868 5296 4870
rect 5352 4868 5376 4870
rect 5432 4868 5456 4870
rect 5512 4868 5518 4870
rect 5210 4859 5518 4868
rect 5210 3836 5518 3845
rect 5210 3834 5216 3836
rect 5272 3834 5296 3836
rect 5352 3834 5376 3836
rect 5432 3834 5456 3836
rect 5512 3834 5518 3836
rect 5272 3782 5274 3834
rect 5454 3782 5456 3834
rect 5210 3780 5216 3782
rect 5272 3780 5296 3782
rect 5352 3780 5376 3782
rect 5432 3780 5456 3782
rect 5512 3780 5518 3782
rect 5210 3771 5518 3780
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5210 2748 5518 2757
rect 5210 2746 5216 2748
rect 5272 2746 5296 2748
rect 5352 2746 5376 2748
rect 5432 2746 5456 2748
rect 5512 2746 5518 2748
rect 5272 2694 5274 2746
rect 5454 2694 5456 2746
rect 5210 2692 5216 2694
rect 5272 2692 5296 2694
rect 5352 2692 5376 2694
rect 5432 2692 5456 2694
rect 5512 2692 5518 2694
rect 5210 2683 5518 2692
rect 5210 1660 5518 1669
rect 5210 1658 5216 1660
rect 5272 1658 5296 1660
rect 5352 1658 5376 1660
rect 5432 1658 5456 1660
rect 5512 1658 5518 1660
rect 5272 1606 5274 1658
rect 5454 1606 5456 1658
rect 5210 1604 5216 1606
rect 5272 1604 5296 1606
rect 5352 1604 5376 1606
rect 5432 1604 5456 1606
rect 5512 1604 5518 1606
rect 5210 1595 5518 1604
rect 5644 1018 5672 15846
rect 5736 3505 5764 19722
rect 5722 3496 5778 3505
rect 5722 3431 5778 3440
rect 5828 3194 5856 23190
rect 5920 22094 5948 25774
rect 6012 23118 6040 25792
rect 6196 25362 6224 25842
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6150 25052 6458 25061
rect 6150 25050 6156 25052
rect 6212 25050 6236 25052
rect 6292 25050 6316 25052
rect 6372 25050 6396 25052
rect 6452 25050 6458 25052
rect 6212 24998 6214 25050
rect 6394 24998 6396 25050
rect 6150 24996 6156 24998
rect 6212 24996 6236 24998
rect 6292 24996 6316 24998
rect 6372 24996 6396 24998
rect 6452 24996 6458 24998
rect 6150 24987 6458 24996
rect 6150 23964 6458 23973
rect 6150 23962 6156 23964
rect 6212 23962 6236 23964
rect 6292 23962 6316 23964
rect 6372 23962 6396 23964
rect 6452 23962 6458 23964
rect 6212 23910 6214 23962
rect 6394 23910 6396 23962
rect 6150 23908 6156 23910
rect 6212 23908 6236 23910
rect 6292 23908 6316 23910
rect 6372 23908 6396 23910
rect 6452 23908 6458 23910
rect 6150 23899 6458 23908
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6150 22876 6458 22885
rect 6150 22874 6156 22876
rect 6212 22874 6236 22876
rect 6292 22874 6316 22876
rect 6372 22874 6396 22876
rect 6452 22874 6458 22876
rect 6212 22822 6214 22874
rect 6394 22822 6396 22874
rect 6150 22820 6156 22822
rect 6212 22820 6236 22822
rect 6292 22820 6316 22822
rect 6372 22820 6396 22822
rect 6452 22820 6458 22822
rect 6150 22811 6458 22820
rect 6564 22710 6592 26166
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6552 22704 6604 22710
rect 6552 22646 6604 22652
rect 5920 22066 6592 22094
rect 5908 21956 5960 21962
rect 5908 21898 5960 21904
rect 5920 3641 5948 21898
rect 6150 21788 6458 21797
rect 6150 21786 6156 21788
rect 6212 21786 6236 21788
rect 6292 21786 6316 21788
rect 6372 21786 6396 21788
rect 6452 21786 6458 21788
rect 6212 21734 6214 21786
rect 6394 21734 6396 21786
rect 6150 21732 6156 21734
rect 6212 21732 6236 21734
rect 6292 21732 6316 21734
rect 6372 21732 6396 21734
rect 6452 21732 6458 21734
rect 6150 21723 6458 21732
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5906 3632 5962 3641
rect 5906 3567 5962 3576
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6012 2650 6040 20810
rect 6150 20700 6458 20709
rect 6150 20698 6156 20700
rect 6212 20698 6236 20700
rect 6292 20698 6316 20700
rect 6372 20698 6396 20700
rect 6452 20698 6458 20700
rect 6212 20646 6214 20698
rect 6394 20646 6396 20698
rect 6150 20644 6156 20646
rect 6212 20644 6236 20646
rect 6292 20644 6316 20646
rect 6372 20644 6396 20646
rect 6452 20644 6458 20646
rect 6150 20635 6458 20644
rect 6150 19612 6458 19621
rect 6150 19610 6156 19612
rect 6212 19610 6236 19612
rect 6292 19610 6316 19612
rect 6372 19610 6396 19612
rect 6452 19610 6458 19612
rect 6212 19558 6214 19610
rect 6394 19558 6396 19610
rect 6150 19556 6156 19558
rect 6212 19556 6236 19558
rect 6292 19556 6316 19558
rect 6372 19556 6396 19558
rect 6452 19556 6458 19558
rect 6150 19547 6458 19556
rect 6150 18524 6458 18533
rect 6150 18522 6156 18524
rect 6212 18522 6236 18524
rect 6292 18522 6316 18524
rect 6372 18522 6396 18524
rect 6452 18522 6458 18524
rect 6212 18470 6214 18522
rect 6394 18470 6396 18522
rect 6150 18468 6156 18470
rect 6212 18468 6236 18470
rect 6292 18468 6316 18470
rect 6372 18468 6396 18470
rect 6452 18468 6458 18470
rect 6150 18459 6458 18468
rect 6150 17436 6458 17445
rect 6150 17434 6156 17436
rect 6212 17434 6236 17436
rect 6292 17434 6316 17436
rect 6372 17434 6396 17436
rect 6452 17434 6458 17436
rect 6212 17382 6214 17434
rect 6394 17382 6396 17434
rect 6150 17380 6156 17382
rect 6212 17380 6236 17382
rect 6292 17380 6316 17382
rect 6372 17380 6396 17382
rect 6452 17380 6458 17382
rect 6150 17371 6458 17380
rect 6150 16348 6458 16357
rect 6150 16346 6156 16348
rect 6212 16346 6236 16348
rect 6292 16346 6316 16348
rect 6372 16346 6396 16348
rect 6452 16346 6458 16348
rect 6212 16294 6214 16346
rect 6394 16294 6396 16346
rect 6150 16292 6156 16294
rect 6212 16292 6236 16294
rect 6292 16292 6316 16294
rect 6372 16292 6396 16294
rect 6452 16292 6458 16294
rect 6150 16283 6458 16292
rect 6150 15260 6458 15269
rect 6150 15258 6156 15260
rect 6212 15258 6236 15260
rect 6292 15258 6316 15260
rect 6372 15258 6396 15260
rect 6452 15258 6458 15260
rect 6212 15206 6214 15258
rect 6394 15206 6396 15258
rect 6150 15204 6156 15206
rect 6212 15204 6236 15206
rect 6292 15204 6316 15206
rect 6372 15204 6396 15206
rect 6452 15204 6458 15206
rect 6150 15195 6458 15204
rect 6150 14172 6458 14181
rect 6150 14170 6156 14172
rect 6212 14170 6236 14172
rect 6292 14170 6316 14172
rect 6372 14170 6396 14172
rect 6452 14170 6458 14172
rect 6212 14118 6214 14170
rect 6394 14118 6396 14170
rect 6150 14116 6156 14118
rect 6212 14116 6236 14118
rect 6292 14116 6316 14118
rect 6372 14116 6396 14118
rect 6452 14116 6458 14118
rect 6150 14107 6458 14116
rect 6150 13084 6458 13093
rect 6150 13082 6156 13084
rect 6212 13082 6236 13084
rect 6292 13082 6316 13084
rect 6372 13082 6396 13084
rect 6452 13082 6458 13084
rect 6212 13030 6214 13082
rect 6394 13030 6396 13082
rect 6150 13028 6156 13030
rect 6212 13028 6236 13030
rect 6292 13028 6316 13030
rect 6372 13028 6396 13030
rect 6452 13028 6458 13030
rect 6150 13019 6458 13028
rect 6150 11996 6458 12005
rect 6150 11994 6156 11996
rect 6212 11994 6236 11996
rect 6292 11994 6316 11996
rect 6372 11994 6396 11996
rect 6452 11994 6458 11996
rect 6212 11942 6214 11994
rect 6394 11942 6396 11994
rect 6150 11940 6156 11942
rect 6212 11940 6236 11942
rect 6292 11940 6316 11942
rect 6372 11940 6396 11942
rect 6452 11940 6458 11942
rect 6150 11931 6458 11940
rect 6150 10908 6458 10917
rect 6150 10906 6156 10908
rect 6212 10906 6236 10908
rect 6292 10906 6316 10908
rect 6372 10906 6396 10908
rect 6452 10906 6458 10908
rect 6212 10854 6214 10906
rect 6394 10854 6396 10906
rect 6150 10852 6156 10854
rect 6212 10852 6236 10854
rect 6292 10852 6316 10854
rect 6372 10852 6396 10854
rect 6452 10852 6458 10854
rect 6150 10843 6458 10852
rect 6150 9820 6458 9829
rect 6150 9818 6156 9820
rect 6212 9818 6236 9820
rect 6292 9818 6316 9820
rect 6372 9818 6396 9820
rect 6452 9818 6458 9820
rect 6212 9766 6214 9818
rect 6394 9766 6396 9818
rect 6150 9764 6156 9766
rect 6212 9764 6236 9766
rect 6292 9764 6316 9766
rect 6372 9764 6396 9766
rect 6452 9764 6458 9766
rect 6150 9755 6458 9764
rect 6150 8732 6458 8741
rect 6150 8730 6156 8732
rect 6212 8730 6236 8732
rect 6292 8730 6316 8732
rect 6372 8730 6396 8732
rect 6452 8730 6458 8732
rect 6212 8678 6214 8730
rect 6394 8678 6396 8730
rect 6150 8676 6156 8678
rect 6212 8676 6236 8678
rect 6292 8676 6316 8678
rect 6372 8676 6396 8678
rect 6452 8676 6458 8678
rect 6150 8667 6458 8676
rect 6150 7644 6458 7653
rect 6150 7642 6156 7644
rect 6212 7642 6236 7644
rect 6292 7642 6316 7644
rect 6372 7642 6396 7644
rect 6452 7642 6458 7644
rect 6212 7590 6214 7642
rect 6394 7590 6396 7642
rect 6150 7588 6156 7590
rect 6212 7588 6236 7590
rect 6292 7588 6316 7590
rect 6372 7588 6396 7590
rect 6452 7588 6458 7590
rect 6150 7579 6458 7588
rect 6150 6556 6458 6565
rect 6150 6554 6156 6556
rect 6212 6554 6236 6556
rect 6292 6554 6316 6556
rect 6372 6554 6396 6556
rect 6452 6554 6458 6556
rect 6212 6502 6214 6554
rect 6394 6502 6396 6554
rect 6150 6500 6156 6502
rect 6212 6500 6236 6502
rect 6292 6500 6316 6502
rect 6372 6500 6396 6502
rect 6452 6500 6458 6502
rect 6150 6491 6458 6500
rect 6150 5468 6458 5477
rect 6150 5466 6156 5468
rect 6212 5466 6236 5468
rect 6292 5466 6316 5468
rect 6372 5466 6396 5468
rect 6452 5466 6458 5468
rect 6212 5414 6214 5466
rect 6394 5414 6396 5466
rect 6150 5412 6156 5414
rect 6212 5412 6236 5414
rect 6292 5412 6316 5414
rect 6372 5412 6396 5414
rect 6452 5412 6458 5414
rect 6150 5403 6458 5412
rect 6150 4380 6458 4389
rect 6150 4378 6156 4380
rect 6212 4378 6236 4380
rect 6292 4378 6316 4380
rect 6372 4378 6396 4380
rect 6452 4378 6458 4380
rect 6212 4326 6214 4378
rect 6394 4326 6396 4378
rect 6150 4324 6156 4326
rect 6212 4324 6236 4326
rect 6292 4324 6316 4326
rect 6372 4324 6396 4326
rect 6452 4324 6458 4326
rect 6150 4315 6458 4324
rect 6150 3292 6458 3301
rect 6150 3290 6156 3292
rect 6212 3290 6236 3292
rect 6292 3290 6316 3292
rect 6372 3290 6396 3292
rect 6452 3290 6458 3292
rect 6212 3238 6214 3290
rect 6394 3238 6396 3290
rect 6150 3236 6156 3238
rect 6212 3236 6236 3238
rect 6292 3236 6316 3238
rect 6372 3236 6396 3238
rect 6452 3236 6458 3238
rect 6150 3227 6458 3236
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6150 2204 6458 2213
rect 6150 2202 6156 2204
rect 6212 2202 6236 2204
rect 6292 2202 6316 2204
rect 6372 2202 6396 2204
rect 6452 2202 6458 2204
rect 6212 2150 6214 2202
rect 6394 2150 6396 2202
rect 6150 2148 6156 2150
rect 6212 2148 6236 2150
rect 6292 2148 6316 2150
rect 6372 2148 6396 2150
rect 6452 2148 6458 2150
rect 6150 2139 6458 2148
rect 6564 2106 6592 22066
rect 6656 3466 6684 24754
rect 6748 21894 6776 26846
rect 6840 26790 6868 27526
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 6932 26926 6960 27338
rect 7116 26994 7144 27628
rect 7194 27568 7250 27577
rect 7194 27503 7250 27512
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6810 26684 7118 26693
rect 6810 26682 6816 26684
rect 6872 26682 6896 26684
rect 6952 26682 6976 26684
rect 7032 26682 7056 26684
rect 7112 26682 7118 26684
rect 6872 26630 6874 26682
rect 7054 26630 7056 26682
rect 6810 26628 6816 26630
rect 6872 26628 6896 26630
rect 6952 26628 6976 26630
rect 7032 26628 7056 26630
rect 7112 26628 7118 26630
rect 6810 26619 7118 26628
rect 7208 26568 7236 27503
rect 6932 26540 7236 26568
rect 6932 26382 6960 26540
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 6932 25974 6960 26318
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 7024 25906 7052 26318
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7116 25838 7144 26386
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7104 25832 7156 25838
rect 7104 25774 7156 25780
rect 6810 25596 7118 25605
rect 6810 25594 6816 25596
rect 6872 25594 6896 25596
rect 6952 25594 6976 25596
rect 7032 25594 7056 25596
rect 7112 25594 7118 25596
rect 6872 25542 6874 25594
rect 7054 25542 7056 25594
rect 6810 25540 6816 25542
rect 6872 25540 6896 25542
rect 6952 25540 6976 25542
rect 7032 25540 7056 25542
rect 7112 25540 7118 25542
rect 6810 25531 7118 25540
rect 7208 25498 7236 26318
rect 7300 25770 7328 29106
rect 7392 27402 7420 31146
rect 7472 31136 7524 31142
rect 7472 31078 7524 31084
rect 7484 28558 7512 31078
rect 7472 28552 7524 28558
rect 7472 28494 7524 28500
rect 7470 28384 7526 28393
rect 7470 28319 7526 28328
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7288 25764 7340 25770
rect 7288 25706 7340 25712
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7300 25378 7328 25706
rect 7208 25350 7328 25378
rect 6810 24508 7118 24517
rect 6810 24506 6816 24508
rect 6872 24506 6896 24508
rect 6952 24506 6976 24508
rect 7032 24506 7056 24508
rect 7112 24506 7118 24508
rect 6872 24454 6874 24506
rect 7054 24454 7056 24506
rect 6810 24452 6816 24454
rect 6872 24452 6896 24454
rect 6952 24452 6976 24454
rect 7032 24452 7056 24454
rect 7112 24452 7118 24454
rect 6810 24443 7118 24452
rect 6810 23420 7118 23429
rect 6810 23418 6816 23420
rect 6872 23418 6896 23420
rect 6952 23418 6976 23420
rect 7032 23418 7056 23420
rect 7112 23418 7118 23420
rect 6872 23366 6874 23418
rect 7054 23366 7056 23418
rect 6810 23364 6816 23366
rect 6872 23364 6896 23366
rect 6952 23364 6976 23366
rect 7032 23364 7056 23366
rect 7112 23364 7118 23366
rect 6810 23355 7118 23364
rect 7208 22710 7236 25350
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24206 7328 25094
rect 7392 24410 7420 26522
rect 7484 26450 7512 28319
rect 7576 26586 7604 31198
rect 7668 29186 7696 31726
rect 7760 31686 7788 31826
rect 7852 31822 7880 32166
rect 7840 31816 7892 31822
rect 7840 31758 7892 31764
rect 8036 31754 8064 32438
rect 8128 32026 8156 32846
rect 8220 32570 8248 33510
rect 8392 33458 8444 33464
rect 8404 33402 8432 33458
rect 8496 33454 8524 33798
rect 8312 33374 8432 33402
rect 8484 33448 8536 33454
rect 8484 33390 8536 33396
rect 8588 33402 8616 34002
rect 8668 33924 8720 33930
rect 8668 33866 8720 33872
rect 8680 33658 8708 33866
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8772 33538 8800 42350
rect 8852 42016 8904 42022
rect 8852 41958 8904 41964
rect 8864 40594 8892 41958
rect 8852 40588 8904 40594
rect 8852 40530 8904 40536
rect 8956 40186 8984 42520
rect 8944 40180 8996 40186
rect 8944 40122 8996 40128
rect 9048 40050 9076 43590
rect 9140 40730 9168 45290
rect 9232 45286 9260 46974
rect 9350 46812 9658 46821
rect 9350 46810 9356 46812
rect 9412 46810 9436 46812
rect 9492 46810 9516 46812
rect 9572 46810 9596 46812
rect 9652 46810 9658 46812
rect 9412 46758 9414 46810
rect 9594 46758 9596 46810
rect 9350 46756 9356 46758
rect 9412 46756 9436 46758
rect 9492 46756 9516 46758
rect 9572 46756 9596 46758
rect 9652 46756 9658 46758
rect 9350 46747 9658 46756
rect 9692 46628 9720 46974
rect 9310 46608 9366 46617
rect 9310 46543 9366 46552
rect 9600 46600 9720 46628
rect 9324 45898 9352 46543
rect 9312 45892 9364 45898
rect 9312 45834 9364 45840
rect 9600 45812 9628 46600
rect 9600 45784 9720 45812
rect 9350 45724 9658 45733
rect 9350 45722 9356 45724
rect 9412 45722 9436 45724
rect 9492 45722 9516 45724
rect 9572 45722 9596 45724
rect 9652 45722 9658 45724
rect 9412 45670 9414 45722
rect 9594 45670 9596 45722
rect 9350 45668 9356 45670
rect 9412 45668 9436 45670
rect 9492 45668 9516 45670
rect 9572 45668 9596 45670
rect 9652 45668 9658 45670
rect 9350 45659 9658 45668
rect 9692 45506 9720 45784
rect 9600 45478 9720 45506
rect 9220 45280 9272 45286
rect 9220 45222 9272 45228
rect 9600 45014 9628 45478
rect 9220 45008 9272 45014
rect 9220 44950 9272 44956
rect 9588 45008 9640 45014
rect 9588 44950 9640 44956
rect 9128 40724 9180 40730
rect 9128 40666 9180 40672
rect 9140 40050 9168 40666
rect 9036 40044 9088 40050
rect 9036 39986 9088 39992
rect 9128 40044 9180 40050
rect 9128 39986 9180 39992
rect 8852 39840 8904 39846
rect 8852 39782 8904 39788
rect 8864 37398 8892 39782
rect 9232 39114 9260 44950
rect 9350 44636 9658 44645
rect 9350 44634 9356 44636
rect 9412 44634 9436 44636
rect 9492 44634 9516 44636
rect 9572 44634 9596 44636
rect 9652 44634 9658 44636
rect 9412 44582 9414 44634
rect 9594 44582 9596 44634
rect 9350 44580 9356 44582
rect 9412 44580 9436 44582
rect 9492 44580 9516 44582
rect 9572 44580 9596 44582
rect 9652 44580 9658 44582
rect 9350 44571 9658 44580
rect 9350 43548 9658 43557
rect 9350 43546 9356 43548
rect 9412 43546 9436 43548
rect 9492 43546 9516 43548
rect 9572 43546 9596 43548
rect 9652 43546 9658 43548
rect 9412 43494 9414 43546
rect 9594 43494 9596 43546
rect 9350 43492 9356 43494
rect 9412 43492 9436 43494
rect 9492 43492 9516 43494
rect 9572 43492 9596 43494
rect 9652 43492 9658 43494
rect 9350 43483 9658 43492
rect 9350 42460 9658 42469
rect 9350 42458 9356 42460
rect 9412 42458 9436 42460
rect 9492 42458 9516 42460
rect 9572 42458 9596 42460
rect 9652 42458 9658 42460
rect 9412 42406 9414 42458
rect 9594 42406 9596 42458
rect 9350 42404 9356 42406
rect 9412 42404 9436 42406
rect 9492 42404 9516 42406
rect 9572 42404 9596 42406
rect 9652 42404 9658 42406
rect 9350 42395 9658 42404
rect 9350 41372 9658 41381
rect 9350 41370 9356 41372
rect 9412 41370 9436 41372
rect 9492 41370 9516 41372
rect 9572 41370 9596 41372
rect 9652 41370 9658 41372
rect 9412 41318 9414 41370
rect 9594 41318 9596 41370
rect 9350 41316 9356 41318
rect 9412 41316 9436 41318
rect 9492 41316 9516 41318
rect 9572 41316 9596 41318
rect 9652 41316 9658 41318
rect 9350 41307 9658 41316
rect 9350 40284 9658 40293
rect 9350 40282 9356 40284
rect 9412 40282 9436 40284
rect 9492 40282 9516 40284
rect 9572 40282 9596 40284
rect 9652 40282 9658 40284
rect 9412 40230 9414 40282
rect 9594 40230 9596 40282
rect 9350 40228 9356 40230
rect 9412 40228 9436 40230
rect 9492 40228 9516 40230
rect 9572 40228 9596 40230
rect 9652 40228 9658 40230
rect 9350 40219 9658 40228
rect 9350 39196 9658 39205
rect 9350 39194 9356 39196
rect 9412 39194 9436 39196
rect 9492 39194 9516 39196
rect 9572 39194 9596 39196
rect 9652 39194 9658 39196
rect 9412 39142 9414 39194
rect 9594 39142 9596 39194
rect 9350 39140 9356 39142
rect 9412 39140 9436 39142
rect 9492 39140 9516 39142
rect 9572 39140 9596 39142
rect 9652 39140 9658 39142
rect 9350 39131 9658 39140
rect 8956 39086 9260 39114
rect 8956 38654 8984 39086
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 8956 38626 9076 38654
rect 8852 37392 8904 37398
rect 8852 37334 8904 37340
rect 8852 36712 8904 36718
rect 8852 36654 8904 36660
rect 8864 36564 8892 36654
rect 8864 36536 8984 36564
rect 8850 36408 8906 36417
rect 8850 36343 8906 36352
rect 8864 36242 8892 36343
rect 8852 36236 8904 36242
rect 8852 36178 8904 36184
rect 8852 36100 8904 36106
rect 8956 36088 8984 36536
rect 8904 36060 8984 36088
rect 8852 36042 8904 36048
rect 8864 34542 8892 36042
rect 9048 34762 9076 38626
rect 9140 36904 9168 38694
rect 9350 38108 9658 38117
rect 9350 38106 9356 38108
rect 9412 38106 9436 38108
rect 9492 38106 9516 38108
rect 9572 38106 9596 38108
rect 9652 38106 9658 38108
rect 9412 38054 9414 38106
rect 9594 38054 9596 38106
rect 9350 38052 9356 38054
rect 9412 38052 9436 38054
rect 9492 38052 9516 38054
rect 9572 38052 9596 38054
rect 9652 38052 9658 38054
rect 9350 38043 9658 38052
rect 9784 37369 9812 53110
rect 9770 37360 9826 37369
rect 9770 37295 9826 37304
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9350 37020 9658 37029
rect 9350 37018 9356 37020
rect 9412 37018 9436 37020
rect 9492 37018 9516 37020
rect 9572 37018 9596 37020
rect 9652 37018 9658 37020
rect 9412 36966 9414 37018
rect 9594 36966 9596 37018
rect 9350 36964 9356 36966
rect 9412 36964 9436 36966
rect 9492 36964 9516 36966
rect 9572 36964 9596 36966
rect 9652 36964 9658 36966
rect 9350 36955 9658 36964
rect 9140 36876 9628 36904
rect 9220 36644 9272 36650
rect 9220 36586 9272 36592
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 8956 34734 9076 34762
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8864 33930 8892 34478
rect 8852 33924 8904 33930
rect 8852 33866 8904 33872
rect 8956 33862 8984 34734
rect 9036 34604 9088 34610
rect 9036 34546 9088 34552
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8772 33510 8892 33538
rect 8588 33374 8800 33402
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 8208 32360 8260 32366
rect 8208 32302 8260 32308
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 8128 31890 8156 31962
rect 8116 31884 8168 31890
rect 8116 31826 8168 31832
rect 8220 31754 8248 32302
rect 8036 31726 8156 31754
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 8128 31634 8156 31726
rect 8208 31748 8260 31754
rect 8208 31690 8260 31696
rect 8128 31606 8248 31634
rect 7750 31580 8058 31589
rect 7750 31578 7756 31580
rect 7812 31578 7836 31580
rect 7892 31578 7916 31580
rect 7972 31578 7996 31580
rect 8052 31578 8058 31580
rect 7812 31526 7814 31578
rect 7994 31526 7996 31578
rect 7750 31524 7756 31526
rect 7812 31524 7836 31526
rect 7892 31524 7916 31526
rect 7972 31524 7996 31526
rect 8052 31524 8058 31526
rect 7750 31515 8058 31524
rect 8116 31476 8168 31482
rect 8116 31418 8168 31424
rect 7750 30492 8058 30501
rect 7750 30490 7756 30492
rect 7812 30490 7836 30492
rect 7892 30490 7916 30492
rect 7972 30490 7996 30492
rect 8052 30490 8058 30492
rect 7812 30438 7814 30490
rect 7994 30438 7996 30490
rect 7750 30436 7756 30438
rect 7812 30436 7836 30438
rect 7892 30436 7916 30438
rect 7972 30436 7996 30438
rect 8052 30436 8058 30438
rect 7750 30427 8058 30436
rect 7750 29404 8058 29413
rect 7750 29402 7756 29404
rect 7812 29402 7836 29404
rect 7892 29402 7916 29404
rect 7972 29402 7996 29404
rect 8052 29402 8058 29404
rect 7812 29350 7814 29402
rect 7994 29350 7996 29402
rect 7750 29348 7756 29350
rect 7812 29348 7836 29350
rect 7892 29348 7916 29350
rect 7972 29348 7996 29350
rect 8052 29348 8058 29350
rect 7750 29339 8058 29348
rect 8128 29288 8156 31418
rect 8036 29260 8156 29288
rect 7668 29158 7788 29186
rect 7656 28620 7708 28626
rect 7656 28562 7708 28568
rect 7668 27674 7696 28562
rect 7760 28422 7788 29158
rect 8036 28994 8064 29260
rect 8220 29186 8248 31606
rect 7944 28966 8064 28994
rect 8128 29158 8248 29186
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7852 28694 7880 28902
rect 7840 28688 7892 28694
rect 7840 28630 7892 28636
rect 7944 28529 7972 28966
rect 7930 28520 7986 28529
rect 8128 28506 8156 29158
rect 8312 29050 8340 33374
rect 8410 33212 8718 33221
rect 8410 33210 8416 33212
rect 8472 33210 8496 33212
rect 8552 33210 8576 33212
rect 8632 33210 8656 33212
rect 8712 33210 8718 33212
rect 8472 33158 8474 33210
rect 8654 33158 8656 33210
rect 8410 33156 8416 33158
rect 8472 33156 8496 33158
rect 8552 33156 8576 33158
rect 8632 33156 8656 33158
rect 8712 33156 8718 33158
rect 8410 33147 8718 33156
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8680 32570 8708 33050
rect 8668 32564 8720 32570
rect 8668 32506 8720 32512
rect 8410 32124 8718 32133
rect 8410 32122 8416 32124
rect 8472 32122 8496 32124
rect 8552 32122 8576 32124
rect 8632 32122 8656 32124
rect 8712 32122 8718 32124
rect 8472 32070 8474 32122
rect 8654 32070 8656 32122
rect 8410 32068 8416 32070
rect 8472 32068 8496 32070
rect 8552 32068 8576 32070
rect 8632 32068 8656 32070
rect 8712 32068 8718 32070
rect 8410 32059 8718 32068
rect 8410 31036 8718 31045
rect 8410 31034 8416 31036
rect 8472 31034 8496 31036
rect 8552 31034 8576 31036
rect 8632 31034 8656 31036
rect 8712 31034 8718 31036
rect 8472 30982 8474 31034
rect 8654 30982 8656 31034
rect 8410 30980 8416 30982
rect 8472 30980 8496 30982
rect 8552 30980 8576 30982
rect 8632 30980 8656 30982
rect 8712 30980 8718 30982
rect 8410 30971 8718 30980
rect 8410 29948 8718 29957
rect 8410 29946 8416 29948
rect 8472 29946 8496 29948
rect 8552 29946 8576 29948
rect 8632 29946 8656 29948
rect 8712 29946 8718 29948
rect 8472 29894 8474 29946
rect 8654 29894 8656 29946
rect 8410 29892 8416 29894
rect 8472 29892 8496 29894
rect 8552 29892 8576 29894
rect 8632 29892 8656 29894
rect 8712 29892 8718 29894
rect 8410 29883 8718 29892
rect 8772 29050 8800 33374
rect 8864 32366 8892 33510
rect 8944 33516 8996 33522
rect 8944 33458 8996 33464
rect 8956 32978 8984 33458
rect 8944 32972 8996 32978
rect 8944 32914 8996 32920
rect 8852 32360 8904 32366
rect 8852 32302 8904 32308
rect 8956 31906 8984 32914
rect 8864 31878 8984 31906
rect 8864 29238 8892 31878
rect 8942 31784 8998 31793
rect 8942 31719 8998 31728
rect 8956 29238 8984 31719
rect 8852 29232 8904 29238
rect 8852 29174 8904 29180
rect 8944 29232 8996 29238
rect 8944 29174 8996 29180
rect 8220 29022 8340 29050
rect 8496 29022 8800 29050
rect 8220 28626 8248 29022
rect 8496 28994 8524 29022
rect 8312 28966 8524 28994
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 8128 28478 8248 28506
rect 7930 28455 7986 28464
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 8116 28416 8168 28422
rect 8116 28358 8168 28364
rect 7750 28316 8058 28325
rect 7750 28314 7756 28316
rect 7812 28314 7836 28316
rect 7892 28314 7916 28316
rect 7972 28314 7996 28316
rect 8052 28314 8058 28316
rect 7812 28262 7814 28314
rect 7994 28262 7996 28314
rect 7750 28260 7756 28262
rect 7812 28260 7836 28262
rect 7892 28260 7916 28262
rect 7972 28260 7996 28262
rect 8052 28260 8058 28262
rect 7750 28251 8058 28260
rect 7656 27668 7708 27674
rect 7656 27610 7708 27616
rect 7668 26926 7696 27610
rect 7750 27228 8058 27237
rect 7750 27226 7756 27228
rect 7812 27226 7836 27228
rect 7892 27226 7916 27228
rect 7972 27226 7996 27228
rect 8052 27226 8058 27228
rect 7812 27174 7814 27226
rect 7994 27174 7996 27226
rect 7750 27172 7756 27174
rect 7812 27172 7836 27174
rect 7892 27172 7916 27174
rect 7972 27172 7996 27174
rect 8052 27172 8058 27174
rect 7750 27163 8058 27172
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7668 26450 7696 26862
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 7668 26042 7696 26386
rect 7750 26140 8058 26149
rect 7750 26138 7756 26140
rect 7812 26138 7836 26140
rect 7892 26138 7916 26140
rect 7972 26138 7996 26140
rect 8052 26138 8058 26140
rect 7812 26086 7814 26138
rect 7994 26086 7996 26138
rect 7750 26084 7756 26086
rect 7812 26084 7836 26086
rect 7892 26084 7916 26086
rect 7972 26084 7996 26086
rect 8052 26084 8058 26086
rect 7750 26075 8058 26084
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 8128 25974 8156 28358
rect 8220 27130 8248 28478
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 8116 25968 8168 25974
rect 8116 25910 8168 25916
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 8024 25900 8076 25906
rect 8024 25842 8076 25848
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7196 22704 7248 22710
rect 7196 22646 7248 22652
rect 6810 22332 7118 22341
rect 6810 22330 6816 22332
rect 6872 22330 6896 22332
rect 6952 22330 6976 22332
rect 7032 22330 7056 22332
rect 7112 22330 7118 22332
rect 6872 22278 6874 22330
rect 7054 22278 7056 22330
rect 6810 22276 6816 22278
rect 6872 22276 6896 22278
rect 6952 22276 6976 22278
rect 7032 22276 7056 22278
rect 7112 22276 7118 22278
rect 6810 22267 7118 22276
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 20806 6776 21830
rect 7300 21554 7328 24142
rect 7392 22982 7420 24346
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7484 23866 7512 24278
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7576 22794 7604 25842
rect 7656 25832 7708 25838
rect 7654 25800 7656 25809
rect 7840 25832 7892 25838
rect 7708 25800 7710 25809
rect 7840 25774 7892 25780
rect 7654 25735 7710 25744
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7392 22766 7604 22794
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7392 21434 7420 22766
rect 7668 22098 7696 25638
rect 7852 25430 7880 25774
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 8036 25140 8064 25842
rect 8036 25112 8156 25140
rect 7750 25052 8058 25061
rect 7750 25050 7756 25052
rect 7812 25050 7836 25052
rect 7892 25050 7916 25052
rect 7972 25050 7996 25052
rect 8052 25050 8058 25052
rect 7812 24998 7814 25050
rect 7994 24998 7996 25050
rect 7750 24996 7756 24998
rect 7812 24996 7836 24998
rect 7892 24996 7916 24998
rect 7972 24996 7996 24998
rect 8052 24996 8058 24998
rect 7750 24987 8058 24996
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7760 24206 7788 24686
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7748 24200 7800 24206
rect 7748 24142 7800 24148
rect 7760 24070 7788 24142
rect 7852 24138 7880 24346
rect 7944 24274 7972 24890
rect 8128 24750 8156 25112
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 7932 24268 7984 24274
rect 7932 24210 7984 24216
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7750 23964 8058 23973
rect 7750 23962 7756 23964
rect 7812 23962 7836 23964
rect 7892 23962 7916 23964
rect 7972 23962 7996 23964
rect 8052 23962 8058 23964
rect 7812 23910 7814 23962
rect 7994 23910 7996 23962
rect 7750 23908 7756 23910
rect 7812 23908 7836 23910
rect 7892 23908 7916 23910
rect 7972 23908 7996 23910
rect 8052 23908 8058 23910
rect 7750 23899 8058 23908
rect 7750 22876 8058 22885
rect 7750 22874 7756 22876
rect 7812 22874 7836 22876
rect 7892 22874 7916 22876
rect 7972 22874 7996 22876
rect 8052 22874 8058 22876
rect 7812 22822 7814 22874
rect 7994 22822 7996 22874
rect 7750 22820 7756 22822
rect 7812 22820 7836 22822
rect 7892 22820 7916 22822
rect 7972 22820 7996 22822
rect 8052 22820 8058 22822
rect 7750 22811 8058 22820
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7656 22092 7708 22098
rect 7852 22094 7880 22374
rect 7656 22034 7708 22040
rect 7760 22066 7880 22094
rect 7760 21978 7788 22066
rect 7668 21950 7788 21978
rect 7300 21406 7420 21434
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 6810 21244 7118 21253
rect 6810 21242 6816 21244
rect 6872 21242 6896 21244
rect 6952 21242 6976 21244
rect 7032 21242 7056 21244
rect 7112 21242 7118 21244
rect 6872 21190 6874 21242
rect 7054 21190 7056 21242
rect 6810 21188 6816 21190
rect 6872 21188 6896 21190
rect 6952 21188 6976 21190
rect 7032 21188 7056 21190
rect 7112 21188 7118 21190
rect 6810 21179 7118 21188
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6810 20156 7118 20165
rect 6810 20154 6816 20156
rect 6872 20154 6896 20156
rect 6952 20154 6976 20156
rect 7032 20154 7056 20156
rect 7112 20154 7118 20156
rect 6872 20102 6874 20154
rect 7054 20102 7056 20154
rect 6810 20100 6816 20102
rect 6872 20100 6896 20102
rect 6952 20100 6976 20102
rect 7032 20100 7056 20102
rect 7112 20100 7118 20102
rect 6810 20091 7118 20100
rect 6810 19068 7118 19077
rect 6810 19066 6816 19068
rect 6872 19066 6896 19068
rect 6952 19066 6976 19068
rect 7032 19066 7056 19068
rect 7112 19066 7118 19068
rect 6872 19014 6874 19066
rect 7054 19014 7056 19066
rect 6810 19012 6816 19014
rect 6872 19012 6896 19014
rect 6952 19012 6976 19014
rect 7032 19012 7056 19014
rect 7112 19012 7118 19014
rect 6810 19003 7118 19012
rect 7300 18970 7328 21406
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 11898 6776 18566
rect 6810 17980 7118 17989
rect 6810 17978 6816 17980
rect 6872 17978 6896 17980
rect 6952 17978 6976 17980
rect 7032 17978 7056 17980
rect 7112 17978 7118 17980
rect 6872 17926 6874 17978
rect 7054 17926 7056 17978
rect 6810 17924 6816 17926
rect 6872 17924 6896 17926
rect 6952 17924 6976 17926
rect 7032 17924 7056 17926
rect 7112 17924 7118 17926
rect 6810 17915 7118 17924
rect 6810 16892 7118 16901
rect 6810 16890 6816 16892
rect 6872 16890 6896 16892
rect 6952 16890 6976 16892
rect 7032 16890 7056 16892
rect 7112 16890 7118 16892
rect 6872 16838 6874 16890
rect 7054 16838 7056 16890
rect 6810 16836 6816 16838
rect 6872 16836 6896 16838
rect 6952 16836 6976 16838
rect 7032 16836 7056 16838
rect 7112 16836 7118 16838
rect 6810 16827 7118 16836
rect 7208 16794 7236 18838
rect 7300 18834 7328 18906
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7300 17746 7328 18634
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7300 16454 7328 17682
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 6810 15804 7118 15813
rect 6810 15802 6816 15804
rect 6872 15802 6896 15804
rect 6952 15802 6976 15804
rect 7032 15802 7056 15804
rect 7112 15802 7118 15804
rect 6872 15750 6874 15802
rect 7054 15750 7056 15802
rect 6810 15748 6816 15750
rect 6872 15748 6896 15750
rect 6952 15748 6976 15750
rect 7032 15748 7056 15750
rect 7112 15748 7118 15750
rect 6810 15739 7118 15748
rect 6810 14716 7118 14725
rect 6810 14714 6816 14716
rect 6872 14714 6896 14716
rect 6952 14714 6976 14716
rect 7032 14714 7056 14716
rect 7112 14714 7118 14716
rect 6872 14662 6874 14714
rect 7054 14662 7056 14714
rect 6810 14660 6816 14662
rect 6872 14660 6896 14662
rect 6952 14660 6976 14662
rect 7032 14660 7056 14662
rect 7112 14660 7118 14662
rect 6810 14651 7118 14660
rect 7300 14346 7328 16390
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7392 14226 7420 20742
rect 7484 17746 7512 21422
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7576 17338 7604 21286
rect 7668 19334 7696 21950
rect 7750 21788 8058 21797
rect 7750 21786 7756 21788
rect 7812 21786 7836 21788
rect 7892 21786 7916 21788
rect 7972 21786 7996 21788
rect 8052 21786 8058 21788
rect 7812 21734 7814 21786
rect 7994 21734 7996 21786
rect 7750 21732 7756 21734
rect 7812 21732 7836 21734
rect 7892 21732 7916 21734
rect 7972 21732 7996 21734
rect 8052 21732 8058 21734
rect 7750 21723 8058 21732
rect 7750 20700 8058 20709
rect 7750 20698 7756 20700
rect 7812 20698 7836 20700
rect 7892 20698 7916 20700
rect 7972 20698 7996 20700
rect 8052 20698 8058 20700
rect 7812 20646 7814 20698
rect 7994 20646 7996 20698
rect 7750 20644 7756 20646
rect 7812 20644 7836 20646
rect 7892 20644 7916 20646
rect 7972 20644 7996 20646
rect 8052 20644 8058 20646
rect 7750 20635 8058 20644
rect 7750 19612 8058 19621
rect 7750 19610 7756 19612
rect 7812 19610 7836 19612
rect 7892 19610 7916 19612
rect 7972 19610 7996 19612
rect 8052 19610 8058 19612
rect 7812 19558 7814 19610
rect 7994 19558 7996 19610
rect 7750 19556 7756 19558
rect 7812 19556 7836 19558
rect 7892 19556 7916 19558
rect 7972 19556 7996 19558
rect 8052 19556 8058 19558
rect 7750 19547 8058 19556
rect 7668 19306 7788 19334
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7300 14198 7420 14226
rect 6810 13628 7118 13637
rect 6810 13626 6816 13628
rect 6872 13626 6896 13628
rect 6952 13626 6976 13628
rect 7032 13626 7056 13628
rect 7112 13626 7118 13628
rect 6872 13574 6874 13626
rect 7054 13574 7056 13626
rect 6810 13572 6816 13574
rect 6872 13572 6896 13574
rect 6952 13572 6976 13574
rect 7032 13572 7056 13574
rect 7112 13572 7118 13574
rect 6810 13563 7118 13572
rect 7300 13258 7328 14198
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 6810 12540 7118 12549
rect 6810 12538 6816 12540
rect 6872 12538 6896 12540
rect 6952 12538 6976 12540
rect 7032 12538 7056 12540
rect 7112 12538 7118 12540
rect 6872 12486 6874 12538
rect 7054 12486 7056 12538
rect 6810 12484 6816 12486
rect 6872 12484 6896 12486
rect 6952 12484 6976 12486
rect 7032 12484 7056 12486
rect 7112 12484 7118 12486
rect 6810 12475 7118 12484
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 7392 11762 7420 13330
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 6810 11452 7118 11461
rect 6810 11450 6816 11452
rect 6872 11450 6896 11452
rect 6952 11450 6976 11452
rect 7032 11450 7056 11452
rect 7112 11450 7118 11452
rect 6872 11398 6874 11450
rect 7054 11398 7056 11450
rect 6810 11396 6816 11398
rect 6872 11396 6896 11398
rect 6952 11396 6976 11398
rect 7032 11396 7056 11398
rect 7112 11396 7118 11398
rect 6810 11387 7118 11396
rect 7392 11218 7420 11698
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 6810 10364 7118 10373
rect 6810 10362 6816 10364
rect 6872 10362 6896 10364
rect 6952 10362 6976 10364
rect 7032 10362 7056 10364
rect 7112 10362 7118 10364
rect 6872 10310 6874 10362
rect 7054 10310 7056 10362
rect 6810 10308 6816 10310
rect 6872 10308 6896 10310
rect 6952 10308 6976 10310
rect 7032 10308 7056 10310
rect 7112 10308 7118 10310
rect 6810 10299 7118 10308
rect 7392 9518 7420 11154
rect 7484 11082 7512 16390
rect 7576 13394 7604 16934
rect 7668 16590 7696 18906
rect 7760 18902 7788 19306
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7750 18524 8058 18533
rect 7750 18522 7756 18524
rect 7812 18522 7836 18524
rect 7892 18522 7916 18524
rect 7972 18522 7996 18524
rect 8052 18522 8058 18524
rect 7812 18470 7814 18522
rect 7994 18470 7996 18522
rect 7750 18468 7756 18470
rect 7812 18468 7836 18470
rect 7892 18468 7916 18470
rect 7972 18468 7996 18470
rect 8052 18468 8058 18470
rect 7750 18459 8058 18468
rect 7750 17436 8058 17445
rect 7750 17434 7756 17436
rect 7812 17434 7836 17436
rect 7892 17434 7916 17436
rect 7972 17434 7996 17436
rect 8052 17434 8058 17436
rect 7812 17382 7814 17434
rect 7994 17382 7996 17434
rect 7750 17380 7756 17382
rect 7812 17380 7836 17382
rect 7892 17380 7916 17382
rect 7972 17380 7996 17382
rect 8052 17380 8058 17382
rect 7750 17371 8058 17380
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7668 16250 7696 16526
rect 7750 16348 8058 16357
rect 7750 16346 7756 16348
rect 7812 16346 7836 16348
rect 7892 16346 7916 16348
rect 7972 16346 7996 16348
rect 8052 16346 8058 16348
rect 7812 16294 7814 16346
rect 7994 16294 7996 16346
rect 7750 16292 7756 16294
rect 7812 16292 7836 16294
rect 7892 16292 7916 16294
rect 7972 16292 7996 16294
rect 8052 16292 8058 16294
rect 7750 16283 8058 16292
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7750 15260 8058 15269
rect 7750 15258 7756 15260
rect 7812 15258 7836 15260
rect 7892 15258 7916 15260
rect 7972 15258 7996 15260
rect 8052 15258 8058 15260
rect 7812 15206 7814 15258
rect 7994 15206 7996 15258
rect 7750 15204 7756 15206
rect 7812 15204 7836 15206
rect 7892 15204 7916 15206
rect 7972 15204 7996 15206
rect 8052 15204 8058 15206
rect 7750 15195 8058 15204
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 6810 9276 7118 9285
rect 6810 9274 6816 9276
rect 6872 9274 6896 9276
rect 6952 9274 6976 9276
rect 7032 9274 7056 9276
rect 7112 9274 7118 9276
rect 6872 9222 6874 9274
rect 7054 9222 7056 9274
rect 6810 9220 6816 9222
rect 6872 9220 6896 9222
rect 6952 9220 6976 9222
rect 7032 9220 7056 9222
rect 7112 9220 7118 9222
rect 6810 9211 7118 9220
rect 6810 8188 7118 8197
rect 6810 8186 6816 8188
rect 6872 8186 6896 8188
rect 6952 8186 6976 8188
rect 7032 8186 7056 8188
rect 7112 8186 7118 8188
rect 6872 8134 6874 8186
rect 7054 8134 7056 8186
rect 6810 8132 6816 8134
rect 6872 8132 6896 8134
rect 6952 8132 6976 8134
rect 7032 8132 7056 8134
rect 7112 8132 7118 8134
rect 6810 8123 7118 8132
rect 6810 7100 7118 7109
rect 6810 7098 6816 7100
rect 6872 7098 6896 7100
rect 6952 7098 6976 7100
rect 7032 7098 7056 7100
rect 7112 7098 7118 7100
rect 6872 7046 6874 7098
rect 7054 7046 7056 7098
rect 6810 7044 6816 7046
rect 6872 7044 6896 7046
rect 6952 7044 6976 7046
rect 7032 7044 7056 7046
rect 7112 7044 7118 7046
rect 6810 7035 7118 7044
rect 6810 6012 7118 6021
rect 6810 6010 6816 6012
rect 6872 6010 6896 6012
rect 6952 6010 6976 6012
rect 7032 6010 7056 6012
rect 7112 6010 7118 6012
rect 6872 5958 6874 6010
rect 7054 5958 7056 6010
rect 6810 5956 6816 5958
rect 6872 5956 6896 5958
rect 6952 5956 6976 5958
rect 7032 5956 7056 5958
rect 7112 5956 7118 5958
rect 6810 5947 7118 5956
rect 6810 4924 7118 4933
rect 6810 4922 6816 4924
rect 6872 4922 6896 4924
rect 6952 4922 6976 4924
rect 7032 4922 7056 4924
rect 7112 4922 7118 4924
rect 6872 4870 6874 4922
rect 7054 4870 7056 4922
rect 6810 4868 6816 4870
rect 6872 4868 6896 4870
rect 6952 4868 6976 4870
rect 7032 4868 7056 4870
rect 7112 4868 7118 4870
rect 6810 4859 7118 4868
rect 6810 3836 7118 3845
rect 6810 3834 6816 3836
rect 6872 3834 6896 3836
rect 6952 3834 6976 3836
rect 7032 3834 7056 3836
rect 7112 3834 7118 3836
rect 6872 3782 6874 3834
rect 7054 3782 7056 3834
rect 6810 3780 6816 3782
rect 6872 3780 6896 3782
rect 6952 3780 6976 3782
rect 7032 3780 7056 3782
rect 7112 3780 7118 3782
rect 6810 3771 7118 3780
rect 7576 3670 7604 13194
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6810 2748 7118 2757
rect 6810 2746 6816 2748
rect 6872 2746 6896 2748
rect 6952 2746 6976 2748
rect 7032 2746 7056 2748
rect 7112 2746 7118 2748
rect 6872 2694 6874 2746
rect 7054 2694 7056 2746
rect 6810 2692 6816 2694
rect 6872 2692 6896 2694
rect 6952 2692 6976 2694
rect 7032 2692 7056 2694
rect 7112 2692 7118 2694
rect 6810 2683 7118 2692
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6810 1660 7118 1669
rect 6810 1658 6816 1660
rect 6872 1658 6896 1660
rect 6952 1658 6976 1660
rect 7032 1658 7056 1660
rect 7112 1658 7118 1660
rect 6872 1606 6874 1658
rect 7054 1606 7056 1658
rect 6810 1604 6816 1606
rect 6872 1604 6896 1606
rect 6952 1604 6976 1606
rect 7032 1604 7056 1606
rect 7112 1604 7118 1606
rect 6810 1595 7118 1604
rect 6150 1116 6458 1125
rect 6150 1114 6156 1116
rect 6212 1114 6236 1116
rect 6292 1114 6316 1116
rect 6372 1114 6396 1116
rect 6452 1114 6458 1116
rect 6212 1062 6214 1114
rect 6394 1062 6396 1114
rect 6150 1060 6156 1062
rect 6212 1060 6236 1062
rect 6292 1060 6316 1062
rect 6372 1060 6396 1062
rect 6452 1060 6458 1062
rect 6150 1051 6458 1060
rect 5632 1012 5684 1018
rect 5632 954 5684 960
rect 4986 776 5042 785
rect 4986 711 5042 720
rect 7668 542 7696 14486
rect 7750 14172 8058 14181
rect 7750 14170 7756 14172
rect 7812 14170 7836 14172
rect 7892 14170 7916 14172
rect 7972 14170 7996 14172
rect 8052 14170 8058 14172
rect 7812 14118 7814 14170
rect 7994 14118 7996 14170
rect 7750 14116 7756 14118
rect 7812 14116 7836 14118
rect 7892 14116 7916 14118
rect 7972 14116 7996 14118
rect 8052 14116 8058 14118
rect 7750 14107 8058 14116
rect 8128 13954 8156 24278
rect 8220 23118 8248 26726
rect 8312 24410 8340 28966
rect 8410 28860 8718 28869
rect 8410 28858 8416 28860
rect 8472 28858 8496 28860
rect 8552 28858 8576 28860
rect 8632 28858 8656 28860
rect 8712 28858 8718 28860
rect 8472 28806 8474 28858
rect 8654 28806 8656 28858
rect 8410 28804 8416 28806
rect 8472 28804 8496 28806
rect 8552 28804 8576 28806
rect 8632 28804 8656 28806
rect 8712 28804 8718 28806
rect 8410 28795 8718 28804
rect 8864 28778 8892 29174
rect 9048 29050 9076 34546
rect 8772 28750 8892 28778
rect 8956 29022 9076 29050
rect 8484 28620 8536 28626
rect 8536 28580 8708 28608
rect 8484 28562 8536 28568
rect 8680 27962 8708 28580
rect 8772 28558 8800 28750
rect 8852 28620 8904 28626
rect 8852 28562 8904 28568
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 8680 27934 8800 27962
rect 8410 27772 8718 27781
rect 8410 27770 8416 27772
rect 8472 27770 8496 27772
rect 8552 27770 8576 27772
rect 8632 27770 8656 27772
rect 8712 27770 8718 27772
rect 8472 27718 8474 27770
rect 8654 27718 8656 27770
rect 8410 27716 8416 27718
rect 8472 27716 8496 27718
rect 8552 27716 8576 27718
rect 8632 27716 8656 27718
rect 8712 27716 8718 27718
rect 8410 27707 8718 27716
rect 8410 26684 8718 26693
rect 8410 26682 8416 26684
rect 8472 26682 8496 26684
rect 8552 26682 8576 26684
rect 8632 26682 8656 26684
rect 8712 26682 8718 26684
rect 8472 26630 8474 26682
rect 8654 26630 8656 26682
rect 8410 26628 8416 26630
rect 8472 26628 8496 26630
rect 8552 26628 8576 26630
rect 8632 26628 8656 26630
rect 8712 26628 8718 26630
rect 8410 26619 8718 26628
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8404 26042 8432 26182
rect 8392 26036 8444 26042
rect 8392 25978 8444 25984
rect 8772 25838 8800 27934
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8410 25596 8718 25605
rect 8410 25594 8416 25596
rect 8472 25594 8496 25596
rect 8552 25594 8576 25596
rect 8632 25594 8656 25596
rect 8712 25594 8718 25596
rect 8472 25542 8474 25594
rect 8654 25542 8656 25594
rect 8410 25540 8416 25542
rect 8472 25540 8496 25542
rect 8552 25540 8576 25542
rect 8632 25540 8656 25542
rect 8712 25540 8718 25542
rect 8410 25531 8718 25540
rect 8410 24508 8718 24517
rect 8410 24506 8416 24508
rect 8472 24506 8496 24508
rect 8552 24506 8576 24508
rect 8632 24506 8656 24508
rect 8712 24506 8718 24508
rect 8472 24454 8474 24506
rect 8654 24454 8656 24506
rect 8410 24452 8416 24454
rect 8472 24452 8496 24454
rect 8552 24452 8576 24454
rect 8632 24452 8656 24454
rect 8712 24452 8718 24454
rect 8410 24443 8718 24452
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8220 18766 8248 22918
rect 8312 19854 8340 23802
rect 8404 23662 8432 24006
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8410 23420 8718 23429
rect 8410 23418 8416 23420
rect 8472 23418 8496 23420
rect 8552 23418 8576 23420
rect 8632 23418 8656 23420
rect 8712 23418 8718 23420
rect 8472 23366 8474 23418
rect 8654 23366 8656 23418
rect 8410 23364 8416 23366
rect 8472 23364 8496 23366
rect 8552 23364 8576 23366
rect 8632 23364 8656 23366
rect 8712 23364 8718 23366
rect 8410 23355 8718 23364
rect 8410 22332 8718 22341
rect 8410 22330 8416 22332
rect 8472 22330 8496 22332
rect 8552 22330 8576 22332
rect 8632 22330 8656 22332
rect 8712 22330 8718 22332
rect 8472 22278 8474 22330
rect 8654 22278 8656 22330
rect 8410 22276 8416 22278
rect 8472 22276 8496 22278
rect 8552 22276 8576 22278
rect 8632 22276 8656 22278
rect 8712 22276 8718 22278
rect 8410 22267 8718 22276
rect 8410 21244 8718 21253
rect 8410 21242 8416 21244
rect 8472 21242 8496 21244
rect 8552 21242 8576 21244
rect 8632 21242 8656 21244
rect 8712 21242 8718 21244
rect 8472 21190 8474 21242
rect 8654 21190 8656 21242
rect 8410 21188 8416 21190
rect 8472 21188 8496 21190
rect 8552 21188 8576 21190
rect 8632 21188 8656 21190
rect 8712 21188 8718 21190
rect 8410 21179 8718 21188
rect 8772 20466 8800 25638
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8864 20262 8892 28562
rect 8956 26790 8984 29022
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8944 26512 8996 26518
rect 8944 26454 8996 26460
rect 8956 23118 8984 26454
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8410 20156 8718 20165
rect 8410 20154 8416 20156
rect 8472 20154 8496 20156
rect 8552 20154 8576 20156
rect 8632 20154 8656 20156
rect 8712 20154 8718 20156
rect 8472 20102 8474 20154
rect 8654 20102 8656 20154
rect 8410 20100 8416 20102
rect 8472 20100 8496 20102
rect 8552 20100 8576 20102
rect 8632 20100 8656 20102
rect 8712 20100 8718 20102
rect 8410 20091 8718 20100
rect 8956 20074 8984 22918
rect 8864 20046 8984 20074
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8410 19068 8718 19077
rect 8410 19066 8416 19068
rect 8472 19066 8496 19068
rect 8552 19066 8576 19068
rect 8632 19066 8656 19068
rect 8712 19066 8718 19068
rect 8472 19014 8474 19066
rect 8654 19014 8656 19066
rect 8410 19012 8416 19014
rect 8472 19012 8496 19014
rect 8552 19012 8576 19014
rect 8632 19012 8656 19014
rect 8712 19012 8718 19014
rect 8410 19003 8718 19012
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8410 17980 8718 17989
rect 8410 17978 8416 17980
rect 8472 17978 8496 17980
rect 8552 17978 8576 17980
rect 8632 17978 8656 17980
rect 8712 17978 8718 17980
rect 8472 17926 8474 17978
rect 8654 17926 8656 17978
rect 8410 17924 8416 17926
rect 8472 17924 8496 17926
rect 8552 17924 8576 17926
rect 8632 17924 8656 17926
rect 8712 17924 8718 17926
rect 8410 17915 8718 17924
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8220 16046 8248 16662
rect 8312 16590 8340 17478
rect 8410 16892 8718 16901
rect 8410 16890 8416 16892
rect 8472 16890 8496 16892
rect 8552 16890 8576 16892
rect 8632 16890 8656 16892
rect 8712 16890 8718 16892
rect 8472 16838 8474 16890
rect 8654 16838 8656 16890
rect 8410 16836 8416 16838
rect 8472 16836 8496 16838
rect 8552 16836 8576 16838
rect 8632 16836 8656 16838
rect 8712 16836 8718 16838
rect 8410 16827 8718 16836
rect 8864 16708 8892 20046
rect 9048 19718 9076 28902
rect 9140 26042 9168 36110
rect 9232 32026 9260 36586
rect 9600 36122 9628 36876
rect 9600 36094 9720 36122
rect 9350 35932 9658 35941
rect 9350 35930 9356 35932
rect 9412 35930 9436 35932
rect 9492 35930 9516 35932
rect 9572 35930 9596 35932
rect 9652 35930 9658 35932
rect 9412 35878 9414 35930
rect 9594 35878 9596 35930
rect 9350 35876 9356 35878
rect 9412 35876 9436 35878
rect 9492 35876 9516 35878
rect 9572 35876 9596 35878
rect 9652 35876 9658 35878
rect 9350 35867 9658 35876
rect 9692 35714 9720 36094
rect 9600 35686 9720 35714
rect 9600 35034 9628 35686
rect 9600 35006 9720 35034
rect 9350 34844 9658 34853
rect 9350 34842 9356 34844
rect 9412 34842 9436 34844
rect 9492 34842 9516 34844
rect 9572 34842 9596 34844
rect 9652 34842 9658 34844
rect 9412 34790 9414 34842
rect 9594 34790 9596 34842
rect 9350 34788 9356 34790
rect 9412 34788 9436 34790
rect 9492 34788 9516 34790
rect 9572 34788 9596 34790
rect 9652 34788 9658 34790
rect 9350 34779 9658 34788
rect 9692 34626 9720 35006
rect 9600 34598 9720 34626
rect 9600 33946 9628 34598
rect 9600 33918 9720 33946
rect 9350 33756 9658 33765
rect 9350 33754 9356 33756
rect 9412 33754 9436 33756
rect 9492 33754 9516 33756
rect 9572 33754 9596 33756
rect 9652 33754 9658 33756
rect 9412 33702 9414 33754
rect 9594 33702 9596 33754
rect 9350 33700 9356 33702
rect 9412 33700 9436 33702
rect 9492 33700 9516 33702
rect 9572 33700 9596 33702
rect 9652 33700 9658 33702
rect 9350 33691 9658 33700
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9324 33114 9352 33594
rect 9692 33538 9720 33918
rect 9600 33510 9720 33538
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9600 32858 9628 33510
rect 9600 32830 9720 32858
rect 9350 32668 9658 32677
rect 9350 32666 9356 32668
rect 9412 32666 9436 32668
rect 9492 32666 9516 32668
rect 9572 32666 9596 32668
rect 9652 32666 9658 32668
rect 9412 32614 9414 32666
rect 9594 32614 9596 32666
rect 9350 32612 9356 32614
rect 9412 32612 9436 32614
rect 9492 32612 9516 32614
rect 9572 32612 9596 32614
rect 9652 32612 9658 32614
rect 9350 32603 9658 32612
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9220 32020 9272 32026
rect 9220 31962 9272 31968
rect 9324 31906 9352 32506
rect 9692 32476 9720 32830
rect 9232 31878 9352 31906
rect 9508 32448 9720 32476
rect 9232 30326 9260 31878
rect 9508 31793 9536 32448
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9494 31784 9550 31793
rect 9494 31719 9550 31728
rect 9600 31754 9628 31894
rect 9600 31726 9720 31754
rect 9350 31580 9658 31589
rect 9350 31578 9356 31580
rect 9412 31578 9436 31580
rect 9492 31578 9516 31580
rect 9572 31578 9596 31580
rect 9652 31578 9658 31580
rect 9412 31526 9414 31578
rect 9594 31526 9596 31578
rect 9350 31524 9356 31526
rect 9412 31524 9436 31526
rect 9492 31524 9516 31526
rect 9572 31524 9596 31526
rect 9652 31524 9658 31526
rect 9350 31515 9658 31524
rect 9692 31362 9720 31726
rect 9600 31334 9720 31362
rect 9600 30682 9628 31334
rect 9600 30654 9720 30682
rect 9350 30492 9658 30501
rect 9350 30490 9356 30492
rect 9412 30490 9436 30492
rect 9492 30490 9516 30492
rect 9572 30490 9596 30492
rect 9652 30490 9658 30492
rect 9412 30438 9414 30490
rect 9594 30438 9596 30490
rect 9350 30436 9356 30438
rect 9412 30436 9436 30438
rect 9492 30436 9516 30438
rect 9572 30436 9596 30438
rect 9652 30436 9658 30438
rect 9350 30427 9658 30436
rect 9220 30320 9272 30326
rect 9692 30274 9720 30654
rect 9220 30262 9272 30268
rect 9600 30246 9720 30274
rect 9600 29594 9628 30246
rect 9600 29566 9720 29594
rect 9350 29404 9658 29413
rect 9350 29402 9356 29404
rect 9412 29402 9436 29404
rect 9492 29402 9516 29404
rect 9572 29402 9596 29404
rect 9652 29402 9658 29404
rect 9412 29350 9414 29402
rect 9594 29350 9596 29402
rect 9350 29348 9356 29350
rect 9412 29348 9436 29350
rect 9492 29348 9516 29350
rect 9572 29348 9596 29350
rect 9652 29348 9658 29350
rect 9350 29339 9658 29348
rect 9692 29186 9720 29566
rect 9600 29158 9720 29186
rect 9220 28756 9272 28762
rect 9220 28698 9272 28704
rect 9128 26036 9180 26042
rect 9128 25978 9180 25984
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9048 19334 9076 19654
rect 8772 16680 8892 16708
rect 8956 19306 9076 19334
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 14482 8248 15982
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8036 13926 8156 13954
rect 8036 13326 8064 13926
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7750 13084 8058 13093
rect 7750 13082 7756 13084
rect 7812 13082 7836 13084
rect 7892 13082 7916 13084
rect 7972 13082 7996 13084
rect 8052 13082 8058 13084
rect 7812 13030 7814 13082
rect 7994 13030 7996 13082
rect 7750 13028 7756 13030
rect 7812 13028 7836 13030
rect 7892 13028 7916 13030
rect 7972 13028 7996 13030
rect 8052 13028 8058 13030
rect 7750 13019 8058 13028
rect 7750 11996 8058 12005
rect 7750 11994 7756 11996
rect 7812 11994 7836 11996
rect 7892 11994 7916 11996
rect 7972 11994 7996 11996
rect 8052 11994 8058 11996
rect 7812 11942 7814 11994
rect 7994 11942 7996 11994
rect 7750 11940 7756 11942
rect 7812 11940 7836 11942
rect 7892 11940 7916 11942
rect 7972 11940 7996 11942
rect 8052 11940 8058 11942
rect 7750 11931 8058 11940
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7750 10908 8058 10917
rect 7750 10906 7756 10908
rect 7812 10906 7836 10908
rect 7892 10906 7916 10908
rect 7972 10906 7996 10908
rect 8052 10906 8058 10908
rect 7812 10854 7814 10906
rect 7994 10854 7996 10906
rect 7750 10852 7756 10854
rect 7812 10852 7836 10854
rect 7892 10852 7916 10854
rect 7972 10852 7996 10854
rect 8052 10852 8058 10854
rect 7750 10843 8058 10852
rect 7750 9820 8058 9829
rect 7750 9818 7756 9820
rect 7812 9818 7836 9820
rect 7892 9818 7916 9820
rect 7972 9818 7996 9820
rect 8052 9818 8058 9820
rect 7812 9766 7814 9818
rect 7994 9766 7996 9818
rect 7750 9764 7756 9766
rect 7812 9764 7836 9766
rect 7892 9764 7916 9766
rect 7972 9764 7996 9766
rect 8052 9764 8058 9766
rect 7750 9755 8058 9764
rect 7750 8732 8058 8741
rect 7750 8730 7756 8732
rect 7812 8730 7836 8732
rect 7892 8730 7916 8732
rect 7972 8730 7996 8732
rect 8052 8730 8058 8732
rect 7812 8678 7814 8730
rect 7994 8678 7996 8730
rect 7750 8676 7756 8678
rect 7812 8676 7836 8678
rect 7892 8676 7916 8678
rect 7972 8676 7996 8678
rect 8052 8676 8058 8678
rect 7750 8667 8058 8676
rect 7750 7644 8058 7653
rect 7750 7642 7756 7644
rect 7812 7642 7836 7644
rect 7892 7642 7916 7644
rect 7972 7642 7996 7644
rect 8052 7642 8058 7644
rect 7812 7590 7814 7642
rect 7994 7590 7996 7642
rect 7750 7588 7756 7590
rect 7812 7588 7836 7590
rect 7892 7588 7916 7590
rect 7972 7588 7996 7590
rect 8052 7588 8058 7590
rect 7750 7579 8058 7588
rect 7750 6556 8058 6565
rect 7750 6554 7756 6556
rect 7812 6554 7836 6556
rect 7892 6554 7916 6556
rect 7972 6554 7996 6556
rect 8052 6554 8058 6556
rect 7812 6502 7814 6554
rect 7994 6502 7996 6554
rect 7750 6500 7756 6502
rect 7812 6500 7836 6502
rect 7892 6500 7916 6502
rect 7972 6500 7996 6502
rect 8052 6500 8058 6502
rect 7750 6491 8058 6500
rect 7750 5468 8058 5477
rect 7750 5466 7756 5468
rect 7812 5466 7836 5468
rect 7892 5466 7916 5468
rect 7972 5466 7996 5468
rect 8052 5466 8058 5468
rect 7812 5414 7814 5466
rect 7994 5414 7996 5466
rect 7750 5412 7756 5414
rect 7812 5412 7836 5414
rect 7892 5412 7916 5414
rect 7972 5412 7996 5414
rect 8052 5412 8058 5414
rect 7750 5403 8058 5412
rect 7750 4380 8058 4389
rect 7750 4378 7756 4380
rect 7812 4378 7836 4380
rect 7892 4378 7916 4380
rect 7972 4378 7996 4380
rect 8052 4378 8058 4380
rect 7812 4326 7814 4378
rect 7994 4326 7996 4378
rect 7750 4324 7756 4326
rect 7812 4324 7836 4326
rect 7892 4324 7916 4326
rect 7972 4324 7996 4326
rect 8052 4324 8058 4326
rect 7750 4315 8058 4324
rect 7750 3292 8058 3301
rect 7750 3290 7756 3292
rect 7812 3290 7836 3292
rect 7892 3290 7916 3292
rect 7972 3290 7996 3292
rect 8052 3290 8058 3292
rect 7812 3238 7814 3290
rect 7994 3238 7996 3290
rect 7750 3236 7756 3238
rect 7812 3236 7836 3238
rect 7892 3236 7916 3238
rect 7972 3236 7996 3238
rect 8052 3236 8058 3238
rect 7750 3227 8058 3236
rect 8128 2582 8156 11494
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 7750 2204 8058 2213
rect 7750 2202 7756 2204
rect 7812 2202 7836 2204
rect 7892 2202 7916 2204
rect 7972 2202 7996 2204
rect 8052 2202 8058 2204
rect 7812 2150 7814 2202
rect 7994 2150 7996 2202
rect 7750 2148 7756 2150
rect 7812 2148 7836 2150
rect 7892 2148 7916 2150
rect 7972 2148 7996 2150
rect 8052 2148 8058 2150
rect 7750 2139 8058 2148
rect 7750 1116 8058 1125
rect 7750 1114 7756 1116
rect 7812 1114 7836 1116
rect 7892 1114 7916 1116
rect 7972 1114 7996 1116
rect 8052 1114 8058 1116
rect 7812 1062 7814 1114
rect 7994 1062 7996 1114
rect 7750 1060 7756 1062
rect 7812 1060 7836 1062
rect 7892 1060 7916 1062
rect 7972 1060 7996 1062
rect 8052 1060 8058 1062
rect 7750 1051 8058 1060
rect 8220 814 8248 9318
rect 8312 9058 8340 16390
rect 8772 16182 8800 16680
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8410 15804 8718 15813
rect 8410 15802 8416 15804
rect 8472 15802 8496 15804
rect 8552 15802 8576 15804
rect 8632 15802 8656 15804
rect 8712 15802 8718 15804
rect 8472 15750 8474 15802
rect 8654 15750 8656 15802
rect 8410 15748 8416 15750
rect 8472 15748 8496 15750
rect 8552 15748 8576 15750
rect 8632 15748 8656 15750
rect 8712 15748 8718 15750
rect 8410 15739 8718 15748
rect 8410 14716 8718 14725
rect 8410 14714 8416 14716
rect 8472 14714 8496 14716
rect 8552 14714 8576 14716
rect 8632 14714 8656 14716
rect 8712 14714 8718 14716
rect 8472 14662 8474 14714
rect 8654 14662 8656 14714
rect 8410 14660 8416 14662
rect 8472 14660 8496 14662
rect 8552 14660 8576 14662
rect 8632 14660 8656 14662
rect 8712 14660 8718 14662
rect 8410 14651 8718 14660
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8410 13628 8718 13637
rect 8410 13626 8416 13628
rect 8472 13626 8496 13628
rect 8552 13626 8576 13628
rect 8632 13626 8656 13628
rect 8712 13626 8718 13628
rect 8472 13574 8474 13626
rect 8654 13574 8656 13626
rect 8410 13572 8416 13574
rect 8472 13572 8496 13574
rect 8552 13572 8576 13574
rect 8632 13572 8656 13574
rect 8712 13572 8718 13574
rect 8410 13563 8718 13572
rect 8410 12540 8718 12549
rect 8410 12538 8416 12540
rect 8472 12538 8496 12540
rect 8552 12538 8576 12540
rect 8632 12538 8656 12540
rect 8712 12538 8718 12540
rect 8472 12486 8474 12538
rect 8654 12486 8656 12538
rect 8410 12484 8416 12486
rect 8472 12484 8496 12486
rect 8552 12484 8576 12486
rect 8632 12484 8656 12486
rect 8712 12484 8718 12486
rect 8410 12475 8718 12484
rect 8410 11452 8718 11461
rect 8410 11450 8416 11452
rect 8472 11450 8496 11452
rect 8552 11450 8576 11452
rect 8632 11450 8656 11452
rect 8712 11450 8718 11452
rect 8472 11398 8474 11450
rect 8654 11398 8656 11450
rect 8410 11396 8416 11398
rect 8472 11396 8496 11398
rect 8552 11396 8576 11398
rect 8632 11396 8656 11398
rect 8712 11396 8718 11398
rect 8410 11387 8718 11396
rect 8410 10364 8718 10373
rect 8410 10362 8416 10364
rect 8472 10362 8496 10364
rect 8552 10362 8576 10364
rect 8632 10362 8656 10364
rect 8712 10362 8718 10364
rect 8472 10310 8474 10362
rect 8654 10310 8656 10362
rect 8410 10308 8416 10310
rect 8472 10308 8496 10310
rect 8552 10308 8576 10310
rect 8632 10308 8656 10310
rect 8712 10308 8718 10310
rect 8410 10299 8718 10308
rect 8772 9466 8800 14418
rect 8864 9586 8892 16458
rect 8956 12782 8984 19306
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9048 14482 9076 15506
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8772 9438 8892 9466
rect 8410 9276 8718 9285
rect 8410 9274 8416 9276
rect 8472 9274 8496 9276
rect 8552 9274 8576 9276
rect 8632 9274 8656 9276
rect 8712 9274 8718 9276
rect 8472 9222 8474 9274
rect 8654 9222 8656 9274
rect 8410 9220 8416 9222
rect 8472 9220 8496 9222
rect 8552 9220 8576 9222
rect 8632 9220 8656 9222
rect 8712 9220 8718 9222
rect 8410 9211 8718 9220
rect 8312 9030 8800 9058
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 2378 8340 8910
rect 8410 8188 8718 8197
rect 8410 8186 8416 8188
rect 8472 8186 8496 8188
rect 8552 8186 8576 8188
rect 8632 8186 8656 8188
rect 8712 8186 8718 8188
rect 8472 8134 8474 8186
rect 8654 8134 8656 8186
rect 8410 8132 8416 8134
rect 8472 8132 8496 8134
rect 8552 8132 8576 8134
rect 8632 8132 8656 8134
rect 8712 8132 8718 8134
rect 8410 8123 8718 8132
rect 8410 7100 8718 7109
rect 8410 7098 8416 7100
rect 8472 7098 8496 7100
rect 8552 7098 8576 7100
rect 8632 7098 8656 7100
rect 8712 7098 8718 7100
rect 8472 7046 8474 7098
rect 8654 7046 8656 7098
rect 8410 7044 8416 7046
rect 8472 7044 8496 7046
rect 8552 7044 8576 7046
rect 8632 7044 8656 7046
rect 8712 7044 8718 7046
rect 8410 7035 8718 7044
rect 8410 6012 8718 6021
rect 8410 6010 8416 6012
rect 8472 6010 8496 6012
rect 8552 6010 8576 6012
rect 8632 6010 8656 6012
rect 8712 6010 8718 6012
rect 8472 5958 8474 6010
rect 8654 5958 8656 6010
rect 8410 5956 8416 5958
rect 8472 5956 8496 5958
rect 8552 5956 8576 5958
rect 8632 5956 8656 5958
rect 8712 5956 8718 5958
rect 8410 5947 8718 5956
rect 8410 4924 8718 4933
rect 8410 4922 8416 4924
rect 8472 4922 8496 4924
rect 8552 4922 8576 4924
rect 8632 4922 8656 4924
rect 8712 4922 8718 4924
rect 8472 4870 8474 4922
rect 8654 4870 8656 4922
rect 8410 4868 8416 4870
rect 8472 4868 8496 4870
rect 8552 4868 8576 4870
rect 8632 4868 8656 4870
rect 8712 4868 8718 4870
rect 8410 4859 8718 4868
rect 8410 3836 8718 3845
rect 8410 3834 8416 3836
rect 8472 3834 8496 3836
rect 8552 3834 8576 3836
rect 8632 3834 8656 3836
rect 8712 3834 8718 3836
rect 8472 3782 8474 3834
rect 8654 3782 8656 3834
rect 8410 3780 8416 3782
rect 8472 3780 8496 3782
rect 8552 3780 8576 3782
rect 8632 3780 8656 3782
rect 8712 3780 8718 3782
rect 8410 3771 8718 3780
rect 8410 2748 8718 2757
rect 8410 2746 8416 2748
rect 8472 2746 8496 2748
rect 8552 2746 8576 2748
rect 8632 2746 8656 2748
rect 8712 2746 8718 2748
rect 8472 2694 8474 2746
rect 8654 2694 8656 2746
rect 8410 2692 8416 2694
rect 8472 2692 8496 2694
rect 8552 2692 8576 2694
rect 8632 2692 8656 2694
rect 8712 2692 8718 2694
rect 8410 2683 8718 2692
rect 8772 2446 8800 9030
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8410 1660 8718 1669
rect 8410 1658 8416 1660
rect 8472 1658 8496 1660
rect 8552 1658 8576 1660
rect 8632 1658 8656 1660
rect 8712 1658 8718 1660
rect 8472 1606 8474 1658
rect 8654 1606 8656 1658
rect 8410 1604 8416 1606
rect 8472 1604 8496 1606
rect 8552 1604 8576 1606
rect 8632 1604 8656 1606
rect 8712 1604 8718 1606
rect 8410 1595 8718 1604
rect 8208 808 8260 814
rect 8208 750 8260 756
rect 8864 610 8892 9438
rect 8956 2514 8984 12582
rect 9048 3942 9076 14214
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9140 3738 9168 25978
rect 9232 24342 9260 28698
rect 9600 28506 9628 29158
rect 9600 28478 9720 28506
rect 9350 28316 9658 28325
rect 9350 28314 9356 28316
rect 9412 28314 9436 28316
rect 9492 28314 9516 28316
rect 9572 28314 9596 28316
rect 9652 28314 9658 28316
rect 9412 28262 9414 28314
rect 9594 28262 9596 28314
rect 9350 28260 9356 28262
rect 9412 28260 9436 28262
rect 9492 28260 9516 28262
rect 9572 28260 9596 28262
rect 9652 28260 9658 28262
rect 9350 28251 9658 28260
rect 9350 27228 9658 27237
rect 9350 27226 9356 27228
rect 9412 27226 9436 27228
rect 9492 27226 9516 27228
rect 9572 27226 9596 27228
rect 9652 27226 9658 27228
rect 9412 27174 9414 27226
rect 9594 27174 9596 27226
rect 9350 27172 9356 27174
rect 9412 27172 9436 27174
rect 9492 27172 9516 27174
rect 9572 27172 9596 27174
rect 9652 27172 9658 27174
rect 9350 27163 9658 27172
rect 9692 27010 9720 28478
rect 9600 26982 9720 27010
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 9508 26586 9536 26794
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9600 26314 9628 26982
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9350 26140 9658 26149
rect 9350 26138 9356 26140
rect 9412 26138 9436 26140
rect 9492 26138 9516 26140
rect 9572 26138 9596 26140
rect 9652 26138 9658 26140
rect 9412 26086 9414 26138
rect 9594 26086 9596 26138
rect 9350 26084 9356 26086
rect 9412 26084 9436 26086
rect 9492 26084 9516 26086
rect 9572 26084 9596 26086
rect 9652 26084 9658 26086
rect 9350 26075 9658 26084
rect 9588 25424 9640 25430
rect 9588 25366 9640 25372
rect 9600 25242 9628 25366
rect 9600 25214 9720 25242
rect 9350 25052 9658 25061
rect 9350 25050 9356 25052
rect 9412 25050 9436 25052
rect 9492 25050 9516 25052
rect 9572 25050 9596 25052
rect 9652 25050 9658 25052
rect 9412 24998 9414 25050
rect 9594 24998 9596 25050
rect 9350 24996 9356 24998
rect 9412 24996 9436 24998
rect 9492 24996 9516 24998
rect 9572 24996 9596 24998
rect 9652 24996 9658 24998
rect 9350 24987 9658 24996
rect 9692 24834 9720 25214
rect 9600 24806 9720 24834
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 9324 24052 9352 24686
rect 9600 24154 9628 24806
rect 9600 24126 9720 24154
rect 9232 24024 9352 24052
rect 9232 23322 9260 24024
rect 9350 23964 9658 23973
rect 9350 23962 9356 23964
rect 9412 23962 9436 23964
rect 9492 23962 9516 23964
rect 9572 23962 9596 23964
rect 9652 23962 9658 23964
rect 9412 23910 9414 23962
rect 9594 23910 9596 23962
rect 9350 23908 9356 23910
rect 9412 23908 9436 23910
rect 9492 23908 9516 23910
rect 9572 23908 9596 23910
rect 9652 23908 9658 23910
rect 9350 23899 9658 23908
rect 9692 23746 9720 24126
rect 9600 23718 9720 23746
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9324 23202 9352 23598
rect 9232 23174 9352 23202
rect 9232 15570 9260 23174
rect 9600 23050 9628 23718
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9350 22876 9658 22885
rect 9350 22874 9356 22876
rect 9412 22874 9436 22876
rect 9492 22874 9516 22876
rect 9572 22874 9596 22876
rect 9652 22874 9658 22876
rect 9412 22822 9414 22874
rect 9594 22822 9596 22874
rect 9350 22820 9356 22822
rect 9412 22820 9436 22822
rect 9492 22820 9516 22822
rect 9572 22820 9596 22822
rect 9652 22820 9658 22822
rect 9350 22811 9658 22820
rect 9350 21788 9658 21797
rect 9350 21786 9356 21788
rect 9412 21786 9436 21788
rect 9492 21786 9516 21788
rect 9572 21786 9596 21788
rect 9652 21786 9658 21788
rect 9412 21734 9414 21786
rect 9594 21734 9596 21786
rect 9350 21732 9356 21734
rect 9412 21732 9436 21734
rect 9492 21732 9516 21734
rect 9572 21732 9596 21734
rect 9652 21732 9658 21734
rect 9350 21723 9658 21732
rect 9350 20700 9658 20709
rect 9350 20698 9356 20700
rect 9412 20698 9436 20700
rect 9492 20698 9516 20700
rect 9572 20698 9596 20700
rect 9652 20698 9658 20700
rect 9412 20646 9414 20698
rect 9594 20646 9596 20698
rect 9350 20644 9356 20646
rect 9412 20644 9436 20646
rect 9492 20644 9516 20646
rect 9572 20644 9596 20646
rect 9652 20644 9658 20646
rect 9350 20635 9658 20644
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9600 19802 9628 20198
rect 9600 19774 9720 19802
rect 9350 19612 9658 19621
rect 9350 19610 9356 19612
rect 9412 19610 9436 19612
rect 9492 19610 9516 19612
rect 9572 19610 9596 19612
rect 9652 19610 9658 19612
rect 9412 19558 9414 19610
rect 9594 19558 9596 19610
rect 9350 19556 9356 19558
rect 9412 19556 9436 19558
rect 9492 19556 9516 19558
rect 9572 19556 9596 19558
rect 9652 19556 9658 19558
rect 9350 19547 9658 19556
rect 9692 19394 9720 19774
rect 9600 19366 9720 19394
rect 9600 18714 9628 19366
rect 9600 18686 9720 18714
rect 9350 18524 9658 18533
rect 9350 18522 9356 18524
rect 9412 18522 9436 18524
rect 9492 18522 9516 18524
rect 9572 18522 9596 18524
rect 9652 18522 9658 18524
rect 9412 18470 9414 18522
rect 9594 18470 9596 18522
rect 9350 18468 9356 18470
rect 9412 18468 9436 18470
rect 9492 18468 9516 18470
rect 9572 18468 9596 18470
rect 9652 18468 9658 18470
rect 9350 18459 9658 18468
rect 9692 18340 9720 18686
rect 9600 18312 9720 18340
rect 9600 17626 9628 18312
rect 9600 17598 9720 17626
rect 9350 17436 9658 17445
rect 9350 17434 9356 17436
rect 9412 17434 9436 17436
rect 9492 17434 9516 17436
rect 9572 17434 9596 17436
rect 9652 17434 9658 17436
rect 9412 17382 9414 17434
rect 9594 17382 9596 17434
rect 9350 17380 9356 17382
rect 9412 17380 9436 17382
rect 9492 17380 9516 17382
rect 9572 17380 9596 17382
rect 9652 17380 9658 17382
rect 9350 17371 9658 17380
rect 9692 17218 9720 17598
rect 9600 17190 9720 17218
rect 9600 16538 9628 17190
rect 9600 16510 9720 16538
rect 9350 16348 9658 16357
rect 9350 16346 9356 16348
rect 9412 16346 9436 16348
rect 9492 16346 9516 16348
rect 9572 16346 9596 16348
rect 9652 16346 9658 16348
rect 9412 16294 9414 16346
rect 9594 16294 9596 16346
rect 9350 16292 9356 16294
rect 9412 16292 9436 16294
rect 9492 16292 9516 16294
rect 9572 16292 9596 16294
rect 9652 16292 9658 16294
rect 9350 16283 9658 16292
rect 9692 16130 9720 16510
rect 9600 16102 9720 16130
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9600 15450 9628 16102
rect 9600 15422 9720 15450
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9232 12866 9260 15302
rect 9350 15260 9658 15269
rect 9350 15258 9356 15260
rect 9412 15258 9436 15260
rect 9492 15258 9516 15260
rect 9572 15258 9596 15260
rect 9652 15258 9658 15260
rect 9412 15206 9414 15258
rect 9594 15206 9596 15258
rect 9350 15204 9356 15206
rect 9412 15204 9436 15206
rect 9492 15204 9516 15206
rect 9572 15204 9596 15206
rect 9652 15204 9658 15206
rect 9350 15195 9658 15204
rect 9692 15042 9720 15422
rect 9600 15014 9720 15042
rect 9600 14362 9628 15014
rect 9784 14414 9812 37198
rect 9876 32842 9904 55218
rect 9968 46578 9996 55406
rect 10060 53174 10088 62630
rect 10048 53168 10100 53174
rect 10048 53110 10100 53116
rect 10152 52018 10180 64874
rect 10244 53786 10272 65010
rect 10336 58614 10364 65282
rect 10428 64462 10456 86974
rect 10508 86896 10560 86902
rect 10508 86838 10560 86844
rect 10520 73166 10548 86838
rect 10600 86624 10652 86630
rect 10600 86566 10652 86572
rect 10508 73160 10560 73166
rect 10508 73102 10560 73108
rect 10506 69320 10562 69329
rect 10506 69255 10562 69264
rect 10520 66450 10548 69255
rect 10612 67046 10640 86566
rect 10692 84856 10744 84862
rect 10692 84798 10744 84804
rect 10600 67040 10652 67046
rect 10600 66982 10652 66988
rect 10704 66638 10732 84798
rect 10796 69562 10824 87042
rect 10950 85980 11258 85989
rect 10950 85978 10956 85980
rect 11012 85978 11036 85980
rect 11092 85978 11116 85980
rect 11172 85978 11196 85980
rect 11252 85978 11258 85980
rect 11012 85926 11014 85978
rect 11194 85926 11196 85978
rect 10950 85924 10956 85926
rect 11012 85924 11036 85926
rect 11092 85924 11116 85926
rect 11172 85924 11196 85926
rect 11252 85924 11258 85926
rect 10950 85915 11258 85924
rect 10876 84924 10928 84930
rect 10876 84866 10928 84872
rect 10888 71738 10916 84866
rect 10968 83564 11020 83570
rect 10968 83506 11020 83512
rect 10876 71732 10928 71738
rect 10876 71674 10928 71680
rect 10876 69964 10928 69970
rect 10876 69906 10928 69912
rect 10784 69556 10836 69562
rect 10784 69498 10836 69504
rect 10784 67652 10836 67658
rect 10784 67594 10836 67600
rect 10692 66632 10744 66638
rect 10692 66574 10744 66580
rect 10520 66422 10732 66450
rect 10416 64456 10468 64462
rect 10416 64398 10468 64404
rect 10600 63980 10652 63986
rect 10600 63922 10652 63928
rect 10416 63572 10468 63578
rect 10416 63514 10468 63520
rect 10324 58608 10376 58614
rect 10324 58550 10376 58556
rect 10428 55162 10456 63514
rect 10612 55162 10640 63922
rect 10336 55134 10456 55162
rect 10520 55134 10640 55162
rect 10232 53780 10284 53786
rect 10232 53722 10284 53728
rect 10140 52012 10192 52018
rect 10140 51954 10192 51960
rect 9956 46572 10008 46578
rect 9956 46514 10008 46520
rect 9968 42362 9996 46514
rect 9956 42356 10008 42362
rect 9956 42298 10008 42304
rect 10048 42220 10100 42226
rect 10048 42162 10100 42168
rect 9956 40112 10008 40118
rect 9956 40054 10008 40060
rect 9864 32836 9916 32842
rect 9864 32778 9916 32784
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 9876 16590 9904 29174
rect 9968 22642 9996 40054
rect 10060 31754 10088 42162
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 10060 23254 10088 26726
rect 10152 26586 10180 31962
rect 10336 29753 10364 55134
rect 10520 55026 10548 55134
rect 10428 54998 10548 55026
rect 10428 31521 10456 54998
rect 10704 54890 10732 66422
rect 10520 54862 10732 54890
rect 10520 38185 10548 54862
rect 10796 54262 10824 67594
rect 10888 58546 10916 69906
rect 10980 69766 11008 83506
rect 11348 71738 11376 87246
rect 17316 87236 17368 87242
rect 17316 87178 17368 87184
rect 11428 86964 11480 86970
rect 11428 86906 11480 86912
rect 11336 71732 11388 71738
rect 11336 71674 11388 71680
rect 11152 71528 11204 71534
rect 11152 71470 11204 71476
rect 10968 69760 11020 69766
rect 10968 69702 11020 69708
rect 10980 66230 11008 69702
rect 10968 66224 11020 66230
rect 10968 66166 11020 66172
rect 11164 65006 11192 71470
rect 11244 71392 11296 71398
rect 11244 71334 11296 71340
rect 11152 65000 11204 65006
rect 11152 64942 11204 64948
rect 11152 59424 11204 59430
rect 11152 59366 11204 59372
rect 10876 58540 10928 58546
rect 10876 58482 10928 58488
rect 11060 56772 11112 56778
rect 11060 56714 11112 56720
rect 10784 54256 10836 54262
rect 10784 54198 10836 54204
rect 10506 38176 10562 38185
rect 10506 38111 10562 38120
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10508 33040 10560 33046
rect 10508 32982 10560 32988
rect 10414 31512 10470 31521
rect 10414 31447 10470 31456
rect 10322 29744 10378 29753
rect 10322 29679 10378 29688
rect 10324 28688 10376 28694
rect 10324 28630 10376 28636
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10048 23248 10100 23254
rect 10048 23190 10100 23196
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 14408 9824 14414
rect 9600 14334 9720 14362
rect 9772 14350 9824 14356
rect 9350 14172 9658 14181
rect 9350 14170 9356 14172
rect 9412 14170 9436 14172
rect 9492 14170 9516 14172
rect 9572 14170 9596 14172
rect 9652 14170 9658 14172
rect 9412 14118 9414 14170
rect 9594 14118 9596 14170
rect 9350 14116 9356 14118
rect 9412 14116 9436 14118
rect 9492 14116 9516 14118
rect 9572 14116 9596 14118
rect 9652 14116 9658 14118
rect 9350 14107 9658 14116
rect 9692 13954 9720 14334
rect 9600 13926 9720 13954
rect 9600 13274 9628 13926
rect 9600 13246 9720 13274
rect 9350 13084 9658 13093
rect 9350 13082 9356 13084
rect 9412 13082 9436 13084
rect 9492 13082 9516 13084
rect 9572 13082 9596 13084
rect 9652 13082 9658 13084
rect 9412 13030 9414 13082
rect 9594 13030 9596 13082
rect 9350 13028 9356 13030
rect 9412 13028 9436 13030
rect 9492 13028 9516 13030
rect 9572 13028 9596 13030
rect 9652 13028 9658 13030
rect 9350 13019 9658 13028
rect 9232 12838 9628 12866
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9232 2038 9260 12718
rect 9600 12186 9628 12838
rect 9692 12646 9720 13246
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9600 12158 9720 12186
rect 9350 11996 9658 12005
rect 9350 11994 9356 11996
rect 9412 11994 9436 11996
rect 9492 11994 9516 11996
rect 9572 11994 9596 11996
rect 9652 11994 9658 11996
rect 9412 11942 9414 11994
rect 9594 11942 9596 11994
rect 9350 11940 9356 11942
rect 9412 11940 9436 11942
rect 9492 11940 9516 11942
rect 9572 11940 9596 11942
rect 9652 11940 9658 11942
rect 9350 11931 9658 11940
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9600 11257 9628 11290
rect 9586 11248 9642 11257
rect 9586 11183 9642 11192
rect 9350 10908 9658 10917
rect 9350 10906 9356 10908
rect 9412 10906 9436 10908
rect 9492 10906 9516 10908
rect 9572 10906 9596 10908
rect 9652 10906 9658 10908
rect 9412 10854 9414 10906
rect 9594 10854 9596 10906
rect 9350 10852 9356 10854
rect 9412 10852 9436 10854
rect 9492 10852 9516 10854
rect 9572 10852 9596 10854
rect 9652 10852 9658 10854
rect 9350 10843 9658 10852
rect 9692 10690 9720 12158
rect 9600 10662 9720 10690
rect 9600 10010 9628 10662
rect 9600 9982 9720 10010
rect 9350 9820 9658 9829
rect 9350 9818 9356 9820
rect 9412 9818 9436 9820
rect 9492 9818 9516 9820
rect 9572 9818 9596 9820
rect 9652 9818 9658 9820
rect 9412 9766 9414 9818
rect 9594 9766 9596 9818
rect 9350 9764 9356 9766
rect 9412 9764 9436 9766
rect 9492 9764 9516 9766
rect 9572 9764 9596 9766
rect 9652 9764 9658 9766
rect 9350 9755 9658 9764
rect 9692 9628 9720 9982
rect 9600 9600 9720 9628
rect 9600 8974 9628 9600
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9350 8732 9658 8741
rect 9350 8730 9356 8732
rect 9412 8730 9436 8732
rect 9492 8730 9516 8732
rect 9572 8730 9596 8732
rect 9652 8730 9658 8732
rect 9412 8678 9414 8730
rect 9594 8678 9596 8730
rect 9350 8676 9356 8678
rect 9412 8676 9436 8678
rect 9492 8676 9516 8678
rect 9572 8676 9596 8678
rect 9652 8676 9658 8678
rect 9350 8667 9658 8676
rect 9350 7644 9658 7653
rect 9350 7642 9356 7644
rect 9412 7642 9436 7644
rect 9492 7642 9516 7644
rect 9572 7642 9596 7644
rect 9652 7642 9658 7644
rect 9412 7590 9414 7642
rect 9594 7590 9596 7642
rect 9350 7588 9356 7590
rect 9412 7588 9436 7590
rect 9492 7588 9516 7590
rect 9572 7588 9596 7590
rect 9652 7588 9658 7590
rect 9350 7579 9658 7588
rect 9350 6556 9658 6565
rect 9350 6554 9356 6556
rect 9412 6554 9436 6556
rect 9492 6554 9516 6556
rect 9572 6554 9596 6556
rect 9652 6554 9658 6556
rect 9412 6502 9414 6554
rect 9594 6502 9596 6554
rect 9350 6500 9356 6502
rect 9412 6500 9436 6502
rect 9492 6500 9516 6502
rect 9572 6500 9596 6502
rect 9652 6500 9658 6502
rect 9350 6491 9658 6500
rect 9350 5468 9658 5477
rect 9350 5466 9356 5468
rect 9412 5466 9436 5468
rect 9492 5466 9516 5468
rect 9572 5466 9596 5468
rect 9652 5466 9658 5468
rect 9412 5414 9414 5466
rect 9594 5414 9596 5466
rect 9350 5412 9356 5414
rect 9412 5412 9436 5414
rect 9492 5412 9516 5414
rect 9572 5412 9596 5414
rect 9652 5412 9658 5414
rect 9350 5403 9658 5412
rect 9350 4380 9658 4389
rect 9350 4378 9356 4380
rect 9412 4378 9436 4380
rect 9492 4378 9516 4380
rect 9572 4378 9596 4380
rect 9652 4378 9658 4380
rect 9412 4326 9414 4378
rect 9594 4326 9596 4378
rect 9350 4324 9356 4326
rect 9412 4324 9436 4326
rect 9492 4324 9516 4326
rect 9572 4324 9596 4326
rect 9652 4324 9658 4326
rect 9350 4315 9658 4324
rect 9350 3292 9658 3301
rect 9350 3290 9356 3292
rect 9412 3290 9436 3292
rect 9492 3290 9516 3292
rect 9572 3290 9596 3292
rect 9652 3290 9658 3292
rect 9412 3238 9414 3290
rect 9594 3238 9596 3290
rect 9350 3236 9356 3238
rect 9412 3236 9436 3238
rect 9492 3236 9516 3238
rect 9572 3236 9596 3238
rect 9652 3236 9658 3238
rect 9350 3227 9658 3236
rect 9350 2204 9658 2213
rect 9350 2202 9356 2204
rect 9412 2202 9436 2204
rect 9492 2202 9516 2204
rect 9572 2202 9596 2204
rect 9652 2202 9658 2204
rect 9412 2150 9414 2202
rect 9594 2150 9596 2202
rect 9350 2148 9356 2150
rect 9412 2148 9436 2150
rect 9492 2148 9516 2150
rect 9572 2148 9596 2150
rect 9652 2148 9658 2150
rect 9350 2139 9658 2148
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9350 1116 9658 1125
rect 9350 1114 9356 1116
rect 9412 1114 9436 1116
rect 9492 1114 9516 1116
rect 9572 1114 9596 1116
rect 9652 1114 9658 1116
rect 9412 1062 9414 1114
rect 9594 1062 9596 1114
rect 9350 1060 9356 1062
rect 9412 1060 9436 1062
rect 9492 1060 9516 1062
rect 9572 1060 9596 1062
rect 9652 1060 9658 1062
rect 9350 1051 9658 1060
rect 8852 604 8904 610
rect 8852 546 8904 552
rect 7656 536 7708 542
rect 7656 478 7708 484
rect 1306 368 1362 377
rect 9876 338 9904 16186
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 3398 10272 11222
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10336 3330 10364 28630
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10324 3324 10376 3330
rect 10324 3266 10376 3272
rect 10010 1660 10318 1669
rect 10010 1658 10016 1660
rect 10072 1658 10096 1660
rect 10152 1658 10176 1660
rect 10232 1658 10256 1660
rect 10312 1658 10318 1660
rect 10072 1606 10074 1658
rect 10254 1606 10256 1658
rect 10010 1604 10016 1606
rect 10072 1604 10096 1606
rect 10152 1604 10176 1606
rect 10232 1604 10256 1606
rect 10312 1604 10318 1606
rect 10010 1595 10318 1604
rect 10428 678 10456 26250
rect 10416 672 10468 678
rect 10416 614 10468 620
rect 10520 474 10548 32982
rect 10600 32360 10652 32366
rect 10600 32302 10652 32308
rect 10612 513 10640 32302
rect 10704 3369 10732 34682
rect 10784 32224 10836 32230
rect 10784 32166 10836 32172
rect 10796 3806 10824 32166
rect 11072 24818 11100 56714
rect 11164 46646 11192 59366
rect 11256 57934 11284 71334
rect 11348 70514 11376 71674
rect 11440 70582 11468 86906
rect 11520 86692 11572 86698
rect 11520 86634 11572 86640
rect 11428 70576 11480 70582
rect 11428 70518 11480 70524
rect 11336 70508 11388 70514
rect 11336 70450 11388 70456
rect 11532 70378 11560 86634
rect 11610 86524 11918 86533
rect 11610 86522 11616 86524
rect 11672 86522 11696 86524
rect 11752 86522 11776 86524
rect 11832 86522 11856 86524
rect 11912 86522 11918 86524
rect 11672 86470 11674 86522
rect 11854 86470 11856 86522
rect 11610 86468 11616 86470
rect 11672 86468 11696 86470
rect 11752 86468 11776 86470
rect 11832 86468 11856 86470
rect 11912 86468 11918 86470
rect 11610 86459 11918 86468
rect 13210 86524 13518 86533
rect 13210 86522 13216 86524
rect 13272 86522 13296 86524
rect 13352 86522 13376 86524
rect 13432 86522 13456 86524
rect 13512 86522 13518 86524
rect 13272 86470 13274 86522
rect 13454 86470 13456 86522
rect 13210 86468 13216 86470
rect 13272 86468 13296 86470
rect 13352 86468 13376 86470
rect 13432 86468 13456 86470
rect 13512 86468 13518 86470
rect 13210 86459 13518 86468
rect 14810 86524 15118 86533
rect 14810 86522 14816 86524
rect 14872 86522 14896 86524
rect 14952 86522 14976 86524
rect 15032 86522 15056 86524
rect 15112 86522 15118 86524
rect 14872 86470 14874 86522
rect 15054 86470 15056 86522
rect 14810 86468 14816 86470
rect 14872 86468 14896 86470
rect 14952 86468 14976 86470
rect 15032 86468 15056 86470
rect 15112 86468 15118 86470
rect 14810 86459 15118 86468
rect 16410 86524 16718 86533
rect 16410 86522 16416 86524
rect 16472 86522 16496 86524
rect 16552 86522 16576 86524
rect 16632 86522 16656 86524
rect 16712 86522 16718 86524
rect 16472 86470 16474 86522
rect 16654 86470 16656 86522
rect 16410 86468 16416 86470
rect 16472 86468 16496 86470
rect 16552 86468 16576 86470
rect 16632 86468 16656 86470
rect 16712 86468 16718 86470
rect 16410 86459 16718 86468
rect 13728 86420 13780 86426
rect 13728 86362 13780 86368
rect 11980 86148 12032 86154
rect 11980 86090 12032 86096
rect 11704 85400 11756 85406
rect 11704 85342 11756 85348
rect 11520 70372 11572 70378
rect 11520 70314 11572 70320
rect 11520 68196 11572 68202
rect 11520 68138 11572 68144
rect 11428 66496 11480 66502
rect 11428 66438 11480 66444
rect 11336 62144 11388 62150
rect 11336 62086 11388 62092
rect 11244 57928 11296 57934
rect 11244 57870 11296 57876
rect 11348 49230 11376 62086
rect 11440 53786 11468 66438
rect 11532 54058 11560 68138
rect 11716 64122 11744 85342
rect 11796 84788 11848 84794
rect 11796 84730 11848 84736
rect 11808 68270 11836 84730
rect 11888 84720 11940 84726
rect 11888 84662 11940 84668
rect 11900 68338 11928 84662
rect 11888 68332 11940 68338
rect 11888 68274 11940 68280
rect 11796 68264 11848 68270
rect 11796 68206 11848 68212
rect 11886 65104 11942 65113
rect 11886 65039 11942 65048
rect 11704 64116 11756 64122
rect 11704 64058 11756 64064
rect 11612 59696 11664 59702
rect 11612 59638 11664 59644
rect 11520 54052 11572 54058
rect 11520 53994 11572 54000
rect 11428 53780 11480 53786
rect 11428 53722 11480 53728
rect 11336 49224 11388 49230
rect 11336 49166 11388 49172
rect 11152 46640 11204 46646
rect 11152 46582 11204 46588
rect 11520 38480 11572 38486
rect 11520 38422 11572 38428
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10784 3800 10836 3806
rect 10784 3742 10836 3748
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 10888 2174 10916 24346
rect 11428 23316 11480 23322
rect 11428 23258 11480 23264
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 3534 11008 13126
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 11348 9625 11376 11183
rect 11334 9616 11390 9625
rect 11334 9551 11390 9560
rect 11440 3874 11468 23258
rect 11428 3868 11480 3874
rect 11428 3810 11480 3816
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10876 2168 10928 2174
rect 10876 2110 10928 2116
rect 11532 1358 11560 38422
rect 11624 36922 11652 59638
rect 11900 41414 11928 65039
rect 11992 59430 12020 86090
rect 12550 85980 12858 85989
rect 12550 85978 12556 85980
rect 12612 85978 12636 85980
rect 12692 85978 12716 85980
rect 12772 85978 12796 85980
rect 12852 85978 12858 85980
rect 12612 85926 12614 85978
rect 12794 85926 12796 85978
rect 12550 85924 12556 85926
rect 12612 85924 12636 85926
rect 12692 85924 12716 85926
rect 12772 85924 12796 85926
rect 12852 85924 12858 85926
rect 12550 85915 12858 85924
rect 13740 85678 13768 86362
rect 16960 86290 17264 86306
rect 16948 86284 17276 86290
rect 17000 86278 17224 86284
rect 16948 86226 17000 86232
rect 17224 86226 17276 86232
rect 17328 86154 17356 87178
rect 24768 87168 24820 87174
rect 24768 87110 24820 87116
rect 18010 86524 18318 86533
rect 18010 86522 18016 86524
rect 18072 86522 18096 86524
rect 18152 86522 18176 86524
rect 18232 86522 18256 86524
rect 18312 86522 18318 86524
rect 18072 86470 18074 86522
rect 18254 86470 18256 86522
rect 18010 86468 18016 86470
rect 18072 86468 18096 86470
rect 18152 86468 18176 86470
rect 18232 86468 18256 86470
rect 18312 86468 18318 86470
rect 18010 86459 18318 86468
rect 19610 86524 19918 86533
rect 19610 86522 19616 86524
rect 19672 86522 19696 86524
rect 19752 86522 19776 86524
rect 19832 86522 19856 86524
rect 19912 86522 19918 86524
rect 19672 86470 19674 86522
rect 19854 86470 19856 86522
rect 19610 86468 19616 86470
rect 19672 86468 19696 86470
rect 19752 86468 19776 86470
rect 19832 86468 19856 86470
rect 19912 86468 19918 86470
rect 19610 86459 19918 86468
rect 21210 86524 21518 86533
rect 21210 86522 21216 86524
rect 21272 86522 21296 86524
rect 21352 86522 21376 86524
rect 21432 86522 21456 86524
rect 21512 86522 21518 86524
rect 21272 86470 21274 86522
rect 21454 86470 21456 86522
rect 21210 86468 21216 86470
rect 21272 86468 21296 86470
rect 21352 86468 21376 86470
rect 21432 86468 21456 86470
rect 21512 86468 21518 86470
rect 21210 86459 21518 86468
rect 22810 86524 23118 86533
rect 22810 86522 22816 86524
rect 22872 86522 22896 86524
rect 22952 86522 22976 86524
rect 23032 86522 23056 86524
rect 23112 86522 23118 86524
rect 22872 86470 22874 86522
rect 23054 86470 23056 86522
rect 22810 86468 22816 86470
rect 22872 86468 22896 86470
rect 22952 86468 22976 86470
rect 23032 86468 23056 86470
rect 23112 86468 23118 86470
rect 22810 86459 23118 86468
rect 24410 86524 24718 86533
rect 24410 86522 24416 86524
rect 24472 86522 24496 86524
rect 24552 86522 24576 86524
rect 24632 86522 24656 86524
rect 24712 86522 24718 86524
rect 24472 86470 24474 86522
rect 24654 86470 24656 86522
rect 24410 86468 24416 86470
rect 24472 86468 24496 86470
rect 24552 86468 24576 86470
rect 24632 86468 24656 86470
rect 24712 86468 24718 86470
rect 24410 86459 24718 86468
rect 24780 86154 24808 87110
rect 26010 86524 26318 86533
rect 26010 86522 26016 86524
rect 26072 86522 26096 86524
rect 26152 86522 26176 86524
rect 26232 86522 26256 86524
rect 26312 86522 26318 86524
rect 26072 86470 26074 86522
rect 26254 86470 26256 86522
rect 26010 86468 26016 86470
rect 26072 86468 26096 86470
rect 26152 86468 26176 86470
rect 26232 86468 26256 86470
rect 26312 86468 26318 86470
rect 26010 86459 26318 86468
rect 25044 86284 25096 86290
rect 25044 86226 25096 86232
rect 27160 86284 27212 86290
rect 27160 86226 27212 86232
rect 17316 86148 17368 86154
rect 17316 86090 17368 86096
rect 19708 86148 19760 86154
rect 19708 86090 19760 86096
rect 19800 86148 19852 86154
rect 19800 86090 19852 86096
rect 19984 86148 20036 86154
rect 19984 86090 20036 86096
rect 24768 86148 24820 86154
rect 24768 86090 24820 86096
rect 14150 85980 14458 85989
rect 14150 85978 14156 85980
rect 14212 85978 14236 85980
rect 14292 85978 14316 85980
rect 14372 85978 14396 85980
rect 14452 85978 14458 85980
rect 14212 85926 14214 85978
rect 14394 85926 14396 85978
rect 14150 85924 14156 85926
rect 14212 85924 14236 85926
rect 14292 85924 14316 85926
rect 14372 85924 14396 85926
rect 14452 85924 14458 85926
rect 14150 85915 14458 85924
rect 15750 85980 16058 85989
rect 15750 85978 15756 85980
rect 15812 85978 15836 85980
rect 15892 85978 15916 85980
rect 15972 85978 15996 85980
rect 16052 85978 16058 85980
rect 15812 85926 15814 85978
rect 15994 85926 15996 85978
rect 15750 85924 15756 85926
rect 15812 85924 15836 85926
rect 15892 85924 15916 85926
rect 15972 85924 15996 85926
rect 16052 85924 16058 85926
rect 15750 85915 16058 85924
rect 17350 85980 17658 85989
rect 17350 85978 17356 85980
rect 17412 85978 17436 85980
rect 17492 85978 17516 85980
rect 17572 85978 17596 85980
rect 17652 85978 17658 85980
rect 17412 85926 17414 85978
rect 17594 85926 17596 85978
rect 17350 85924 17356 85926
rect 17412 85924 17436 85926
rect 17492 85924 17516 85926
rect 17572 85924 17596 85926
rect 17652 85924 17658 85926
rect 17350 85915 17658 85924
rect 18950 85980 19258 85989
rect 18950 85978 18956 85980
rect 19012 85978 19036 85980
rect 19092 85978 19116 85980
rect 19172 85978 19196 85980
rect 19252 85978 19258 85980
rect 19012 85926 19014 85978
rect 19194 85926 19196 85978
rect 18950 85924 18956 85926
rect 19012 85924 19036 85926
rect 19092 85924 19116 85926
rect 19172 85924 19196 85926
rect 19252 85924 19258 85926
rect 18950 85915 19258 85924
rect 19720 85678 19748 86090
rect 19812 85814 19840 86090
rect 19800 85808 19852 85814
rect 19800 85750 19852 85756
rect 19996 85746 20024 86090
rect 24952 86080 25004 86086
rect 24952 86022 25004 86028
rect 20550 85980 20858 85989
rect 20550 85978 20556 85980
rect 20612 85978 20636 85980
rect 20692 85978 20716 85980
rect 20772 85978 20796 85980
rect 20852 85978 20858 85980
rect 20612 85926 20614 85978
rect 20794 85926 20796 85978
rect 20550 85924 20556 85926
rect 20612 85924 20636 85926
rect 20692 85924 20716 85926
rect 20772 85924 20796 85926
rect 20852 85924 20858 85926
rect 20550 85915 20858 85924
rect 22150 85980 22458 85989
rect 22150 85978 22156 85980
rect 22212 85978 22236 85980
rect 22292 85978 22316 85980
rect 22372 85978 22396 85980
rect 22452 85978 22458 85980
rect 22212 85926 22214 85978
rect 22394 85926 22396 85978
rect 22150 85924 22156 85926
rect 22212 85924 22236 85926
rect 22292 85924 22316 85926
rect 22372 85924 22396 85926
rect 22452 85924 22458 85926
rect 22150 85915 22458 85924
rect 23750 85980 24058 85989
rect 23750 85978 23756 85980
rect 23812 85978 23836 85980
rect 23892 85978 23916 85980
rect 23972 85978 23996 85980
rect 24052 85978 24058 85980
rect 23812 85926 23814 85978
rect 23994 85926 23996 85978
rect 23750 85924 23756 85926
rect 23812 85924 23836 85926
rect 23892 85924 23916 85926
rect 23972 85924 23996 85926
rect 24052 85924 24058 85926
rect 23750 85915 24058 85924
rect 24964 85746 24992 86022
rect 25056 85882 25084 86226
rect 26792 86216 26844 86222
rect 27172 86170 27200 86226
rect 26844 86164 27200 86170
rect 26792 86158 27200 86164
rect 26804 86142 27200 86158
rect 27264 86142 27384 86170
rect 27264 86086 27292 86142
rect 26792 86080 26844 86086
rect 26792 86022 26844 86028
rect 27252 86080 27304 86086
rect 27252 86022 27304 86028
rect 25350 85980 25658 85989
rect 25350 85978 25356 85980
rect 25412 85978 25436 85980
rect 25492 85978 25516 85980
rect 25572 85978 25596 85980
rect 25652 85978 25658 85980
rect 25412 85926 25414 85978
rect 25594 85926 25596 85978
rect 25350 85924 25356 85926
rect 25412 85924 25436 85926
rect 25492 85924 25516 85926
rect 25572 85924 25596 85926
rect 25652 85924 25658 85926
rect 25350 85915 25658 85924
rect 25044 85876 25096 85882
rect 25044 85818 25096 85824
rect 19984 85740 20036 85746
rect 19984 85682 20036 85688
rect 24952 85740 25004 85746
rect 24952 85682 25004 85688
rect 13728 85672 13780 85678
rect 13728 85614 13780 85620
rect 19708 85672 19760 85678
rect 19708 85614 19760 85620
rect 26804 85626 26832 86022
rect 26950 85980 27258 85989
rect 26950 85978 26956 85980
rect 27012 85978 27036 85980
rect 27092 85978 27116 85980
rect 27172 85978 27196 85980
rect 27252 85978 27258 85980
rect 27012 85926 27014 85978
rect 27194 85926 27196 85978
rect 26950 85924 26956 85926
rect 27012 85924 27036 85926
rect 27092 85924 27116 85926
rect 27172 85924 27196 85926
rect 27252 85924 27258 85926
rect 26950 85915 27258 85924
rect 26976 85672 27028 85678
rect 26804 85620 26976 85626
rect 26804 85614 27028 85620
rect 26804 85610 27016 85614
rect 26792 85604 27016 85610
rect 26844 85598 27016 85604
rect 26792 85546 26844 85552
rect 27356 84658 27384 86142
rect 27540 86086 27568 87518
rect 33876 87508 33928 87514
rect 33876 87450 33928 87456
rect 30196 87304 30248 87310
rect 30196 87246 30248 87252
rect 30380 87304 30432 87310
rect 30380 87246 30432 87252
rect 27610 86524 27918 86533
rect 27610 86522 27616 86524
rect 27672 86522 27696 86524
rect 27752 86522 27776 86524
rect 27832 86522 27856 86524
rect 27912 86522 27918 86524
rect 27672 86470 27674 86522
rect 27854 86470 27856 86522
rect 27610 86468 27616 86470
rect 27672 86468 27696 86470
rect 27752 86468 27776 86470
rect 27832 86468 27856 86470
rect 27912 86468 27918 86470
rect 27610 86459 27918 86468
rect 29210 86524 29518 86533
rect 29210 86522 29216 86524
rect 29272 86522 29296 86524
rect 29352 86522 29376 86524
rect 29432 86522 29456 86524
rect 29512 86522 29518 86524
rect 29272 86470 29274 86522
rect 29454 86470 29456 86522
rect 29210 86468 29216 86470
rect 29272 86468 29296 86470
rect 29352 86468 29376 86470
rect 29432 86468 29456 86470
rect 29512 86468 29518 86470
rect 29210 86459 29518 86468
rect 27620 86216 27672 86222
rect 27620 86158 27672 86164
rect 30012 86216 30064 86222
rect 30012 86158 30064 86164
rect 27632 86086 27660 86158
rect 27528 86080 27580 86086
rect 27528 86022 27580 86028
rect 27620 86080 27672 86086
rect 27620 86022 27672 86028
rect 27632 85882 27660 86022
rect 28550 85980 28858 85989
rect 28550 85978 28556 85980
rect 28612 85978 28636 85980
rect 28692 85978 28716 85980
rect 28772 85978 28796 85980
rect 28852 85978 28858 85980
rect 28612 85926 28614 85978
rect 28794 85926 28796 85978
rect 28550 85924 28556 85926
rect 28612 85924 28636 85926
rect 28692 85924 28716 85926
rect 28772 85924 28796 85926
rect 28852 85924 28858 85926
rect 28550 85915 28858 85924
rect 30024 85882 30052 86158
rect 30208 86154 30236 87246
rect 30196 86148 30248 86154
rect 30196 86090 30248 86096
rect 30392 86086 30420 87246
rect 30810 86524 31118 86533
rect 30810 86522 30816 86524
rect 30872 86522 30896 86524
rect 30952 86522 30976 86524
rect 31032 86522 31056 86524
rect 31112 86522 31118 86524
rect 30872 86470 30874 86522
rect 31054 86470 31056 86522
rect 30810 86468 30816 86470
rect 30872 86468 30896 86470
rect 30952 86468 30976 86470
rect 31032 86468 31056 86470
rect 31112 86468 31118 86470
rect 30810 86459 31118 86468
rect 32410 86524 32718 86533
rect 32410 86522 32416 86524
rect 32472 86522 32496 86524
rect 32552 86522 32576 86524
rect 32632 86522 32656 86524
rect 32712 86522 32718 86524
rect 32472 86470 32474 86522
rect 32654 86470 32656 86522
rect 32410 86468 32416 86470
rect 32472 86468 32496 86470
rect 32552 86468 32576 86470
rect 32632 86468 32656 86470
rect 32712 86468 32718 86470
rect 32410 86459 32718 86468
rect 33888 86340 33916 87450
rect 35348 87168 35400 87174
rect 35348 87110 35400 87116
rect 34010 86524 34318 86533
rect 34010 86522 34016 86524
rect 34072 86522 34096 86524
rect 34152 86522 34176 86524
rect 34232 86522 34256 86524
rect 34312 86522 34318 86524
rect 34072 86470 34074 86522
rect 34254 86470 34256 86522
rect 34010 86468 34016 86470
rect 34072 86468 34096 86470
rect 34152 86468 34176 86470
rect 34232 86468 34256 86470
rect 34312 86468 34318 86470
rect 34010 86459 34318 86468
rect 34796 86352 34848 86358
rect 33888 86312 34008 86340
rect 33980 86154 34008 86312
rect 34796 86294 34848 86300
rect 34808 86222 34836 86294
rect 34796 86216 34848 86222
rect 34796 86158 34848 86164
rect 33876 86148 33928 86154
rect 33876 86090 33928 86096
rect 33968 86148 34020 86154
rect 33968 86090 34020 86096
rect 30380 86080 30432 86086
rect 30380 86022 30432 86028
rect 30150 85980 30458 85989
rect 30150 85978 30156 85980
rect 30212 85978 30236 85980
rect 30292 85978 30316 85980
rect 30372 85978 30396 85980
rect 30452 85978 30458 85980
rect 30212 85926 30214 85978
rect 30394 85926 30396 85978
rect 30150 85924 30156 85926
rect 30212 85924 30236 85926
rect 30292 85924 30316 85926
rect 30372 85924 30396 85926
rect 30452 85924 30458 85926
rect 30150 85915 30458 85924
rect 31750 85980 32058 85989
rect 31750 85978 31756 85980
rect 31812 85978 31836 85980
rect 31892 85978 31916 85980
rect 31972 85978 31996 85980
rect 32052 85978 32058 85980
rect 31812 85926 31814 85978
rect 31994 85926 31996 85978
rect 31750 85924 31756 85926
rect 31812 85924 31836 85926
rect 31892 85924 31916 85926
rect 31972 85924 31996 85926
rect 32052 85924 32058 85926
rect 31750 85915 32058 85924
rect 33350 85980 33658 85989
rect 33350 85978 33356 85980
rect 33412 85978 33436 85980
rect 33492 85978 33516 85980
rect 33572 85978 33596 85980
rect 33652 85978 33658 85980
rect 33412 85926 33414 85978
rect 33594 85926 33596 85978
rect 33350 85924 33356 85926
rect 33412 85924 33436 85926
rect 33492 85924 33516 85926
rect 33572 85924 33596 85926
rect 33652 85924 33658 85926
rect 33350 85915 33658 85924
rect 33888 85882 33916 86090
rect 27620 85876 27672 85882
rect 27620 85818 27672 85824
rect 30012 85876 30064 85882
rect 30012 85818 30064 85824
rect 33876 85876 33928 85882
rect 33876 85818 33928 85824
rect 34808 84998 34836 86158
rect 35360 86154 35388 87110
rect 36556 87038 36584 87586
rect 41696 87576 41748 87582
rect 41696 87518 41748 87524
rect 37648 87440 37700 87446
rect 37648 87382 37700 87388
rect 36544 87032 36596 87038
rect 36544 86974 36596 86980
rect 35610 86524 35918 86533
rect 35610 86522 35616 86524
rect 35672 86522 35696 86524
rect 35752 86522 35776 86524
rect 35832 86522 35856 86524
rect 35912 86522 35918 86524
rect 35672 86470 35674 86522
rect 35854 86470 35856 86522
rect 35610 86468 35616 86470
rect 35672 86468 35696 86470
rect 35752 86468 35776 86470
rect 35832 86468 35856 86470
rect 35912 86468 35918 86470
rect 35610 86459 35918 86468
rect 37210 86524 37518 86533
rect 37210 86522 37216 86524
rect 37272 86522 37296 86524
rect 37352 86522 37376 86524
rect 37432 86522 37456 86524
rect 37512 86522 37518 86524
rect 37272 86470 37274 86522
rect 37454 86470 37456 86522
rect 37210 86468 37216 86470
rect 37272 86468 37296 86470
rect 37352 86468 37376 86470
rect 37432 86468 37456 86470
rect 37512 86468 37518 86470
rect 37210 86459 37518 86468
rect 37372 86352 37424 86358
rect 37372 86294 37424 86300
rect 36084 86284 36136 86290
rect 36084 86226 36136 86232
rect 35348 86148 35400 86154
rect 35348 86090 35400 86096
rect 34950 85980 35258 85989
rect 34950 85978 34956 85980
rect 35012 85978 35036 85980
rect 35092 85978 35116 85980
rect 35172 85978 35196 85980
rect 35252 85978 35258 85980
rect 35012 85926 35014 85978
rect 35194 85926 35196 85978
rect 34950 85924 34956 85926
rect 35012 85924 35036 85926
rect 35092 85924 35116 85926
rect 35172 85924 35196 85926
rect 35252 85924 35258 85926
rect 34950 85915 35258 85924
rect 36096 85882 36124 86226
rect 36452 86080 36504 86086
rect 36452 86022 36504 86028
rect 36084 85876 36136 85882
rect 36084 85818 36136 85824
rect 36464 85746 36492 86022
rect 36550 85980 36858 85989
rect 36550 85978 36556 85980
rect 36612 85978 36636 85980
rect 36692 85978 36716 85980
rect 36772 85978 36796 85980
rect 36852 85978 36858 85980
rect 36612 85926 36614 85978
rect 36794 85926 36796 85978
rect 36550 85924 36556 85926
rect 36612 85924 36636 85926
rect 36692 85924 36716 85926
rect 36772 85924 36796 85926
rect 36852 85924 36858 85926
rect 36550 85915 36858 85924
rect 36452 85740 36504 85746
rect 36452 85682 36504 85688
rect 34796 84992 34848 84998
rect 34796 84934 34848 84940
rect 27344 84652 27396 84658
rect 27344 84594 27396 84600
rect 37384 83910 37412 86294
rect 37660 86154 37688 87382
rect 38810 86524 39118 86533
rect 38810 86522 38816 86524
rect 38872 86522 38896 86524
rect 38952 86522 38976 86524
rect 39032 86522 39056 86524
rect 39112 86522 39118 86524
rect 38872 86470 38874 86522
rect 39054 86470 39056 86522
rect 38810 86468 38816 86470
rect 38872 86468 38896 86470
rect 38952 86468 38976 86470
rect 39032 86468 39056 86470
rect 39112 86468 39118 86470
rect 38810 86459 39118 86468
rect 40410 86524 40718 86533
rect 40410 86522 40416 86524
rect 40472 86522 40496 86524
rect 40552 86522 40576 86524
rect 40632 86522 40656 86524
rect 40712 86522 40718 86524
rect 40472 86470 40474 86522
rect 40654 86470 40656 86522
rect 40410 86468 40416 86470
rect 40472 86468 40496 86470
rect 40552 86468 40576 86470
rect 40632 86468 40656 86470
rect 40712 86468 40718 86470
rect 40410 86459 40718 86468
rect 41708 86426 41736 87518
rect 44824 87304 44876 87310
rect 44824 87246 44876 87252
rect 41788 87100 41840 87106
rect 41788 87042 41840 87048
rect 40776 86420 40828 86426
rect 40776 86362 40828 86368
rect 41696 86420 41748 86426
rect 41696 86362 41748 86368
rect 40408 86284 40460 86290
rect 40408 86226 40460 86232
rect 38842 86184 38898 86193
rect 37648 86148 37700 86154
rect 38842 86119 38844 86128
rect 37648 86090 37700 86096
rect 38896 86119 38898 86128
rect 38844 86090 38896 86096
rect 37660 85814 37688 86090
rect 37832 86080 37884 86086
rect 37832 86022 37884 86028
rect 37648 85808 37700 85814
rect 37648 85750 37700 85756
rect 37844 85746 37872 86022
rect 38150 85980 38458 85989
rect 38150 85978 38156 85980
rect 38212 85978 38236 85980
rect 38292 85978 38316 85980
rect 38372 85978 38396 85980
rect 38452 85978 38458 85980
rect 38212 85926 38214 85978
rect 38394 85926 38396 85978
rect 38150 85924 38156 85926
rect 38212 85924 38236 85926
rect 38292 85924 38316 85926
rect 38372 85924 38396 85926
rect 38452 85924 38458 85926
rect 38150 85915 38458 85924
rect 37832 85740 37884 85746
rect 37832 85682 37884 85688
rect 38856 85610 38884 86090
rect 39750 85980 40058 85989
rect 39750 85978 39756 85980
rect 39812 85978 39836 85980
rect 39892 85978 39916 85980
rect 39972 85978 39996 85980
rect 40052 85978 40058 85980
rect 39812 85926 39814 85978
rect 39994 85926 39996 85978
rect 39750 85924 39756 85926
rect 39812 85924 39836 85926
rect 39892 85924 39916 85926
rect 39972 85924 39996 85926
rect 40052 85924 40058 85926
rect 39750 85915 40058 85924
rect 40420 85882 40448 86226
rect 40408 85876 40460 85882
rect 40408 85818 40460 85824
rect 40788 85678 40816 86362
rect 40868 86148 40920 86154
rect 40868 86090 40920 86096
rect 40880 85814 40908 86090
rect 41350 85980 41658 85989
rect 41350 85978 41356 85980
rect 41412 85978 41436 85980
rect 41492 85978 41516 85980
rect 41572 85978 41596 85980
rect 41652 85978 41658 85980
rect 41412 85926 41414 85978
rect 41594 85926 41596 85978
rect 41350 85924 41356 85926
rect 41412 85924 41436 85926
rect 41492 85924 41516 85926
rect 41572 85924 41596 85926
rect 41652 85924 41658 85926
rect 41350 85915 41658 85924
rect 40868 85808 40920 85814
rect 40868 85750 40920 85756
rect 40776 85672 40828 85678
rect 40038 85640 40094 85649
rect 38844 85604 38896 85610
rect 41800 85649 41828 87042
rect 42010 86524 42318 86533
rect 42010 86522 42016 86524
rect 42072 86522 42096 86524
rect 42152 86522 42176 86524
rect 42232 86522 42256 86524
rect 42312 86522 42318 86524
rect 42072 86470 42074 86522
rect 42254 86470 42256 86522
rect 42010 86468 42016 86470
rect 42072 86468 42096 86470
rect 42152 86468 42176 86470
rect 42232 86468 42256 86470
rect 42312 86468 42318 86470
rect 42010 86459 42318 86468
rect 43610 86524 43918 86533
rect 43610 86522 43616 86524
rect 43672 86522 43696 86524
rect 43752 86522 43776 86524
rect 43832 86522 43856 86524
rect 43912 86522 43918 86524
rect 43672 86470 43674 86522
rect 43854 86470 43856 86522
rect 43610 86468 43616 86470
rect 43672 86468 43696 86470
rect 43752 86468 43776 86470
rect 43832 86468 43856 86470
rect 43912 86468 43918 86470
rect 43610 86459 43918 86468
rect 44836 86358 44864 87246
rect 44916 87236 44968 87242
rect 44916 87178 44968 87184
rect 45100 87236 45152 87242
rect 45100 87178 45152 87184
rect 44928 87038 44956 87178
rect 44916 87032 44968 87038
rect 44916 86974 44968 86980
rect 44824 86352 44876 86358
rect 44824 86294 44876 86300
rect 42708 86284 42760 86290
rect 42708 86226 42760 86232
rect 42800 86284 42852 86290
rect 42800 86226 42852 86232
rect 42720 85678 42748 86226
rect 42812 86086 42840 86226
rect 44928 86154 44956 86974
rect 44916 86148 44968 86154
rect 44916 86090 44968 86096
rect 42800 86080 42852 86086
rect 42800 86022 42852 86028
rect 42812 85882 42840 86022
rect 42950 85980 43258 85989
rect 42950 85978 42956 85980
rect 43012 85978 43036 85980
rect 43092 85978 43116 85980
rect 43172 85978 43196 85980
rect 43252 85978 43258 85980
rect 43012 85926 43014 85978
rect 43194 85926 43196 85978
rect 42950 85924 42956 85926
rect 43012 85924 43036 85926
rect 43092 85924 43116 85926
rect 43172 85924 43196 85926
rect 43252 85924 43258 85926
rect 42950 85915 43258 85924
rect 44550 85980 44858 85989
rect 44550 85978 44556 85980
rect 44612 85978 44636 85980
rect 44692 85978 44716 85980
rect 44772 85978 44796 85980
rect 44852 85978 44858 85980
rect 44612 85926 44614 85978
rect 44794 85926 44796 85978
rect 44550 85924 44556 85926
rect 44612 85924 44636 85926
rect 44692 85924 44716 85926
rect 44772 85924 44796 85926
rect 44852 85924 44858 85926
rect 44550 85915 44858 85924
rect 42800 85876 42852 85882
rect 42800 85818 42852 85824
rect 42708 85672 42760 85678
rect 40776 85614 40828 85620
rect 41786 85640 41842 85649
rect 40038 85575 40094 85584
rect 42708 85614 42760 85620
rect 42798 85640 42854 85649
rect 41786 85575 41842 85584
rect 42798 85575 42800 85584
rect 38844 85546 38896 85552
rect 40052 85542 40080 85575
rect 42852 85575 42854 85584
rect 42800 85546 42852 85552
rect 40040 85536 40092 85542
rect 40040 85478 40092 85484
rect 44732 84788 44784 84794
rect 44732 84730 44784 84736
rect 42524 84720 42576 84726
rect 42524 84662 42576 84668
rect 42536 84425 42564 84662
rect 44744 84425 44772 84730
rect 42522 84416 42578 84425
rect 42522 84351 42578 84360
rect 44730 84416 44786 84425
rect 44730 84351 44786 84360
rect 37372 83904 37424 83910
rect 37372 83846 37424 83852
rect 45112 83706 45140 87178
rect 45210 86524 45518 86533
rect 45210 86522 45216 86524
rect 45272 86522 45296 86524
rect 45352 86522 45376 86524
rect 45432 86522 45456 86524
rect 45512 86522 45518 86524
rect 45272 86470 45274 86522
rect 45454 86470 45456 86522
rect 45210 86468 45216 86470
rect 45272 86468 45296 86470
rect 45352 86468 45376 86470
rect 45432 86468 45456 86470
rect 45512 86468 45518 86470
rect 45210 86459 45518 86468
rect 46810 86524 47118 86533
rect 46810 86522 46816 86524
rect 46872 86522 46896 86524
rect 46952 86522 46976 86524
rect 47032 86522 47056 86524
rect 47112 86522 47118 86524
rect 46872 86470 46874 86522
rect 47054 86470 47056 86522
rect 46810 86468 46816 86470
rect 46872 86468 46896 86470
rect 46952 86468 46976 86470
rect 47032 86468 47056 86470
rect 47112 86468 47118 86470
rect 46810 86459 47118 86468
rect 46150 85980 46458 85989
rect 46150 85978 46156 85980
rect 46212 85978 46236 85980
rect 46292 85978 46316 85980
rect 46372 85978 46396 85980
rect 46452 85978 46458 85980
rect 46212 85926 46214 85978
rect 46394 85926 46396 85978
rect 46150 85924 46156 85926
rect 46212 85924 46236 85926
rect 46292 85924 46316 85926
rect 46372 85924 46396 85926
rect 46452 85924 46458 85926
rect 46150 85915 46458 85924
rect 46572 85808 46624 85814
rect 46572 85750 46624 85756
rect 46584 85649 46612 85750
rect 47320 85649 47348 87586
rect 47860 87508 47912 87514
rect 47860 87450 47912 87456
rect 47872 86358 47900 87450
rect 53564 87440 53616 87446
rect 53564 87382 53616 87388
rect 50804 86964 50856 86970
rect 50804 86906 50856 86912
rect 48410 86524 48718 86533
rect 48410 86522 48416 86524
rect 48472 86522 48496 86524
rect 48552 86522 48576 86524
rect 48632 86522 48656 86524
rect 48712 86522 48718 86524
rect 48472 86470 48474 86522
rect 48654 86470 48656 86522
rect 48410 86468 48416 86470
rect 48472 86468 48496 86470
rect 48552 86468 48576 86470
rect 48632 86468 48656 86470
rect 48712 86468 48718 86470
rect 48410 86459 48718 86468
rect 50010 86524 50318 86533
rect 50010 86522 50016 86524
rect 50072 86522 50096 86524
rect 50152 86522 50176 86524
rect 50232 86522 50256 86524
rect 50312 86522 50318 86524
rect 50072 86470 50074 86522
rect 50254 86470 50256 86522
rect 50010 86468 50016 86470
rect 50072 86468 50096 86470
rect 50152 86468 50176 86470
rect 50232 86468 50256 86470
rect 50312 86468 50318 86470
rect 50010 86459 50318 86468
rect 50816 86426 50844 86906
rect 51610 86524 51918 86533
rect 51610 86522 51616 86524
rect 51672 86522 51696 86524
rect 51752 86522 51776 86524
rect 51832 86522 51856 86524
rect 51912 86522 51918 86524
rect 51672 86470 51674 86522
rect 51854 86470 51856 86522
rect 51610 86468 51616 86470
rect 51672 86468 51696 86470
rect 51752 86468 51776 86470
rect 51832 86468 51856 86470
rect 51912 86468 51918 86470
rect 51610 86459 51918 86468
rect 53210 86524 53518 86533
rect 53210 86522 53216 86524
rect 53272 86522 53296 86524
rect 53352 86522 53376 86524
rect 53432 86522 53456 86524
rect 53512 86522 53518 86524
rect 53272 86470 53274 86522
rect 53454 86470 53456 86522
rect 53210 86468 53216 86470
rect 53272 86468 53296 86470
rect 53352 86468 53376 86470
rect 53432 86468 53456 86470
rect 53512 86468 53518 86470
rect 53210 86459 53518 86468
rect 48964 86420 49016 86426
rect 48964 86362 49016 86368
rect 50712 86420 50764 86426
rect 50712 86362 50764 86368
rect 50804 86420 50856 86426
rect 50804 86362 50856 86368
rect 47860 86352 47912 86358
rect 47860 86294 47912 86300
rect 48870 86184 48926 86193
rect 48976 86154 49004 86362
rect 50724 86154 50752 86362
rect 48870 86119 48872 86128
rect 48924 86119 48926 86128
rect 48964 86148 49016 86154
rect 48872 86090 48924 86096
rect 48964 86090 49016 86096
rect 50712 86148 50764 86154
rect 50712 86090 50764 86096
rect 49240 86080 49292 86086
rect 49240 86022 49292 86028
rect 49884 86080 49936 86086
rect 49884 86022 49936 86028
rect 47750 85980 48058 85989
rect 47750 85978 47756 85980
rect 47812 85978 47836 85980
rect 47892 85978 47916 85980
rect 47972 85978 47996 85980
rect 48052 85978 48058 85980
rect 47812 85926 47814 85978
rect 47994 85926 47996 85978
rect 47750 85924 47756 85926
rect 47812 85924 47836 85926
rect 47892 85924 47916 85926
rect 47972 85924 47996 85926
rect 48052 85924 48058 85926
rect 47750 85915 48058 85924
rect 49252 85649 49280 86022
rect 49350 85980 49658 85989
rect 49350 85978 49356 85980
rect 49412 85978 49436 85980
rect 49492 85978 49516 85980
rect 49572 85978 49596 85980
rect 49652 85978 49658 85980
rect 49412 85926 49414 85978
rect 49594 85926 49596 85978
rect 49350 85924 49356 85926
rect 49412 85924 49436 85926
rect 49492 85924 49516 85926
rect 49572 85924 49596 85926
rect 49652 85924 49658 85926
rect 49350 85915 49658 85924
rect 49896 85814 49924 86022
rect 49884 85808 49936 85814
rect 49884 85750 49936 85756
rect 50816 85649 50844 86362
rect 53576 86154 53604 87382
rect 91284 87372 91336 87378
rect 91284 87314 91336 87320
rect 63500 87236 63552 87242
rect 63500 87178 63552 87184
rect 62488 86896 62540 86902
rect 62488 86838 62540 86844
rect 58348 86828 58400 86834
rect 58348 86770 58400 86776
rect 54810 86524 55118 86533
rect 54810 86522 54816 86524
rect 54872 86522 54896 86524
rect 54952 86522 54976 86524
rect 55032 86522 55056 86524
rect 55112 86522 55118 86524
rect 54872 86470 54874 86522
rect 55054 86470 55056 86522
rect 54810 86468 54816 86470
rect 54872 86468 54896 86470
rect 54952 86468 54976 86470
rect 55032 86468 55056 86470
rect 55112 86468 55118 86470
rect 54810 86459 55118 86468
rect 56410 86524 56718 86533
rect 56410 86522 56416 86524
rect 56472 86522 56496 86524
rect 56552 86522 56576 86524
rect 56632 86522 56656 86524
rect 56712 86522 56718 86524
rect 56472 86470 56474 86522
rect 56654 86470 56656 86522
rect 56410 86468 56416 86470
rect 56472 86468 56496 86470
rect 56552 86468 56576 86470
rect 56632 86468 56656 86470
rect 56712 86468 56718 86470
rect 56410 86459 56718 86468
rect 58010 86524 58318 86533
rect 58010 86522 58016 86524
rect 58072 86522 58096 86524
rect 58152 86522 58176 86524
rect 58232 86522 58256 86524
rect 58312 86522 58318 86524
rect 58072 86470 58074 86522
rect 58254 86470 58256 86522
rect 58010 86468 58016 86470
rect 58072 86468 58096 86470
rect 58152 86468 58176 86470
rect 58232 86468 58256 86470
rect 58312 86468 58318 86470
rect 58010 86459 58318 86468
rect 58360 86426 58388 86770
rect 61016 86760 61068 86766
rect 61016 86702 61068 86708
rect 59610 86524 59918 86533
rect 59610 86522 59616 86524
rect 59672 86522 59696 86524
rect 59752 86522 59776 86524
rect 59832 86522 59856 86524
rect 59912 86522 59918 86524
rect 59672 86470 59674 86522
rect 59854 86470 59856 86522
rect 59610 86468 59616 86470
rect 59672 86468 59696 86470
rect 59752 86468 59776 86470
rect 59832 86468 59856 86470
rect 59912 86468 59918 86470
rect 59610 86459 59918 86468
rect 58348 86420 58400 86426
rect 58348 86362 58400 86368
rect 55312 86216 55364 86222
rect 55310 86184 55312 86193
rect 55364 86184 55366 86193
rect 53564 86148 53616 86154
rect 55310 86119 55366 86128
rect 53564 86090 53616 86096
rect 52000 86080 52052 86086
rect 52000 86022 52052 86028
rect 53012 86080 53064 86086
rect 53012 86022 53064 86028
rect 56692 86080 56744 86086
rect 56692 86022 56744 86028
rect 50950 85980 51258 85989
rect 50950 85978 50956 85980
rect 51012 85978 51036 85980
rect 51092 85978 51116 85980
rect 51172 85978 51196 85980
rect 51252 85978 51258 85980
rect 51012 85926 51014 85978
rect 51194 85926 51196 85978
rect 50950 85924 50956 85926
rect 51012 85924 51036 85926
rect 51092 85924 51116 85926
rect 51172 85924 51196 85926
rect 51252 85924 51258 85926
rect 50950 85915 51258 85924
rect 52012 85746 52040 86022
rect 52550 85980 52858 85989
rect 52550 85978 52556 85980
rect 52612 85978 52636 85980
rect 52692 85978 52716 85980
rect 52772 85978 52796 85980
rect 52852 85978 52858 85980
rect 52612 85926 52614 85978
rect 52794 85926 52796 85978
rect 52550 85924 52556 85926
rect 52612 85924 52636 85926
rect 52692 85924 52716 85926
rect 52772 85924 52796 85926
rect 52852 85924 52858 85926
rect 52550 85915 52858 85924
rect 52000 85740 52052 85746
rect 52000 85682 52052 85688
rect 46570 85640 46626 85649
rect 47306 85640 47362 85649
rect 46570 85575 46626 85584
rect 46940 85604 46992 85610
rect 46584 85474 46612 85575
rect 47306 85575 47362 85584
rect 49238 85640 49294 85649
rect 49238 85575 49294 85584
rect 50802 85640 50858 85649
rect 50802 85575 50858 85584
rect 46940 85546 46992 85552
rect 46572 85468 46624 85474
rect 46572 85410 46624 85416
rect 45100 83700 45152 83706
rect 45100 83642 45152 83648
rect 46952 83638 46980 85546
rect 49252 85406 49280 85575
rect 49240 85400 49292 85406
rect 49240 85342 49292 85348
rect 52460 85332 52512 85338
rect 52460 85274 52512 85280
rect 51172 85196 51224 85202
rect 51172 85138 51224 85144
rect 51184 84697 51212 85138
rect 52472 84833 52500 85274
rect 53024 85105 53052 86022
rect 54150 85980 54458 85989
rect 54150 85978 54156 85980
rect 54212 85978 54236 85980
rect 54292 85978 54316 85980
rect 54372 85978 54396 85980
rect 54452 85978 54458 85980
rect 54212 85926 54214 85978
rect 54394 85926 54396 85978
rect 54150 85924 54156 85926
rect 54212 85924 54236 85926
rect 54292 85924 54316 85926
rect 54372 85924 54396 85926
rect 54452 85924 54458 85926
rect 54150 85915 54458 85924
rect 55750 85980 56058 85989
rect 55750 85978 55756 85980
rect 55812 85978 55836 85980
rect 55892 85978 55916 85980
rect 55972 85978 55996 85980
rect 56052 85978 56058 85980
rect 55812 85926 55814 85978
rect 55994 85926 55996 85978
rect 55750 85924 55756 85926
rect 55812 85924 55836 85926
rect 55892 85924 55916 85926
rect 55972 85924 55996 85926
rect 56052 85924 56058 85926
rect 55750 85915 56058 85924
rect 56704 85814 56732 86022
rect 57350 85980 57658 85989
rect 57350 85978 57356 85980
rect 57412 85978 57436 85980
rect 57492 85978 57516 85980
rect 57572 85978 57596 85980
rect 57652 85978 57658 85980
rect 57412 85926 57414 85978
rect 57594 85926 57596 85978
rect 57350 85924 57356 85926
rect 57412 85924 57436 85926
rect 57492 85924 57516 85926
rect 57572 85924 57596 85926
rect 57652 85924 57658 85926
rect 57350 85915 57658 85924
rect 56692 85808 56744 85814
rect 56692 85750 56744 85756
rect 55220 85672 55272 85678
rect 55218 85640 55220 85649
rect 58360 85649 58388 86362
rect 58950 85980 59258 85989
rect 58950 85978 58956 85980
rect 59012 85978 59036 85980
rect 59092 85978 59116 85980
rect 59172 85978 59196 85980
rect 59252 85978 59258 85980
rect 59012 85926 59014 85978
rect 59194 85926 59196 85978
rect 58950 85924 58956 85926
rect 59012 85924 59036 85926
rect 59092 85924 59116 85926
rect 59172 85924 59196 85926
rect 59252 85924 59258 85926
rect 58950 85915 59258 85924
rect 60550 85980 60858 85989
rect 60550 85978 60556 85980
rect 60612 85978 60636 85980
rect 60692 85978 60716 85980
rect 60772 85978 60796 85980
rect 60852 85978 60858 85980
rect 60612 85926 60614 85978
rect 60794 85926 60796 85978
rect 60550 85924 60556 85926
rect 60612 85924 60636 85926
rect 60692 85924 60716 85926
rect 60772 85924 60796 85926
rect 60852 85924 60858 85926
rect 60550 85915 60858 85924
rect 61028 85921 61056 86702
rect 61210 86524 61518 86533
rect 61210 86522 61216 86524
rect 61272 86522 61296 86524
rect 61352 86522 61376 86524
rect 61432 86522 61456 86524
rect 61512 86522 61518 86524
rect 61272 86470 61274 86522
rect 61454 86470 61456 86522
rect 61210 86468 61216 86470
rect 61272 86468 61296 86470
rect 61352 86468 61376 86470
rect 61432 86468 61456 86470
rect 61512 86468 61518 86470
rect 61210 86459 61518 86468
rect 62150 85980 62458 85989
rect 62150 85978 62156 85980
rect 62212 85978 62236 85980
rect 62292 85978 62316 85980
rect 62372 85978 62396 85980
rect 62452 85978 62458 85980
rect 62212 85926 62214 85978
rect 62394 85926 62396 85978
rect 62150 85924 62156 85926
rect 62212 85924 62236 85926
rect 62292 85924 62316 85926
rect 62372 85924 62396 85926
rect 62452 85924 62458 85926
rect 61014 85912 61070 85921
rect 62150 85915 62458 85924
rect 61014 85847 61070 85856
rect 62500 85649 62528 86838
rect 62810 86524 63118 86533
rect 62810 86522 62816 86524
rect 62872 86522 62896 86524
rect 62952 86522 62976 86524
rect 63032 86522 63056 86524
rect 63112 86522 63118 86524
rect 62872 86470 62874 86522
rect 63054 86470 63056 86522
rect 62810 86468 62816 86470
rect 62872 86468 62896 86470
rect 62952 86468 62976 86470
rect 63032 86468 63056 86470
rect 63112 86468 63118 86470
rect 62810 86459 63118 86468
rect 63512 85921 63540 87178
rect 72148 87168 72200 87174
rect 72148 87110 72200 87116
rect 68100 86692 68152 86698
rect 68100 86634 68152 86640
rect 68008 86624 68060 86630
rect 68008 86566 68060 86572
rect 64410 86524 64718 86533
rect 64410 86522 64416 86524
rect 64472 86522 64496 86524
rect 64552 86522 64576 86524
rect 64632 86522 64656 86524
rect 64712 86522 64718 86524
rect 64472 86470 64474 86522
rect 64654 86470 64656 86522
rect 64410 86468 64416 86470
rect 64472 86468 64496 86470
rect 64552 86468 64576 86470
rect 64632 86468 64656 86470
rect 64712 86468 64718 86470
rect 64410 86459 64718 86468
rect 66010 86524 66318 86533
rect 66010 86522 66016 86524
rect 66072 86522 66096 86524
rect 66152 86522 66176 86524
rect 66232 86522 66256 86524
rect 66312 86522 66318 86524
rect 66072 86470 66074 86522
rect 66254 86470 66256 86522
rect 66010 86468 66016 86470
rect 66072 86468 66096 86470
rect 66152 86468 66176 86470
rect 66232 86468 66256 86470
rect 66312 86468 66318 86470
rect 66010 86459 66318 86468
rect 67610 86524 67918 86533
rect 67610 86522 67616 86524
rect 67672 86522 67696 86524
rect 67752 86522 67776 86524
rect 67832 86522 67856 86524
rect 67912 86522 67918 86524
rect 67672 86470 67674 86522
rect 67854 86470 67856 86522
rect 67610 86468 67616 86470
rect 67672 86468 67696 86470
rect 67752 86468 67776 86470
rect 67832 86468 67856 86470
rect 67912 86468 67918 86470
rect 67610 86459 67918 86468
rect 63750 85980 64058 85989
rect 63750 85978 63756 85980
rect 63812 85978 63836 85980
rect 63892 85978 63916 85980
rect 63972 85978 63996 85980
rect 64052 85978 64058 85980
rect 63812 85926 63814 85978
rect 63994 85926 63996 85978
rect 63750 85924 63756 85926
rect 63812 85924 63836 85926
rect 63892 85924 63916 85926
rect 63972 85924 63996 85926
rect 64052 85924 64058 85926
rect 63498 85912 63554 85921
rect 63750 85915 64058 85924
rect 65350 85980 65658 85989
rect 65350 85978 65356 85980
rect 65412 85978 65436 85980
rect 65492 85978 65516 85980
rect 65572 85978 65596 85980
rect 65652 85978 65658 85980
rect 65412 85926 65414 85978
rect 65594 85926 65596 85978
rect 65350 85924 65356 85926
rect 65412 85924 65436 85926
rect 65492 85924 65516 85926
rect 65572 85924 65596 85926
rect 65652 85924 65658 85926
rect 65350 85915 65658 85924
rect 66950 85980 67258 85989
rect 66950 85978 66956 85980
rect 67012 85978 67036 85980
rect 67092 85978 67116 85980
rect 67172 85978 67196 85980
rect 67252 85978 67258 85980
rect 67012 85926 67014 85978
rect 67194 85926 67196 85978
rect 66950 85924 66956 85926
rect 67012 85924 67036 85926
rect 67092 85924 67116 85926
rect 67172 85924 67196 85926
rect 67252 85924 67258 85926
rect 66950 85915 67258 85924
rect 63498 85847 63554 85856
rect 68020 85785 68048 86566
rect 68112 85921 68140 86634
rect 69210 86524 69518 86533
rect 69210 86522 69216 86524
rect 69272 86522 69296 86524
rect 69352 86522 69376 86524
rect 69432 86522 69456 86524
rect 69512 86522 69518 86524
rect 69272 86470 69274 86522
rect 69454 86470 69456 86522
rect 69210 86468 69216 86470
rect 69272 86468 69296 86470
rect 69352 86468 69376 86470
rect 69432 86468 69456 86470
rect 69512 86468 69518 86470
rect 69210 86459 69518 86468
rect 70810 86524 71118 86533
rect 70810 86522 70816 86524
rect 70872 86522 70896 86524
rect 70952 86522 70976 86524
rect 71032 86522 71056 86524
rect 71112 86522 71118 86524
rect 70872 86470 70874 86522
rect 71054 86470 71056 86522
rect 70810 86468 70816 86470
rect 70872 86468 70896 86470
rect 70952 86468 70976 86470
rect 71032 86468 71056 86470
rect 71112 86468 71118 86470
rect 70810 86459 71118 86468
rect 68550 85980 68858 85989
rect 68550 85978 68556 85980
rect 68612 85978 68636 85980
rect 68692 85978 68716 85980
rect 68772 85978 68796 85980
rect 68852 85978 68858 85980
rect 68612 85926 68614 85978
rect 68794 85926 68796 85978
rect 68550 85924 68556 85926
rect 68612 85924 68636 85926
rect 68692 85924 68716 85926
rect 68772 85924 68796 85926
rect 68852 85924 68858 85926
rect 68098 85912 68154 85921
rect 68550 85915 68858 85924
rect 70150 85980 70458 85989
rect 70150 85978 70156 85980
rect 70212 85978 70236 85980
rect 70292 85978 70316 85980
rect 70372 85978 70396 85980
rect 70452 85978 70458 85980
rect 70212 85926 70214 85978
rect 70394 85926 70396 85978
rect 70150 85924 70156 85926
rect 70212 85924 70236 85926
rect 70292 85924 70316 85926
rect 70372 85924 70396 85926
rect 70452 85924 70458 85926
rect 70150 85915 70458 85924
rect 71750 85980 72058 85989
rect 71750 85978 71756 85980
rect 71812 85978 71836 85980
rect 71892 85978 71916 85980
rect 71972 85978 71996 85980
rect 72052 85978 72058 85980
rect 71812 85926 71814 85978
rect 71994 85926 71996 85978
rect 71750 85924 71756 85926
rect 71812 85924 71836 85926
rect 71892 85924 71916 85926
rect 71972 85924 71996 85926
rect 72052 85924 72058 85926
rect 71750 85915 72058 85924
rect 72160 85921 72188 87110
rect 77668 87100 77720 87106
rect 77668 87042 77720 87048
rect 72410 86524 72718 86533
rect 72410 86522 72416 86524
rect 72472 86522 72496 86524
rect 72552 86522 72576 86524
rect 72632 86522 72656 86524
rect 72712 86522 72718 86524
rect 72472 86470 72474 86522
rect 72654 86470 72656 86522
rect 72410 86468 72416 86470
rect 72472 86468 72496 86470
rect 72552 86468 72576 86470
rect 72632 86468 72656 86470
rect 72712 86468 72718 86470
rect 72410 86459 72718 86468
rect 74010 86524 74318 86533
rect 74010 86522 74016 86524
rect 74072 86522 74096 86524
rect 74152 86522 74176 86524
rect 74232 86522 74256 86524
rect 74312 86522 74318 86524
rect 74072 86470 74074 86522
rect 74254 86470 74256 86522
rect 74010 86468 74016 86470
rect 74072 86468 74096 86470
rect 74152 86468 74176 86470
rect 74232 86468 74256 86470
rect 74312 86468 74318 86470
rect 74010 86459 74318 86468
rect 75610 86524 75918 86533
rect 75610 86522 75616 86524
rect 75672 86522 75696 86524
rect 75752 86522 75776 86524
rect 75832 86522 75856 86524
rect 75912 86522 75918 86524
rect 75672 86470 75674 86522
rect 75854 86470 75856 86522
rect 75610 86468 75616 86470
rect 75672 86468 75696 86470
rect 75752 86468 75776 86470
rect 75832 86468 75856 86470
rect 75912 86468 75918 86470
rect 75610 86459 75918 86468
rect 77210 86524 77518 86533
rect 77210 86522 77216 86524
rect 77272 86522 77296 86524
rect 77352 86522 77376 86524
rect 77432 86522 77456 86524
rect 77512 86522 77518 86524
rect 77272 86470 77274 86522
rect 77454 86470 77456 86522
rect 77210 86468 77216 86470
rect 77272 86468 77296 86470
rect 77352 86468 77376 86470
rect 77432 86468 77456 86470
rect 77512 86468 77518 86470
rect 77210 86459 77518 86468
rect 74632 86148 74684 86154
rect 74632 86090 74684 86096
rect 73350 85980 73658 85989
rect 73350 85978 73356 85980
rect 73412 85978 73436 85980
rect 73492 85978 73516 85980
rect 73572 85978 73596 85980
rect 73652 85978 73658 85980
rect 73412 85926 73414 85978
rect 73594 85926 73596 85978
rect 73350 85924 73356 85926
rect 73412 85924 73436 85926
rect 73492 85924 73516 85926
rect 73572 85924 73596 85926
rect 73652 85924 73658 85926
rect 68098 85847 68154 85856
rect 72146 85912 72202 85921
rect 73350 85915 73658 85924
rect 72146 85847 72202 85856
rect 68006 85776 68062 85785
rect 68006 85711 68062 85720
rect 73160 85740 73212 85746
rect 73160 85682 73212 85688
rect 73172 85649 73200 85682
rect 74644 85649 74672 86090
rect 74950 85980 75258 85989
rect 74950 85978 74956 85980
rect 75012 85978 75036 85980
rect 75092 85978 75116 85980
rect 75172 85978 75196 85980
rect 75252 85978 75258 85980
rect 75012 85926 75014 85978
rect 75194 85926 75196 85978
rect 74950 85924 74956 85926
rect 75012 85924 75036 85926
rect 75092 85924 75116 85926
rect 75172 85924 75196 85926
rect 75252 85924 75258 85926
rect 74950 85915 75258 85924
rect 76550 85980 76858 85989
rect 76550 85978 76556 85980
rect 76612 85978 76636 85980
rect 76692 85978 76716 85980
rect 76772 85978 76796 85980
rect 76852 85978 76858 85980
rect 76612 85926 76614 85978
rect 76794 85926 76796 85978
rect 76550 85924 76556 85926
rect 76612 85924 76636 85926
rect 76692 85924 76716 85926
rect 76772 85924 76796 85926
rect 76852 85924 76858 85926
rect 76550 85915 76858 85924
rect 75920 85876 75972 85882
rect 75920 85818 75972 85824
rect 75932 85649 75960 85818
rect 77680 85649 77708 87042
rect 78810 86524 79118 86533
rect 78810 86522 78816 86524
rect 78872 86522 78896 86524
rect 78952 86522 78976 86524
rect 79032 86522 79056 86524
rect 79112 86522 79118 86524
rect 78872 86470 78874 86522
rect 79054 86470 79056 86522
rect 78810 86468 78816 86470
rect 78872 86468 78896 86470
rect 78952 86468 78976 86470
rect 79032 86468 79056 86470
rect 79112 86468 79118 86470
rect 78810 86459 79118 86468
rect 80410 86524 80718 86533
rect 80410 86522 80416 86524
rect 80472 86522 80496 86524
rect 80552 86522 80576 86524
rect 80632 86522 80656 86524
rect 80712 86522 80718 86524
rect 80472 86470 80474 86522
rect 80654 86470 80656 86522
rect 80410 86468 80416 86470
rect 80472 86468 80496 86470
rect 80552 86468 80576 86470
rect 80632 86468 80656 86470
rect 80712 86468 80718 86470
rect 80410 86459 80718 86468
rect 82010 86524 82318 86533
rect 82010 86522 82016 86524
rect 82072 86522 82096 86524
rect 82152 86522 82176 86524
rect 82232 86522 82256 86524
rect 82312 86522 82318 86524
rect 82072 86470 82074 86522
rect 82254 86470 82256 86522
rect 82010 86468 82016 86470
rect 82072 86468 82096 86470
rect 82152 86468 82176 86470
rect 82232 86468 82256 86470
rect 82312 86468 82318 86470
rect 82010 86459 82318 86468
rect 83610 86524 83918 86533
rect 83610 86522 83616 86524
rect 83672 86522 83696 86524
rect 83752 86522 83776 86524
rect 83832 86522 83856 86524
rect 83912 86522 83918 86524
rect 83672 86470 83674 86522
rect 83854 86470 83856 86522
rect 83610 86468 83616 86470
rect 83672 86468 83696 86470
rect 83752 86468 83776 86470
rect 83832 86468 83856 86470
rect 83912 86468 83918 86470
rect 83610 86459 83918 86468
rect 85210 86524 85518 86533
rect 85210 86522 85216 86524
rect 85272 86522 85296 86524
rect 85352 86522 85376 86524
rect 85432 86522 85456 86524
rect 85512 86522 85518 86524
rect 85272 86470 85274 86522
rect 85454 86470 85456 86522
rect 85210 86468 85216 86470
rect 85272 86468 85296 86470
rect 85352 86468 85376 86470
rect 85432 86468 85456 86470
rect 85512 86468 85518 86470
rect 85210 86459 85518 86468
rect 86810 86524 87118 86533
rect 86810 86522 86816 86524
rect 86872 86522 86896 86524
rect 86952 86522 86976 86524
rect 87032 86522 87056 86524
rect 87112 86522 87118 86524
rect 86872 86470 86874 86522
rect 87054 86470 87056 86522
rect 86810 86468 86816 86470
rect 86872 86468 86896 86470
rect 86952 86468 86976 86470
rect 87032 86468 87056 86470
rect 87112 86468 87118 86470
rect 86810 86459 87118 86468
rect 88410 86524 88718 86533
rect 88410 86522 88416 86524
rect 88472 86522 88496 86524
rect 88552 86522 88576 86524
rect 88632 86522 88656 86524
rect 88712 86522 88718 86524
rect 88472 86470 88474 86522
rect 88654 86470 88656 86522
rect 88410 86468 88416 86470
rect 88472 86468 88496 86470
rect 88552 86468 88576 86470
rect 88632 86468 88656 86470
rect 88712 86468 88718 86470
rect 88410 86459 88718 86468
rect 90010 86524 90318 86533
rect 90010 86522 90016 86524
rect 90072 86522 90096 86524
rect 90152 86522 90176 86524
rect 90232 86522 90256 86524
rect 90312 86522 90318 86524
rect 90072 86470 90074 86522
rect 90254 86470 90256 86522
rect 90010 86468 90016 86470
rect 90072 86468 90096 86470
rect 90152 86468 90176 86470
rect 90232 86468 90256 86470
rect 90312 86468 90318 86470
rect 90010 86459 90318 86468
rect 78150 85980 78458 85989
rect 78150 85978 78156 85980
rect 78212 85978 78236 85980
rect 78292 85978 78316 85980
rect 78372 85978 78396 85980
rect 78452 85978 78458 85980
rect 78212 85926 78214 85978
rect 78394 85926 78396 85978
rect 78150 85924 78156 85926
rect 78212 85924 78236 85926
rect 78292 85924 78316 85926
rect 78372 85924 78396 85926
rect 78452 85924 78458 85926
rect 78150 85915 78458 85924
rect 79750 85980 80058 85989
rect 79750 85978 79756 85980
rect 79812 85978 79836 85980
rect 79892 85978 79916 85980
rect 79972 85978 79996 85980
rect 80052 85978 80058 85980
rect 79812 85926 79814 85978
rect 79994 85926 79996 85978
rect 79750 85924 79756 85926
rect 79812 85924 79836 85926
rect 79892 85924 79916 85926
rect 79972 85924 79996 85926
rect 80052 85924 80058 85926
rect 79750 85915 80058 85924
rect 81350 85980 81658 85989
rect 81350 85978 81356 85980
rect 81412 85978 81436 85980
rect 81492 85978 81516 85980
rect 81572 85978 81596 85980
rect 81652 85978 81658 85980
rect 81412 85926 81414 85978
rect 81594 85926 81596 85978
rect 81350 85924 81356 85926
rect 81412 85924 81436 85926
rect 81492 85924 81516 85926
rect 81572 85924 81596 85926
rect 81652 85924 81658 85926
rect 81350 85915 81658 85924
rect 82950 85980 83258 85989
rect 82950 85978 82956 85980
rect 83012 85978 83036 85980
rect 83092 85978 83116 85980
rect 83172 85978 83196 85980
rect 83252 85978 83258 85980
rect 83012 85926 83014 85978
rect 83194 85926 83196 85978
rect 82950 85924 82956 85926
rect 83012 85924 83036 85926
rect 83092 85924 83116 85926
rect 83172 85924 83196 85926
rect 83252 85924 83258 85926
rect 82950 85915 83258 85924
rect 84550 85980 84858 85989
rect 84550 85978 84556 85980
rect 84612 85978 84636 85980
rect 84692 85978 84716 85980
rect 84772 85978 84796 85980
rect 84852 85978 84858 85980
rect 84612 85926 84614 85978
rect 84794 85926 84796 85978
rect 84550 85924 84556 85926
rect 84612 85924 84636 85926
rect 84692 85924 84716 85926
rect 84772 85924 84796 85926
rect 84852 85924 84858 85926
rect 84550 85915 84858 85924
rect 86150 85980 86458 85989
rect 86150 85978 86156 85980
rect 86212 85978 86236 85980
rect 86292 85978 86316 85980
rect 86372 85978 86396 85980
rect 86452 85978 86458 85980
rect 86212 85926 86214 85978
rect 86394 85926 86396 85978
rect 86150 85924 86156 85926
rect 86212 85924 86236 85926
rect 86292 85924 86316 85926
rect 86372 85924 86396 85926
rect 86452 85924 86458 85926
rect 86150 85915 86458 85924
rect 87750 85980 88058 85989
rect 87750 85978 87756 85980
rect 87812 85978 87836 85980
rect 87892 85978 87916 85980
rect 87972 85978 87996 85980
rect 88052 85978 88058 85980
rect 87812 85926 87814 85978
rect 87994 85926 87996 85978
rect 87750 85924 87756 85926
rect 87812 85924 87836 85926
rect 87892 85924 87916 85926
rect 87972 85924 87996 85926
rect 88052 85924 88058 85926
rect 87750 85915 88058 85924
rect 89350 85980 89658 85989
rect 89350 85978 89356 85980
rect 89412 85978 89436 85980
rect 89492 85978 89516 85980
rect 89572 85978 89596 85980
rect 89652 85978 89658 85980
rect 89412 85926 89414 85978
rect 89594 85926 89596 85978
rect 89350 85924 89356 85926
rect 89412 85924 89436 85926
rect 89492 85924 89516 85926
rect 89572 85924 89596 85926
rect 89652 85924 89658 85926
rect 89350 85915 89658 85924
rect 90950 85980 91258 85989
rect 90950 85978 90956 85980
rect 91012 85978 91036 85980
rect 91092 85978 91116 85980
rect 91172 85978 91196 85980
rect 91252 85978 91258 85980
rect 91012 85926 91014 85978
rect 91194 85926 91196 85978
rect 90950 85924 90956 85926
rect 91012 85924 91036 85926
rect 91092 85924 91116 85926
rect 91172 85924 91196 85926
rect 91252 85924 91258 85926
rect 90950 85915 91258 85924
rect 91296 85649 91324 87314
rect 91610 86524 91918 86533
rect 91610 86522 91616 86524
rect 91672 86522 91696 86524
rect 91752 86522 91776 86524
rect 91832 86522 91856 86524
rect 91912 86522 91918 86524
rect 91672 86470 91674 86522
rect 91854 86470 91856 86522
rect 91610 86468 91616 86470
rect 91672 86468 91696 86470
rect 91752 86468 91776 86470
rect 91832 86468 91856 86470
rect 91912 86468 91918 86470
rect 91610 86459 91918 86468
rect 93210 86524 93518 86533
rect 93210 86522 93216 86524
rect 93272 86522 93296 86524
rect 93352 86522 93376 86524
rect 93432 86522 93456 86524
rect 93512 86522 93518 86524
rect 93272 86470 93274 86522
rect 93454 86470 93456 86522
rect 93210 86468 93216 86470
rect 93272 86468 93296 86470
rect 93352 86468 93376 86470
rect 93432 86468 93456 86470
rect 93512 86468 93518 86470
rect 93210 86459 93518 86468
rect 94810 86524 95118 86533
rect 94810 86522 94816 86524
rect 94872 86522 94896 86524
rect 94952 86522 94976 86524
rect 95032 86522 95056 86524
rect 95112 86522 95118 86524
rect 94872 86470 94874 86522
rect 95054 86470 95056 86522
rect 94810 86468 94816 86470
rect 94872 86468 94896 86470
rect 94952 86468 94976 86470
rect 95032 86468 95056 86470
rect 95112 86468 95118 86470
rect 94810 86459 95118 86468
rect 96410 86524 96718 86533
rect 96410 86522 96416 86524
rect 96472 86522 96496 86524
rect 96552 86522 96576 86524
rect 96632 86522 96656 86524
rect 96712 86522 96718 86524
rect 96472 86470 96474 86522
rect 96654 86470 96656 86522
rect 96410 86468 96416 86470
rect 96472 86468 96496 86470
rect 96552 86468 96576 86470
rect 96632 86468 96656 86470
rect 96712 86468 96718 86470
rect 96410 86459 96718 86468
rect 98010 86524 98318 86533
rect 98010 86522 98016 86524
rect 98072 86522 98096 86524
rect 98152 86522 98176 86524
rect 98232 86522 98256 86524
rect 98312 86522 98318 86524
rect 98072 86470 98074 86522
rect 98254 86470 98256 86522
rect 98010 86468 98016 86470
rect 98072 86468 98096 86470
rect 98152 86468 98176 86470
rect 98232 86468 98256 86470
rect 98312 86468 98318 86470
rect 98010 86459 98318 86468
rect 99610 86524 99918 86533
rect 99610 86522 99616 86524
rect 99672 86522 99696 86524
rect 99752 86522 99776 86524
rect 99832 86522 99856 86524
rect 99912 86522 99918 86524
rect 99672 86470 99674 86522
rect 99854 86470 99856 86522
rect 99610 86468 99616 86470
rect 99672 86468 99696 86470
rect 99752 86468 99776 86470
rect 99832 86468 99856 86470
rect 99912 86468 99918 86470
rect 99610 86459 99918 86468
rect 101210 86524 101518 86533
rect 101210 86522 101216 86524
rect 101272 86522 101296 86524
rect 101352 86522 101376 86524
rect 101432 86522 101456 86524
rect 101512 86522 101518 86524
rect 101272 86470 101274 86522
rect 101454 86470 101456 86522
rect 101210 86468 101216 86470
rect 101272 86468 101296 86470
rect 101352 86468 101376 86470
rect 101432 86468 101456 86470
rect 101512 86468 101518 86470
rect 101210 86459 101518 86468
rect 102810 86524 103118 86533
rect 102810 86522 102816 86524
rect 102872 86522 102896 86524
rect 102952 86522 102976 86524
rect 103032 86522 103056 86524
rect 103112 86522 103118 86524
rect 102872 86470 102874 86522
rect 103054 86470 103056 86522
rect 102810 86468 102816 86470
rect 102872 86468 102896 86470
rect 102952 86468 102976 86470
rect 103032 86468 103056 86470
rect 103112 86468 103118 86470
rect 102810 86459 103118 86468
rect 104410 86524 104718 86533
rect 104410 86522 104416 86524
rect 104472 86522 104496 86524
rect 104552 86522 104576 86524
rect 104632 86522 104656 86524
rect 104712 86522 104718 86524
rect 104472 86470 104474 86522
rect 104654 86470 104656 86522
rect 104410 86468 104416 86470
rect 104472 86468 104496 86470
rect 104552 86468 104576 86470
rect 104632 86468 104656 86470
rect 104712 86468 104718 86470
rect 104410 86459 104718 86468
rect 106010 86524 106318 86533
rect 106010 86522 106016 86524
rect 106072 86522 106096 86524
rect 106152 86522 106176 86524
rect 106232 86522 106256 86524
rect 106312 86522 106318 86524
rect 106072 86470 106074 86522
rect 106254 86470 106256 86522
rect 106010 86468 106016 86470
rect 106072 86468 106096 86470
rect 106152 86468 106176 86470
rect 106232 86468 106256 86470
rect 106312 86468 106318 86470
rect 106010 86459 106318 86468
rect 107610 86524 107918 86533
rect 107610 86522 107616 86524
rect 107672 86522 107696 86524
rect 107752 86522 107776 86524
rect 107832 86522 107856 86524
rect 107912 86522 107918 86524
rect 107672 86470 107674 86522
rect 107854 86470 107856 86522
rect 107610 86468 107616 86470
rect 107672 86468 107696 86470
rect 107752 86468 107776 86470
rect 107832 86468 107856 86470
rect 107912 86468 107918 86470
rect 107610 86459 107918 86468
rect 100944 86216 100996 86222
rect 100944 86158 100996 86164
rect 108028 86216 108080 86222
rect 108028 86158 108080 86164
rect 92550 85980 92858 85989
rect 92550 85978 92556 85980
rect 92612 85978 92636 85980
rect 92692 85978 92716 85980
rect 92772 85978 92796 85980
rect 92852 85978 92858 85980
rect 92612 85926 92614 85978
rect 92794 85926 92796 85978
rect 92550 85924 92556 85926
rect 92612 85924 92636 85926
rect 92692 85924 92716 85926
rect 92772 85924 92796 85926
rect 92852 85924 92858 85926
rect 92550 85915 92858 85924
rect 94150 85980 94458 85989
rect 94150 85978 94156 85980
rect 94212 85978 94236 85980
rect 94292 85978 94316 85980
rect 94372 85978 94396 85980
rect 94452 85978 94458 85980
rect 94212 85926 94214 85978
rect 94394 85926 94396 85978
rect 94150 85924 94156 85926
rect 94212 85924 94236 85926
rect 94292 85924 94316 85926
rect 94372 85924 94396 85926
rect 94452 85924 94458 85926
rect 94150 85915 94458 85924
rect 95750 85980 96058 85989
rect 95750 85978 95756 85980
rect 95812 85978 95836 85980
rect 95892 85978 95916 85980
rect 95972 85978 95996 85980
rect 96052 85978 96058 85980
rect 95812 85926 95814 85978
rect 95994 85926 95996 85978
rect 95750 85924 95756 85926
rect 95812 85924 95836 85926
rect 95892 85924 95916 85926
rect 95972 85924 95996 85926
rect 96052 85924 96058 85926
rect 95750 85915 96058 85924
rect 97350 85980 97658 85989
rect 97350 85978 97356 85980
rect 97412 85978 97436 85980
rect 97492 85978 97516 85980
rect 97572 85978 97596 85980
rect 97652 85978 97658 85980
rect 97412 85926 97414 85978
rect 97594 85926 97596 85978
rect 97350 85924 97356 85926
rect 97412 85924 97436 85926
rect 97492 85924 97516 85926
rect 97572 85924 97596 85926
rect 97652 85924 97658 85926
rect 97350 85915 97658 85924
rect 98950 85980 99258 85989
rect 98950 85978 98956 85980
rect 99012 85978 99036 85980
rect 99092 85978 99116 85980
rect 99172 85978 99196 85980
rect 99252 85978 99258 85980
rect 99012 85926 99014 85978
rect 99194 85926 99196 85978
rect 98950 85924 98956 85926
rect 99012 85924 99036 85926
rect 99092 85924 99116 85926
rect 99172 85924 99196 85926
rect 99252 85924 99258 85926
rect 98950 85915 99258 85924
rect 100550 85980 100858 85989
rect 100550 85978 100556 85980
rect 100612 85978 100636 85980
rect 100692 85978 100716 85980
rect 100772 85978 100796 85980
rect 100852 85978 100858 85980
rect 100612 85926 100614 85978
rect 100794 85926 100796 85978
rect 100550 85924 100556 85926
rect 100612 85924 100636 85926
rect 100692 85924 100716 85926
rect 100772 85924 100796 85926
rect 100852 85924 100858 85926
rect 100550 85915 100858 85924
rect 100956 85649 100984 86158
rect 102150 85980 102458 85989
rect 102150 85978 102156 85980
rect 102212 85978 102236 85980
rect 102292 85978 102316 85980
rect 102372 85978 102396 85980
rect 102452 85978 102458 85980
rect 102212 85926 102214 85978
rect 102394 85926 102396 85978
rect 102150 85924 102156 85926
rect 102212 85924 102236 85926
rect 102292 85924 102316 85926
rect 102372 85924 102396 85926
rect 102452 85924 102458 85926
rect 102150 85915 102458 85924
rect 103750 85980 104058 85989
rect 103750 85978 103756 85980
rect 103812 85978 103836 85980
rect 103892 85978 103916 85980
rect 103972 85978 103996 85980
rect 104052 85978 104058 85980
rect 103812 85926 103814 85978
rect 103994 85926 103996 85978
rect 103750 85924 103756 85926
rect 103812 85924 103836 85926
rect 103892 85924 103916 85926
rect 103972 85924 103996 85926
rect 104052 85924 104058 85926
rect 103750 85915 104058 85924
rect 105350 85980 105658 85989
rect 105350 85978 105356 85980
rect 105412 85978 105436 85980
rect 105492 85978 105516 85980
rect 105572 85978 105596 85980
rect 105652 85978 105658 85980
rect 105412 85926 105414 85978
rect 105594 85926 105596 85978
rect 105350 85924 105356 85926
rect 105412 85924 105436 85926
rect 105492 85924 105516 85926
rect 105572 85924 105596 85926
rect 105652 85924 105658 85926
rect 105350 85915 105658 85924
rect 106950 85980 107258 85989
rect 106950 85978 106956 85980
rect 107012 85978 107036 85980
rect 107092 85978 107116 85980
rect 107172 85978 107196 85980
rect 107252 85978 107258 85980
rect 107012 85926 107014 85978
rect 107194 85926 107196 85978
rect 106950 85924 106956 85926
rect 107012 85924 107036 85926
rect 107092 85924 107116 85926
rect 107172 85924 107196 85926
rect 107252 85924 107258 85926
rect 106950 85915 107258 85924
rect 55272 85640 55274 85649
rect 55218 85575 55274 85584
rect 55678 85640 55734 85649
rect 55678 85575 55680 85584
rect 55732 85575 55734 85584
rect 58346 85640 58402 85649
rect 58346 85575 58402 85584
rect 62486 85640 62542 85649
rect 62486 85575 62542 85584
rect 73158 85640 73214 85649
rect 73158 85575 73214 85584
rect 74630 85640 74686 85649
rect 74630 85575 74686 85584
rect 75918 85640 75974 85649
rect 75918 85575 75974 85584
rect 77666 85640 77722 85649
rect 77666 85575 77722 85584
rect 91282 85640 91338 85649
rect 91282 85575 91338 85584
rect 100942 85640 100998 85649
rect 100942 85575 100998 85584
rect 55680 85546 55732 85552
rect 53840 85264 53892 85270
rect 53840 85206 53892 85212
rect 53010 85096 53066 85105
rect 53010 85031 53066 85040
rect 52458 84824 52514 84833
rect 52458 84759 52514 84768
rect 53852 84697 53880 85206
rect 66260 85128 66312 85134
rect 66260 85070 66312 85076
rect 57612 84924 57664 84930
rect 57612 84866 57664 84872
rect 51170 84688 51226 84697
rect 51170 84623 51226 84632
rect 53838 84688 53894 84697
rect 53838 84623 53894 84632
rect 57624 84561 57652 84866
rect 66272 84697 66300 85070
rect 71228 85060 71280 85066
rect 71228 85002 71280 85008
rect 71240 84697 71268 85002
rect 78680 84856 78732 84862
rect 78680 84798 78732 84804
rect 66258 84688 66314 84697
rect 66258 84623 66314 84632
rect 71226 84688 71282 84697
rect 71226 84623 71282 84632
rect 78692 84561 78720 84798
rect 57610 84552 57666 84561
rect 57610 84487 57666 84496
rect 78678 84552 78734 84561
rect 78678 84487 78734 84496
rect 59910 83736 59966 83745
rect 59910 83671 59966 83680
rect 70214 83736 70270 83745
rect 70214 83671 70270 83680
rect 46940 83632 46992 83638
rect 46940 83574 46992 83580
rect 59924 83570 59952 83671
rect 59912 83564 59964 83570
rect 59912 83506 59964 83512
rect 70228 83502 70256 83671
rect 70216 83496 70268 83502
rect 70216 83438 70268 83444
rect 108040 80507 108068 86158
rect 108550 85980 108858 85989
rect 108550 85978 108556 85980
rect 108612 85978 108636 85980
rect 108692 85978 108716 85980
rect 108772 85978 108796 85980
rect 108852 85978 108858 85980
rect 108612 85926 108614 85978
rect 108794 85926 108796 85978
rect 108550 85924 108556 85926
rect 108612 85924 108636 85926
rect 108692 85924 108716 85926
rect 108772 85924 108796 85926
rect 108852 85924 108858 85926
rect 108550 85915 108858 85924
rect 108026 80498 108082 80507
rect 108026 80433 108082 80442
rect 11980 59424 12032 59430
rect 11980 59366 12032 59372
rect 11808 41386 11928 41414
rect 11704 38752 11756 38758
rect 11704 38694 11756 38700
rect 11612 36916 11664 36922
rect 11612 36858 11664 36864
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11624 2242 11652 27066
rect 11716 4010 11744 38694
rect 11808 32499 11836 41386
rect 11980 37664 12032 37670
rect 11980 37606 12032 37612
rect 11888 34128 11940 34134
rect 11888 34070 11940 34076
rect 11794 32490 11850 32499
rect 11794 32425 11850 32434
rect 11900 31754 11928 34070
rect 11808 31726 11928 31754
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11808 2718 11836 31726
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11900 2786 11928 29106
rect 11888 2780 11940 2786
rect 11888 2722 11940 2728
rect 11796 2712 11848 2718
rect 11796 2654 11848 2660
rect 11612 2236 11664 2242
rect 11612 2178 11664 2184
rect 11610 1660 11918 1669
rect 11610 1658 11616 1660
rect 11672 1658 11696 1660
rect 11752 1658 11776 1660
rect 11832 1658 11856 1660
rect 11912 1658 11918 1660
rect 11672 1606 11674 1658
rect 11854 1606 11856 1658
rect 11610 1604 11616 1606
rect 11672 1604 11696 1606
rect 11752 1604 11776 1606
rect 11832 1604 11856 1606
rect 11912 1604 11918 1606
rect 11610 1595 11918 1604
rect 11520 1352 11572 1358
rect 11520 1294 11572 1300
rect 10950 1116 11258 1125
rect 10950 1114 10956 1116
rect 11012 1114 11036 1116
rect 11092 1114 11116 1116
rect 11172 1114 11196 1116
rect 11252 1114 11258 1116
rect 11012 1062 11014 1114
rect 11194 1062 11196 1114
rect 10950 1060 10956 1062
rect 11012 1060 11036 1062
rect 11092 1060 11116 1062
rect 11172 1060 11196 1062
rect 11252 1060 11258 1062
rect 10950 1051 11258 1060
rect 11992 746 12020 37606
rect 108026 20658 108082 20667
rect 108026 20593 108082 20602
rect 107934 18456 107990 18465
rect 107934 18391 107990 18400
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17880 3913 17908 3946
rect 54392 3936 54444 3942
rect 17866 3904 17922 3913
rect 17866 3839 17922 3848
rect 39210 3904 39266 3913
rect 39210 3839 39266 3848
rect 40314 3904 40370 3913
rect 40314 3839 40370 3848
rect 45006 3904 45062 3913
rect 45006 3839 45062 3848
rect 46110 3904 46166 3913
rect 46110 3839 46112 3848
rect 28722 3768 28778 3777
rect 28722 3703 28778 3712
rect 29826 3768 29882 3777
rect 29826 3703 29882 3712
rect 28736 3398 28764 3703
rect 29840 3534 29868 3703
rect 39224 3602 39252 3839
rect 40328 3806 40356 3839
rect 40316 3800 40368 3806
rect 40316 3742 40368 3748
rect 45020 3670 45048 3839
rect 46164 3839 46166 3848
rect 50894 3904 50950 3913
rect 50894 3839 50950 3848
rect 54390 3904 54392 3913
rect 54444 3904 54446 3913
rect 54390 3839 54446 3848
rect 46112 3810 46164 3816
rect 47490 3768 47546 3777
rect 50908 3738 50936 3839
rect 47490 3703 47546 3712
rect 50896 3732 50948 3738
rect 45008 3664 45060 3670
rect 45008 3606 45060 3612
rect 39212 3596 39264 3602
rect 39212 3538 39264 3544
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 28724 3392 28776 3398
rect 28724 3334 28776 3340
rect 29642 3360 29698 3369
rect 29642 3295 29698 3304
rect 32128 3324 32180 3330
rect 27528 2780 27580 2786
rect 27528 2722 27580 2728
rect 13210 1660 13518 1669
rect 13210 1658 13216 1660
rect 13272 1658 13296 1660
rect 13352 1658 13376 1660
rect 13432 1658 13456 1660
rect 13512 1658 13518 1660
rect 13272 1606 13274 1658
rect 13454 1606 13456 1658
rect 13210 1604 13216 1606
rect 13272 1604 13296 1606
rect 13352 1604 13376 1606
rect 13432 1604 13456 1606
rect 13512 1604 13518 1606
rect 13210 1595 13518 1604
rect 14810 1660 15118 1669
rect 14810 1658 14816 1660
rect 14872 1658 14896 1660
rect 14952 1658 14976 1660
rect 15032 1658 15056 1660
rect 15112 1658 15118 1660
rect 14872 1606 14874 1658
rect 15054 1606 15056 1658
rect 14810 1604 14816 1606
rect 14872 1604 14896 1606
rect 14952 1604 14976 1606
rect 15032 1604 15056 1606
rect 15112 1604 15118 1606
rect 14810 1595 15118 1604
rect 16410 1660 16718 1669
rect 16410 1658 16416 1660
rect 16472 1658 16496 1660
rect 16552 1658 16576 1660
rect 16632 1658 16656 1660
rect 16712 1658 16718 1660
rect 16472 1606 16474 1658
rect 16654 1606 16656 1658
rect 16410 1604 16416 1606
rect 16472 1604 16496 1606
rect 16552 1604 16576 1606
rect 16632 1604 16656 1606
rect 16712 1604 16718 1606
rect 16410 1595 16718 1604
rect 18010 1660 18318 1669
rect 18010 1658 18016 1660
rect 18072 1658 18096 1660
rect 18152 1658 18176 1660
rect 18232 1658 18256 1660
rect 18312 1658 18318 1660
rect 18072 1606 18074 1658
rect 18254 1606 18256 1658
rect 18010 1604 18016 1606
rect 18072 1604 18096 1606
rect 18152 1604 18176 1606
rect 18232 1604 18256 1606
rect 18312 1604 18318 1606
rect 18010 1595 18318 1604
rect 19610 1660 19918 1669
rect 19610 1658 19616 1660
rect 19672 1658 19696 1660
rect 19752 1658 19776 1660
rect 19832 1658 19856 1660
rect 19912 1658 19918 1660
rect 19672 1606 19674 1658
rect 19854 1606 19856 1658
rect 19610 1604 19616 1606
rect 19672 1604 19696 1606
rect 19752 1604 19776 1606
rect 19832 1604 19856 1606
rect 19912 1604 19918 1606
rect 19610 1595 19918 1604
rect 21210 1660 21518 1669
rect 21210 1658 21216 1660
rect 21272 1658 21296 1660
rect 21352 1658 21376 1660
rect 21432 1658 21456 1660
rect 21512 1658 21518 1660
rect 21272 1606 21274 1658
rect 21454 1606 21456 1658
rect 21210 1604 21216 1606
rect 21272 1604 21296 1606
rect 21352 1604 21376 1606
rect 21432 1604 21456 1606
rect 21512 1604 21518 1606
rect 21210 1595 21518 1604
rect 22810 1660 23118 1669
rect 22810 1658 22816 1660
rect 22872 1658 22896 1660
rect 22952 1658 22976 1660
rect 23032 1658 23056 1660
rect 23112 1658 23118 1660
rect 22872 1606 22874 1658
rect 23054 1606 23056 1658
rect 22810 1604 22816 1606
rect 22872 1604 22896 1606
rect 22952 1604 22976 1606
rect 23032 1604 23056 1606
rect 23112 1604 23118 1606
rect 22810 1595 23118 1604
rect 24410 1660 24718 1669
rect 24410 1658 24416 1660
rect 24472 1658 24496 1660
rect 24552 1658 24576 1660
rect 24632 1658 24656 1660
rect 24712 1658 24718 1660
rect 24472 1606 24474 1658
rect 24654 1606 24656 1658
rect 24410 1604 24416 1606
rect 24472 1604 24496 1606
rect 24552 1604 24576 1606
rect 24632 1604 24656 1606
rect 24712 1604 24718 1606
rect 24410 1595 24718 1604
rect 26010 1660 26318 1669
rect 26010 1658 26016 1660
rect 26072 1658 26096 1660
rect 26152 1658 26176 1660
rect 26232 1658 26256 1660
rect 26312 1658 26318 1660
rect 26072 1606 26074 1658
rect 26254 1606 26256 1658
rect 26010 1604 26016 1606
rect 26072 1604 26096 1606
rect 26152 1604 26176 1606
rect 26232 1604 26256 1606
rect 26312 1604 26318 1606
rect 26010 1595 26318 1604
rect 23664 1488 23716 1494
rect 23664 1430 23716 1436
rect 23204 1420 23256 1426
rect 23204 1362 23256 1368
rect 17224 1216 17276 1222
rect 17224 1158 17276 1164
rect 22928 1216 22980 1222
rect 22928 1158 22980 1164
rect 12550 1116 12858 1125
rect 12550 1114 12556 1116
rect 12612 1114 12636 1116
rect 12692 1114 12716 1116
rect 12772 1114 12796 1116
rect 12852 1114 12858 1116
rect 12612 1062 12614 1114
rect 12794 1062 12796 1114
rect 12550 1060 12556 1062
rect 12612 1060 12636 1062
rect 12692 1060 12716 1062
rect 12772 1060 12796 1062
rect 12852 1060 12858 1062
rect 12550 1051 12858 1060
rect 14150 1116 14458 1125
rect 14150 1114 14156 1116
rect 14212 1114 14236 1116
rect 14292 1114 14316 1116
rect 14372 1114 14396 1116
rect 14452 1114 14458 1116
rect 14212 1062 14214 1114
rect 14394 1062 14396 1114
rect 14150 1060 14156 1062
rect 14212 1060 14236 1062
rect 14292 1060 14316 1062
rect 14372 1060 14396 1062
rect 14452 1060 14458 1062
rect 14150 1051 14458 1060
rect 15750 1116 16058 1125
rect 15750 1114 15756 1116
rect 15812 1114 15836 1116
rect 15892 1114 15916 1116
rect 15972 1114 15996 1116
rect 16052 1114 16058 1116
rect 15812 1062 15814 1114
rect 15994 1062 15996 1114
rect 15750 1060 15756 1062
rect 15812 1060 15836 1062
rect 15892 1060 15916 1062
rect 15972 1060 15996 1062
rect 16052 1060 16058 1062
rect 15750 1051 16058 1060
rect 17236 1018 17264 1158
rect 17350 1116 17658 1125
rect 17350 1114 17356 1116
rect 17412 1114 17436 1116
rect 17492 1114 17516 1116
rect 17572 1114 17596 1116
rect 17652 1114 17658 1116
rect 17412 1062 17414 1114
rect 17594 1062 17596 1114
rect 17350 1060 17356 1062
rect 17412 1060 17436 1062
rect 17492 1060 17516 1062
rect 17572 1060 17596 1062
rect 17652 1060 17658 1062
rect 17350 1051 17658 1060
rect 18950 1116 19258 1125
rect 18950 1114 18956 1116
rect 19012 1114 19036 1116
rect 19092 1114 19116 1116
rect 19172 1114 19196 1116
rect 19252 1114 19258 1116
rect 19012 1062 19014 1114
rect 19194 1062 19196 1114
rect 18950 1060 18956 1062
rect 19012 1060 19036 1062
rect 19092 1060 19116 1062
rect 19172 1060 19196 1062
rect 19252 1060 19258 1062
rect 18950 1051 19258 1060
rect 20550 1116 20858 1125
rect 20550 1114 20556 1116
rect 20612 1114 20636 1116
rect 20692 1114 20716 1116
rect 20772 1114 20796 1116
rect 20852 1114 20858 1116
rect 20612 1062 20614 1114
rect 20794 1062 20796 1114
rect 20550 1060 20556 1062
rect 20612 1060 20636 1062
rect 20692 1060 20716 1062
rect 20772 1060 20796 1062
rect 20852 1060 20858 1062
rect 20550 1051 20858 1060
rect 22150 1116 22458 1125
rect 22150 1114 22156 1116
rect 22212 1114 22236 1116
rect 22292 1114 22316 1116
rect 22372 1114 22396 1116
rect 22452 1114 22458 1116
rect 22212 1062 22214 1114
rect 22394 1062 22396 1114
rect 22150 1060 22156 1062
rect 22212 1060 22236 1062
rect 22292 1060 22316 1062
rect 22372 1060 22396 1062
rect 22452 1060 22458 1062
rect 22150 1051 22458 1060
rect 17224 1012 17276 1018
rect 17224 954 17276 960
rect 11980 740 12032 746
rect 11980 682 12032 688
rect 10598 504 10654 513
rect 10508 468 10560 474
rect 10598 439 10654 448
rect 10508 410 10560 416
rect 1306 303 1362 312
rect 9864 332 9916 338
rect 9864 274 9916 280
rect 22940 134 22968 1158
rect 23216 474 23244 1362
rect 23480 1284 23532 1290
rect 23480 1226 23532 1232
rect 23492 746 23520 1226
rect 23480 740 23532 746
rect 23480 682 23532 688
rect 23676 542 23704 1430
rect 27540 1426 27568 2722
rect 27610 1660 27918 1669
rect 27610 1658 27616 1660
rect 27672 1658 27696 1660
rect 27752 1658 27776 1660
rect 27832 1658 27856 1660
rect 27912 1658 27918 1660
rect 27672 1606 27674 1658
rect 27854 1606 27856 1658
rect 27610 1604 27616 1606
rect 27672 1604 27696 1606
rect 27752 1604 27776 1606
rect 27832 1604 27856 1606
rect 27912 1604 27918 1606
rect 27610 1595 27918 1604
rect 29210 1660 29518 1669
rect 29210 1658 29216 1660
rect 29272 1658 29296 1660
rect 29352 1658 29376 1660
rect 29432 1658 29456 1660
rect 29512 1658 29518 1660
rect 29272 1606 29274 1658
rect 29454 1606 29456 1658
rect 29210 1604 29216 1606
rect 29272 1604 29296 1606
rect 29352 1604 29376 1606
rect 29432 1604 29456 1606
rect 29512 1604 29518 1606
rect 29210 1595 29518 1604
rect 27528 1420 27580 1426
rect 27528 1362 27580 1368
rect 29656 1358 29684 3295
rect 32128 3266 32180 3272
rect 32036 2576 32088 2582
rect 32036 2518 32088 2524
rect 32048 2417 32076 2518
rect 32034 2408 32090 2417
rect 32034 2343 32090 2352
rect 30810 1660 31118 1669
rect 30810 1658 30816 1660
rect 30872 1658 30896 1660
rect 30952 1658 30976 1660
rect 31032 1658 31056 1660
rect 31112 1658 31118 1660
rect 30872 1606 30874 1658
rect 31054 1606 31056 1658
rect 30810 1604 30816 1606
rect 30872 1604 30896 1606
rect 30952 1604 30976 1606
rect 31032 1604 31056 1606
rect 31112 1604 31118 1606
rect 30810 1595 31118 1604
rect 32140 1358 32168 3266
rect 47504 3194 47532 3703
rect 50896 3674 50948 3680
rect 54576 3460 54628 3466
rect 54576 3402 54628 3408
rect 47492 3188 47544 3194
rect 47492 3130 47544 3136
rect 34704 2712 34756 2718
rect 34704 2654 34756 2660
rect 37002 2680 37058 2689
rect 32410 1660 32718 1669
rect 32410 1658 32416 1660
rect 32472 1658 32496 1660
rect 32552 1658 32576 1660
rect 32632 1658 32656 1660
rect 32712 1658 32718 1660
rect 32472 1606 32474 1658
rect 32654 1606 32656 1658
rect 32410 1604 32416 1606
rect 32472 1604 32496 1606
rect 32552 1604 32576 1606
rect 32632 1604 32656 1606
rect 32712 1604 32718 1606
rect 32410 1595 32718 1604
rect 34010 1660 34318 1669
rect 34010 1658 34016 1660
rect 34072 1658 34096 1660
rect 34152 1658 34176 1660
rect 34232 1658 34256 1660
rect 34312 1658 34318 1660
rect 34072 1606 34074 1658
rect 34254 1606 34256 1658
rect 34010 1604 34016 1606
rect 34072 1604 34096 1606
rect 34152 1604 34176 1606
rect 34232 1604 34256 1606
rect 34312 1604 34318 1606
rect 34010 1595 34318 1604
rect 34716 1426 34744 2654
rect 37002 2615 37058 2624
rect 49698 2680 49754 2689
rect 49698 2615 49754 2624
rect 37016 2242 37044 2615
rect 43812 2508 43864 2514
rect 43812 2450 43864 2456
rect 43824 2417 43852 2450
rect 42798 2408 42854 2417
rect 42798 2343 42854 2352
rect 43810 2408 43866 2417
rect 43810 2343 43866 2352
rect 48594 2408 48650 2417
rect 48594 2343 48650 2352
rect 37004 2236 37056 2242
rect 37004 2178 37056 2184
rect 37462 2136 37518 2145
rect 37518 2094 37596 2122
rect 37462 2071 37518 2080
rect 35610 1660 35918 1669
rect 35610 1658 35616 1660
rect 35672 1658 35696 1660
rect 35752 1658 35776 1660
rect 35832 1658 35856 1660
rect 35912 1658 35918 1660
rect 35672 1606 35674 1658
rect 35854 1606 35856 1658
rect 35610 1604 35616 1606
rect 35672 1604 35696 1606
rect 35752 1604 35776 1606
rect 35832 1604 35856 1606
rect 35912 1604 35918 1606
rect 35610 1595 35918 1604
rect 37210 1660 37518 1669
rect 37210 1658 37216 1660
rect 37272 1658 37296 1660
rect 37352 1658 37376 1660
rect 37432 1658 37456 1660
rect 37512 1658 37518 1660
rect 37272 1606 37274 1658
rect 37454 1606 37456 1658
rect 37210 1604 37216 1606
rect 37272 1604 37296 1606
rect 37352 1604 37376 1606
rect 37432 1604 37456 1606
rect 37512 1604 37518 1606
rect 37210 1595 37518 1604
rect 34704 1420 34756 1426
rect 34704 1362 34756 1368
rect 37568 1358 37596 2094
rect 42812 2038 42840 2343
rect 48608 2174 48636 2343
rect 49712 2310 49740 2615
rect 49700 2304 49752 2310
rect 49700 2246 49752 2252
rect 48596 2168 48648 2174
rect 48596 2110 48648 2116
rect 42800 2032 42852 2038
rect 42800 1974 42852 1980
rect 38810 1660 39118 1669
rect 38810 1658 38816 1660
rect 38872 1658 38896 1660
rect 38952 1658 38976 1660
rect 39032 1658 39056 1660
rect 39112 1658 39118 1660
rect 38872 1606 38874 1658
rect 39054 1606 39056 1658
rect 38810 1604 38816 1606
rect 38872 1604 38896 1606
rect 38952 1604 38976 1606
rect 39032 1604 39056 1606
rect 39112 1604 39118 1606
rect 38810 1595 39118 1604
rect 40410 1660 40718 1669
rect 40410 1658 40416 1660
rect 40472 1658 40496 1660
rect 40552 1658 40576 1660
rect 40632 1658 40656 1660
rect 40712 1658 40718 1660
rect 40472 1606 40474 1658
rect 40654 1606 40656 1658
rect 40410 1604 40416 1606
rect 40472 1604 40496 1606
rect 40552 1604 40576 1606
rect 40632 1604 40656 1606
rect 40712 1604 40718 1606
rect 40410 1595 40718 1604
rect 42010 1660 42318 1669
rect 42010 1658 42016 1660
rect 42072 1658 42096 1660
rect 42152 1658 42176 1660
rect 42232 1658 42256 1660
rect 42312 1658 42318 1660
rect 42072 1606 42074 1658
rect 42254 1606 42256 1658
rect 42010 1604 42016 1606
rect 42072 1604 42096 1606
rect 42152 1604 42176 1606
rect 42232 1604 42256 1606
rect 42312 1604 42318 1606
rect 42010 1595 42318 1604
rect 43610 1660 43918 1669
rect 43610 1658 43616 1660
rect 43672 1658 43696 1660
rect 43752 1658 43776 1660
rect 43832 1658 43856 1660
rect 43912 1658 43918 1660
rect 43672 1606 43674 1658
rect 43854 1606 43856 1658
rect 43610 1604 43616 1606
rect 43672 1604 43696 1606
rect 43752 1604 43776 1606
rect 43832 1604 43856 1606
rect 43912 1604 43918 1606
rect 43610 1595 43918 1604
rect 45210 1660 45518 1669
rect 45210 1658 45216 1660
rect 45272 1658 45296 1660
rect 45352 1658 45376 1660
rect 45432 1658 45456 1660
rect 45512 1658 45518 1660
rect 45272 1606 45274 1658
rect 45454 1606 45456 1658
rect 45210 1604 45216 1606
rect 45272 1604 45296 1606
rect 45352 1604 45376 1606
rect 45432 1604 45456 1606
rect 45512 1604 45518 1606
rect 45210 1595 45518 1604
rect 46810 1660 47118 1669
rect 46810 1658 46816 1660
rect 46872 1658 46896 1660
rect 46952 1658 46976 1660
rect 47032 1658 47056 1660
rect 47112 1658 47118 1660
rect 46872 1606 46874 1658
rect 47054 1606 47056 1658
rect 46810 1604 46816 1606
rect 46872 1604 46896 1606
rect 46952 1604 46976 1606
rect 47032 1604 47056 1606
rect 47112 1604 47118 1606
rect 46810 1595 47118 1604
rect 48410 1660 48718 1669
rect 48410 1658 48416 1660
rect 48472 1658 48496 1660
rect 48552 1658 48576 1660
rect 48632 1658 48656 1660
rect 48712 1658 48718 1660
rect 48472 1606 48474 1658
rect 48654 1606 48656 1658
rect 48410 1604 48416 1606
rect 48472 1604 48496 1606
rect 48552 1604 48576 1606
rect 48632 1604 48656 1606
rect 48712 1604 48718 1606
rect 48410 1595 48718 1604
rect 50010 1660 50318 1669
rect 50010 1658 50016 1660
rect 50072 1658 50096 1660
rect 50152 1658 50176 1660
rect 50232 1658 50256 1660
rect 50312 1658 50318 1660
rect 50072 1606 50074 1658
rect 50254 1606 50256 1658
rect 50010 1604 50016 1606
rect 50072 1604 50096 1606
rect 50152 1604 50176 1606
rect 50232 1604 50256 1606
rect 50312 1604 50318 1606
rect 50010 1595 50318 1604
rect 51610 1660 51918 1669
rect 51610 1658 51616 1660
rect 51672 1658 51696 1660
rect 51752 1658 51776 1660
rect 51832 1658 51856 1660
rect 51912 1658 51918 1660
rect 51672 1606 51674 1658
rect 51854 1606 51856 1658
rect 51610 1604 51616 1606
rect 51672 1604 51696 1606
rect 51752 1604 51776 1606
rect 51832 1604 51856 1606
rect 51912 1604 51918 1606
rect 51610 1595 51918 1604
rect 53210 1660 53518 1669
rect 53210 1658 53216 1660
rect 53272 1658 53296 1660
rect 53352 1658 53376 1660
rect 53432 1658 53456 1660
rect 53512 1658 53518 1660
rect 53272 1606 53274 1658
rect 53454 1606 53456 1658
rect 53210 1604 53216 1606
rect 53272 1604 53296 1606
rect 53352 1604 53376 1606
rect 53432 1604 53456 1606
rect 53512 1604 53518 1606
rect 53210 1595 53518 1604
rect 24124 1352 24176 1358
rect 24124 1294 24176 1300
rect 27804 1352 27856 1358
rect 27804 1294 27856 1300
rect 29644 1352 29696 1358
rect 32128 1352 32180 1358
rect 29644 1294 29696 1300
rect 30562 1320 30618 1329
rect 23750 1116 24058 1125
rect 23750 1114 23756 1116
rect 23812 1114 23836 1116
rect 23892 1114 23916 1116
rect 23972 1114 23996 1116
rect 24052 1114 24058 1116
rect 23812 1062 23814 1114
rect 23994 1062 23996 1114
rect 23750 1060 23756 1062
rect 23812 1060 23836 1062
rect 23892 1060 23916 1062
rect 23972 1060 23996 1062
rect 24052 1060 24058 1062
rect 23750 1051 24058 1060
rect 24136 950 24164 1294
rect 27344 1284 27396 1290
rect 27344 1226 27396 1232
rect 26240 1216 26292 1222
rect 26240 1158 26292 1164
rect 26332 1216 26384 1222
rect 26332 1158 26384 1164
rect 25350 1116 25658 1125
rect 25350 1114 25356 1116
rect 25412 1114 25436 1116
rect 25492 1114 25516 1116
rect 25572 1114 25596 1116
rect 25652 1114 25658 1116
rect 25412 1062 25414 1114
rect 25594 1062 25596 1114
rect 25350 1060 25356 1062
rect 25412 1060 25436 1062
rect 25492 1060 25516 1062
rect 25572 1060 25596 1062
rect 25652 1060 25658 1062
rect 25350 1051 25658 1060
rect 26252 1018 26280 1158
rect 26240 1012 26292 1018
rect 26240 954 26292 960
rect 24124 944 24176 950
rect 26344 921 26372 1158
rect 26950 1116 27258 1125
rect 26950 1114 26956 1116
rect 27012 1114 27036 1116
rect 27092 1114 27116 1116
rect 27172 1114 27196 1116
rect 27252 1114 27258 1116
rect 27012 1062 27014 1114
rect 27194 1062 27196 1114
rect 26950 1060 26956 1062
rect 27012 1060 27036 1062
rect 27092 1060 27116 1062
rect 27172 1060 27196 1062
rect 27252 1060 27258 1062
rect 26950 1051 27258 1060
rect 24124 886 24176 892
rect 26330 912 26386 921
rect 26330 847 26386 856
rect 24400 808 24452 814
rect 24400 750 24452 756
rect 23664 536 23716 542
rect 23664 478 23716 484
rect 23204 468 23256 474
rect 23204 410 23256 416
rect 24412 270 24440 750
rect 27356 610 27384 1226
rect 27816 610 27844 1294
rect 32128 1294 32180 1300
rect 32404 1352 32456 1358
rect 32404 1294 32456 1300
rect 33140 1352 33192 1358
rect 33876 1352 33928 1358
rect 33140 1294 33192 1300
rect 33230 1320 33286 1329
rect 30562 1255 30618 1264
rect 29460 1216 29512 1222
rect 29460 1158 29512 1164
rect 29736 1216 29788 1222
rect 29736 1158 29788 1164
rect 29828 1216 29880 1222
rect 29828 1158 29880 1164
rect 28550 1116 28858 1125
rect 28550 1114 28556 1116
rect 28612 1114 28636 1116
rect 28692 1114 28716 1116
rect 28772 1114 28796 1116
rect 28852 1114 28858 1116
rect 28612 1062 28614 1114
rect 28794 1062 28796 1114
rect 28550 1060 28556 1062
rect 28612 1060 28636 1062
rect 28692 1060 28716 1062
rect 28772 1060 28796 1062
rect 28852 1060 28858 1062
rect 28550 1051 28858 1060
rect 29472 746 29500 1158
rect 29748 1018 29776 1158
rect 29736 1012 29788 1018
rect 29736 954 29788 960
rect 29840 898 29868 1158
rect 30150 1116 30458 1125
rect 30150 1114 30156 1116
rect 30212 1114 30236 1116
rect 30292 1114 30316 1116
rect 30372 1114 30396 1116
rect 30452 1114 30458 1116
rect 30212 1062 30214 1114
rect 30394 1062 30396 1114
rect 30150 1060 30156 1062
rect 30212 1060 30236 1062
rect 30292 1060 30316 1062
rect 30372 1060 30396 1062
rect 30452 1060 30458 1062
rect 30150 1051 30458 1060
rect 29564 870 29868 898
rect 29564 814 29592 870
rect 29552 808 29604 814
rect 29552 750 29604 756
rect 29460 740 29512 746
rect 29460 682 29512 688
rect 27344 604 27396 610
rect 27344 546 27396 552
rect 27804 604 27856 610
rect 27804 546 27856 552
rect 30576 270 30604 1255
rect 30656 1216 30708 1222
rect 30656 1158 30708 1164
rect 32312 1216 32364 1222
rect 32312 1158 32364 1164
rect 30668 814 30696 1158
rect 31750 1116 32058 1125
rect 31750 1114 31756 1116
rect 31812 1114 31836 1116
rect 31892 1114 31916 1116
rect 31972 1114 31996 1116
rect 32052 1114 32058 1116
rect 31812 1062 31814 1114
rect 31994 1062 31996 1114
rect 31750 1060 31756 1062
rect 31812 1060 31836 1062
rect 31892 1060 31916 1062
rect 31972 1060 31996 1062
rect 32052 1060 32058 1062
rect 31750 1051 32058 1060
rect 30656 808 30708 814
rect 30656 750 30708 756
rect 32324 746 32352 1158
rect 32220 740 32272 746
rect 32220 682 32272 688
rect 32312 740 32364 746
rect 32312 682 32364 688
rect 32232 649 32260 682
rect 32218 640 32274 649
rect 32218 575 32274 584
rect 32416 542 32444 1294
rect 32404 536 32456 542
rect 32404 478 32456 484
rect 33152 377 33180 1294
rect 37372 1352 37424 1358
rect 33876 1294 33928 1300
rect 34518 1320 34574 1329
rect 33230 1255 33286 1264
rect 33138 368 33194 377
rect 33244 338 33272 1255
rect 33350 1116 33658 1125
rect 33350 1114 33356 1116
rect 33412 1114 33436 1116
rect 33492 1114 33516 1116
rect 33572 1114 33596 1116
rect 33652 1114 33658 1116
rect 33412 1062 33414 1114
rect 33594 1062 33596 1114
rect 33350 1060 33356 1062
rect 33412 1060 33436 1062
rect 33492 1060 33516 1062
rect 33572 1060 33596 1062
rect 33652 1060 33658 1062
rect 33350 1051 33658 1060
rect 33888 950 33916 1294
rect 34518 1255 34574 1264
rect 37278 1320 37334 1329
rect 37372 1294 37424 1300
rect 37556 1352 37608 1358
rect 37556 1294 37608 1300
rect 37740 1352 37792 1358
rect 37740 1294 37792 1300
rect 37278 1255 37334 1264
rect 33876 944 33928 950
rect 33876 886 33928 892
rect 34532 338 34560 1255
rect 37292 1222 37320 1255
rect 37280 1216 37332 1222
rect 37280 1158 37332 1164
rect 34950 1116 35258 1125
rect 34950 1114 34956 1116
rect 35012 1114 35036 1116
rect 35092 1114 35116 1116
rect 35172 1114 35196 1116
rect 35252 1114 35258 1116
rect 35012 1062 35014 1114
rect 35194 1062 35196 1114
rect 34950 1060 34956 1062
rect 35012 1060 35036 1062
rect 35092 1060 35116 1062
rect 35172 1060 35196 1062
rect 35252 1060 35258 1062
rect 34950 1051 35258 1060
rect 36550 1116 36858 1125
rect 36550 1114 36556 1116
rect 36612 1114 36636 1116
rect 36692 1114 36716 1116
rect 36772 1114 36796 1116
rect 36852 1114 36858 1116
rect 36612 1062 36614 1114
rect 36794 1062 36796 1114
rect 36550 1060 36556 1062
rect 36612 1060 36636 1062
rect 36692 1060 36716 1062
rect 36772 1060 36796 1062
rect 36852 1060 36858 1062
rect 36550 1051 36858 1060
rect 37384 610 37412 1294
rect 37568 1222 37596 1294
rect 37556 1216 37608 1222
rect 37556 1158 37608 1164
rect 37752 678 37780 1294
rect 38150 1116 38458 1125
rect 38150 1114 38156 1116
rect 38212 1114 38236 1116
rect 38292 1114 38316 1116
rect 38372 1114 38396 1116
rect 38452 1114 38458 1116
rect 38212 1062 38214 1114
rect 38394 1062 38396 1114
rect 38150 1060 38156 1062
rect 38212 1060 38236 1062
rect 38292 1060 38316 1062
rect 38372 1060 38396 1062
rect 38452 1060 38458 1062
rect 38150 1051 38458 1060
rect 39750 1116 40058 1125
rect 39750 1114 39756 1116
rect 39812 1114 39836 1116
rect 39892 1114 39916 1116
rect 39972 1114 39996 1116
rect 40052 1114 40058 1116
rect 39812 1062 39814 1114
rect 39994 1062 39996 1114
rect 39750 1060 39756 1062
rect 39812 1060 39836 1062
rect 39892 1060 39916 1062
rect 39972 1060 39996 1062
rect 40052 1060 40058 1062
rect 39750 1051 40058 1060
rect 41350 1116 41658 1125
rect 41350 1114 41356 1116
rect 41412 1114 41436 1116
rect 41492 1114 41516 1116
rect 41572 1114 41596 1116
rect 41652 1114 41658 1116
rect 41412 1062 41414 1114
rect 41594 1062 41596 1114
rect 41350 1060 41356 1062
rect 41412 1060 41436 1062
rect 41492 1060 41516 1062
rect 41572 1060 41596 1062
rect 41652 1060 41658 1062
rect 41350 1051 41658 1060
rect 42950 1116 43258 1125
rect 42950 1114 42956 1116
rect 43012 1114 43036 1116
rect 43092 1114 43116 1116
rect 43172 1114 43196 1116
rect 43252 1114 43258 1116
rect 43012 1062 43014 1114
rect 43194 1062 43196 1114
rect 42950 1060 42956 1062
rect 43012 1060 43036 1062
rect 43092 1060 43116 1062
rect 43172 1060 43196 1062
rect 43252 1060 43258 1062
rect 42950 1051 43258 1060
rect 44550 1116 44858 1125
rect 44550 1114 44556 1116
rect 44612 1114 44636 1116
rect 44692 1114 44716 1116
rect 44772 1114 44796 1116
rect 44852 1114 44858 1116
rect 44612 1062 44614 1114
rect 44794 1062 44796 1114
rect 44550 1060 44556 1062
rect 44612 1060 44636 1062
rect 44692 1060 44716 1062
rect 44772 1060 44796 1062
rect 44852 1060 44858 1062
rect 44550 1051 44858 1060
rect 46150 1116 46458 1125
rect 46150 1114 46156 1116
rect 46212 1114 46236 1116
rect 46292 1114 46316 1116
rect 46372 1114 46396 1116
rect 46452 1114 46458 1116
rect 46212 1062 46214 1114
rect 46394 1062 46396 1114
rect 46150 1060 46156 1062
rect 46212 1060 46236 1062
rect 46292 1060 46316 1062
rect 46372 1060 46396 1062
rect 46452 1060 46458 1062
rect 46150 1051 46458 1060
rect 47750 1116 48058 1125
rect 47750 1114 47756 1116
rect 47812 1114 47836 1116
rect 47892 1114 47916 1116
rect 47972 1114 47996 1116
rect 48052 1114 48058 1116
rect 47812 1062 47814 1114
rect 47994 1062 47996 1114
rect 47750 1060 47756 1062
rect 47812 1060 47836 1062
rect 47892 1060 47916 1062
rect 47972 1060 47996 1062
rect 48052 1060 48058 1062
rect 47750 1051 48058 1060
rect 49350 1116 49658 1125
rect 49350 1114 49356 1116
rect 49412 1114 49436 1116
rect 49492 1114 49516 1116
rect 49572 1114 49596 1116
rect 49652 1114 49658 1116
rect 49412 1062 49414 1114
rect 49594 1062 49596 1114
rect 49350 1060 49356 1062
rect 49412 1060 49436 1062
rect 49492 1060 49516 1062
rect 49572 1060 49596 1062
rect 49652 1060 49658 1062
rect 49350 1051 49658 1060
rect 50950 1116 51258 1125
rect 50950 1114 50956 1116
rect 51012 1114 51036 1116
rect 51092 1114 51116 1116
rect 51172 1114 51196 1116
rect 51252 1114 51258 1116
rect 51012 1062 51014 1114
rect 51194 1062 51196 1114
rect 50950 1060 50956 1062
rect 51012 1060 51036 1062
rect 51092 1060 51116 1062
rect 51172 1060 51196 1062
rect 51252 1060 51258 1062
rect 50950 1051 51258 1060
rect 52550 1116 52858 1125
rect 52550 1114 52556 1116
rect 52612 1114 52636 1116
rect 52692 1114 52716 1116
rect 52772 1114 52796 1116
rect 52852 1114 52858 1116
rect 52612 1062 52614 1114
rect 52794 1062 52796 1114
rect 52550 1060 52556 1062
rect 52612 1060 52636 1062
rect 52692 1060 52716 1062
rect 52772 1060 52796 1062
rect 52852 1060 52858 1062
rect 52550 1051 52858 1060
rect 54150 1116 54458 1125
rect 54150 1114 54156 1116
rect 54212 1114 54236 1116
rect 54292 1114 54316 1116
rect 54372 1114 54396 1116
rect 54452 1114 54458 1116
rect 54212 1062 54214 1114
rect 54394 1062 54396 1114
rect 54150 1060 54156 1062
rect 54212 1060 54236 1062
rect 54292 1060 54316 1062
rect 54372 1060 54396 1062
rect 54452 1060 54458 1062
rect 54150 1051 54458 1060
rect 54588 762 54616 3402
rect 55402 2680 55458 2689
rect 55402 2615 55458 2624
rect 57978 2680 58034 2689
rect 107948 2650 107976 18391
rect 108040 3505 108068 20593
rect 108118 17666 108174 17675
rect 108118 17601 108174 17610
rect 108132 3641 108160 17601
rect 108118 3632 108174 3641
rect 108118 3567 108174 3576
rect 108026 3496 108082 3505
rect 108026 3431 108082 3440
rect 57978 2615 58034 2624
rect 107936 2644 107988 2650
rect 55416 2446 55444 2615
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 57992 2378 58020 2615
rect 107936 2586 107988 2592
rect 94962 2544 95018 2553
rect 94962 2479 95018 2488
rect 57980 2372 58032 2378
rect 57980 2314 58032 2320
rect 94976 2106 95004 2479
rect 94964 2100 95016 2106
rect 94964 2042 95016 2048
rect 54810 1660 55118 1669
rect 54810 1658 54816 1660
rect 54872 1658 54896 1660
rect 54952 1658 54976 1660
rect 55032 1658 55056 1660
rect 55112 1658 55118 1660
rect 54872 1606 54874 1658
rect 55054 1606 55056 1658
rect 54810 1604 54816 1606
rect 54872 1604 54896 1606
rect 54952 1604 54976 1606
rect 55032 1604 55056 1606
rect 55112 1604 55118 1606
rect 54810 1595 55118 1604
rect 56410 1660 56718 1669
rect 56410 1658 56416 1660
rect 56472 1658 56496 1660
rect 56552 1658 56576 1660
rect 56632 1658 56656 1660
rect 56712 1658 56718 1660
rect 56472 1606 56474 1658
rect 56654 1606 56656 1658
rect 56410 1604 56416 1606
rect 56472 1604 56496 1606
rect 56552 1604 56576 1606
rect 56632 1604 56656 1606
rect 56712 1604 56718 1606
rect 56410 1595 56718 1604
rect 58010 1660 58318 1669
rect 58010 1658 58016 1660
rect 58072 1658 58096 1660
rect 58152 1658 58176 1660
rect 58232 1658 58256 1660
rect 58312 1658 58318 1660
rect 58072 1606 58074 1658
rect 58254 1606 58256 1658
rect 58010 1604 58016 1606
rect 58072 1604 58096 1606
rect 58152 1604 58176 1606
rect 58232 1604 58256 1606
rect 58312 1604 58318 1606
rect 58010 1595 58318 1604
rect 59610 1660 59918 1669
rect 59610 1658 59616 1660
rect 59672 1658 59696 1660
rect 59752 1658 59776 1660
rect 59832 1658 59856 1660
rect 59912 1658 59918 1660
rect 59672 1606 59674 1658
rect 59854 1606 59856 1658
rect 59610 1604 59616 1606
rect 59672 1604 59696 1606
rect 59752 1604 59776 1606
rect 59832 1604 59856 1606
rect 59912 1604 59918 1606
rect 59610 1595 59918 1604
rect 61210 1660 61518 1669
rect 61210 1658 61216 1660
rect 61272 1658 61296 1660
rect 61352 1658 61376 1660
rect 61432 1658 61456 1660
rect 61512 1658 61518 1660
rect 61272 1606 61274 1658
rect 61454 1606 61456 1658
rect 61210 1604 61216 1606
rect 61272 1604 61296 1606
rect 61352 1604 61376 1606
rect 61432 1604 61456 1606
rect 61512 1604 61518 1606
rect 61210 1595 61518 1604
rect 62810 1660 63118 1669
rect 62810 1658 62816 1660
rect 62872 1658 62896 1660
rect 62952 1658 62976 1660
rect 63032 1658 63056 1660
rect 63112 1658 63118 1660
rect 62872 1606 62874 1658
rect 63054 1606 63056 1658
rect 62810 1604 62816 1606
rect 62872 1604 62896 1606
rect 62952 1604 62976 1606
rect 63032 1604 63056 1606
rect 63112 1604 63118 1606
rect 62810 1595 63118 1604
rect 64410 1660 64718 1669
rect 64410 1658 64416 1660
rect 64472 1658 64496 1660
rect 64552 1658 64576 1660
rect 64632 1658 64656 1660
rect 64712 1658 64718 1660
rect 64472 1606 64474 1658
rect 64654 1606 64656 1658
rect 64410 1604 64416 1606
rect 64472 1604 64496 1606
rect 64552 1604 64576 1606
rect 64632 1604 64656 1606
rect 64712 1604 64718 1606
rect 64410 1595 64718 1604
rect 66010 1660 66318 1669
rect 66010 1658 66016 1660
rect 66072 1658 66096 1660
rect 66152 1658 66176 1660
rect 66232 1658 66256 1660
rect 66312 1658 66318 1660
rect 66072 1606 66074 1658
rect 66254 1606 66256 1658
rect 66010 1604 66016 1606
rect 66072 1604 66096 1606
rect 66152 1604 66176 1606
rect 66232 1604 66256 1606
rect 66312 1604 66318 1606
rect 66010 1595 66318 1604
rect 67610 1660 67918 1669
rect 67610 1658 67616 1660
rect 67672 1658 67696 1660
rect 67752 1658 67776 1660
rect 67832 1658 67856 1660
rect 67912 1658 67918 1660
rect 67672 1606 67674 1658
rect 67854 1606 67856 1658
rect 67610 1604 67616 1606
rect 67672 1604 67696 1606
rect 67752 1604 67776 1606
rect 67832 1604 67856 1606
rect 67912 1604 67918 1606
rect 67610 1595 67918 1604
rect 69210 1660 69518 1669
rect 69210 1658 69216 1660
rect 69272 1658 69296 1660
rect 69352 1658 69376 1660
rect 69432 1658 69456 1660
rect 69512 1658 69518 1660
rect 69272 1606 69274 1658
rect 69454 1606 69456 1658
rect 69210 1604 69216 1606
rect 69272 1604 69296 1606
rect 69352 1604 69376 1606
rect 69432 1604 69456 1606
rect 69512 1604 69518 1606
rect 69210 1595 69518 1604
rect 70810 1660 71118 1669
rect 70810 1658 70816 1660
rect 70872 1658 70896 1660
rect 70952 1658 70976 1660
rect 71032 1658 71056 1660
rect 71112 1658 71118 1660
rect 70872 1606 70874 1658
rect 71054 1606 71056 1658
rect 70810 1604 70816 1606
rect 70872 1604 70896 1606
rect 70952 1604 70976 1606
rect 71032 1604 71056 1606
rect 71112 1604 71118 1606
rect 70810 1595 71118 1604
rect 72410 1660 72718 1669
rect 72410 1658 72416 1660
rect 72472 1658 72496 1660
rect 72552 1658 72576 1660
rect 72632 1658 72656 1660
rect 72712 1658 72718 1660
rect 72472 1606 72474 1658
rect 72654 1606 72656 1658
rect 72410 1604 72416 1606
rect 72472 1604 72496 1606
rect 72552 1604 72576 1606
rect 72632 1604 72656 1606
rect 72712 1604 72718 1606
rect 72410 1595 72718 1604
rect 74010 1660 74318 1669
rect 74010 1658 74016 1660
rect 74072 1658 74096 1660
rect 74152 1658 74176 1660
rect 74232 1658 74256 1660
rect 74312 1658 74318 1660
rect 74072 1606 74074 1658
rect 74254 1606 74256 1658
rect 74010 1604 74016 1606
rect 74072 1604 74096 1606
rect 74152 1604 74176 1606
rect 74232 1604 74256 1606
rect 74312 1604 74318 1606
rect 74010 1595 74318 1604
rect 75610 1660 75918 1669
rect 75610 1658 75616 1660
rect 75672 1658 75696 1660
rect 75752 1658 75776 1660
rect 75832 1658 75856 1660
rect 75912 1658 75918 1660
rect 75672 1606 75674 1658
rect 75854 1606 75856 1658
rect 75610 1604 75616 1606
rect 75672 1604 75696 1606
rect 75752 1604 75776 1606
rect 75832 1604 75856 1606
rect 75912 1604 75918 1606
rect 75610 1595 75918 1604
rect 77210 1660 77518 1669
rect 77210 1658 77216 1660
rect 77272 1658 77296 1660
rect 77352 1658 77376 1660
rect 77432 1658 77456 1660
rect 77512 1658 77518 1660
rect 77272 1606 77274 1658
rect 77454 1606 77456 1658
rect 77210 1604 77216 1606
rect 77272 1604 77296 1606
rect 77352 1604 77376 1606
rect 77432 1604 77456 1606
rect 77512 1604 77518 1606
rect 77210 1595 77518 1604
rect 78810 1660 79118 1669
rect 78810 1658 78816 1660
rect 78872 1658 78896 1660
rect 78952 1658 78976 1660
rect 79032 1658 79056 1660
rect 79112 1658 79118 1660
rect 78872 1606 78874 1658
rect 79054 1606 79056 1658
rect 78810 1604 78816 1606
rect 78872 1604 78896 1606
rect 78952 1604 78976 1606
rect 79032 1604 79056 1606
rect 79112 1604 79118 1606
rect 78810 1595 79118 1604
rect 80410 1660 80718 1669
rect 80410 1658 80416 1660
rect 80472 1658 80496 1660
rect 80552 1658 80576 1660
rect 80632 1658 80656 1660
rect 80712 1658 80718 1660
rect 80472 1606 80474 1658
rect 80654 1606 80656 1658
rect 80410 1604 80416 1606
rect 80472 1604 80496 1606
rect 80552 1604 80576 1606
rect 80632 1604 80656 1606
rect 80712 1604 80718 1606
rect 80410 1595 80718 1604
rect 82010 1660 82318 1669
rect 82010 1658 82016 1660
rect 82072 1658 82096 1660
rect 82152 1658 82176 1660
rect 82232 1658 82256 1660
rect 82312 1658 82318 1660
rect 82072 1606 82074 1658
rect 82254 1606 82256 1658
rect 82010 1604 82016 1606
rect 82072 1604 82096 1606
rect 82152 1604 82176 1606
rect 82232 1604 82256 1606
rect 82312 1604 82318 1606
rect 82010 1595 82318 1604
rect 83610 1660 83918 1669
rect 83610 1658 83616 1660
rect 83672 1658 83696 1660
rect 83752 1658 83776 1660
rect 83832 1658 83856 1660
rect 83912 1658 83918 1660
rect 83672 1606 83674 1658
rect 83854 1606 83856 1658
rect 83610 1604 83616 1606
rect 83672 1604 83696 1606
rect 83752 1604 83776 1606
rect 83832 1604 83856 1606
rect 83912 1604 83918 1606
rect 83610 1595 83918 1604
rect 85210 1660 85518 1669
rect 85210 1658 85216 1660
rect 85272 1658 85296 1660
rect 85352 1658 85376 1660
rect 85432 1658 85456 1660
rect 85512 1658 85518 1660
rect 85272 1606 85274 1658
rect 85454 1606 85456 1658
rect 85210 1604 85216 1606
rect 85272 1604 85296 1606
rect 85352 1604 85376 1606
rect 85432 1604 85456 1606
rect 85512 1604 85518 1606
rect 85210 1595 85518 1604
rect 86810 1660 87118 1669
rect 86810 1658 86816 1660
rect 86872 1658 86896 1660
rect 86952 1658 86976 1660
rect 87032 1658 87056 1660
rect 87112 1658 87118 1660
rect 86872 1606 86874 1658
rect 87054 1606 87056 1658
rect 86810 1604 86816 1606
rect 86872 1604 86896 1606
rect 86952 1604 86976 1606
rect 87032 1604 87056 1606
rect 87112 1604 87118 1606
rect 86810 1595 87118 1604
rect 88410 1660 88718 1669
rect 88410 1658 88416 1660
rect 88472 1658 88496 1660
rect 88552 1658 88576 1660
rect 88632 1658 88656 1660
rect 88712 1658 88718 1660
rect 88472 1606 88474 1658
rect 88654 1606 88656 1658
rect 88410 1604 88416 1606
rect 88472 1604 88496 1606
rect 88552 1604 88576 1606
rect 88632 1604 88656 1606
rect 88712 1604 88718 1606
rect 88410 1595 88718 1604
rect 90010 1660 90318 1669
rect 90010 1658 90016 1660
rect 90072 1658 90096 1660
rect 90152 1658 90176 1660
rect 90232 1658 90256 1660
rect 90312 1658 90318 1660
rect 90072 1606 90074 1658
rect 90254 1606 90256 1658
rect 90010 1604 90016 1606
rect 90072 1604 90096 1606
rect 90152 1604 90176 1606
rect 90232 1604 90256 1606
rect 90312 1604 90318 1606
rect 90010 1595 90318 1604
rect 91610 1660 91918 1669
rect 91610 1658 91616 1660
rect 91672 1658 91696 1660
rect 91752 1658 91776 1660
rect 91832 1658 91856 1660
rect 91912 1658 91918 1660
rect 91672 1606 91674 1658
rect 91854 1606 91856 1658
rect 91610 1604 91616 1606
rect 91672 1604 91696 1606
rect 91752 1604 91776 1606
rect 91832 1604 91856 1606
rect 91912 1604 91918 1606
rect 91610 1595 91918 1604
rect 93210 1660 93518 1669
rect 93210 1658 93216 1660
rect 93272 1658 93296 1660
rect 93352 1658 93376 1660
rect 93432 1658 93456 1660
rect 93512 1658 93518 1660
rect 93272 1606 93274 1658
rect 93454 1606 93456 1658
rect 93210 1604 93216 1606
rect 93272 1604 93296 1606
rect 93352 1604 93376 1606
rect 93432 1604 93456 1606
rect 93512 1604 93518 1606
rect 93210 1595 93518 1604
rect 94810 1660 95118 1669
rect 94810 1658 94816 1660
rect 94872 1658 94896 1660
rect 94952 1658 94976 1660
rect 95032 1658 95056 1660
rect 95112 1658 95118 1660
rect 94872 1606 94874 1658
rect 95054 1606 95056 1658
rect 94810 1604 94816 1606
rect 94872 1604 94896 1606
rect 94952 1604 94976 1606
rect 95032 1604 95056 1606
rect 95112 1604 95118 1606
rect 94810 1595 95118 1604
rect 96410 1660 96718 1669
rect 96410 1658 96416 1660
rect 96472 1658 96496 1660
rect 96552 1658 96576 1660
rect 96632 1658 96656 1660
rect 96712 1658 96718 1660
rect 96472 1606 96474 1658
rect 96654 1606 96656 1658
rect 96410 1604 96416 1606
rect 96472 1604 96496 1606
rect 96552 1604 96576 1606
rect 96632 1604 96656 1606
rect 96712 1604 96718 1606
rect 96410 1595 96718 1604
rect 98010 1660 98318 1669
rect 98010 1658 98016 1660
rect 98072 1658 98096 1660
rect 98152 1658 98176 1660
rect 98232 1658 98256 1660
rect 98312 1658 98318 1660
rect 98072 1606 98074 1658
rect 98254 1606 98256 1658
rect 98010 1604 98016 1606
rect 98072 1604 98096 1606
rect 98152 1604 98176 1606
rect 98232 1604 98256 1606
rect 98312 1604 98318 1606
rect 98010 1595 98318 1604
rect 99610 1660 99918 1669
rect 99610 1658 99616 1660
rect 99672 1658 99696 1660
rect 99752 1658 99776 1660
rect 99832 1658 99856 1660
rect 99912 1658 99918 1660
rect 99672 1606 99674 1658
rect 99854 1606 99856 1658
rect 99610 1604 99616 1606
rect 99672 1604 99696 1606
rect 99752 1604 99776 1606
rect 99832 1604 99856 1606
rect 99912 1604 99918 1606
rect 99610 1595 99918 1604
rect 101210 1660 101518 1669
rect 101210 1658 101216 1660
rect 101272 1658 101296 1660
rect 101352 1658 101376 1660
rect 101432 1658 101456 1660
rect 101512 1658 101518 1660
rect 101272 1606 101274 1658
rect 101454 1606 101456 1658
rect 101210 1604 101216 1606
rect 101272 1604 101296 1606
rect 101352 1604 101376 1606
rect 101432 1604 101456 1606
rect 101512 1604 101518 1606
rect 101210 1595 101518 1604
rect 102810 1660 103118 1669
rect 102810 1658 102816 1660
rect 102872 1658 102896 1660
rect 102952 1658 102976 1660
rect 103032 1658 103056 1660
rect 103112 1658 103118 1660
rect 102872 1606 102874 1658
rect 103054 1606 103056 1658
rect 102810 1604 102816 1606
rect 102872 1604 102896 1606
rect 102952 1604 102976 1606
rect 103032 1604 103056 1606
rect 103112 1604 103118 1606
rect 102810 1595 103118 1604
rect 104410 1660 104718 1669
rect 104410 1658 104416 1660
rect 104472 1658 104496 1660
rect 104552 1658 104576 1660
rect 104632 1658 104656 1660
rect 104712 1658 104718 1660
rect 104472 1606 104474 1658
rect 104654 1606 104656 1658
rect 104410 1604 104416 1606
rect 104472 1604 104496 1606
rect 104552 1604 104576 1606
rect 104632 1604 104656 1606
rect 104712 1604 104718 1606
rect 104410 1595 104718 1604
rect 106010 1660 106318 1669
rect 106010 1658 106016 1660
rect 106072 1658 106096 1660
rect 106152 1658 106176 1660
rect 106232 1658 106256 1660
rect 106312 1658 106318 1660
rect 106072 1606 106074 1658
rect 106254 1606 106256 1658
rect 106010 1604 106016 1606
rect 106072 1604 106096 1606
rect 106152 1604 106176 1606
rect 106232 1604 106256 1606
rect 106312 1604 106318 1606
rect 106010 1595 106318 1604
rect 107610 1660 107918 1669
rect 107610 1658 107616 1660
rect 107672 1658 107696 1660
rect 107752 1658 107776 1660
rect 107832 1658 107856 1660
rect 107912 1658 107918 1660
rect 107672 1606 107674 1658
rect 107854 1606 107856 1658
rect 107610 1604 107616 1606
rect 107672 1604 107696 1606
rect 107752 1604 107776 1606
rect 107832 1604 107856 1606
rect 107912 1604 107918 1606
rect 107610 1595 107918 1604
rect 56598 1320 56654 1329
rect 56598 1255 56654 1264
rect 57978 1320 58034 1329
rect 57978 1255 58034 1264
rect 59358 1320 59414 1329
rect 59358 1255 59360 1264
rect 55750 1116 56058 1125
rect 55750 1114 55756 1116
rect 55812 1114 55836 1116
rect 55892 1114 55916 1116
rect 55972 1114 55996 1116
rect 56052 1114 56058 1116
rect 55812 1062 55814 1114
rect 55994 1062 55996 1114
rect 55750 1060 55756 1062
rect 55812 1060 55836 1062
rect 55892 1060 55916 1062
rect 55972 1060 55996 1062
rect 56052 1060 56058 1062
rect 55750 1051 56058 1060
rect 54864 870 54984 898
rect 56612 882 56640 1255
rect 57350 1116 57658 1125
rect 57350 1114 57356 1116
rect 57412 1114 57436 1116
rect 57492 1114 57516 1116
rect 57572 1114 57596 1116
rect 57652 1114 57658 1116
rect 57412 1062 57414 1114
rect 57594 1062 57596 1114
rect 57350 1060 57356 1062
rect 57412 1060 57436 1062
rect 57492 1060 57516 1062
rect 57572 1060 57596 1062
rect 57652 1060 57658 1062
rect 57350 1051 57658 1060
rect 54864 762 54892 870
rect 54588 734 54892 762
rect 37740 672 37792 678
rect 37740 614 37792 620
rect 37372 604 37424 610
rect 37372 546 37424 552
rect 33138 303 33194 312
rect 33232 332 33284 338
rect 33232 274 33284 280
rect 34520 332 34572 338
rect 34520 274 34572 280
rect 24400 264 24452 270
rect 24400 206 24452 212
rect 30564 264 30616 270
rect 30564 206 30616 212
rect 22928 128 22980 134
rect 22928 70 22980 76
rect 54956 0 54984 870
rect 56600 876 56652 882
rect 56600 818 56652 824
rect 57992 270 58020 1255
rect 59412 1255 59414 1264
rect 60922 1320 60978 1329
rect 60922 1255 60978 1264
rect 62486 1320 62542 1329
rect 62486 1255 62542 1264
rect 63498 1320 63554 1329
rect 63498 1255 63554 1264
rect 64878 1320 64934 1329
rect 64878 1255 64934 1264
rect 65154 1320 65210 1329
rect 65154 1255 65210 1264
rect 66258 1320 66314 1329
rect 66258 1255 66314 1264
rect 67638 1320 67694 1329
rect 67638 1255 67694 1264
rect 69018 1320 69074 1329
rect 69018 1255 69074 1264
rect 59360 1226 59412 1232
rect 58950 1116 59258 1125
rect 58950 1114 58956 1116
rect 59012 1114 59036 1116
rect 59092 1114 59116 1116
rect 59172 1114 59196 1116
rect 59252 1114 59258 1116
rect 59012 1062 59014 1114
rect 59194 1062 59196 1114
rect 58950 1060 58956 1062
rect 59012 1060 59036 1062
rect 59092 1060 59116 1062
rect 59172 1060 59196 1062
rect 59252 1060 59258 1062
rect 58950 1051 59258 1060
rect 60550 1116 60858 1125
rect 60550 1114 60556 1116
rect 60612 1114 60636 1116
rect 60692 1114 60716 1116
rect 60772 1114 60796 1116
rect 60852 1114 60858 1116
rect 60612 1062 60614 1114
rect 60794 1062 60796 1114
rect 60550 1060 60556 1062
rect 60612 1060 60636 1062
rect 60692 1060 60716 1062
rect 60772 1060 60796 1062
rect 60852 1060 60858 1062
rect 60550 1051 60858 1060
rect 60936 746 60964 1255
rect 62150 1116 62458 1125
rect 62150 1114 62156 1116
rect 62212 1114 62236 1116
rect 62292 1114 62316 1116
rect 62372 1114 62396 1116
rect 62452 1114 62458 1116
rect 62212 1062 62214 1114
rect 62394 1062 62396 1114
rect 62150 1060 62156 1062
rect 62212 1060 62236 1062
rect 62292 1060 62316 1062
rect 62372 1060 62396 1062
rect 62452 1060 62458 1062
rect 62150 1051 62458 1060
rect 60924 740 60976 746
rect 60924 682 60976 688
rect 62500 542 62528 1255
rect 62488 536 62540 542
rect 62488 478 62540 484
rect 63512 406 63540 1255
rect 63750 1116 64058 1125
rect 63750 1114 63756 1116
rect 63812 1114 63836 1116
rect 63892 1114 63916 1116
rect 63972 1114 63996 1116
rect 64052 1114 64058 1116
rect 63812 1062 63814 1114
rect 63994 1062 63996 1114
rect 63750 1060 63756 1062
rect 63812 1060 63836 1062
rect 63892 1060 63916 1062
rect 63972 1060 63996 1062
rect 64052 1060 64058 1062
rect 63750 1051 64058 1060
rect 64892 814 64920 1255
rect 65168 1018 65196 1255
rect 65350 1116 65658 1125
rect 65350 1114 65356 1116
rect 65412 1114 65436 1116
rect 65492 1114 65516 1116
rect 65572 1114 65596 1116
rect 65652 1114 65658 1116
rect 65412 1062 65414 1114
rect 65594 1062 65596 1114
rect 65350 1060 65356 1062
rect 65412 1060 65436 1062
rect 65492 1060 65516 1062
rect 65572 1060 65596 1062
rect 65652 1060 65658 1062
rect 65350 1051 65658 1060
rect 65156 1012 65208 1018
rect 65156 954 65208 960
rect 64880 808 64932 814
rect 64880 750 64932 756
rect 66272 610 66300 1255
rect 66950 1116 67258 1125
rect 66950 1114 66956 1116
rect 67012 1114 67036 1116
rect 67092 1114 67116 1116
rect 67172 1114 67196 1116
rect 67252 1114 67258 1116
rect 67012 1062 67014 1114
rect 67194 1062 67196 1114
rect 66950 1060 66956 1062
rect 67012 1060 67036 1062
rect 67092 1060 67116 1062
rect 67172 1060 67196 1062
rect 67252 1060 67258 1062
rect 66950 1051 67258 1060
rect 67652 950 67680 1255
rect 68550 1116 68858 1125
rect 68550 1114 68556 1116
rect 68612 1114 68636 1116
rect 68692 1114 68716 1116
rect 68772 1114 68796 1116
rect 68852 1114 68858 1116
rect 68612 1062 68614 1114
rect 68794 1062 68796 1114
rect 68550 1060 68556 1062
rect 68612 1060 68636 1062
rect 68692 1060 68716 1062
rect 68772 1060 68796 1062
rect 68852 1060 68858 1062
rect 68550 1051 68858 1060
rect 67640 944 67692 950
rect 67640 886 67692 892
rect 69032 678 69060 1255
rect 70150 1116 70458 1125
rect 70150 1114 70156 1116
rect 70212 1114 70236 1116
rect 70292 1114 70316 1116
rect 70372 1114 70396 1116
rect 70452 1114 70458 1116
rect 70212 1062 70214 1114
rect 70394 1062 70396 1114
rect 70150 1060 70156 1062
rect 70212 1060 70236 1062
rect 70292 1060 70316 1062
rect 70372 1060 70396 1062
rect 70452 1060 70458 1062
rect 70150 1051 70458 1060
rect 71750 1116 72058 1125
rect 71750 1114 71756 1116
rect 71812 1114 71836 1116
rect 71892 1114 71916 1116
rect 71972 1114 71996 1116
rect 72052 1114 72058 1116
rect 71812 1062 71814 1114
rect 71994 1062 71996 1114
rect 71750 1060 71756 1062
rect 71812 1060 71836 1062
rect 71892 1060 71916 1062
rect 71972 1060 71996 1062
rect 72052 1060 72058 1062
rect 71750 1051 72058 1060
rect 73350 1116 73658 1125
rect 73350 1114 73356 1116
rect 73412 1114 73436 1116
rect 73492 1114 73516 1116
rect 73572 1114 73596 1116
rect 73652 1114 73658 1116
rect 73412 1062 73414 1114
rect 73594 1062 73596 1114
rect 73350 1060 73356 1062
rect 73412 1060 73436 1062
rect 73492 1060 73516 1062
rect 73572 1060 73596 1062
rect 73652 1060 73658 1062
rect 73350 1051 73658 1060
rect 74950 1116 75258 1125
rect 74950 1114 74956 1116
rect 75012 1114 75036 1116
rect 75092 1114 75116 1116
rect 75172 1114 75196 1116
rect 75252 1114 75258 1116
rect 75012 1062 75014 1114
rect 75194 1062 75196 1114
rect 74950 1060 74956 1062
rect 75012 1060 75036 1062
rect 75092 1060 75116 1062
rect 75172 1060 75196 1062
rect 75252 1060 75258 1062
rect 74950 1051 75258 1060
rect 76550 1116 76858 1125
rect 76550 1114 76556 1116
rect 76612 1114 76636 1116
rect 76692 1114 76716 1116
rect 76772 1114 76796 1116
rect 76852 1114 76858 1116
rect 76612 1062 76614 1114
rect 76794 1062 76796 1114
rect 76550 1060 76556 1062
rect 76612 1060 76636 1062
rect 76692 1060 76716 1062
rect 76772 1060 76796 1062
rect 76852 1060 76858 1062
rect 76550 1051 76858 1060
rect 78150 1116 78458 1125
rect 78150 1114 78156 1116
rect 78212 1114 78236 1116
rect 78292 1114 78316 1116
rect 78372 1114 78396 1116
rect 78452 1114 78458 1116
rect 78212 1062 78214 1114
rect 78394 1062 78396 1114
rect 78150 1060 78156 1062
rect 78212 1060 78236 1062
rect 78292 1060 78316 1062
rect 78372 1060 78396 1062
rect 78452 1060 78458 1062
rect 78150 1051 78458 1060
rect 79750 1116 80058 1125
rect 79750 1114 79756 1116
rect 79812 1114 79836 1116
rect 79892 1114 79916 1116
rect 79972 1114 79996 1116
rect 80052 1114 80058 1116
rect 79812 1062 79814 1114
rect 79994 1062 79996 1114
rect 79750 1060 79756 1062
rect 79812 1060 79836 1062
rect 79892 1060 79916 1062
rect 79972 1060 79996 1062
rect 80052 1060 80058 1062
rect 79750 1051 80058 1060
rect 81350 1116 81658 1125
rect 81350 1114 81356 1116
rect 81412 1114 81436 1116
rect 81492 1114 81516 1116
rect 81572 1114 81596 1116
rect 81652 1114 81658 1116
rect 81412 1062 81414 1114
rect 81594 1062 81596 1114
rect 81350 1060 81356 1062
rect 81412 1060 81436 1062
rect 81492 1060 81516 1062
rect 81572 1060 81596 1062
rect 81652 1060 81658 1062
rect 81350 1051 81658 1060
rect 82950 1116 83258 1125
rect 82950 1114 82956 1116
rect 83012 1114 83036 1116
rect 83092 1114 83116 1116
rect 83172 1114 83196 1116
rect 83252 1114 83258 1116
rect 83012 1062 83014 1114
rect 83194 1062 83196 1114
rect 82950 1060 82956 1062
rect 83012 1060 83036 1062
rect 83092 1060 83116 1062
rect 83172 1060 83196 1062
rect 83252 1060 83258 1062
rect 82950 1051 83258 1060
rect 84550 1116 84858 1125
rect 84550 1114 84556 1116
rect 84612 1114 84636 1116
rect 84692 1114 84716 1116
rect 84772 1114 84796 1116
rect 84852 1114 84858 1116
rect 84612 1062 84614 1114
rect 84794 1062 84796 1114
rect 84550 1060 84556 1062
rect 84612 1060 84636 1062
rect 84692 1060 84716 1062
rect 84772 1060 84796 1062
rect 84852 1060 84858 1062
rect 84550 1051 84858 1060
rect 86150 1116 86458 1125
rect 86150 1114 86156 1116
rect 86212 1114 86236 1116
rect 86292 1114 86316 1116
rect 86372 1114 86396 1116
rect 86452 1114 86458 1116
rect 86212 1062 86214 1114
rect 86394 1062 86396 1114
rect 86150 1060 86156 1062
rect 86212 1060 86236 1062
rect 86292 1060 86316 1062
rect 86372 1060 86396 1062
rect 86452 1060 86458 1062
rect 86150 1051 86458 1060
rect 87750 1116 88058 1125
rect 87750 1114 87756 1116
rect 87812 1114 87836 1116
rect 87892 1114 87916 1116
rect 87972 1114 87996 1116
rect 88052 1114 88058 1116
rect 87812 1062 87814 1114
rect 87994 1062 87996 1114
rect 87750 1060 87756 1062
rect 87812 1060 87836 1062
rect 87892 1060 87916 1062
rect 87972 1060 87996 1062
rect 88052 1060 88058 1062
rect 87750 1051 88058 1060
rect 89350 1116 89658 1125
rect 89350 1114 89356 1116
rect 89412 1114 89436 1116
rect 89492 1114 89516 1116
rect 89572 1114 89596 1116
rect 89652 1114 89658 1116
rect 89412 1062 89414 1114
rect 89594 1062 89596 1114
rect 89350 1060 89356 1062
rect 89412 1060 89436 1062
rect 89492 1060 89516 1062
rect 89572 1060 89596 1062
rect 89652 1060 89658 1062
rect 89350 1051 89658 1060
rect 90950 1116 91258 1125
rect 90950 1114 90956 1116
rect 91012 1114 91036 1116
rect 91092 1114 91116 1116
rect 91172 1114 91196 1116
rect 91252 1114 91258 1116
rect 91012 1062 91014 1114
rect 91194 1062 91196 1114
rect 90950 1060 90956 1062
rect 91012 1060 91036 1062
rect 91092 1060 91116 1062
rect 91172 1060 91196 1062
rect 91252 1060 91258 1062
rect 90950 1051 91258 1060
rect 92550 1116 92858 1125
rect 92550 1114 92556 1116
rect 92612 1114 92636 1116
rect 92692 1114 92716 1116
rect 92772 1114 92796 1116
rect 92852 1114 92858 1116
rect 92612 1062 92614 1114
rect 92794 1062 92796 1114
rect 92550 1060 92556 1062
rect 92612 1060 92636 1062
rect 92692 1060 92716 1062
rect 92772 1060 92796 1062
rect 92852 1060 92858 1062
rect 92550 1051 92858 1060
rect 94150 1116 94458 1125
rect 94150 1114 94156 1116
rect 94212 1114 94236 1116
rect 94292 1114 94316 1116
rect 94372 1114 94396 1116
rect 94452 1114 94458 1116
rect 94212 1062 94214 1114
rect 94394 1062 94396 1114
rect 94150 1060 94156 1062
rect 94212 1060 94236 1062
rect 94292 1060 94316 1062
rect 94372 1060 94396 1062
rect 94452 1060 94458 1062
rect 94150 1051 94458 1060
rect 95750 1116 96058 1125
rect 95750 1114 95756 1116
rect 95812 1114 95836 1116
rect 95892 1114 95916 1116
rect 95972 1114 95996 1116
rect 96052 1114 96058 1116
rect 95812 1062 95814 1114
rect 95994 1062 95996 1114
rect 95750 1060 95756 1062
rect 95812 1060 95836 1062
rect 95892 1060 95916 1062
rect 95972 1060 95996 1062
rect 96052 1060 96058 1062
rect 95750 1051 96058 1060
rect 97350 1116 97658 1125
rect 97350 1114 97356 1116
rect 97412 1114 97436 1116
rect 97492 1114 97516 1116
rect 97572 1114 97596 1116
rect 97652 1114 97658 1116
rect 97412 1062 97414 1114
rect 97594 1062 97596 1114
rect 97350 1060 97356 1062
rect 97412 1060 97436 1062
rect 97492 1060 97516 1062
rect 97572 1060 97596 1062
rect 97652 1060 97658 1062
rect 97350 1051 97658 1060
rect 98950 1116 99258 1125
rect 98950 1114 98956 1116
rect 99012 1114 99036 1116
rect 99092 1114 99116 1116
rect 99172 1114 99196 1116
rect 99252 1114 99258 1116
rect 99012 1062 99014 1114
rect 99194 1062 99196 1114
rect 98950 1060 98956 1062
rect 99012 1060 99036 1062
rect 99092 1060 99116 1062
rect 99172 1060 99196 1062
rect 99252 1060 99258 1062
rect 98950 1051 99258 1060
rect 100550 1116 100858 1125
rect 100550 1114 100556 1116
rect 100612 1114 100636 1116
rect 100692 1114 100716 1116
rect 100772 1114 100796 1116
rect 100852 1114 100858 1116
rect 100612 1062 100614 1114
rect 100794 1062 100796 1114
rect 100550 1060 100556 1062
rect 100612 1060 100636 1062
rect 100692 1060 100716 1062
rect 100772 1060 100796 1062
rect 100852 1060 100858 1062
rect 100550 1051 100858 1060
rect 102150 1116 102458 1125
rect 102150 1114 102156 1116
rect 102212 1114 102236 1116
rect 102292 1114 102316 1116
rect 102372 1114 102396 1116
rect 102452 1114 102458 1116
rect 102212 1062 102214 1114
rect 102394 1062 102396 1114
rect 102150 1060 102156 1062
rect 102212 1060 102236 1062
rect 102292 1060 102316 1062
rect 102372 1060 102396 1062
rect 102452 1060 102458 1062
rect 102150 1051 102458 1060
rect 103750 1116 104058 1125
rect 103750 1114 103756 1116
rect 103812 1114 103836 1116
rect 103892 1114 103916 1116
rect 103972 1114 103996 1116
rect 104052 1114 104058 1116
rect 103812 1062 103814 1114
rect 103994 1062 103996 1114
rect 103750 1060 103756 1062
rect 103812 1060 103836 1062
rect 103892 1060 103916 1062
rect 103972 1060 103996 1062
rect 104052 1060 104058 1062
rect 103750 1051 104058 1060
rect 105350 1116 105658 1125
rect 105350 1114 105356 1116
rect 105412 1114 105436 1116
rect 105492 1114 105516 1116
rect 105572 1114 105596 1116
rect 105652 1114 105658 1116
rect 105412 1062 105414 1114
rect 105594 1062 105596 1114
rect 105350 1060 105356 1062
rect 105412 1060 105436 1062
rect 105492 1060 105516 1062
rect 105572 1060 105596 1062
rect 105652 1060 105658 1062
rect 105350 1051 105658 1060
rect 106950 1116 107258 1125
rect 106950 1114 106956 1116
rect 107012 1114 107036 1116
rect 107092 1114 107116 1116
rect 107172 1114 107196 1116
rect 107252 1114 107258 1116
rect 107012 1062 107014 1114
rect 107194 1062 107196 1114
rect 106950 1060 106956 1062
rect 107012 1060 107036 1062
rect 107092 1060 107116 1062
rect 107172 1060 107196 1062
rect 107252 1060 107258 1062
rect 106950 1051 107258 1060
rect 108550 1116 108858 1125
rect 108550 1114 108556 1116
rect 108612 1114 108636 1116
rect 108692 1114 108716 1116
rect 108772 1114 108796 1116
rect 108852 1114 108858 1116
rect 108612 1062 108614 1114
rect 108794 1062 108796 1114
rect 108550 1060 108556 1062
rect 108612 1060 108636 1062
rect 108692 1060 108716 1062
rect 108772 1060 108796 1062
rect 108852 1060 108858 1062
rect 108550 1051 108858 1060
rect 69020 672 69072 678
rect 69020 614 69072 620
rect 66260 604 66312 610
rect 66260 546 66312 552
rect 63500 400 63552 406
rect 63500 342 63552 348
rect 57980 264 58032 270
rect 57980 206 58032 212
<< via2 >>
rect 938 84360 994 84416
rect 938 83408 994 83464
rect 938 81504 994 81560
rect 938 80552 994 80608
rect 938 79620 994 79656
rect 938 79600 940 79620
rect 940 79600 992 79620
rect 992 79600 994 79620
rect 938 78648 994 78704
rect 938 77696 994 77752
rect 938 76744 994 76800
rect 938 74840 994 74896
rect 938 73888 994 73944
rect 938 72936 994 72992
rect 938 72004 994 72040
rect 938 71984 940 72004
rect 940 71984 992 72004
rect 992 71984 994 72004
rect 938 71032 994 71088
rect 938 69128 994 69184
rect 938 68176 994 68232
rect 938 66272 994 66328
rect 938 65320 994 65376
rect 2956 85978 3012 85980
rect 3036 85978 3092 85980
rect 3116 85978 3172 85980
rect 3196 85978 3252 85980
rect 2956 85926 3002 85978
rect 3002 85926 3012 85978
rect 3036 85926 3066 85978
rect 3066 85926 3078 85978
rect 3078 85926 3092 85978
rect 3116 85926 3130 85978
rect 3130 85926 3142 85978
rect 3142 85926 3172 85978
rect 3196 85926 3206 85978
rect 3206 85926 3252 85978
rect 2956 85924 3012 85926
rect 3036 85924 3092 85926
rect 3116 85924 3172 85926
rect 3196 85924 3252 85926
rect 2956 84890 3012 84892
rect 3036 84890 3092 84892
rect 3116 84890 3172 84892
rect 3196 84890 3252 84892
rect 2956 84838 3002 84890
rect 3002 84838 3012 84890
rect 3036 84838 3066 84890
rect 3066 84838 3078 84890
rect 3078 84838 3092 84890
rect 3116 84838 3130 84890
rect 3130 84838 3142 84890
rect 3142 84838 3172 84890
rect 3196 84838 3206 84890
rect 3206 84838 3252 84890
rect 2956 84836 3012 84838
rect 3036 84836 3092 84838
rect 3116 84836 3172 84838
rect 3196 84836 3252 84838
rect 1490 82728 1546 82784
rect 1490 75792 1546 75848
rect 1398 70352 1454 70408
rect 938 64388 994 64424
rect 938 64368 940 64388
rect 940 64368 992 64388
rect 992 64368 994 64388
rect 1122 65048 1178 65104
rect 938 62464 994 62520
rect 938 61512 994 61568
rect 938 60560 994 60616
rect 938 59608 994 59664
rect 938 58656 994 58712
rect 938 56752 994 56808
rect 938 55800 994 55856
rect 938 54848 994 54904
rect 938 53932 940 53952
rect 940 53932 992 53952
rect 992 53932 994 53952
rect 938 53896 994 53932
rect 938 52944 994 53000
rect 938 51040 994 51096
rect 1582 71884 1584 71904
rect 1584 71884 1636 71904
rect 1636 71884 1638 71904
rect 1582 71848 1638 71884
rect 1490 67496 1546 67552
rect 1582 65048 1638 65104
rect 1490 63416 1546 63472
rect 938 50124 940 50144
rect 940 50124 992 50144
rect 992 50124 994 50144
rect 938 50088 994 50124
rect 938 49136 994 49192
rect 938 47232 994 47288
rect 938 46316 940 46336
rect 940 46316 992 46336
rect 992 46316 994 46336
rect 938 46280 994 46316
rect 938 45328 994 45384
rect 938 44376 994 44432
rect 938 43424 994 43480
rect 938 42472 994 42528
rect 938 41540 994 41576
rect 938 41520 940 41540
rect 940 41520 992 41540
rect 992 41520 994 41540
rect 1030 40568 1086 40624
rect 1030 38664 1086 38720
rect 1030 37712 1086 37768
rect 1030 36760 1086 36816
rect 1582 57740 1584 57760
rect 1584 57740 1636 57760
rect 1636 57740 1638 57760
rect 1582 57704 1638 57740
rect 1582 52300 1584 52320
rect 1584 52300 1636 52320
rect 1636 52300 1638 52320
rect 1582 52264 1638 52300
rect 1582 48184 1638 48240
rect 1490 39888 1546 39944
rect 2956 83802 3012 83804
rect 3036 83802 3092 83804
rect 3116 83802 3172 83804
rect 3196 83802 3252 83804
rect 2956 83750 3002 83802
rect 3002 83750 3012 83802
rect 3036 83750 3066 83802
rect 3066 83750 3078 83802
rect 3078 83750 3092 83802
rect 3116 83750 3130 83802
rect 3130 83750 3142 83802
rect 3142 83750 3172 83802
rect 3196 83750 3206 83802
rect 3206 83750 3252 83802
rect 2956 83748 3012 83750
rect 3036 83748 3092 83750
rect 3116 83748 3172 83750
rect 3196 83748 3252 83750
rect 938 34856 994 34912
rect 938 33940 940 33960
rect 940 33940 992 33960
rect 992 33940 994 33960
rect 938 33904 994 33940
rect 938 32000 994 32056
rect 938 31048 994 31104
rect 938 30096 994 30152
rect 938 29144 994 29200
rect 938 28192 994 28248
rect 938 27240 994 27296
rect 938 26324 940 26344
rect 940 26324 992 26344
rect 992 26324 994 26344
rect 938 26288 994 26324
rect 938 25336 994 25392
rect 938 24384 994 24440
rect 938 23432 994 23488
rect 938 22480 994 22536
rect 938 21528 994 21584
rect 938 19624 994 19680
rect 938 18692 994 18728
rect 938 18672 940 18692
rect 940 18672 992 18692
rect 992 18672 994 18692
rect 938 16768 994 16824
rect 938 15852 940 15872
rect 940 15852 992 15872
rect 992 15852 994 15872
rect 938 15816 994 15852
rect 938 14864 994 14920
rect 938 13912 994 13968
rect 938 12960 994 13016
rect 938 12044 940 12064
rect 940 12044 992 12064
rect 992 12044 994 12064
rect 938 12008 994 12044
rect 938 11056 994 11112
rect 938 10104 994 10160
rect 938 9152 994 9208
rect 938 7248 994 7304
rect 938 6296 994 6352
rect 938 4428 940 4448
rect 940 4428 992 4448
rect 992 4428 994 4448
rect 938 4392 994 4428
rect 938 3440 994 3496
rect 1398 35808 1454 35864
rect 1214 2488 1270 2544
rect 2134 69284 2190 69320
rect 2134 69264 2136 69284
rect 2136 69264 2188 69284
rect 2188 69264 2190 69284
rect 2134 65048 2190 65104
rect 2956 82714 3012 82716
rect 3036 82714 3092 82716
rect 3116 82714 3172 82716
rect 3196 82714 3252 82716
rect 2956 82662 3002 82714
rect 3002 82662 3012 82714
rect 3036 82662 3066 82714
rect 3066 82662 3078 82714
rect 3078 82662 3092 82714
rect 3116 82662 3130 82714
rect 3130 82662 3142 82714
rect 3142 82662 3172 82714
rect 3196 82662 3206 82714
rect 3206 82662 3252 82714
rect 2956 82660 3012 82662
rect 3036 82660 3092 82662
rect 3116 82660 3172 82662
rect 3196 82660 3252 82662
rect 2956 81626 3012 81628
rect 3036 81626 3092 81628
rect 3116 81626 3172 81628
rect 3196 81626 3252 81628
rect 2956 81574 3002 81626
rect 3002 81574 3012 81626
rect 3036 81574 3066 81626
rect 3066 81574 3078 81626
rect 3078 81574 3092 81626
rect 3116 81574 3130 81626
rect 3130 81574 3142 81626
rect 3142 81574 3172 81626
rect 3196 81574 3206 81626
rect 3206 81574 3252 81626
rect 2956 81572 3012 81574
rect 3036 81572 3092 81574
rect 3116 81572 3172 81574
rect 3196 81572 3252 81574
rect 2956 80538 3012 80540
rect 3036 80538 3092 80540
rect 3116 80538 3172 80540
rect 3196 80538 3252 80540
rect 2956 80486 3002 80538
rect 3002 80486 3012 80538
rect 3036 80486 3066 80538
rect 3066 80486 3078 80538
rect 3078 80486 3092 80538
rect 3116 80486 3130 80538
rect 3130 80486 3142 80538
rect 3142 80486 3172 80538
rect 3196 80486 3206 80538
rect 3206 80486 3252 80538
rect 2956 80484 3012 80486
rect 3036 80484 3092 80486
rect 3116 80484 3172 80486
rect 3196 80484 3252 80486
rect 2956 79450 3012 79452
rect 3036 79450 3092 79452
rect 3116 79450 3172 79452
rect 3196 79450 3252 79452
rect 2956 79398 3002 79450
rect 3002 79398 3012 79450
rect 3036 79398 3066 79450
rect 3066 79398 3078 79450
rect 3078 79398 3092 79450
rect 3116 79398 3130 79450
rect 3130 79398 3142 79450
rect 3142 79398 3172 79450
rect 3196 79398 3206 79450
rect 3206 79398 3252 79450
rect 2956 79396 3012 79398
rect 3036 79396 3092 79398
rect 3116 79396 3172 79398
rect 3196 79396 3252 79398
rect 2956 78362 3012 78364
rect 3036 78362 3092 78364
rect 3116 78362 3172 78364
rect 3196 78362 3252 78364
rect 2956 78310 3002 78362
rect 3002 78310 3012 78362
rect 3036 78310 3066 78362
rect 3066 78310 3078 78362
rect 3078 78310 3092 78362
rect 3116 78310 3130 78362
rect 3130 78310 3142 78362
rect 3142 78310 3172 78362
rect 3196 78310 3206 78362
rect 3206 78310 3252 78362
rect 2956 78308 3012 78310
rect 3036 78308 3092 78310
rect 3116 78308 3172 78310
rect 3196 78308 3252 78310
rect 2956 77274 3012 77276
rect 3036 77274 3092 77276
rect 3116 77274 3172 77276
rect 3196 77274 3252 77276
rect 2956 77222 3002 77274
rect 3002 77222 3012 77274
rect 3036 77222 3066 77274
rect 3066 77222 3078 77274
rect 3078 77222 3092 77274
rect 3116 77222 3130 77274
rect 3130 77222 3142 77274
rect 3142 77222 3172 77274
rect 3196 77222 3206 77274
rect 3206 77222 3252 77274
rect 2956 77220 3012 77222
rect 3036 77220 3092 77222
rect 3116 77220 3172 77222
rect 3196 77220 3252 77222
rect 2956 76186 3012 76188
rect 3036 76186 3092 76188
rect 3116 76186 3172 76188
rect 3196 76186 3252 76188
rect 2956 76134 3002 76186
rect 3002 76134 3012 76186
rect 3036 76134 3066 76186
rect 3066 76134 3078 76186
rect 3078 76134 3092 76186
rect 3116 76134 3130 76186
rect 3130 76134 3142 76186
rect 3142 76134 3172 76186
rect 3196 76134 3206 76186
rect 3206 76134 3252 76186
rect 2956 76132 3012 76134
rect 3036 76132 3092 76134
rect 3116 76132 3172 76134
rect 3196 76132 3252 76134
rect 2956 75098 3012 75100
rect 3036 75098 3092 75100
rect 3116 75098 3172 75100
rect 3196 75098 3252 75100
rect 2956 75046 3002 75098
rect 3002 75046 3012 75098
rect 3036 75046 3066 75098
rect 3066 75046 3078 75098
rect 3078 75046 3092 75098
rect 3116 75046 3130 75098
rect 3130 75046 3142 75098
rect 3142 75046 3172 75098
rect 3196 75046 3206 75098
rect 3206 75046 3252 75098
rect 2956 75044 3012 75046
rect 3036 75044 3092 75046
rect 3116 75044 3172 75046
rect 3196 75044 3252 75046
rect 2956 74010 3012 74012
rect 3036 74010 3092 74012
rect 3116 74010 3172 74012
rect 3196 74010 3252 74012
rect 2956 73958 3002 74010
rect 3002 73958 3012 74010
rect 3036 73958 3066 74010
rect 3066 73958 3078 74010
rect 3078 73958 3092 74010
rect 3116 73958 3130 74010
rect 3130 73958 3142 74010
rect 3142 73958 3172 74010
rect 3196 73958 3206 74010
rect 3206 73958 3252 74010
rect 2956 73956 3012 73958
rect 3036 73956 3092 73958
rect 3116 73956 3172 73958
rect 3196 73956 3252 73958
rect 2956 72922 3012 72924
rect 3036 72922 3092 72924
rect 3116 72922 3172 72924
rect 3196 72922 3252 72924
rect 2956 72870 3002 72922
rect 3002 72870 3012 72922
rect 3036 72870 3066 72922
rect 3066 72870 3078 72922
rect 3078 72870 3092 72922
rect 3116 72870 3130 72922
rect 3130 72870 3142 72922
rect 3142 72870 3172 72922
rect 3196 72870 3206 72922
rect 3206 72870 3252 72922
rect 2956 72868 3012 72870
rect 3036 72868 3092 72870
rect 3116 72868 3172 72870
rect 3196 72868 3252 72870
rect 2956 71834 3012 71836
rect 3036 71834 3092 71836
rect 3116 71834 3172 71836
rect 3196 71834 3252 71836
rect 2956 71782 3002 71834
rect 3002 71782 3012 71834
rect 3036 71782 3066 71834
rect 3066 71782 3078 71834
rect 3078 71782 3092 71834
rect 3116 71782 3130 71834
rect 3130 71782 3142 71834
rect 3142 71782 3172 71834
rect 3196 71782 3206 71834
rect 3206 71782 3252 71834
rect 2956 71780 3012 71782
rect 3036 71780 3092 71782
rect 3116 71780 3172 71782
rect 3196 71780 3252 71782
rect 2870 71440 2926 71496
rect 2686 69944 2742 70000
rect 2594 69808 2650 69864
rect 2778 68176 2834 68232
rect 2956 70746 3012 70748
rect 3036 70746 3092 70748
rect 3116 70746 3172 70748
rect 3196 70746 3252 70748
rect 2956 70694 3002 70746
rect 3002 70694 3012 70746
rect 3036 70694 3066 70746
rect 3066 70694 3078 70746
rect 3078 70694 3092 70746
rect 3116 70694 3130 70746
rect 3130 70694 3142 70746
rect 3142 70694 3172 70746
rect 3196 70694 3206 70746
rect 3206 70694 3252 70746
rect 2956 70692 3012 70694
rect 3036 70692 3092 70694
rect 3116 70692 3172 70694
rect 3196 70692 3252 70694
rect 2956 69658 3012 69660
rect 3036 69658 3092 69660
rect 3116 69658 3172 69660
rect 3196 69658 3252 69660
rect 2956 69606 3002 69658
rect 3002 69606 3012 69658
rect 3036 69606 3066 69658
rect 3066 69606 3078 69658
rect 3078 69606 3092 69658
rect 3116 69606 3130 69658
rect 3130 69606 3142 69658
rect 3142 69606 3172 69658
rect 3196 69606 3206 69658
rect 3206 69606 3252 69658
rect 2956 69604 3012 69606
rect 3036 69604 3092 69606
rect 3116 69604 3172 69606
rect 3196 69604 3252 69606
rect 2956 68570 3012 68572
rect 3036 68570 3092 68572
rect 3116 68570 3172 68572
rect 3196 68570 3252 68572
rect 2956 68518 3002 68570
rect 3002 68518 3012 68570
rect 3036 68518 3066 68570
rect 3066 68518 3078 68570
rect 3078 68518 3092 68570
rect 3116 68518 3130 68570
rect 3130 68518 3142 68570
rect 3142 68518 3172 68570
rect 3196 68518 3206 68570
rect 3206 68518 3252 68570
rect 2956 68516 3012 68518
rect 3036 68516 3092 68518
rect 3116 68516 3172 68518
rect 3196 68516 3252 68518
rect 2956 67482 3012 67484
rect 3036 67482 3092 67484
rect 3116 67482 3172 67484
rect 3196 67482 3252 67484
rect 2956 67430 3002 67482
rect 3002 67430 3012 67482
rect 3036 67430 3066 67482
rect 3066 67430 3078 67482
rect 3078 67430 3092 67482
rect 3116 67430 3130 67482
rect 3130 67430 3142 67482
rect 3142 67430 3172 67482
rect 3196 67430 3206 67482
rect 3206 67430 3252 67482
rect 2956 67428 3012 67430
rect 3036 67428 3092 67430
rect 3116 67428 3172 67430
rect 3196 67428 3252 67430
rect 2956 66394 3012 66396
rect 3036 66394 3092 66396
rect 3116 66394 3172 66396
rect 3196 66394 3252 66396
rect 2956 66342 3002 66394
rect 3002 66342 3012 66394
rect 3036 66342 3066 66394
rect 3066 66342 3078 66394
rect 3078 66342 3092 66394
rect 3116 66342 3130 66394
rect 3130 66342 3142 66394
rect 3142 66342 3172 66394
rect 3196 66342 3206 66394
rect 3206 66342 3252 66394
rect 2956 66340 3012 66342
rect 3036 66340 3092 66342
rect 3116 66340 3172 66342
rect 3196 66340 3252 66342
rect 2778 65728 2834 65784
rect 2778 65320 2834 65376
rect 2956 65306 3012 65308
rect 3036 65306 3092 65308
rect 3116 65306 3172 65308
rect 3196 65306 3252 65308
rect 2956 65254 3002 65306
rect 3002 65254 3012 65306
rect 3036 65254 3066 65306
rect 3066 65254 3078 65306
rect 3078 65254 3092 65306
rect 3116 65254 3130 65306
rect 3130 65254 3142 65306
rect 3142 65254 3172 65306
rect 3196 65254 3206 65306
rect 3206 65254 3252 65306
rect 2956 65252 3012 65254
rect 3036 65252 3092 65254
rect 3116 65252 3172 65254
rect 3196 65252 3252 65254
rect 1490 33088 1546 33144
rect 1398 20576 1454 20632
rect 1582 17720 1638 17776
rect 1398 8200 1454 8256
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 2956 64218 3012 64220
rect 3036 64218 3092 64220
rect 3116 64218 3172 64220
rect 3196 64218 3252 64220
rect 2956 64166 3002 64218
rect 3002 64166 3012 64218
rect 3036 64166 3066 64218
rect 3066 64166 3078 64218
rect 3078 64166 3092 64218
rect 3116 64166 3130 64218
rect 3130 64166 3142 64218
rect 3142 64166 3172 64218
rect 3196 64166 3206 64218
rect 3206 64166 3252 64218
rect 2956 64164 3012 64166
rect 3036 64164 3092 64166
rect 3116 64164 3172 64166
rect 3196 64164 3252 64166
rect 2956 63130 3012 63132
rect 3036 63130 3092 63132
rect 3116 63130 3172 63132
rect 3196 63130 3252 63132
rect 2956 63078 3002 63130
rect 3002 63078 3012 63130
rect 3036 63078 3066 63130
rect 3066 63078 3078 63130
rect 3078 63078 3092 63130
rect 3116 63078 3130 63130
rect 3130 63078 3142 63130
rect 3142 63078 3172 63130
rect 3196 63078 3206 63130
rect 3206 63078 3252 63130
rect 2956 63076 3012 63078
rect 3036 63076 3092 63078
rect 3116 63076 3172 63078
rect 3196 63076 3252 63078
rect 2956 62042 3012 62044
rect 3036 62042 3092 62044
rect 3116 62042 3172 62044
rect 3196 62042 3252 62044
rect 2956 61990 3002 62042
rect 3002 61990 3012 62042
rect 3036 61990 3066 62042
rect 3066 61990 3078 62042
rect 3078 61990 3092 62042
rect 3116 61990 3130 62042
rect 3130 61990 3142 62042
rect 3142 61990 3172 62042
rect 3196 61990 3206 62042
rect 3206 61990 3252 62042
rect 2956 61988 3012 61990
rect 3036 61988 3092 61990
rect 3116 61988 3172 61990
rect 3196 61988 3252 61990
rect 2956 60954 3012 60956
rect 3036 60954 3092 60956
rect 3116 60954 3172 60956
rect 3196 60954 3252 60956
rect 2956 60902 3002 60954
rect 3002 60902 3012 60954
rect 3036 60902 3066 60954
rect 3066 60902 3078 60954
rect 3078 60902 3092 60954
rect 3116 60902 3130 60954
rect 3130 60902 3142 60954
rect 3142 60902 3172 60954
rect 3196 60902 3206 60954
rect 3206 60902 3252 60954
rect 2956 60900 3012 60902
rect 3036 60900 3092 60902
rect 3116 60900 3172 60902
rect 3196 60900 3252 60902
rect 2956 59866 3012 59868
rect 3036 59866 3092 59868
rect 3116 59866 3172 59868
rect 3196 59866 3252 59868
rect 2956 59814 3002 59866
rect 3002 59814 3012 59866
rect 3036 59814 3066 59866
rect 3066 59814 3078 59866
rect 3078 59814 3092 59866
rect 3116 59814 3130 59866
rect 3130 59814 3142 59866
rect 3142 59814 3172 59866
rect 3196 59814 3206 59866
rect 3206 59814 3252 59866
rect 2956 59812 3012 59814
rect 3036 59812 3092 59814
rect 3116 59812 3172 59814
rect 3196 59812 3252 59814
rect 2956 58778 3012 58780
rect 3036 58778 3092 58780
rect 3116 58778 3172 58780
rect 3196 58778 3252 58780
rect 2956 58726 3002 58778
rect 3002 58726 3012 58778
rect 3036 58726 3066 58778
rect 3066 58726 3078 58778
rect 3078 58726 3092 58778
rect 3116 58726 3130 58778
rect 3130 58726 3142 58778
rect 3142 58726 3172 58778
rect 3196 58726 3206 58778
rect 3206 58726 3252 58778
rect 2956 58724 3012 58726
rect 3036 58724 3092 58726
rect 3116 58724 3172 58726
rect 3196 58724 3252 58726
rect 2956 57690 3012 57692
rect 3036 57690 3092 57692
rect 3116 57690 3172 57692
rect 3196 57690 3252 57692
rect 2956 57638 3002 57690
rect 3002 57638 3012 57690
rect 3036 57638 3066 57690
rect 3066 57638 3078 57690
rect 3078 57638 3092 57690
rect 3116 57638 3130 57690
rect 3130 57638 3142 57690
rect 3142 57638 3172 57690
rect 3196 57638 3206 57690
rect 3206 57638 3252 57690
rect 2956 57636 3012 57638
rect 3036 57636 3092 57638
rect 3116 57636 3172 57638
rect 3196 57636 3252 57638
rect 2956 56602 3012 56604
rect 3036 56602 3092 56604
rect 3116 56602 3172 56604
rect 3196 56602 3252 56604
rect 2956 56550 3002 56602
rect 3002 56550 3012 56602
rect 3036 56550 3066 56602
rect 3066 56550 3078 56602
rect 3078 56550 3092 56602
rect 3116 56550 3130 56602
rect 3130 56550 3142 56602
rect 3142 56550 3172 56602
rect 3196 56550 3206 56602
rect 3206 56550 3252 56602
rect 2956 56548 3012 56550
rect 3036 56548 3092 56550
rect 3116 56548 3172 56550
rect 3196 56548 3252 56550
rect 2956 55514 3012 55516
rect 3036 55514 3092 55516
rect 3116 55514 3172 55516
rect 3196 55514 3252 55516
rect 2956 55462 3002 55514
rect 3002 55462 3012 55514
rect 3036 55462 3066 55514
rect 3066 55462 3078 55514
rect 3078 55462 3092 55514
rect 3116 55462 3130 55514
rect 3130 55462 3142 55514
rect 3142 55462 3172 55514
rect 3196 55462 3206 55514
rect 3206 55462 3252 55514
rect 2956 55460 3012 55462
rect 3036 55460 3092 55462
rect 3116 55460 3172 55462
rect 3196 55460 3252 55462
rect 2956 54426 3012 54428
rect 3036 54426 3092 54428
rect 3116 54426 3172 54428
rect 3196 54426 3252 54428
rect 2956 54374 3002 54426
rect 3002 54374 3012 54426
rect 3036 54374 3066 54426
rect 3066 54374 3078 54426
rect 3078 54374 3092 54426
rect 3116 54374 3130 54426
rect 3130 54374 3142 54426
rect 3142 54374 3172 54426
rect 3196 54374 3206 54426
rect 3206 54374 3252 54426
rect 2956 54372 3012 54374
rect 3036 54372 3092 54374
rect 3116 54372 3172 54374
rect 3196 54372 3252 54374
rect 2956 53338 3012 53340
rect 3036 53338 3092 53340
rect 3116 53338 3172 53340
rect 3196 53338 3252 53340
rect 2956 53286 3002 53338
rect 3002 53286 3012 53338
rect 3036 53286 3066 53338
rect 3066 53286 3078 53338
rect 3078 53286 3092 53338
rect 3116 53286 3130 53338
rect 3130 53286 3142 53338
rect 3142 53286 3172 53338
rect 3196 53286 3206 53338
rect 3206 53286 3252 53338
rect 2956 53284 3012 53286
rect 3036 53284 3092 53286
rect 3116 53284 3172 53286
rect 3196 53284 3252 53286
rect 2956 52250 3012 52252
rect 3036 52250 3092 52252
rect 3116 52250 3172 52252
rect 3196 52250 3252 52252
rect 2956 52198 3002 52250
rect 3002 52198 3012 52250
rect 3036 52198 3066 52250
rect 3066 52198 3078 52250
rect 3078 52198 3092 52250
rect 3116 52198 3130 52250
rect 3130 52198 3142 52250
rect 3142 52198 3172 52250
rect 3196 52198 3206 52250
rect 3206 52198 3252 52250
rect 2956 52196 3012 52198
rect 3036 52196 3092 52198
rect 3116 52196 3172 52198
rect 3196 52196 3252 52198
rect 2956 51162 3012 51164
rect 3036 51162 3092 51164
rect 3116 51162 3172 51164
rect 3196 51162 3252 51164
rect 2956 51110 3002 51162
rect 3002 51110 3012 51162
rect 3036 51110 3066 51162
rect 3066 51110 3078 51162
rect 3078 51110 3092 51162
rect 3116 51110 3130 51162
rect 3130 51110 3142 51162
rect 3142 51110 3172 51162
rect 3196 51110 3206 51162
rect 3206 51110 3252 51162
rect 2956 51108 3012 51110
rect 3036 51108 3092 51110
rect 3116 51108 3172 51110
rect 3196 51108 3252 51110
rect 2956 50074 3012 50076
rect 3036 50074 3092 50076
rect 3116 50074 3172 50076
rect 3196 50074 3252 50076
rect 2956 50022 3002 50074
rect 3002 50022 3012 50074
rect 3036 50022 3066 50074
rect 3066 50022 3078 50074
rect 3078 50022 3092 50074
rect 3116 50022 3130 50074
rect 3130 50022 3142 50074
rect 3142 50022 3172 50074
rect 3196 50022 3206 50074
rect 3206 50022 3252 50074
rect 2956 50020 3012 50022
rect 3036 50020 3092 50022
rect 3116 50020 3172 50022
rect 3196 50020 3252 50022
rect 2956 48986 3012 48988
rect 3036 48986 3092 48988
rect 3116 48986 3172 48988
rect 3196 48986 3252 48988
rect 2956 48934 3002 48986
rect 3002 48934 3012 48986
rect 3036 48934 3066 48986
rect 3066 48934 3078 48986
rect 3078 48934 3092 48986
rect 3116 48934 3130 48986
rect 3130 48934 3142 48986
rect 3142 48934 3172 48986
rect 3196 48934 3206 48986
rect 3206 48934 3252 48986
rect 2956 48932 3012 48934
rect 3036 48932 3092 48934
rect 3116 48932 3172 48934
rect 3196 48932 3252 48934
rect 2956 47898 3012 47900
rect 3036 47898 3092 47900
rect 3116 47898 3172 47900
rect 3196 47898 3252 47900
rect 2956 47846 3002 47898
rect 3002 47846 3012 47898
rect 3036 47846 3066 47898
rect 3066 47846 3078 47898
rect 3078 47846 3092 47898
rect 3116 47846 3130 47898
rect 3130 47846 3142 47898
rect 3142 47846 3172 47898
rect 3196 47846 3206 47898
rect 3206 47846 3252 47898
rect 2956 47844 3012 47846
rect 3036 47844 3092 47846
rect 3116 47844 3172 47846
rect 3196 47844 3252 47846
rect 2956 46810 3012 46812
rect 3036 46810 3092 46812
rect 3116 46810 3172 46812
rect 3196 46810 3252 46812
rect 2956 46758 3002 46810
rect 3002 46758 3012 46810
rect 3036 46758 3066 46810
rect 3066 46758 3078 46810
rect 3078 46758 3092 46810
rect 3116 46758 3130 46810
rect 3130 46758 3142 46810
rect 3142 46758 3172 46810
rect 3196 46758 3206 46810
rect 3206 46758 3252 46810
rect 2956 46756 3012 46758
rect 3036 46756 3092 46758
rect 3116 46756 3172 46758
rect 3196 46756 3252 46758
rect 2956 45722 3012 45724
rect 3036 45722 3092 45724
rect 3116 45722 3172 45724
rect 3196 45722 3252 45724
rect 2956 45670 3002 45722
rect 3002 45670 3012 45722
rect 3036 45670 3066 45722
rect 3066 45670 3078 45722
rect 3078 45670 3092 45722
rect 3116 45670 3130 45722
rect 3130 45670 3142 45722
rect 3142 45670 3172 45722
rect 3196 45670 3206 45722
rect 3206 45670 3252 45722
rect 2956 45668 3012 45670
rect 3036 45668 3092 45670
rect 3116 45668 3172 45670
rect 3196 45668 3252 45670
rect 2956 44634 3012 44636
rect 3036 44634 3092 44636
rect 3116 44634 3172 44636
rect 3196 44634 3252 44636
rect 2956 44582 3002 44634
rect 3002 44582 3012 44634
rect 3036 44582 3066 44634
rect 3066 44582 3078 44634
rect 3078 44582 3092 44634
rect 3116 44582 3130 44634
rect 3130 44582 3142 44634
rect 3142 44582 3172 44634
rect 3196 44582 3206 44634
rect 3206 44582 3252 44634
rect 2956 44580 3012 44582
rect 3036 44580 3092 44582
rect 3116 44580 3172 44582
rect 3196 44580 3252 44582
rect 2956 43546 3012 43548
rect 3036 43546 3092 43548
rect 3116 43546 3172 43548
rect 3196 43546 3252 43548
rect 2956 43494 3002 43546
rect 3002 43494 3012 43546
rect 3036 43494 3066 43546
rect 3066 43494 3078 43546
rect 3078 43494 3092 43546
rect 3116 43494 3130 43546
rect 3130 43494 3142 43546
rect 3142 43494 3172 43546
rect 3196 43494 3206 43546
rect 3206 43494 3252 43546
rect 2956 43492 3012 43494
rect 3036 43492 3092 43494
rect 3116 43492 3172 43494
rect 3196 43492 3252 43494
rect 2956 42458 3012 42460
rect 3036 42458 3092 42460
rect 3116 42458 3172 42460
rect 3196 42458 3252 42460
rect 2956 42406 3002 42458
rect 3002 42406 3012 42458
rect 3036 42406 3066 42458
rect 3066 42406 3078 42458
rect 3078 42406 3092 42458
rect 3116 42406 3130 42458
rect 3130 42406 3142 42458
rect 3142 42406 3172 42458
rect 3196 42406 3206 42458
rect 3206 42406 3252 42458
rect 2956 42404 3012 42406
rect 3036 42404 3092 42406
rect 3116 42404 3172 42406
rect 3196 42404 3252 42406
rect 2956 41370 3012 41372
rect 3036 41370 3092 41372
rect 3116 41370 3172 41372
rect 3196 41370 3252 41372
rect 2956 41318 3002 41370
rect 3002 41318 3012 41370
rect 3036 41318 3066 41370
rect 3066 41318 3078 41370
rect 3078 41318 3092 41370
rect 3116 41318 3130 41370
rect 3130 41318 3142 41370
rect 3142 41318 3172 41370
rect 3196 41318 3206 41370
rect 3206 41318 3252 41370
rect 2956 41316 3012 41318
rect 3036 41316 3092 41318
rect 3116 41316 3172 41318
rect 3196 41316 3252 41318
rect 2956 40282 3012 40284
rect 3036 40282 3092 40284
rect 3116 40282 3172 40284
rect 3196 40282 3252 40284
rect 2956 40230 3002 40282
rect 3002 40230 3012 40282
rect 3036 40230 3066 40282
rect 3066 40230 3078 40282
rect 3078 40230 3092 40282
rect 3116 40230 3130 40282
rect 3130 40230 3142 40282
rect 3142 40230 3172 40282
rect 3196 40230 3206 40282
rect 3206 40230 3252 40282
rect 2956 40228 3012 40230
rect 3036 40228 3092 40230
rect 3116 40228 3172 40230
rect 3196 40228 3252 40230
rect 2956 39194 3012 39196
rect 3036 39194 3092 39196
rect 3116 39194 3172 39196
rect 3196 39194 3252 39196
rect 2956 39142 3002 39194
rect 3002 39142 3012 39194
rect 3036 39142 3066 39194
rect 3066 39142 3078 39194
rect 3078 39142 3092 39194
rect 3116 39142 3130 39194
rect 3130 39142 3142 39194
rect 3142 39142 3172 39194
rect 3196 39142 3206 39194
rect 3206 39142 3252 39194
rect 2956 39140 3012 39142
rect 3036 39140 3092 39142
rect 3116 39140 3172 39142
rect 3196 39140 3252 39142
rect 2956 38106 3012 38108
rect 3036 38106 3092 38108
rect 3116 38106 3172 38108
rect 3196 38106 3252 38108
rect 2956 38054 3002 38106
rect 3002 38054 3012 38106
rect 3036 38054 3066 38106
rect 3066 38054 3078 38106
rect 3078 38054 3092 38106
rect 3116 38054 3130 38106
rect 3130 38054 3142 38106
rect 3142 38054 3172 38106
rect 3196 38054 3206 38106
rect 3206 38054 3252 38106
rect 2956 38052 3012 38054
rect 3036 38052 3092 38054
rect 3116 38052 3172 38054
rect 3196 38052 3252 38054
rect 2956 37018 3012 37020
rect 3036 37018 3092 37020
rect 3116 37018 3172 37020
rect 3196 37018 3252 37020
rect 2956 36966 3002 37018
rect 3002 36966 3012 37018
rect 3036 36966 3066 37018
rect 3066 36966 3078 37018
rect 3078 36966 3092 37018
rect 3116 36966 3130 37018
rect 3130 36966 3142 37018
rect 3142 36966 3172 37018
rect 3196 36966 3206 37018
rect 3206 36966 3252 37018
rect 2956 36964 3012 36966
rect 3036 36964 3092 36966
rect 3116 36964 3172 36966
rect 3196 36964 3252 36966
rect 2956 35930 3012 35932
rect 3036 35930 3092 35932
rect 3116 35930 3172 35932
rect 3196 35930 3252 35932
rect 2956 35878 3002 35930
rect 3002 35878 3012 35930
rect 3036 35878 3066 35930
rect 3066 35878 3078 35930
rect 3078 35878 3092 35930
rect 3116 35878 3130 35930
rect 3130 35878 3142 35930
rect 3142 35878 3172 35930
rect 3196 35878 3206 35930
rect 3206 35878 3252 35930
rect 2956 35876 3012 35878
rect 3036 35876 3092 35878
rect 3116 35876 3172 35878
rect 3196 35876 3252 35878
rect 2956 34842 3012 34844
rect 3036 34842 3092 34844
rect 3116 34842 3172 34844
rect 3196 34842 3252 34844
rect 2956 34790 3002 34842
rect 3002 34790 3012 34842
rect 3036 34790 3066 34842
rect 3066 34790 3078 34842
rect 3078 34790 3092 34842
rect 3116 34790 3130 34842
rect 3130 34790 3142 34842
rect 3142 34790 3172 34842
rect 3196 34790 3206 34842
rect 3206 34790 3252 34842
rect 2956 34788 3012 34790
rect 3036 34788 3092 34790
rect 3116 34788 3172 34790
rect 3196 34788 3252 34790
rect 2956 33754 3012 33756
rect 3036 33754 3092 33756
rect 3116 33754 3172 33756
rect 3196 33754 3252 33756
rect 2956 33702 3002 33754
rect 3002 33702 3012 33754
rect 3036 33702 3066 33754
rect 3066 33702 3078 33754
rect 3078 33702 3092 33754
rect 3116 33702 3130 33754
rect 3130 33702 3142 33754
rect 3142 33702 3172 33754
rect 3196 33702 3206 33754
rect 3206 33702 3252 33754
rect 2956 33700 3012 33702
rect 3036 33700 3092 33702
rect 3116 33700 3172 33702
rect 3196 33700 3252 33702
rect 2956 32666 3012 32668
rect 3036 32666 3092 32668
rect 3116 32666 3172 32668
rect 3196 32666 3252 32668
rect 2956 32614 3002 32666
rect 3002 32614 3012 32666
rect 3036 32614 3066 32666
rect 3066 32614 3078 32666
rect 3078 32614 3092 32666
rect 3116 32614 3130 32666
rect 3130 32614 3142 32666
rect 3142 32614 3172 32666
rect 3196 32614 3206 32666
rect 3206 32614 3252 32666
rect 2956 32612 3012 32614
rect 3036 32612 3092 32614
rect 3116 32612 3172 32614
rect 3196 32612 3252 32614
rect 2956 31578 3012 31580
rect 3036 31578 3092 31580
rect 3116 31578 3172 31580
rect 3196 31578 3252 31580
rect 2956 31526 3002 31578
rect 3002 31526 3012 31578
rect 3036 31526 3066 31578
rect 3066 31526 3078 31578
rect 3078 31526 3092 31578
rect 3116 31526 3130 31578
rect 3130 31526 3142 31578
rect 3142 31526 3172 31578
rect 3196 31526 3206 31578
rect 3206 31526 3252 31578
rect 2956 31524 3012 31526
rect 3036 31524 3092 31526
rect 3116 31524 3172 31526
rect 3196 31524 3252 31526
rect 2956 30490 3012 30492
rect 3036 30490 3092 30492
rect 3116 30490 3172 30492
rect 3196 30490 3252 30492
rect 2956 30438 3002 30490
rect 3002 30438 3012 30490
rect 3036 30438 3066 30490
rect 3066 30438 3078 30490
rect 3078 30438 3092 30490
rect 3116 30438 3130 30490
rect 3130 30438 3142 30490
rect 3142 30438 3172 30490
rect 3196 30438 3206 30490
rect 3206 30438 3252 30490
rect 2956 30436 3012 30438
rect 3036 30436 3092 30438
rect 3116 30436 3172 30438
rect 3196 30436 3252 30438
rect 2956 29402 3012 29404
rect 3036 29402 3092 29404
rect 3116 29402 3172 29404
rect 3196 29402 3252 29404
rect 2956 29350 3002 29402
rect 3002 29350 3012 29402
rect 3036 29350 3066 29402
rect 3066 29350 3078 29402
rect 3078 29350 3092 29402
rect 3116 29350 3130 29402
rect 3130 29350 3142 29402
rect 3142 29350 3172 29402
rect 3196 29350 3206 29402
rect 3206 29350 3252 29402
rect 2956 29348 3012 29350
rect 3036 29348 3092 29350
rect 3116 29348 3172 29350
rect 3196 29348 3252 29350
rect 2956 28314 3012 28316
rect 3036 28314 3092 28316
rect 3116 28314 3172 28316
rect 3196 28314 3252 28316
rect 2956 28262 3002 28314
rect 3002 28262 3012 28314
rect 3036 28262 3066 28314
rect 3066 28262 3078 28314
rect 3078 28262 3092 28314
rect 3116 28262 3130 28314
rect 3130 28262 3142 28314
rect 3142 28262 3172 28314
rect 3196 28262 3206 28314
rect 3206 28262 3252 28314
rect 2956 28260 3012 28262
rect 3036 28260 3092 28262
rect 3116 28260 3172 28262
rect 3196 28260 3252 28262
rect 2956 27226 3012 27228
rect 3036 27226 3092 27228
rect 3116 27226 3172 27228
rect 3196 27226 3252 27228
rect 2956 27174 3002 27226
rect 3002 27174 3012 27226
rect 3036 27174 3066 27226
rect 3066 27174 3078 27226
rect 3078 27174 3092 27226
rect 3116 27174 3130 27226
rect 3130 27174 3142 27226
rect 3142 27174 3172 27226
rect 3196 27174 3206 27226
rect 3206 27174 3252 27226
rect 2956 27172 3012 27174
rect 3036 27172 3092 27174
rect 3116 27172 3172 27174
rect 3196 27172 3252 27174
rect 2956 26138 3012 26140
rect 3036 26138 3092 26140
rect 3116 26138 3172 26140
rect 3196 26138 3252 26140
rect 2956 26086 3002 26138
rect 3002 26086 3012 26138
rect 3036 26086 3066 26138
rect 3066 26086 3078 26138
rect 3078 26086 3092 26138
rect 3116 26086 3130 26138
rect 3130 26086 3142 26138
rect 3142 26086 3172 26138
rect 3196 26086 3206 26138
rect 3206 26086 3252 26138
rect 2956 26084 3012 26086
rect 3036 26084 3092 26086
rect 3116 26084 3172 26086
rect 3196 26084 3252 26086
rect 2956 25050 3012 25052
rect 3036 25050 3092 25052
rect 3116 25050 3172 25052
rect 3196 25050 3252 25052
rect 2956 24998 3002 25050
rect 3002 24998 3012 25050
rect 3036 24998 3066 25050
rect 3066 24998 3078 25050
rect 3078 24998 3092 25050
rect 3116 24998 3130 25050
rect 3130 24998 3142 25050
rect 3142 24998 3172 25050
rect 3196 24998 3206 25050
rect 3206 24998 3252 25050
rect 2956 24996 3012 24998
rect 3036 24996 3092 24998
rect 3116 24996 3172 24998
rect 3196 24996 3252 24998
rect 2956 23962 3012 23964
rect 3036 23962 3092 23964
rect 3116 23962 3172 23964
rect 3196 23962 3252 23964
rect 2956 23910 3002 23962
rect 3002 23910 3012 23962
rect 3036 23910 3066 23962
rect 3066 23910 3078 23962
rect 3078 23910 3092 23962
rect 3116 23910 3130 23962
rect 3130 23910 3142 23962
rect 3142 23910 3172 23962
rect 3196 23910 3206 23962
rect 3206 23910 3252 23962
rect 2956 23908 3012 23910
rect 3036 23908 3092 23910
rect 3116 23908 3172 23910
rect 3196 23908 3252 23910
rect 2956 22874 3012 22876
rect 3036 22874 3092 22876
rect 3116 22874 3172 22876
rect 3196 22874 3252 22876
rect 2956 22822 3002 22874
rect 3002 22822 3012 22874
rect 3036 22822 3066 22874
rect 3066 22822 3078 22874
rect 3078 22822 3092 22874
rect 3116 22822 3130 22874
rect 3130 22822 3142 22874
rect 3142 22822 3172 22874
rect 3196 22822 3206 22874
rect 3206 22822 3252 22874
rect 2956 22820 3012 22822
rect 3036 22820 3092 22822
rect 3116 22820 3172 22822
rect 3196 22820 3252 22822
rect 2956 21786 3012 21788
rect 3036 21786 3092 21788
rect 3116 21786 3172 21788
rect 3196 21786 3252 21788
rect 2956 21734 3002 21786
rect 3002 21734 3012 21786
rect 3036 21734 3066 21786
rect 3066 21734 3078 21786
rect 3078 21734 3092 21786
rect 3116 21734 3130 21786
rect 3130 21734 3142 21786
rect 3142 21734 3172 21786
rect 3196 21734 3206 21786
rect 3206 21734 3252 21786
rect 2956 21732 3012 21734
rect 3036 21732 3092 21734
rect 3116 21732 3172 21734
rect 3196 21732 3252 21734
rect 2956 20698 3012 20700
rect 3036 20698 3092 20700
rect 3116 20698 3172 20700
rect 3196 20698 3252 20700
rect 2956 20646 3002 20698
rect 3002 20646 3012 20698
rect 3036 20646 3066 20698
rect 3066 20646 3078 20698
rect 3078 20646 3092 20698
rect 3116 20646 3130 20698
rect 3130 20646 3142 20698
rect 3142 20646 3172 20698
rect 3196 20646 3206 20698
rect 3206 20646 3252 20698
rect 2956 20644 3012 20646
rect 3036 20644 3092 20646
rect 3116 20644 3172 20646
rect 3196 20644 3252 20646
rect 2956 19610 3012 19612
rect 3036 19610 3092 19612
rect 3116 19610 3172 19612
rect 3196 19610 3252 19612
rect 2956 19558 3002 19610
rect 3002 19558 3012 19610
rect 3036 19558 3066 19610
rect 3066 19558 3078 19610
rect 3078 19558 3092 19610
rect 3116 19558 3130 19610
rect 3130 19558 3142 19610
rect 3142 19558 3172 19610
rect 3196 19558 3206 19610
rect 3206 19558 3252 19610
rect 2956 19556 3012 19558
rect 3036 19556 3092 19558
rect 3116 19556 3172 19558
rect 3196 19556 3252 19558
rect 2956 18522 3012 18524
rect 3036 18522 3092 18524
rect 3116 18522 3172 18524
rect 3196 18522 3252 18524
rect 2956 18470 3002 18522
rect 3002 18470 3012 18522
rect 3036 18470 3066 18522
rect 3066 18470 3078 18522
rect 3078 18470 3092 18522
rect 3116 18470 3130 18522
rect 3130 18470 3142 18522
rect 3142 18470 3172 18522
rect 3196 18470 3206 18522
rect 3206 18470 3252 18522
rect 2956 18468 3012 18470
rect 3036 18468 3092 18470
rect 3116 18468 3172 18470
rect 3196 18468 3252 18470
rect 2956 17434 3012 17436
rect 3036 17434 3092 17436
rect 3116 17434 3172 17436
rect 3196 17434 3252 17436
rect 2956 17382 3002 17434
rect 3002 17382 3012 17434
rect 3036 17382 3066 17434
rect 3066 17382 3078 17434
rect 3078 17382 3092 17434
rect 3116 17382 3130 17434
rect 3130 17382 3142 17434
rect 3142 17382 3172 17434
rect 3196 17382 3206 17434
rect 3206 17382 3252 17434
rect 2956 17380 3012 17382
rect 3036 17380 3092 17382
rect 3116 17380 3172 17382
rect 3196 17380 3252 17382
rect 2956 16346 3012 16348
rect 3036 16346 3092 16348
rect 3116 16346 3172 16348
rect 3196 16346 3252 16348
rect 2956 16294 3002 16346
rect 3002 16294 3012 16346
rect 3036 16294 3066 16346
rect 3066 16294 3078 16346
rect 3078 16294 3092 16346
rect 3116 16294 3130 16346
rect 3130 16294 3142 16346
rect 3142 16294 3172 16346
rect 3196 16294 3206 16346
rect 3206 16294 3252 16346
rect 2956 16292 3012 16294
rect 3036 16292 3092 16294
rect 3116 16292 3172 16294
rect 3196 16292 3252 16294
rect 2956 15258 3012 15260
rect 3036 15258 3092 15260
rect 3116 15258 3172 15260
rect 3196 15258 3252 15260
rect 2956 15206 3002 15258
rect 3002 15206 3012 15258
rect 3036 15206 3066 15258
rect 3066 15206 3078 15258
rect 3078 15206 3092 15258
rect 3116 15206 3130 15258
rect 3130 15206 3142 15258
rect 3142 15206 3172 15258
rect 3196 15206 3206 15258
rect 3206 15206 3252 15258
rect 2956 15204 3012 15206
rect 3036 15204 3092 15206
rect 3116 15204 3172 15206
rect 3196 15204 3252 15206
rect 2956 14170 3012 14172
rect 3036 14170 3092 14172
rect 3116 14170 3172 14172
rect 3196 14170 3252 14172
rect 2956 14118 3002 14170
rect 3002 14118 3012 14170
rect 3036 14118 3066 14170
rect 3066 14118 3078 14170
rect 3078 14118 3092 14170
rect 3116 14118 3130 14170
rect 3130 14118 3142 14170
rect 3142 14118 3172 14170
rect 3196 14118 3206 14170
rect 3206 14118 3252 14170
rect 2956 14116 3012 14118
rect 3036 14116 3092 14118
rect 3116 14116 3172 14118
rect 3196 14116 3252 14118
rect 2956 13082 3012 13084
rect 3036 13082 3092 13084
rect 3116 13082 3172 13084
rect 3196 13082 3252 13084
rect 2956 13030 3002 13082
rect 3002 13030 3012 13082
rect 3036 13030 3066 13082
rect 3066 13030 3078 13082
rect 3078 13030 3092 13082
rect 3116 13030 3130 13082
rect 3130 13030 3142 13082
rect 3142 13030 3172 13082
rect 3196 13030 3206 13082
rect 3206 13030 3252 13082
rect 2956 13028 3012 13030
rect 3036 13028 3092 13030
rect 3116 13028 3172 13030
rect 3196 13028 3252 13030
rect 2956 11994 3012 11996
rect 3036 11994 3092 11996
rect 3116 11994 3172 11996
rect 3196 11994 3252 11996
rect 2956 11942 3002 11994
rect 3002 11942 3012 11994
rect 3036 11942 3066 11994
rect 3066 11942 3078 11994
rect 3078 11942 3092 11994
rect 3116 11942 3130 11994
rect 3130 11942 3142 11994
rect 3142 11942 3172 11994
rect 3196 11942 3206 11994
rect 3206 11942 3252 11994
rect 2956 11940 3012 11942
rect 3036 11940 3092 11942
rect 3116 11940 3172 11942
rect 3196 11940 3252 11942
rect 2956 10906 3012 10908
rect 3036 10906 3092 10908
rect 3116 10906 3172 10908
rect 3196 10906 3252 10908
rect 2956 10854 3002 10906
rect 3002 10854 3012 10906
rect 3036 10854 3066 10906
rect 3066 10854 3078 10906
rect 3078 10854 3092 10906
rect 3116 10854 3130 10906
rect 3130 10854 3142 10906
rect 3142 10854 3172 10906
rect 3196 10854 3206 10906
rect 3206 10854 3252 10906
rect 2956 10852 3012 10854
rect 3036 10852 3092 10854
rect 3116 10852 3172 10854
rect 3196 10852 3252 10854
rect 2956 9818 3012 9820
rect 3036 9818 3092 9820
rect 3116 9818 3172 9820
rect 3196 9818 3252 9820
rect 2956 9766 3002 9818
rect 3002 9766 3012 9818
rect 3036 9766 3066 9818
rect 3066 9766 3078 9818
rect 3078 9766 3092 9818
rect 3116 9766 3130 9818
rect 3130 9766 3142 9818
rect 3142 9766 3172 9818
rect 3196 9766 3206 9818
rect 3206 9766 3252 9818
rect 2956 9764 3012 9766
rect 3036 9764 3092 9766
rect 3116 9764 3172 9766
rect 3196 9764 3252 9766
rect 2956 8730 3012 8732
rect 3036 8730 3092 8732
rect 3116 8730 3172 8732
rect 3196 8730 3252 8732
rect 2956 8678 3002 8730
rect 3002 8678 3012 8730
rect 3036 8678 3066 8730
rect 3066 8678 3078 8730
rect 3078 8678 3092 8730
rect 3116 8678 3130 8730
rect 3130 8678 3142 8730
rect 3142 8678 3172 8730
rect 3196 8678 3206 8730
rect 3206 8678 3252 8730
rect 2956 8676 3012 8678
rect 3036 8676 3092 8678
rect 3116 8676 3172 8678
rect 3196 8676 3252 8678
rect 2956 7642 3012 7644
rect 3036 7642 3092 7644
rect 3116 7642 3172 7644
rect 3196 7642 3252 7644
rect 2956 7590 3002 7642
rect 3002 7590 3012 7642
rect 3036 7590 3066 7642
rect 3066 7590 3078 7642
rect 3078 7590 3092 7642
rect 3116 7590 3130 7642
rect 3130 7590 3142 7642
rect 3142 7590 3172 7642
rect 3196 7590 3206 7642
rect 3206 7590 3252 7642
rect 2956 7588 3012 7590
rect 3036 7588 3092 7590
rect 3116 7588 3172 7590
rect 3196 7588 3252 7590
rect 3616 86522 3672 86524
rect 3696 86522 3752 86524
rect 3776 86522 3832 86524
rect 3856 86522 3912 86524
rect 3616 86470 3662 86522
rect 3662 86470 3672 86522
rect 3696 86470 3726 86522
rect 3726 86470 3738 86522
rect 3738 86470 3752 86522
rect 3776 86470 3790 86522
rect 3790 86470 3802 86522
rect 3802 86470 3832 86522
rect 3856 86470 3866 86522
rect 3866 86470 3912 86522
rect 3616 86468 3672 86470
rect 3696 86468 3752 86470
rect 3776 86468 3832 86470
rect 3856 86468 3912 86470
rect 3616 85434 3672 85436
rect 3696 85434 3752 85436
rect 3776 85434 3832 85436
rect 3856 85434 3912 85436
rect 3616 85382 3662 85434
rect 3662 85382 3672 85434
rect 3696 85382 3726 85434
rect 3726 85382 3738 85434
rect 3738 85382 3752 85434
rect 3776 85382 3790 85434
rect 3790 85382 3802 85434
rect 3802 85382 3832 85434
rect 3856 85382 3866 85434
rect 3866 85382 3912 85434
rect 3616 85380 3672 85382
rect 3696 85380 3752 85382
rect 3776 85380 3832 85382
rect 3856 85380 3912 85382
rect 3616 84346 3672 84348
rect 3696 84346 3752 84348
rect 3776 84346 3832 84348
rect 3856 84346 3912 84348
rect 3616 84294 3662 84346
rect 3662 84294 3672 84346
rect 3696 84294 3726 84346
rect 3726 84294 3738 84346
rect 3738 84294 3752 84346
rect 3776 84294 3790 84346
rect 3790 84294 3802 84346
rect 3802 84294 3832 84346
rect 3856 84294 3866 84346
rect 3866 84294 3912 84346
rect 3616 84292 3672 84294
rect 3696 84292 3752 84294
rect 3776 84292 3832 84294
rect 3856 84292 3912 84294
rect 3616 83258 3672 83260
rect 3696 83258 3752 83260
rect 3776 83258 3832 83260
rect 3856 83258 3912 83260
rect 3616 83206 3662 83258
rect 3662 83206 3672 83258
rect 3696 83206 3726 83258
rect 3726 83206 3738 83258
rect 3738 83206 3752 83258
rect 3776 83206 3790 83258
rect 3790 83206 3802 83258
rect 3802 83206 3832 83258
rect 3856 83206 3866 83258
rect 3866 83206 3912 83258
rect 3616 83204 3672 83206
rect 3696 83204 3752 83206
rect 3776 83204 3832 83206
rect 3856 83204 3912 83206
rect 3616 82170 3672 82172
rect 3696 82170 3752 82172
rect 3776 82170 3832 82172
rect 3856 82170 3912 82172
rect 3616 82118 3662 82170
rect 3662 82118 3672 82170
rect 3696 82118 3726 82170
rect 3726 82118 3738 82170
rect 3738 82118 3752 82170
rect 3776 82118 3790 82170
rect 3790 82118 3802 82170
rect 3802 82118 3832 82170
rect 3856 82118 3866 82170
rect 3866 82118 3912 82170
rect 3616 82116 3672 82118
rect 3696 82116 3752 82118
rect 3776 82116 3832 82118
rect 3856 82116 3912 82118
rect 3616 81082 3672 81084
rect 3696 81082 3752 81084
rect 3776 81082 3832 81084
rect 3856 81082 3912 81084
rect 3616 81030 3662 81082
rect 3662 81030 3672 81082
rect 3696 81030 3726 81082
rect 3726 81030 3738 81082
rect 3738 81030 3752 81082
rect 3776 81030 3790 81082
rect 3790 81030 3802 81082
rect 3802 81030 3832 81082
rect 3856 81030 3866 81082
rect 3866 81030 3912 81082
rect 3616 81028 3672 81030
rect 3696 81028 3752 81030
rect 3776 81028 3832 81030
rect 3856 81028 3912 81030
rect 3616 79994 3672 79996
rect 3696 79994 3752 79996
rect 3776 79994 3832 79996
rect 3856 79994 3912 79996
rect 3616 79942 3662 79994
rect 3662 79942 3672 79994
rect 3696 79942 3726 79994
rect 3726 79942 3738 79994
rect 3738 79942 3752 79994
rect 3776 79942 3790 79994
rect 3790 79942 3802 79994
rect 3802 79942 3832 79994
rect 3856 79942 3866 79994
rect 3866 79942 3912 79994
rect 3616 79940 3672 79942
rect 3696 79940 3752 79942
rect 3776 79940 3832 79942
rect 3856 79940 3912 79942
rect 3616 78906 3672 78908
rect 3696 78906 3752 78908
rect 3776 78906 3832 78908
rect 3856 78906 3912 78908
rect 3616 78854 3662 78906
rect 3662 78854 3672 78906
rect 3696 78854 3726 78906
rect 3726 78854 3738 78906
rect 3738 78854 3752 78906
rect 3776 78854 3790 78906
rect 3790 78854 3802 78906
rect 3802 78854 3832 78906
rect 3856 78854 3866 78906
rect 3866 78854 3912 78906
rect 3616 78852 3672 78854
rect 3696 78852 3752 78854
rect 3776 78852 3832 78854
rect 3856 78852 3912 78854
rect 3616 77818 3672 77820
rect 3696 77818 3752 77820
rect 3776 77818 3832 77820
rect 3856 77818 3912 77820
rect 3616 77766 3662 77818
rect 3662 77766 3672 77818
rect 3696 77766 3726 77818
rect 3726 77766 3738 77818
rect 3738 77766 3752 77818
rect 3776 77766 3790 77818
rect 3790 77766 3802 77818
rect 3802 77766 3832 77818
rect 3856 77766 3866 77818
rect 3866 77766 3912 77818
rect 3616 77764 3672 77766
rect 3696 77764 3752 77766
rect 3776 77764 3832 77766
rect 3856 77764 3912 77766
rect 3616 76730 3672 76732
rect 3696 76730 3752 76732
rect 3776 76730 3832 76732
rect 3856 76730 3912 76732
rect 3616 76678 3662 76730
rect 3662 76678 3672 76730
rect 3696 76678 3726 76730
rect 3726 76678 3738 76730
rect 3738 76678 3752 76730
rect 3776 76678 3790 76730
rect 3790 76678 3802 76730
rect 3802 76678 3832 76730
rect 3856 76678 3866 76730
rect 3866 76678 3912 76730
rect 3616 76676 3672 76678
rect 3696 76676 3752 76678
rect 3776 76676 3832 76678
rect 3856 76676 3912 76678
rect 3616 75642 3672 75644
rect 3696 75642 3752 75644
rect 3776 75642 3832 75644
rect 3856 75642 3912 75644
rect 3616 75590 3662 75642
rect 3662 75590 3672 75642
rect 3696 75590 3726 75642
rect 3726 75590 3738 75642
rect 3738 75590 3752 75642
rect 3776 75590 3790 75642
rect 3790 75590 3802 75642
rect 3802 75590 3832 75642
rect 3856 75590 3866 75642
rect 3866 75590 3912 75642
rect 3616 75588 3672 75590
rect 3696 75588 3752 75590
rect 3776 75588 3832 75590
rect 3856 75588 3912 75590
rect 3616 74554 3672 74556
rect 3696 74554 3752 74556
rect 3776 74554 3832 74556
rect 3856 74554 3912 74556
rect 3616 74502 3662 74554
rect 3662 74502 3672 74554
rect 3696 74502 3726 74554
rect 3726 74502 3738 74554
rect 3738 74502 3752 74554
rect 3776 74502 3790 74554
rect 3790 74502 3802 74554
rect 3802 74502 3832 74554
rect 3856 74502 3866 74554
rect 3866 74502 3912 74554
rect 3616 74500 3672 74502
rect 3696 74500 3752 74502
rect 3776 74500 3832 74502
rect 3856 74500 3912 74502
rect 3616 73466 3672 73468
rect 3696 73466 3752 73468
rect 3776 73466 3832 73468
rect 3856 73466 3912 73468
rect 3616 73414 3662 73466
rect 3662 73414 3672 73466
rect 3696 73414 3726 73466
rect 3726 73414 3738 73466
rect 3738 73414 3752 73466
rect 3776 73414 3790 73466
rect 3790 73414 3802 73466
rect 3802 73414 3832 73466
rect 3856 73414 3866 73466
rect 3866 73414 3912 73466
rect 3616 73412 3672 73414
rect 3696 73412 3752 73414
rect 3776 73412 3832 73414
rect 3856 73412 3912 73414
rect 3616 72378 3672 72380
rect 3696 72378 3752 72380
rect 3776 72378 3832 72380
rect 3856 72378 3912 72380
rect 3616 72326 3662 72378
rect 3662 72326 3672 72378
rect 3696 72326 3726 72378
rect 3726 72326 3738 72378
rect 3738 72326 3752 72378
rect 3776 72326 3790 72378
rect 3790 72326 3802 72378
rect 3802 72326 3832 72378
rect 3856 72326 3866 72378
rect 3866 72326 3912 72378
rect 3616 72324 3672 72326
rect 3696 72324 3752 72326
rect 3776 72324 3832 72326
rect 3856 72324 3912 72326
rect 3616 71290 3672 71292
rect 3696 71290 3752 71292
rect 3776 71290 3832 71292
rect 3856 71290 3912 71292
rect 3616 71238 3662 71290
rect 3662 71238 3672 71290
rect 3696 71238 3726 71290
rect 3726 71238 3738 71290
rect 3738 71238 3752 71290
rect 3776 71238 3790 71290
rect 3790 71238 3802 71290
rect 3802 71238 3832 71290
rect 3856 71238 3866 71290
rect 3866 71238 3912 71290
rect 3616 71236 3672 71238
rect 3696 71236 3752 71238
rect 3776 71236 3832 71238
rect 3856 71236 3912 71238
rect 3616 70202 3672 70204
rect 3696 70202 3752 70204
rect 3776 70202 3832 70204
rect 3856 70202 3912 70204
rect 3616 70150 3662 70202
rect 3662 70150 3672 70202
rect 3696 70150 3726 70202
rect 3726 70150 3738 70202
rect 3738 70150 3752 70202
rect 3776 70150 3790 70202
rect 3790 70150 3802 70202
rect 3802 70150 3832 70202
rect 3856 70150 3866 70202
rect 3866 70150 3912 70202
rect 3616 70148 3672 70150
rect 3696 70148 3752 70150
rect 3776 70148 3832 70150
rect 3856 70148 3912 70150
rect 3616 69114 3672 69116
rect 3696 69114 3752 69116
rect 3776 69114 3832 69116
rect 3856 69114 3912 69116
rect 3616 69062 3662 69114
rect 3662 69062 3672 69114
rect 3696 69062 3726 69114
rect 3726 69062 3738 69114
rect 3738 69062 3752 69114
rect 3776 69062 3790 69114
rect 3790 69062 3802 69114
rect 3802 69062 3832 69114
rect 3856 69062 3866 69114
rect 3866 69062 3912 69114
rect 3616 69060 3672 69062
rect 3696 69060 3752 69062
rect 3776 69060 3832 69062
rect 3856 69060 3912 69062
rect 3616 68026 3672 68028
rect 3696 68026 3752 68028
rect 3776 68026 3832 68028
rect 3856 68026 3912 68028
rect 3616 67974 3662 68026
rect 3662 67974 3672 68026
rect 3696 67974 3726 68026
rect 3726 67974 3738 68026
rect 3738 67974 3752 68026
rect 3776 67974 3790 68026
rect 3790 67974 3802 68026
rect 3802 67974 3832 68026
rect 3856 67974 3866 68026
rect 3866 67974 3912 68026
rect 3616 67972 3672 67974
rect 3696 67972 3752 67974
rect 3776 67972 3832 67974
rect 3856 67972 3912 67974
rect 3882 67768 3938 67824
rect 3616 66938 3672 66940
rect 3696 66938 3752 66940
rect 3776 66938 3832 66940
rect 3856 66938 3912 66940
rect 3616 66886 3662 66938
rect 3662 66886 3672 66938
rect 3696 66886 3726 66938
rect 3726 66886 3738 66938
rect 3738 66886 3752 66938
rect 3776 66886 3790 66938
rect 3790 66886 3802 66938
rect 3802 66886 3832 66938
rect 3856 66886 3866 66938
rect 3866 66886 3912 66938
rect 3616 66884 3672 66886
rect 3696 66884 3752 66886
rect 3776 66884 3832 66886
rect 3856 66884 3912 66886
rect 3616 65850 3672 65852
rect 3696 65850 3752 65852
rect 3776 65850 3832 65852
rect 3856 65850 3912 65852
rect 3616 65798 3662 65850
rect 3662 65798 3672 65850
rect 3696 65798 3726 65850
rect 3726 65798 3738 65850
rect 3738 65798 3752 65850
rect 3776 65798 3790 65850
rect 3790 65798 3802 65850
rect 3802 65798 3832 65850
rect 3856 65798 3866 65850
rect 3866 65798 3912 65850
rect 3616 65796 3672 65798
rect 3696 65796 3752 65798
rect 3776 65796 3832 65798
rect 3856 65796 3912 65798
rect 3616 64762 3672 64764
rect 3696 64762 3752 64764
rect 3776 64762 3832 64764
rect 3856 64762 3912 64764
rect 3616 64710 3662 64762
rect 3662 64710 3672 64762
rect 3696 64710 3726 64762
rect 3726 64710 3738 64762
rect 3738 64710 3752 64762
rect 3776 64710 3790 64762
rect 3790 64710 3802 64762
rect 3802 64710 3832 64762
rect 3856 64710 3866 64762
rect 3866 64710 3912 64762
rect 3616 64708 3672 64710
rect 3696 64708 3752 64710
rect 3776 64708 3832 64710
rect 3856 64708 3912 64710
rect 3616 63674 3672 63676
rect 3696 63674 3752 63676
rect 3776 63674 3832 63676
rect 3856 63674 3912 63676
rect 3616 63622 3662 63674
rect 3662 63622 3672 63674
rect 3696 63622 3726 63674
rect 3726 63622 3738 63674
rect 3738 63622 3752 63674
rect 3776 63622 3790 63674
rect 3790 63622 3802 63674
rect 3802 63622 3832 63674
rect 3856 63622 3866 63674
rect 3866 63622 3912 63674
rect 3616 63620 3672 63622
rect 3696 63620 3752 63622
rect 3776 63620 3832 63622
rect 3856 63620 3912 63622
rect 3606 62872 3662 62928
rect 3616 62586 3672 62588
rect 3696 62586 3752 62588
rect 3776 62586 3832 62588
rect 3856 62586 3912 62588
rect 3616 62534 3662 62586
rect 3662 62534 3672 62586
rect 3696 62534 3726 62586
rect 3726 62534 3738 62586
rect 3738 62534 3752 62586
rect 3776 62534 3790 62586
rect 3790 62534 3802 62586
rect 3802 62534 3832 62586
rect 3856 62534 3866 62586
rect 3866 62534 3912 62586
rect 3616 62532 3672 62534
rect 3696 62532 3752 62534
rect 3776 62532 3832 62534
rect 3856 62532 3912 62534
rect 3616 61498 3672 61500
rect 3696 61498 3752 61500
rect 3776 61498 3832 61500
rect 3856 61498 3912 61500
rect 3616 61446 3662 61498
rect 3662 61446 3672 61498
rect 3696 61446 3726 61498
rect 3726 61446 3738 61498
rect 3738 61446 3752 61498
rect 3776 61446 3790 61498
rect 3790 61446 3802 61498
rect 3802 61446 3832 61498
rect 3856 61446 3866 61498
rect 3866 61446 3912 61498
rect 3616 61444 3672 61446
rect 3696 61444 3752 61446
rect 3776 61444 3832 61446
rect 3856 61444 3912 61446
rect 3616 60410 3672 60412
rect 3696 60410 3752 60412
rect 3776 60410 3832 60412
rect 3856 60410 3912 60412
rect 3616 60358 3662 60410
rect 3662 60358 3672 60410
rect 3696 60358 3726 60410
rect 3726 60358 3738 60410
rect 3738 60358 3752 60410
rect 3776 60358 3790 60410
rect 3790 60358 3802 60410
rect 3802 60358 3832 60410
rect 3856 60358 3866 60410
rect 3866 60358 3912 60410
rect 3616 60356 3672 60358
rect 3696 60356 3752 60358
rect 3776 60356 3832 60358
rect 3856 60356 3912 60358
rect 3616 59322 3672 59324
rect 3696 59322 3752 59324
rect 3776 59322 3832 59324
rect 3856 59322 3912 59324
rect 3616 59270 3662 59322
rect 3662 59270 3672 59322
rect 3696 59270 3726 59322
rect 3726 59270 3738 59322
rect 3738 59270 3752 59322
rect 3776 59270 3790 59322
rect 3790 59270 3802 59322
rect 3802 59270 3832 59322
rect 3856 59270 3866 59322
rect 3866 59270 3912 59322
rect 3616 59268 3672 59270
rect 3696 59268 3752 59270
rect 3776 59268 3832 59270
rect 3856 59268 3912 59270
rect 3616 58234 3672 58236
rect 3696 58234 3752 58236
rect 3776 58234 3832 58236
rect 3856 58234 3912 58236
rect 3616 58182 3662 58234
rect 3662 58182 3672 58234
rect 3696 58182 3726 58234
rect 3726 58182 3738 58234
rect 3738 58182 3752 58234
rect 3776 58182 3790 58234
rect 3790 58182 3802 58234
rect 3802 58182 3832 58234
rect 3856 58182 3866 58234
rect 3866 58182 3912 58234
rect 3616 58180 3672 58182
rect 3696 58180 3752 58182
rect 3776 58180 3832 58182
rect 3856 58180 3912 58182
rect 3616 57146 3672 57148
rect 3696 57146 3752 57148
rect 3776 57146 3832 57148
rect 3856 57146 3912 57148
rect 3616 57094 3662 57146
rect 3662 57094 3672 57146
rect 3696 57094 3726 57146
rect 3726 57094 3738 57146
rect 3738 57094 3752 57146
rect 3776 57094 3790 57146
rect 3790 57094 3802 57146
rect 3802 57094 3832 57146
rect 3856 57094 3866 57146
rect 3866 57094 3912 57146
rect 3616 57092 3672 57094
rect 3696 57092 3752 57094
rect 3776 57092 3832 57094
rect 3856 57092 3912 57094
rect 3616 56058 3672 56060
rect 3696 56058 3752 56060
rect 3776 56058 3832 56060
rect 3856 56058 3912 56060
rect 3616 56006 3662 56058
rect 3662 56006 3672 56058
rect 3696 56006 3726 56058
rect 3726 56006 3738 56058
rect 3738 56006 3752 56058
rect 3776 56006 3790 56058
rect 3790 56006 3802 56058
rect 3802 56006 3832 56058
rect 3856 56006 3866 56058
rect 3866 56006 3912 56058
rect 3616 56004 3672 56006
rect 3696 56004 3752 56006
rect 3776 56004 3832 56006
rect 3856 56004 3912 56006
rect 3616 54970 3672 54972
rect 3696 54970 3752 54972
rect 3776 54970 3832 54972
rect 3856 54970 3912 54972
rect 3616 54918 3662 54970
rect 3662 54918 3672 54970
rect 3696 54918 3726 54970
rect 3726 54918 3738 54970
rect 3738 54918 3752 54970
rect 3776 54918 3790 54970
rect 3790 54918 3802 54970
rect 3802 54918 3832 54970
rect 3856 54918 3866 54970
rect 3866 54918 3912 54970
rect 3616 54916 3672 54918
rect 3696 54916 3752 54918
rect 3776 54916 3832 54918
rect 3856 54916 3912 54918
rect 3616 53882 3672 53884
rect 3696 53882 3752 53884
rect 3776 53882 3832 53884
rect 3856 53882 3912 53884
rect 3616 53830 3662 53882
rect 3662 53830 3672 53882
rect 3696 53830 3726 53882
rect 3726 53830 3738 53882
rect 3738 53830 3752 53882
rect 3776 53830 3790 53882
rect 3790 53830 3802 53882
rect 3802 53830 3832 53882
rect 3856 53830 3866 53882
rect 3866 53830 3912 53882
rect 3616 53828 3672 53830
rect 3696 53828 3752 53830
rect 3776 53828 3832 53830
rect 3856 53828 3912 53830
rect 3616 52794 3672 52796
rect 3696 52794 3752 52796
rect 3776 52794 3832 52796
rect 3856 52794 3912 52796
rect 3616 52742 3662 52794
rect 3662 52742 3672 52794
rect 3696 52742 3726 52794
rect 3726 52742 3738 52794
rect 3738 52742 3752 52794
rect 3776 52742 3790 52794
rect 3790 52742 3802 52794
rect 3802 52742 3832 52794
rect 3856 52742 3866 52794
rect 3866 52742 3912 52794
rect 3616 52740 3672 52742
rect 3696 52740 3752 52742
rect 3776 52740 3832 52742
rect 3856 52740 3912 52742
rect 3616 51706 3672 51708
rect 3696 51706 3752 51708
rect 3776 51706 3832 51708
rect 3856 51706 3912 51708
rect 3616 51654 3662 51706
rect 3662 51654 3672 51706
rect 3696 51654 3726 51706
rect 3726 51654 3738 51706
rect 3738 51654 3752 51706
rect 3776 51654 3790 51706
rect 3790 51654 3802 51706
rect 3802 51654 3832 51706
rect 3856 51654 3866 51706
rect 3866 51654 3912 51706
rect 3616 51652 3672 51654
rect 3696 51652 3752 51654
rect 3776 51652 3832 51654
rect 3856 51652 3912 51654
rect 3616 50618 3672 50620
rect 3696 50618 3752 50620
rect 3776 50618 3832 50620
rect 3856 50618 3912 50620
rect 3616 50566 3662 50618
rect 3662 50566 3672 50618
rect 3696 50566 3726 50618
rect 3726 50566 3738 50618
rect 3738 50566 3752 50618
rect 3776 50566 3790 50618
rect 3790 50566 3802 50618
rect 3802 50566 3832 50618
rect 3856 50566 3866 50618
rect 3866 50566 3912 50618
rect 3616 50564 3672 50566
rect 3696 50564 3752 50566
rect 3776 50564 3832 50566
rect 3856 50564 3912 50566
rect 3616 49530 3672 49532
rect 3696 49530 3752 49532
rect 3776 49530 3832 49532
rect 3856 49530 3912 49532
rect 3616 49478 3662 49530
rect 3662 49478 3672 49530
rect 3696 49478 3726 49530
rect 3726 49478 3738 49530
rect 3738 49478 3752 49530
rect 3776 49478 3790 49530
rect 3790 49478 3802 49530
rect 3802 49478 3832 49530
rect 3856 49478 3866 49530
rect 3866 49478 3912 49530
rect 3616 49476 3672 49478
rect 3696 49476 3752 49478
rect 3776 49476 3832 49478
rect 3856 49476 3912 49478
rect 3616 48442 3672 48444
rect 3696 48442 3752 48444
rect 3776 48442 3832 48444
rect 3856 48442 3912 48444
rect 3616 48390 3662 48442
rect 3662 48390 3672 48442
rect 3696 48390 3726 48442
rect 3726 48390 3738 48442
rect 3738 48390 3752 48442
rect 3776 48390 3790 48442
rect 3790 48390 3802 48442
rect 3802 48390 3832 48442
rect 3856 48390 3866 48442
rect 3866 48390 3912 48442
rect 3616 48388 3672 48390
rect 3696 48388 3752 48390
rect 3776 48388 3832 48390
rect 3856 48388 3912 48390
rect 3616 47354 3672 47356
rect 3696 47354 3752 47356
rect 3776 47354 3832 47356
rect 3856 47354 3912 47356
rect 3616 47302 3662 47354
rect 3662 47302 3672 47354
rect 3696 47302 3726 47354
rect 3726 47302 3738 47354
rect 3738 47302 3752 47354
rect 3776 47302 3790 47354
rect 3790 47302 3802 47354
rect 3802 47302 3832 47354
rect 3856 47302 3866 47354
rect 3866 47302 3912 47354
rect 3616 47300 3672 47302
rect 3696 47300 3752 47302
rect 3776 47300 3832 47302
rect 3856 47300 3912 47302
rect 3616 46266 3672 46268
rect 3696 46266 3752 46268
rect 3776 46266 3832 46268
rect 3856 46266 3912 46268
rect 3616 46214 3662 46266
rect 3662 46214 3672 46266
rect 3696 46214 3726 46266
rect 3726 46214 3738 46266
rect 3738 46214 3752 46266
rect 3776 46214 3790 46266
rect 3790 46214 3802 46266
rect 3802 46214 3832 46266
rect 3856 46214 3866 46266
rect 3866 46214 3912 46266
rect 3616 46212 3672 46214
rect 3696 46212 3752 46214
rect 3776 46212 3832 46214
rect 3856 46212 3912 46214
rect 3616 45178 3672 45180
rect 3696 45178 3752 45180
rect 3776 45178 3832 45180
rect 3856 45178 3912 45180
rect 3616 45126 3662 45178
rect 3662 45126 3672 45178
rect 3696 45126 3726 45178
rect 3726 45126 3738 45178
rect 3738 45126 3752 45178
rect 3776 45126 3790 45178
rect 3790 45126 3802 45178
rect 3802 45126 3832 45178
rect 3856 45126 3866 45178
rect 3866 45126 3912 45178
rect 3616 45124 3672 45126
rect 3696 45124 3752 45126
rect 3776 45124 3832 45126
rect 3856 45124 3912 45126
rect 4556 85978 4612 85980
rect 4636 85978 4692 85980
rect 4716 85978 4772 85980
rect 4796 85978 4852 85980
rect 4556 85926 4602 85978
rect 4602 85926 4612 85978
rect 4636 85926 4666 85978
rect 4666 85926 4678 85978
rect 4678 85926 4692 85978
rect 4716 85926 4730 85978
rect 4730 85926 4742 85978
rect 4742 85926 4772 85978
rect 4796 85926 4806 85978
rect 4806 85926 4852 85978
rect 4556 85924 4612 85926
rect 4636 85924 4692 85926
rect 4716 85924 4772 85926
rect 4796 85924 4852 85926
rect 4556 84890 4612 84892
rect 4636 84890 4692 84892
rect 4716 84890 4772 84892
rect 4796 84890 4852 84892
rect 4556 84838 4602 84890
rect 4602 84838 4612 84890
rect 4636 84838 4666 84890
rect 4666 84838 4678 84890
rect 4678 84838 4692 84890
rect 4716 84838 4730 84890
rect 4730 84838 4742 84890
rect 4742 84838 4772 84890
rect 4796 84838 4806 84890
rect 4806 84838 4852 84890
rect 4556 84836 4612 84838
rect 4636 84836 4692 84838
rect 4716 84836 4772 84838
rect 4796 84836 4852 84838
rect 4556 83802 4612 83804
rect 4636 83802 4692 83804
rect 4716 83802 4772 83804
rect 4796 83802 4852 83804
rect 4556 83750 4602 83802
rect 4602 83750 4612 83802
rect 4636 83750 4666 83802
rect 4666 83750 4678 83802
rect 4678 83750 4692 83802
rect 4716 83750 4730 83802
rect 4730 83750 4742 83802
rect 4742 83750 4772 83802
rect 4796 83750 4806 83802
rect 4806 83750 4852 83802
rect 4556 83748 4612 83750
rect 4636 83748 4692 83750
rect 4716 83748 4772 83750
rect 4796 83748 4852 83750
rect 4556 82714 4612 82716
rect 4636 82714 4692 82716
rect 4716 82714 4772 82716
rect 4796 82714 4852 82716
rect 4556 82662 4602 82714
rect 4602 82662 4612 82714
rect 4636 82662 4666 82714
rect 4666 82662 4678 82714
rect 4678 82662 4692 82714
rect 4716 82662 4730 82714
rect 4730 82662 4742 82714
rect 4742 82662 4772 82714
rect 4796 82662 4806 82714
rect 4806 82662 4852 82714
rect 4556 82660 4612 82662
rect 4636 82660 4692 82662
rect 4716 82660 4772 82662
rect 4796 82660 4852 82662
rect 4556 81626 4612 81628
rect 4636 81626 4692 81628
rect 4716 81626 4772 81628
rect 4796 81626 4852 81628
rect 4556 81574 4602 81626
rect 4602 81574 4612 81626
rect 4636 81574 4666 81626
rect 4666 81574 4678 81626
rect 4678 81574 4692 81626
rect 4716 81574 4730 81626
rect 4730 81574 4742 81626
rect 4742 81574 4772 81626
rect 4796 81574 4806 81626
rect 4806 81574 4852 81626
rect 4556 81572 4612 81574
rect 4636 81572 4692 81574
rect 4716 81572 4772 81574
rect 4796 81572 4852 81574
rect 4556 80538 4612 80540
rect 4636 80538 4692 80540
rect 4716 80538 4772 80540
rect 4796 80538 4852 80540
rect 4556 80486 4602 80538
rect 4602 80486 4612 80538
rect 4636 80486 4666 80538
rect 4666 80486 4678 80538
rect 4678 80486 4692 80538
rect 4716 80486 4730 80538
rect 4730 80486 4742 80538
rect 4742 80486 4772 80538
rect 4796 80486 4806 80538
rect 4806 80486 4852 80538
rect 4556 80484 4612 80486
rect 4636 80484 4692 80486
rect 4716 80484 4772 80486
rect 4796 80484 4852 80486
rect 4556 79450 4612 79452
rect 4636 79450 4692 79452
rect 4716 79450 4772 79452
rect 4796 79450 4852 79452
rect 4556 79398 4602 79450
rect 4602 79398 4612 79450
rect 4636 79398 4666 79450
rect 4666 79398 4678 79450
rect 4678 79398 4692 79450
rect 4716 79398 4730 79450
rect 4730 79398 4742 79450
rect 4742 79398 4772 79450
rect 4796 79398 4806 79450
rect 4806 79398 4852 79450
rect 4556 79396 4612 79398
rect 4636 79396 4692 79398
rect 4716 79396 4772 79398
rect 4796 79396 4852 79398
rect 4556 78362 4612 78364
rect 4636 78362 4692 78364
rect 4716 78362 4772 78364
rect 4796 78362 4852 78364
rect 4556 78310 4602 78362
rect 4602 78310 4612 78362
rect 4636 78310 4666 78362
rect 4666 78310 4678 78362
rect 4678 78310 4692 78362
rect 4716 78310 4730 78362
rect 4730 78310 4742 78362
rect 4742 78310 4772 78362
rect 4796 78310 4806 78362
rect 4806 78310 4852 78362
rect 4556 78308 4612 78310
rect 4636 78308 4692 78310
rect 4716 78308 4772 78310
rect 4796 78308 4852 78310
rect 4556 77274 4612 77276
rect 4636 77274 4692 77276
rect 4716 77274 4772 77276
rect 4796 77274 4852 77276
rect 4556 77222 4602 77274
rect 4602 77222 4612 77274
rect 4636 77222 4666 77274
rect 4666 77222 4678 77274
rect 4678 77222 4692 77274
rect 4716 77222 4730 77274
rect 4730 77222 4742 77274
rect 4742 77222 4772 77274
rect 4796 77222 4806 77274
rect 4806 77222 4852 77274
rect 4556 77220 4612 77222
rect 4636 77220 4692 77222
rect 4716 77220 4772 77222
rect 4796 77220 4852 77222
rect 4556 76186 4612 76188
rect 4636 76186 4692 76188
rect 4716 76186 4772 76188
rect 4796 76186 4852 76188
rect 4556 76134 4602 76186
rect 4602 76134 4612 76186
rect 4636 76134 4666 76186
rect 4666 76134 4678 76186
rect 4678 76134 4692 76186
rect 4716 76134 4730 76186
rect 4730 76134 4742 76186
rect 4742 76134 4772 76186
rect 4796 76134 4806 76186
rect 4806 76134 4852 76186
rect 4556 76132 4612 76134
rect 4636 76132 4692 76134
rect 4716 76132 4772 76134
rect 4796 76132 4852 76134
rect 5216 86522 5272 86524
rect 5296 86522 5352 86524
rect 5376 86522 5432 86524
rect 5456 86522 5512 86524
rect 5216 86470 5262 86522
rect 5262 86470 5272 86522
rect 5296 86470 5326 86522
rect 5326 86470 5338 86522
rect 5338 86470 5352 86522
rect 5376 86470 5390 86522
rect 5390 86470 5402 86522
rect 5402 86470 5432 86522
rect 5456 86470 5466 86522
rect 5466 86470 5512 86522
rect 5216 86468 5272 86470
rect 5296 86468 5352 86470
rect 5376 86468 5432 86470
rect 5456 86468 5512 86470
rect 5216 85434 5272 85436
rect 5296 85434 5352 85436
rect 5376 85434 5432 85436
rect 5456 85434 5512 85436
rect 5216 85382 5262 85434
rect 5262 85382 5272 85434
rect 5296 85382 5326 85434
rect 5326 85382 5338 85434
rect 5338 85382 5352 85434
rect 5376 85382 5390 85434
rect 5390 85382 5402 85434
rect 5402 85382 5432 85434
rect 5456 85382 5466 85434
rect 5466 85382 5512 85434
rect 5216 85380 5272 85382
rect 5296 85380 5352 85382
rect 5376 85380 5432 85382
rect 5456 85380 5512 85382
rect 5078 85040 5134 85096
rect 4556 75098 4612 75100
rect 4636 75098 4692 75100
rect 4716 75098 4772 75100
rect 4796 75098 4852 75100
rect 4556 75046 4602 75098
rect 4602 75046 4612 75098
rect 4636 75046 4666 75098
rect 4666 75046 4678 75098
rect 4678 75046 4692 75098
rect 4716 75046 4730 75098
rect 4730 75046 4742 75098
rect 4742 75046 4772 75098
rect 4796 75046 4806 75098
rect 4806 75046 4852 75098
rect 4556 75044 4612 75046
rect 4636 75044 4692 75046
rect 4716 75044 4772 75046
rect 4796 75044 4852 75046
rect 4556 74010 4612 74012
rect 4636 74010 4692 74012
rect 4716 74010 4772 74012
rect 4796 74010 4852 74012
rect 4556 73958 4602 74010
rect 4602 73958 4612 74010
rect 4636 73958 4666 74010
rect 4666 73958 4678 74010
rect 4678 73958 4692 74010
rect 4716 73958 4730 74010
rect 4730 73958 4742 74010
rect 4742 73958 4772 74010
rect 4796 73958 4806 74010
rect 4806 73958 4852 74010
rect 4556 73956 4612 73958
rect 4636 73956 4692 73958
rect 4716 73956 4772 73958
rect 4796 73956 4852 73958
rect 4556 72922 4612 72924
rect 4636 72922 4692 72924
rect 4716 72922 4772 72924
rect 4796 72922 4852 72924
rect 4556 72870 4602 72922
rect 4602 72870 4612 72922
rect 4636 72870 4666 72922
rect 4666 72870 4678 72922
rect 4678 72870 4692 72922
rect 4716 72870 4730 72922
rect 4730 72870 4742 72922
rect 4742 72870 4772 72922
rect 4796 72870 4806 72922
rect 4806 72870 4852 72922
rect 4556 72868 4612 72870
rect 4636 72868 4692 72870
rect 4716 72868 4772 72870
rect 4796 72868 4852 72870
rect 4556 71834 4612 71836
rect 4636 71834 4692 71836
rect 4716 71834 4772 71836
rect 4796 71834 4852 71836
rect 4556 71782 4602 71834
rect 4602 71782 4612 71834
rect 4636 71782 4666 71834
rect 4666 71782 4678 71834
rect 4678 71782 4692 71834
rect 4716 71782 4730 71834
rect 4730 71782 4742 71834
rect 4742 71782 4772 71834
rect 4796 71782 4806 71834
rect 4806 71782 4852 71834
rect 4556 71780 4612 71782
rect 4636 71780 4692 71782
rect 4716 71780 4772 71782
rect 4796 71780 4852 71782
rect 4556 70746 4612 70748
rect 4636 70746 4692 70748
rect 4716 70746 4772 70748
rect 4796 70746 4852 70748
rect 4556 70694 4602 70746
rect 4602 70694 4612 70746
rect 4636 70694 4666 70746
rect 4666 70694 4678 70746
rect 4678 70694 4692 70746
rect 4716 70694 4730 70746
rect 4730 70694 4742 70746
rect 4742 70694 4772 70746
rect 4796 70694 4806 70746
rect 4806 70694 4852 70746
rect 4556 70692 4612 70694
rect 4636 70692 4692 70694
rect 4716 70692 4772 70694
rect 4796 70692 4852 70694
rect 4158 68856 4214 68912
rect 4710 70352 4766 70408
rect 4556 69658 4612 69660
rect 4636 69658 4692 69660
rect 4716 69658 4772 69660
rect 4796 69658 4852 69660
rect 4556 69606 4602 69658
rect 4602 69606 4612 69658
rect 4636 69606 4666 69658
rect 4666 69606 4678 69658
rect 4678 69606 4692 69658
rect 4716 69606 4730 69658
rect 4730 69606 4742 69658
rect 4742 69606 4772 69658
rect 4796 69606 4806 69658
rect 4806 69606 4852 69658
rect 4556 69604 4612 69606
rect 4636 69604 4692 69606
rect 4716 69604 4772 69606
rect 4796 69604 4852 69606
rect 4556 68570 4612 68572
rect 4636 68570 4692 68572
rect 4716 68570 4772 68572
rect 4796 68570 4852 68572
rect 4556 68518 4602 68570
rect 4602 68518 4612 68570
rect 4636 68518 4666 68570
rect 4666 68518 4678 68570
rect 4678 68518 4692 68570
rect 4716 68518 4730 68570
rect 4730 68518 4742 68570
rect 4742 68518 4772 68570
rect 4796 68518 4806 68570
rect 4806 68518 4852 68570
rect 4556 68516 4612 68518
rect 4636 68516 4692 68518
rect 4716 68516 4772 68518
rect 4796 68516 4852 68518
rect 4342 67768 4398 67824
rect 4342 67260 4344 67280
rect 4344 67260 4396 67280
rect 4396 67260 4398 67280
rect 4342 67224 4398 67260
rect 4618 67788 4674 67824
rect 4618 67768 4620 67788
rect 4620 67768 4672 67788
rect 4672 67768 4674 67788
rect 4526 67632 4582 67688
rect 5216 84346 5272 84348
rect 5296 84346 5352 84348
rect 5376 84346 5432 84348
rect 5456 84346 5512 84348
rect 5216 84294 5262 84346
rect 5262 84294 5272 84346
rect 5296 84294 5326 84346
rect 5326 84294 5338 84346
rect 5338 84294 5352 84346
rect 5376 84294 5390 84346
rect 5390 84294 5402 84346
rect 5402 84294 5432 84346
rect 5456 84294 5466 84346
rect 5466 84294 5512 84346
rect 5216 84292 5272 84294
rect 5296 84292 5352 84294
rect 5376 84292 5432 84294
rect 5456 84292 5512 84294
rect 5216 83258 5272 83260
rect 5296 83258 5352 83260
rect 5376 83258 5432 83260
rect 5456 83258 5512 83260
rect 5216 83206 5262 83258
rect 5262 83206 5272 83258
rect 5296 83206 5326 83258
rect 5326 83206 5338 83258
rect 5338 83206 5352 83258
rect 5376 83206 5390 83258
rect 5390 83206 5402 83258
rect 5402 83206 5432 83258
rect 5456 83206 5466 83258
rect 5466 83206 5512 83258
rect 5216 83204 5272 83206
rect 5296 83204 5352 83206
rect 5376 83204 5432 83206
rect 5456 83204 5512 83206
rect 5216 82170 5272 82172
rect 5296 82170 5352 82172
rect 5376 82170 5432 82172
rect 5456 82170 5512 82172
rect 5216 82118 5262 82170
rect 5262 82118 5272 82170
rect 5296 82118 5326 82170
rect 5326 82118 5338 82170
rect 5338 82118 5352 82170
rect 5376 82118 5390 82170
rect 5390 82118 5402 82170
rect 5402 82118 5432 82170
rect 5456 82118 5466 82170
rect 5466 82118 5512 82170
rect 5216 82116 5272 82118
rect 5296 82116 5352 82118
rect 5376 82116 5432 82118
rect 5456 82116 5512 82118
rect 5216 81082 5272 81084
rect 5296 81082 5352 81084
rect 5376 81082 5432 81084
rect 5456 81082 5512 81084
rect 5216 81030 5262 81082
rect 5262 81030 5272 81082
rect 5296 81030 5326 81082
rect 5326 81030 5338 81082
rect 5338 81030 5352 81082
rect 5376 81030 5390 81082
rect 5390 81030 5402 81082
rect 5402 81030 5432 81082
rect 5456 81030 5466 81082
rect 5466 81030 5512 81082
rect 5216 81028 5272 81030
rect 5296 81028 5352 81030
rect 5376 81028 5432 81030
rect 5456 81028 5512 81030
rect 5216 79994 5272 79996
rect 5296 79994 5352 79996
rect 5376 79994 5432 79996
rect 5456 79994 5512 79996
rect 5216 79942 5262 79994
rect 5262 79942 5272 79994
rect 5296 79942 5326 79994
rect 5326 79942 5338 79994
rect 5338 79942 5352 79994
rect 5376 79942 5390 79994
rect 5390 79942 5402 79994
rect 5402 79942 5432 79994
rect 5456 79942 5466 79994
rect 5466 79942 5512 79994
rect 5216 79940 5272 79942
rect 5296 79940 5352 79942
rect 5376 79940 5432 79942
rect 5456 79940 5512 79942
rect 5216 78906 5272 78908
rect 5296 78906 5352 78908
rect 5376 78906 5432 78908
rect 5456 78906 5512 78908
rect 5216 78854 5262 78906
rect 5262 78854 5272 78906
rect 5296 78854 5326 78906
rect 5326 78854 5338 78906
rect 5338 78854 5352 78906
rect 5376 78854 5390 78906
rect 5390 78854 5402 78906
rect 5402 78854 5432 78906
rect 5456 78854 5466 78906
rect 5466 78854 5512 78906
rect 5216 78852 5272 78854
rect 5296 78852 5352 78854
rect 5376 78852 5432 78854
rect 5456 78852 5512 78854
rect 5216 77818 5272 77820
rect 5296 77818 5352 77820
rect 5376 77818 5432 77820
rect 5456 77818 5512 77820
rect 5216 77766 5262 77818
rect 5262 77766 5272 77818
rect 5296 77766 5326 77818
rect 5326 77766 5338 77818
rect 5338 77766 5352 77818
rect 5376 77766 5390 77818
rect 5390 77766 5402 77818
rect 5402 77766 5432 77818
rect 5456 77766 5466 77818
rect 5466 77766 5512 77818
rect 5216 77764 5272 77766
rect 5296 77764 5352 77766
rect 5376 77764 5432 77766
rect 5456 77764 5512 77766
rect 5216 76730 5272 76732
rect 5296 76730 5352 76732
rect 5376 76730 5432 76732
rect 5456 76730 5512 76732
rect 5216 76678 5262 76730
rect 5262 76678 5272 76730
rect 5296 76678 5326 76730
rect 5326 76678 5338 76730
rect 5338 76678 5352 76730
rect 5376 76678 5390 76730
rect 5390 76678 5402 76730
rect 5402 76678 5432 76730
rect 5456 76678 5466 76730
rect 5466 76678 5512 76730
rect 5216 76676 5272 76678
rect 5296 76676 5352 76678
rect 5376 76676 5432 76678
rect 5456 76676 5512 76678
rect 5216 75642 5272 75644
rect 5296 75642 5352 75644
rect 5376 75642 5432 75644
rect 5456 75642 5512 75644
rect 5216 75590 5262 75642
rect 5262 75590 5272 75642
rect 5296 75590 5326 75642
rect 5326 75590 5338 75642
rect 5338 75590 5352 75642
rect 5376 75590 5390 75642
rect 5390 75590 5402 75642
rect 5402 75590 5432 75642
rect 5456 75590 5466 75642
rect 5466 75590 5512 75642
rect 5216 75588 5272 75590
rect 5296 75588 5352 75590
rect 5376 75588 5432 75590
rect 5456 75588 5512 75590
rect 5216 74554 5272 74556
rect 5296 74554 5352 74556
rect 5376 74554 5432 74556
rect 5456 74554 5512 74556
rect 5216 74502 5262 74554
rect 5262 74502 5272 74554
rect 5296 74502 5326 74554
rect 5326 74502 5338 74554
rect 5338 74502 5352 74554
rect 5376 74502 5390 74554
rect 5390 74502 5402 74554
rect 5402 74502 5432 74554
rect 5456 74502 5466 74554
rect 5466 74502 5512 74554
rect 5216 74500 5272 74502
rect 5296 74500 5352 74502
rect 5376 74500 5432 74502
rect 5456 74500 5512 74502
rect 5216 73466 5272 73468
rect 5296 73466 5352 73468
rect 5376 73466 5432 73468
rect 5456 73466 5512 73468
rect 5216 73414 5262 73466
rect 5262 73414 5272 73466
rect 5296 73414 5326 73466
rect 5326 73414 5338 73466
rect 5338 73414 5352 73466
rect 5376 73414 5390 73466
rect 5390 73414 5402 73466
rect 5402 73414 5432 73466
rect 5456 73414 5466 73466
rect 5466 73414 5512 73466
rect 5216 73412 5272 73414
rect 5296 73412 5352 73414
rect 5376 73412 5432 73414
rect 5456 73412 5512 73414
rect 5216 72378 5272 72380
rect 5296 72378 5352 72380
rect 5376 72378 5432 72380
rect 5456 72378 5512 72380
rect 5216 72326 5262 72378
rect 5262 72326 5272 72378
rect 5296 72326 5326 72378
rect 5326 72326 5338 72378
rect 5338 72326 5352 72378
rect 5376 72326 5390 72378
rect 5390 72326 5402 72378
rect 5402 72326 5432 72378
rect 5456 72326 5466 72378
rect 5466 72326 5512 72378
rect 5216 72324 5272 72326
rect 5296 72324 5352 72326
rect 5376 72324 5432 72326
rect 5456 72324 5512 72326
rect 6816 86522 6872 86524
rect 6896 86522 6952 86524
rect 6976 86522 7032 86524
rect 7056 86522 7112 86524
rect 6816 86470 6862 86522
rect 6862 86470 6872 86522
rect 6896 86470 6926 86522
rect 6926 86470 6938 86522
rect 6938 86470 6952 86522
rect 6976 86470 6990 86522
rect 6990 86470 7002 86522
rect 7002 86470 7032 86522
rect 7056 86470 7066 86522
rect 7066 86470 7112 86522
rect 6816 86468 6872 86470
rect 6896 86468 6952 86470
rect 6976 86468 7032 86470
rect 7056 86468 7112 86470
rect 8416 86522 8472 86524
rect 8496 86522 8552 86524
rect 8576 86522 8632 86524
rect 8656 86522 8712 86524
rect 8416 86470 8462 86522
rect 8462 86470 8472 86522
rect 8496 86470 8526 86522
rect 8526 86470 8538 86522
rect 8538 86470 8552 86522
rect 8576 86470 8590 86522
rect 8590 86470 8602 86522
rect 8602 86470 8632 86522
rect 8656 86470 8666 86522
rect 8666 86470 8712 86522
rect 8416 86468 8472 86470
rect 8496 86468 8552 86470
rect 8576 86468 8632 86470
rect 8656 86468 8712 86470
rect 5216 71290 5272 71292
rect 5296 71290 5352 71292
rect 5376 71290 5432 71292
rect 5456 71290 5512 71292
rect 5216 71238 5262 71290
rect 5262 71238 5272 71290
rect 5296 71238 5326 71290
rect 5326 71238 5338 71290
rect 5338 71238 5352 71290
rect 5376 71238 5390 71290
rect 5390 71238 5402 71290
rect 5402 71238 5432 71290
rect 5456 71238 5466 71290
rect 5466 71238 5512 71290
rect 5216 71236 5272 71238
rect 5296 71236 5352 71238
rect 5376 71236 5432 71238
rect 5456 71236 5512 71238
rect 5216 70202 5272 70204
rect 5296 70202 5352 70204
rect 5376 70202 5432 70204
rect 5456 70202 5512 70204
rect 5216 70150 5262 70202
rect 5262 70150 5272 70202
rect 5296 70150 5326 70202
rect 5326 70150 5338 70202
rect 5338 70150 5352 70202
rect 5376 70150 5390 70202
rect 5390 70150 5402 70202
rect 5402 70150 5432 70202
rect 5456 70150 5466 70202
rect 5466 70150 5512 70202
rect 5216 70148 5272 70150
rect 5296 70148 5352 70150
rect 5376 70148 5432 70150
rect 5456 70148 5512 70150
rect 5354 69944 5410 70000
rect 5354 69400 5410 69456
rect 5216 69114 5272 69116
rect 5296 69114 5352 69116
rect 5376 69114 5432 69116
rect 5456 69114 5512 69116
rect 5216 69062 5262 69114
rect 5262 69062 5272 69114
rect 5296 69062 5326 69114
rect 5326 69062 5338 69114
rect 5338 69062 5352 69114
rect 5376 69062 5390 69114
rect 5390 69062 5402 69114
rect 5402 69062 5432 69114
rect 5456 69062 5466 69114
rect 5466 69062 5512 69114
rect 5216 69060 5272 69062
rect 5296 69060 5352 69062
rect 5376 69060 5432 69062
rect 5456 69060 5512 69062
rect 4556 67482 4612 67484
rect 4636 67482 4692 67484
rect 4716 67482 4772 67484
rect 4796 67482 4852 67484
rect 4556 67430 4602 67482
rect 4602 67430 4612 67482
rect 4636 67430 4666 67482
rect 4666 67430 4678 67482
rect 4678 67430 4692 67482
rect 4716 67430 4730 67482
rect 4730 67430 4742 67482
rect 4742 67430 4772 67482
rect 4796 67430 4806 67482
rect 4806 67430 4852 67482
rect 4556 67428 4612 67430
rect 4636 67428 4692 67430
rect 4716 67428 4772 67430
rect 4796 67428 4852 67430
rect 4526 66700 4582 66736
rect 4526 66680 4528 66700
rect 4528 66680 4580 66700
rect 4580 66680 4582 66700
rect 4342 66408 4398 66464
rect 4710 66544 4766 66600
rect 4556 66394 4612 66396
rect 4636 66394 4692 66396
rect 4716 66394 4772 66396
rect 4796 66394 4852 66396
rect 4556 66342 4602 66394
rect 4602 66342 4612 66394
rect 4636 66342 4666 66394
rect 4666 66342 4678 66394
rect 4678 66342 4692 66394
rect 4716 66342 4730 66394
rect 4730 66342 4742 66394
rect 4742 66342 4772 66394
rect 4796 66342 4806 66394
rect 4806 66342 4852 66394
rect 4556 66340 4612 66342
rect 4636 66340 4692 66342
rect 4716 66340 4772 66342
rect 4796 66340 4852 66342
rect 4618 66136 4674 66192
rect 5722 72120 5778 72176
rect 5814 70488 5870 70544
rect 6156 85978 6212 85980
rect 6236 85978 6292 85980
rect 6316 85978 6372 85980
rect 6396 85978 6452 85980
rect 6156 85926 6202 85978
rect 6202 85926 6212 85978
rect 6236 85926 6266 85978
rect 6266 85926 6278 85978
rect 6278 85926 6292 85978
rect 6316 85926 6330 85978
rect 6330 85926 6342 85978
rect 6342 85926 6372 85978
rect 6396 85926 6406 85978
rect 6406 85926 6452 85978
rect 6156 85924 6212 85926
rect 6236 85924 6292 85926
rect 6316 85924 6372 85926
rect 6396 85924 6452 85926
rect 7756 85978 7812 85980
rect 7836 85978 7892 85980
rect 7916 85978 7972 85980
rect 7996 85978 8052 85980
rect 7756 85926 7802 85978
rect 7802 85926 7812 85978
rect 7836 85926 7866 85978
rect 7866 85926 7878 85978
rect 7878 85926 7892 85978
rect 7916 85926 7930 85978
rect 7930 85926 7942 85978
rect 7942 85926 7972 85978
rect 7996 85926 8006 85978
rect 8006 85926 8052 85978
rect 7756 85924 7812 85926
rect 7836 85924 7892 85926
rect 7916 85924 7972 85926
rect 7996 85924 8052 85926
rect 6816 85434 6872 85436
rect 6896 85434 6952 85436
rect 6976 85434 7032 85436
rect 7056 85434 7112 85436
rect 6816 85382 6862 85434
rect 6862 85382 6872 85434
rect 6896 85382 6926 85434
rect 6926 85382 6938 85434
rect 6938 85382 6952 85434
rect 6976 85382 6990 85434
rect 6990 85382 7002 85434
rect 7002 85382 7032 85434
rect 7056 85382 7066 85434
rect 7066 85382 7112 85434
rect 6816 85380 6872 85382
rect 6896 85380 6952 85382
rect 6976 85380 7032 85382
rect 7056 85380 7112 85382
rect 8416 85434 8472 85436
rect 8496 85434 8552 85436
rect 8576 85434 8632 85436
rect 8656 85434 8712 85436
rect 8416 85382 8462 85434
rect 8462 85382 8472 85434
rect 8496 85382 8526 85434
rect 8526 85382 8538 85434
rect 8538 85382 8552 85434
rect 8576 85382 8590 85434
rect 8590 85382 8602 85434
rect 8602 85382 8632 85434
rect 8656 85382 8666 85434
rect 8666 85382 8712 85434
rect 8416 85380 8472 85382
rect 8496 85380 8552 85382
rect 8576 85380 8632 85382
rect 8656 85380 8712 85382
rect 6156 84890 6212 84892
rect 6236 84890 6292 84892
rect 6316 84890 6372 84892
rect 6396 84890 6452 84892
rect 6156 84838 6202 84890
rect 6202 84838 6212 84890
rect 6236 84838 6266 84890
rect 6266 84838 6278 84890
rect 6278 84838 6292 84890
rect 6316 84838 6330 84890
rect 6330 84838 6342 84890
rect 6342 84838 6372 84890
rect 6396 84838 6406 84890
rect 6406 84838 6452 84890
rect 6156 84836 6212 84838
rect 6236 84836 6292 84838
rect 6316 84836 6372 84838
rect 6396 84836 6452 84838
rect 6156 83802 6212 83804
rect 6236 83802 6292 83804
rect 6316 83802 6372 83804
rect 6396 83802 6452 83804
rect 6156 83750 6202 83802
rect 6202 83750 6212 83802
rect 6236 83750 6266 83802
rect 6266 83750 6278 83802
rect 6278 83750 6292 83802
rect 6316 83750 6330 83802
rect 6330 83750 6342 83802
rect 6342 83750 6372 83802
rect 6396 83750 6406 83802
rect 6406 83750 6452 83802
rect 6156 83748 6212 83750
rect 6236 83748 6292 83750
rect 6316 83748 6372 83750
rect 6396 83748 6452 83750
rect 6156 82714 6212 82716
rect 6236 82714 6292 82716
rect 6316 82714 6372 82716
rect 6396 82714 6452 82716
rect 6156 82662 6202 82714
rect 6202 82662 6212 82714
rect 6236 82662 6266 82714
rect 6266 82662 6278 82714
rect 6278 82662 6292 82714
rect 6316 82662 6330 82714
rect 6330 82662 6342 82714
rect 6342 82662 6372 82714
rect 6396 82662 6406 82714
rect 6406 82662 6452 82714
rect 6156 82660 6212 82662
rect 6236 82660 6292 82662
rect 6316 82660 6372 82662
rect 6396 82660 6452 82662
rect 6156 81626 6212 81628
rect 6236 81626 6292 81628
rect 6316 81626 6372 81628
rect 6396 81626 6452 81628
rect 6156 81574 6202 81626
rect 6202 81574 6212 81626
rect 6236 81574 6266 81626
rect 6266 81574 6278 81626
rect 6278 81574 6292 81626
rect 6316 81574 6330 81626
rect 6330 81574 6342 81626
rect 6342 81574 6372 81626
rect 6396 81574 6406 81626
rect 6406 81574 6452 81626
rect 6156 81572 6212 81574
rect 6236 81572 6292 81574
rect 6316 81572 6372 81574
rect 6396 81572 6452 81574
rect 6156 80538 6212 80540
rect 6236 80538 6292 80540
rect 6316 80538 6372 80540
rect 6396 80538 6452 80540
rect 6156 80486 6202 80538
rect 6202 80486 6212 80538
rect 6236 80486 6266 80538
rect 6266 80486 6278 80538
rect 6278 80486 6292 80538
rect 6316 80486 6330 80538
rect 6330 80486 6342 80538
rect 6342 80486 6372 80538
rect 6396 80486 6406 80538
rect 6406 80486 6452 80538
rect 6156 80484 6212 80486
rect 6236 80484 6292 80486
rect 6316 80484 6372 80486
rect 6396 80484 6452 80486
rect 6156 79450 6212 79452
rect 6236 79450 6292 79452
rect 6316 79450 6372 79452
rect 6396 79450 6452 79452
rect 6156 79398 6202 79450
rect 6202 79398 6212 79450
rect 6236 79398 6266 79450
rect 6266 79398 6278 79450
rect 6278 79398 6292 79450
rect 6316 79398 6330 79450
rect 6330 79398 6342 79450
rect 6342 79398 6372 79450
rect 6396 79398 6406 79450
rect 6406 79398 6452 79450
rect 6156 79396 6212 79398
rect 6236 79396 6292 79398
rect 6316 79396 6372 79398
rect 6396 79396 6452 79398
rect 6156 78362 6212 78364
rect 6236 78362 6292 78364
rect 6316 78362 6372 78364
rect 6396 78362 6452 78364
rect 6156 78310 6202 78362
rect 6202 78310 6212 78362
rect 6236 78310 6266 78362
rect 6266 78310 6278 78362
rect 6278 78310 6292 78362
rect 6316 78310 6330 78362
rect 6330 78310 6342 78362
rect 6342 78310 6372 78362
rect 6396 78310 6406 78362
rect 6406 78310 6452 78362
rect 6156 78308 6212 78310
rect 6236 78308 6292 78310
rect 6316 78308 6372 78310
rect 6396 78308 6452 78310
rect 6156 77274 6212 77276
rect 6236 77274 6292 77276
rect 6316 77274 6372 77276
rect 6396 77274 6452 77276
rect 6156 77222 6202 77274
rect 6202 77222 6212 77274
rect 6236 77222 6266 77274
rect 6266 77222 6278 77274
rect 6278 77222 6292 77274
rect 6316 77222 6330 77274
rect 6330 77222 6342 77274
rect 6342 77222 6372 77274
rect 6396 77222 6406 77274
rect 6406 77222 6452 77274
rect 6156 77220 6212 77222
rect 6236 77220 6292 77222
rect 6316 77220 6372 77222
rect 6396 77220 6452 77222
rect 6156 76186 6212 76188
rect 6236 76186 6292 76188
rect 6316 76186 6372 76188
rect 6396 76186 6452 76188
rect 6156 76134 6202 76186
rect 6202 76134 6212 76186
rect 6236 76134 6266 76186
rect 6266 76134 6278 76186
rect 6278 76134 6292 76186
rect 6316 76134 6330 76186
rect 6330 76134 6342 76186
rect 6342 76134 6372 76186
rect 6396 76134 6406 76186
rect 6406 76134 6452 76186
rect 6156 76132 6212 76134
rect 6236 76132 6292 76134
rect 6316 76132 6372 76134
rect 6396 76132 6452 76134
rect 6156 75098 6212 75100
rect 6236 75098 6292 75100
rect 6316 75098 6372 75100
rect 6396 75098 6452 75100
rect 6156 75046 6202 75098
rect 6202 75046 6212 75098
rect 6236 75046 6266 75098
rect 6266 75046 6278 75098
rect 6278 75046 6292 75098
rect 6316 75046 6330 75098
rect 6330 75046 6342 75098
rect 6342 75046 6372 75098
rect 6396 75046 6406 75098
rect 6406 75046 6452 75098
rect 6156 75044 6212 75046
rect 6236 75044 6292 75046
rect 6316 75044 6372 75046
rect 6396 75044 6452 75046
rect 6156 74010 6212 74012
rect 6236 74010 6292 74012
rect 6316 74010 6372 74012
rect 6396 74010 6452 74012
rect 6156 73958 6202 74010
rect 6202 73958 6212 74010
rect 6236 73958 6266 74010
rect 6266 73958 6278 74010
rect 6278 73958 6292 74010
rect 6316 73958 6330 74010
rect 6330 73958 6342 74010
rect 6342 73958 6372 74010
rect 6396 73958 6406 74010
rect 6406 73958 6452 74010
rect 6156 73956 6212 73958
rect 6236 73956 6292 73958
rect 6316 73956 6372 73958
rect 6396 73956 6452 73958
rect 6156 72922 6212 72924
rect 6236 72922 6292 72924
rect 6316 72922 6372 72924
rect 6396 72922 6452 72924
rect 6156 72870 6202 72922
rect 6202 72870 6212 72922
rect 6236 72870 6266 72922
rect 6266 72870 6278 72922
rect 6278 72870 6292 72922
rect 6316 72870 6330 72922
rect 6330 72870 6342 72922
rect 6342 72870 6372 72922
rect 6396 72870 6406 72922
rect 6406 72870 6452 72922
rect 6156 72868 6212 72870
rect 6236 72868 6292 72870
rect 6316 72868 6372 72870
rect 6396 72868 6452 72870
rect 6274 72664 6330 72720
rect 6156 71834 6212 71836
rect 6236 71834 6292 71836
rect 6316 71834 6372 71836
rect 6396 71834 6452 71836
rect 6156 71782 6202 71834
rect 6202 71782 6212 71834
rect 6236 71782 6266 71834
rect 6266 71782 6278 71834
rect 6278 71782 6292 71834
rect 6316 71782 6330 71834
rect 6330 71782 6342 71834
rect 6342 71782 6372 71834
rect 6396 71782 6406 71834
rect 6406 71782 6452 71834
rect 6156 71780 6212 71782
rect 6236 71780 6292 71782
rect 6316 71780 6372 71782
rect 6396 71780 6452 71782
rect 6816 84346 6872 84348
rect 6896 84346 6952 84348
rect 6976 84346 7032 84348
rect 7056 84346 7112 84348
rect 6816 84294 6862 84346
rect 6862 84294 6872 84346
rect 6896 84294 6926 84346
rect 6926 84294 6938 84346
rect 6938 84294 6952 84346
rect 6976 84294 6990 84346
rect 6990 84294 7002 84346
rect 7002 84294 7032 84346
rect 7056 84294 7066 84346
rect 7066 84294 7112 84346
rect 6816 84292 6872 84294
rect 6896 84292 6952 84294
rect 6976 84292 7032 84294
rect 7056 84292 7112 84294
rect 6816 83258 6872 83260
rect 6896 83258 6952 83260
rect 6976 83258 7032 83260
rect 7056 83258 7112 83260
rect 6816 83206 6862 83258
rect 6862 83206 6872 83258
rect 6896 83206 6926 83258
rect 6926 83206 6938 83258
rect 6938 83206 6952 83258
rect 6976 83206 6990 83258
rect 6990 83206 7002 83258
rect 7002 83206 7032 83258
rect 7056 83206 7066 83258
rect 7066 83206 7112 83258
rect 6816 83204 6872 83206
rect 6896 83204 6952 83206
rect 6976 83204 7032 83206
rect 7056 83204 7112 83206
rect 6816 82170 6872 82172
rect 6896 82170 6952 82172
rect 6976 82170 7032 82172
rect 7056 82170 7112 82172
rect 6816 82118 6862 82170
rect 6862 82118 6872 82170
rect 6896 82118 6926 82170
rect 6926 82118 6938 82170
rect 6938 82118 6952 82170
rect 6976 82118 6990 82170
rect 6990 82118 7002 82170
rect 7002 82118 7032 82170
rect 7056 82118 7066 82170
rect 7066 82118 7112 82170
rect 6816 82116 6872 82118
rect 6896 82116 6952 82118
rect 6976 82116 7032 82118
rect 7056 82116 7112 82118
rect 6816 81082 6872 81084
rect 6896 81082 6952 81084
rect 6976 81082 7032 81084
rect 7056 81082 7112 81084
rect 6816 81030 6862 81082
rect 6862 81030 6872 81082
rect 6896 81030 6926 81082
rect 6926 81030 6938 81082
rect 6938 81030 6952 81082
rect 6976 81030 6990 81082
rect 6990 81030 7002 81082
rect 7002 81030 7032 81082
rect 7056 81030 7066 81082
rect 7066 81030 7112 81082
rect 6816 81028 6872 81030
rect 6896 81028 6952 81030
rect 6976 81028 7032 81030
rect 7056 81028 7112 81030
rect 6816 79994 6872 79996
rect 6896 79994 6952 79996
rect 6976 79994 7032 79996
rect 7056 79994 7112 79996
rect 6816 79942 6862 79994
rect 6862 79942 6872 79994
rect 6896 79942 6926 79994
rect 6926 79942 6938 79994
rect 6938 79942 6952 79994
rect 6976 79942 6990 79994
rect 6990 79942 7002 79994
rect 7002 79942 7032 79994
rect 7056 79942 7066 79994
rect 7066 79942 7112 79994
rect 6816 79940 6872 79942
rect 6896 79940 6952 79942
rect 6976 79940 7032 79942
rect 7056 79940 7112 79942
rect 6816 78906 6872 78908
rect 6896 78906 6952 78908
rect 6976 78906 7032 78908
rect 7056 78906 7112 78908
rect 6816 78854 6862 78906
rect 6862 78854 6872 78906
rect 6896 78854 6926 78906
rect 6926 78854 6938 78906
rect 6938 78854 6952 78906
rect 6976 78854 6990 78906
rect 6990 78854 7002 78906
rect 7002 78854 7032 78906
rect 7056 78854 7066 78906
rect 7066 78854 7112 78906
rect 6816 78852 6872 78854
rect 6896 78852 6952 78854
rect 6976 78852 7032 78854
rect 7056 78852 7112 78854
rect 6816 77818 6872 77820
rect 6896 77818 6952 77820
rect 6976 77818 7032 77820
rect 7056 77818 7112 77820
rect 6816 77766 6862 77818
rect 6862 77766 6872 77818
rect 6896 77766 6926 77818
rect 6926 77766 6938 77818
rect 6938 77766 6952 77818
rect 6976 77766 6990 77818
rect 6990 77766 7002 77818
rect 7002 77766 7032 77818
rect 7056 77766 7066 77818
rect 7066 77766 7112 77818
rect 6816 77764 6872 77766
rect 6896 77764 6952 77766
rect 6976 77764 7032 77766
rect 7056 77764 7112 77766
rect 6816 76730 6872 76732
rect 6896 76730 6952 76732
rect 6976 76730 7032 76732
rect 7056 76730 7112 76732
rect 6816 76678 6862 76730
rect 6862 76678 6872 76730
rect 6896 76678 6926 76730
rect 6926 76678 6938 76730
rect 6938 76678 6952 76730
rect 6976 76678 6990 76730
rect 6990 76678 7002 76730
rect 7002 76678 7032 76730
rect 7056 76678 7066 76730
rect 7066 76678 7112 76730
rect 6816 76676 6872 76678
rect 6896 76676 6952 76678
rect 6976 76676 7032 76678
rect 7056 76676 7112 76678
rect 6816 75642 6872 75644
rect 6896 75642 6952 75644
rect 6976 75642 7032 75644
rect 7056 75642 7112 75644
rect 6816 75590 6862 75642
rect 6862 75590 6872 75642
rect 6896 75590 6926 75642
rect 6926 75590 6938 75642
rect 6938 75590 6952 75642
rect 6976 75590 6990 75642
rect 6990 75590 7002 75642
rect 7002 75590 7032 75642
rect 7056 75590 7066 75642
rect 7066 75590 7112 75642
rect 6816 75588 6872 75590
rect 6896 75588 6952 75590
rect 6976 75588 7032 75590
rect 7056 75588 7112 75590
rect 6816 74554 6872 74556
rect 6896 74554 6952 74556
rect 6976 74554 7032 74556
rect 7056 74554 7112 74556
rect 6816 74502 6862 74554
rect 6862 74502 6872 74554
rect 6896 74502 6926 74554
rect 6926 74502 6938 74554
rect 6938 74502 6952 74554
rect 6976 74502 6990 74554
rect 6990 74502 7002 74554
rect 7002 74502 7032 74554
rect 7056 74502 7066 74554
rect 7066 74502 7112 74554
rect 6816 74500 6872 74502
rect 6896 74500 6952 74502
rect 6976 74500 7032 74502
rect 7056 74500 7112 74502
rect 7286 74568 7342 74624
rect 6816 73466 6872 73468
rect 6896 73466 6952 73468
rect 6976 73466 7032 73468
rect 7056 73466 7112 73468
rect 6816 73414 6862 73466
rect 6862 73414 6872 73466
rect 6896 73414 6926 73466
rect 6926 73414 6938 73466
rect 6938 73414 6952 73466
rect 6976 73414 6990 73466
rect 6990 73414 7002 73466
rect 7002 73414 7032 73466
rect 7056 73414 7066 73466
rect 7066 73414 7112 73466
rect 6816 73412 6872 73414
rect 6896 73412 6952 73414
rect 6976 73412 7032 73414
rect 7056 73412 7112 73414
rect 7010 73208 7066 73264
rect 6734 73072 6790 73128
rect 6826 72528 6882 72584
rect 7194 72800 7250 72856
rect 6816 72378 6872 72380
rect 6896 72378 6952 72380
rect 6976 72378 7032 72380
rect 7056 72378 7112 72380
rect 6816 72326 6862 72378
rect 6862 72326 6872 72378
rect 6896 72326 6926 72378
rect 6926 72326 6938 72378
rect 6938 72326 6952 72378
rect 6976 72326 6990 72378
rect 6990 72326 7002 72378
rect 7002 72326 7032 72378
rect 7056 72326 7066 72378
rect 7066 72326 7112 72378
rect 6816 72324 6872 72326
rect 6896 72324 6952 72326
rect 6976 72324 7032 72326
rect 7056 72324 7112 72326
rect 7756 84890 7812 84892
rect 7836 84890 7892 84892
rect 7916 84890 7972 84892
rect 7996 84890 8052 84892
rect 7756 84838 7802 84890
rect 7802 84838 7812 84890
rect 7836 84838 7866 84890
rect 7866 84838 7878 84890
rect 7878 84838 7892 84890
rect 7916 84838 7930 84890
rect 7930 84838 7942 84890
rect 7942 84838 7972 84890
rect 7996 84838 8006 84890
rect 8006 84838 8052 84890
rect 7756 84836 7812 84838
rect 7836 84836 7892 84838
rect 7916 84836 7972 84838
rect 7996 84836 8052 84838
rect 7756 83802 7812 83804
rect 7836 83802 7892 83804
rect 7916 83802 7972 83804
rect 7996 83802 8052 83804
rect 7756 83750 7802 83802
rect 7802 83750 7812 83802
rect 7836 83750 7866 83802
rect 7866 83750 7878 83802
rect 7878 83750 7892 83802
rect 7916 83750 7930 83802
rect 7930 83750 7942 83802
rect 7942 83750 7972 83802
rect 7996 83750 8006 83802
rect 8006 83750 8052 83802
rect 7756 83748 7812 83750
rect 7836 83748 7892 83750
rect 7916 83748 7972 83750
rect 7996 83748 8052 83750
rect 7756 82714 7812 82716
rect 7836 82714 7892 82716
rect 7916 82714 7972 82716
rect 7996 82714 8052 82716
rect 7756 82662 7802 82714
rect 7802 82662 7812 82714
rect 7836 82662 7866 82714
rect 7866 82662 7878 82714
rect 7878 82662 7892 82714
rect 7916 82662 7930 82714
rect 7930 82662 7942 82714
rect 7942 82662 7972 82714
rect 7996 82662 8006 82714
rect 8006 82662 8052 82714
rect 7756 82660 7812 82662
rect 7836 82660 7892 82662
rect 7916 82660 7972 82662
rect 7996 82660 8052 82662
rect 7756 81626 7812 81628
rect 7836 81626 7892 81628
rect 7916 81626 7972 81628
rect 7996 81626 8052 81628
rect 7756 81574 7802 81626
rect 7802 81574 7812 81626
rect 7836 81574 7866 81626
rect 7866 81574 7878 81626
rect 7878 81574 7892 81626
rect 7916 81574 7930 81626
rect 7930 81574 7942 81626
rect 7942 81574 7972 81626
rect 7996 81574 8006 81626
rect 8006 81574 8052 81626
rect 7756 81572 7812 81574
rect 7836 81572 7892 81574
rect 7916 81572 7972 81574
rect 7996 81572 8052 81574
rect 7756 80538 7812 80540
rect 7836 80538 7892 80540
rect 7916 80538 7972 80540
rect 7996 80538 8052 80540
rect 7756 80486 7802 80538
rect 7802 80486 7812 80538
rect 7836 80486 7866 80538
rect 7866 80486 7878 80538
rect 7878 80486 7892 80538
rect 7916 80486 7930 80538
rect 7930 80486 7942 80538
rect 7942 80486 7972 80538
rect 7996 80486 8006 80538
rect 8006 80486 8052 80538
rect 7756 80484 7812 80486
rect 7836 80484 7892 80486
rect 7916 80484 7972 80486
rect 7996 80484 8052 80486
rect 7756 79450 7812 79452
rect 7836 79450 7892 79452
rect 7916 79450 7972 79452
rect 7996 79450 8052 79452
rect 7756 79398 7802 79450
rect 7802 79398 7812 79450
rect 7836 79398 7866 79450
rect 7866 79398 7878 79450
rect 7878 79398 7892 79450
rect 7916 79398 7930 79450
rect 7930 79398 7942 79450
rect 7942 79398 7972 79450
rect 7996 79398 8006 79450
rect 8006 79398 8052 79450
rect 7756 79396 7812 79398
rect 7836 79396 7892 79398
rect 7916 79396 7972 79398
rect 7996 79396 8052 79398
rect 7756 78362 7812 78364
rect 7836 78362 7892 78364
rect 7916 78362 7972 78364
rect 7996 78362 8052 78364
rect 7756 78310 7802 78362
rect 7802 78310 7812 78362
rect 7836 78310 7866 78362
rect 7866 78310 7878 78362
rect 7878 78310 7892 78362
rect 7916 78310 7930 78362
rect 7930 78310 7942 78362
rect 7942 78310 7972 78362
rect 7996 78310 8006 78362
rect 8006 78310 8052 78362
rect 7756 78308 7812 78310
rect 7836 78308 7892 78310
rect 7916 78308 7972 78310
rect 7996 78308 8052 78310
rect 7756 77274 7812 77276
rect 7836 77274 7892 77276
rect 7916 77274 7972 77276
rect 7996 77274 8052 77276
rect 7756 77222 7802 77274
rect 7802 77222 7812 77274
rect 7836 77222 7866 77274
rect 7866 77222 7878 77274
rect 7878 77222 7892 77274
rect 7916 77222 7930 77274
rect 7930 77222 7942 77274
rect 7942 77222 7972 77274
rect 7996 77222 8006 77274
rect 8006 77222 8052 77274
rect 7756 77220 7812 77222
rect 7836 77220 7892 77222
rect 7916 77220 7972 77222
rect 7996 77220 8052 77222
rect 7470 73480 7526 73536
rect 7756 76186 7812 76188
rect 7836 76186 7892 76188
rect 7916 76186 7972 76188
rect 7996 76186 8052 76188
rect 7756 76134 7802 76186
rect 7802 76134 7812 76186
rect 7836 76134 7866 76186
rect 7866 76134 7878 76186
rect 7878 76134 7892 76186
rect 7916 76134 7930 76186
rect 7930 76134 7942 76186
rect 7942 76134 7972 76186
rect 7996 76134 8006 76186
rect 8006 76134 8052 76186
rect 7756 76132 7812 76134
rect 7836 76132 7892 76134
rect 7916 76132 7972 76134
rect 7996 76132 8052 76134
rect 7756 75098 7812 75100
rect 7836 75098 7892 75100
rect 7916 75098 7972 75100
rect 7996 75098 8052 75100
rect 7756 75046 7802 75098
rect 7802 75046 7812 75098
rect 7836 75046 7866 75098
rect 7866 75046 7878 75098
rect 7878 75046 7892 75098
rect 7916 75046 7930 75098
rect 7930 75046 7942 75098
rect 7942 75046 7972 75098
rect 7996 75046 8006 75098
rect 8006 75046 8052 75098
rect 7756 75044 7812 75046
rect 7836 75044 7892 75046
rect 7916 75044 7972 75046
rect 7996 75044 8052 75046
rect 7756 74010 7812 74012
rect 7836 74010 7892 74012
rect 7916 74010 7972 74012
rect 7996 74010 8052 74012
rect 7756 73958 7802 74010
rect 7802 73958 7812 74010
rect 7836 73958 7866 74010
rect 7866 73958 7878 74010
rect 7878 73958 7892 74010
rect 7916 73958 7930 74010
rect 7930 73958 7942 74010
rect 7942 73958 7972 74010
rect 7996 73958 8006 74010
rect 8006 73958 8052 74010
rect 7756 73956 7812 73958
rect 7836 73956 7892 73958
rect 7916 73956 7972 73958
rect 7996 73956 8052 73958
rect 8416 84346 8472 84348
rect 8496 84346 8552 84348
rect 8576 84346 8632 84348
rect 8656 84346 8712 84348
rect 8416 84294 8462 84346
rect 8462 84294 8472 84346
rect 8496 84294 8526 84346
rect 8526 84294 8538 84346
rect 8538 84294 8552 84346
rect 8576 84294 8590 84346
rect 8590 84294 8602 84346
rect 8602 84294 8632 84346
rect 8656 84294 8666 84346
rect 8666 84294 8712 84346
rect 8416 84292 8472 84294
rect 8496 84292 8552 84294
rect 8576 84292 8632 84294
rect 8656 84292 8712 84294
rect 8416 83258 8472 83260
rect 8496 83258 8552 83260
rect 8576 83258 8632 83260
rect 8656 83258 8712 83260
rect 8416 83206 8462 83258
rect 8462 83206 8472 83258
rect 8496 83206 8526 83258
rect 8526 83206 8538 83258
rect 8538 83206 8552 83258
rect 8576 83206 8590 83258
rect 8590 83206 8602 83258
rect 8602 83206 8632 83258
rect 8656 83206 8666 83258
rect 8666 83206 8712 83258
rect 8416 83204 8472 83206
rect 8496 83204 8552 83206
rect 8576 83204 8632 83206
rect 8656 83204 8712 83206
rect 8416 82170 8472 82172
rect 8496 82170 8552 82172
rect 8576 82170 8632 82172
rect 8656 82170 8712 82172
rect 8416 82118 8462 82170
rect 8462 82118 8472 82170
rect 8496 82118 8526 82170
rect 8526 82118 8538 82170
rect 8538 82118 8552 82170
rect 8576 82118 8590 82170
rect 8590 82118 8602 82170
rect 8602 82118 8632 82170
rect 8656 82118 8666 82170
rect 8666 82118 8712 82170
rect 8416 82116 8472 82118
rect 8496 82116 8552 82118
rect 8576 82116 8632 82118
rect 8656 82116 8712 82118
rect 8416 81082 8472 81084
rect 8496 81082 8552 81084
rect 8576 81082 8632 81084
rect 8656 81082 8712 81084
rect 8416 81030 8462 81082
rect 8462 81030 8472 81082
rect 8496 81030 8526 81082
rect 8526 81030 8538 81082
rect 8538 81030 8552 81082
rect 8576 81030 8590 81082
rect 8590 81030 8602 81082
rect 8602 81030 8632 81082
rect 8656 81030 8666 81082
rect 8666 81030 8712 81082
rect 8416 81028 8472 81030
rect 8496 81028 8552 81030
rect 8576 81028 8632 81030
rect 8656 81028 8712 81030
rect 8416 79994 8472 79996
rect 8496 79994 8552 79996
rect 8576 79994 8632 79996
rect 8656 79994 8712 79996
rect 8416 79942 8462 79994
rect 8462 79942 8472 79994
rect 8496 79942 8526 79994
rect 8526 79942 8538 79994
rect 8538 79942 8552 79994
rect 8576 79942 8590 79994
rect 8590 79942 8602 79994
rect 8602 79942 8632 79994
rect 8656 79942 8666 79994
rect 8666 79942 8712 79994
rect 8416 79940 8472 79942
rect 8496 79940 8552 79942
rect 8576 79940 8632 79942
rect 8656 79940 8712 79942
rect 8416 78906 8472 78908
rect 8496 78906 8552 78908
rect 8576 78906 8632 78908
rect 8656 78906 8712 78908
rect 8416 78854 8462 78906
rect 8462 78854 8472 78906
rect 8496 78854 8526 78906
rect 8526 78854 8538 78906
rect 8538 78854 8552 78906
rect 8576 78854 8590 78906
rect 8590 78854 8602 78906
rect 8602 78854 8632 78906
rect 8656 78854 8666 78906
rect 8666 78854 8712 78906
rect 8416 78852 8472 78854
rect 8496 78852 8552 78854
rect 8576 78852 8632 78854
rect 8656 78852 8712 78854
rect 8416 77818 8472 77820
rect 8496 77818 8552 77820
rect 8576 77818 8632 77820
rect 8656 77818 8712 77820
rect 8416 77766 8462 77818
rect 8462 77766 8472 77818
rect 8496 77766 8526 77818
rect 8526 77766 8538 77818
rect 8538 77766 8552 77818
rect 8576 77766 8590 77818
rect 8590 77766 8602 77818
rect 8602 77766 8632 77818
rect 8656 77766 8666 77818
rect 8666 77766 8712 77818
rect 8416 77764 8472 77766
rect 8496 77764 8552 77766
rect 8576 77764 8632 77766
rect 8656 77764 8712 77766
rect 8416 76730 8472 76732
rect 8496 76730 8552 76732
rect 8576 76730 8632 76732
rect 8656 76730 8712 76732
rect 8416 76678 8462 76730
rect 8462 76678 8472 76730
rect 8496 76678 8526 76730
rect 8526 76678 8538 76730
rect 8538 76678 8552 76730
rect 8576 76678 8590 76730
rect 8590 76678 8602 76730
rect 8602 76678 8632 76730
rect 8656 76678 8666 76730
rect 8666 76678 8712 76730
rect 8416 76676 8472 76678
rect 8496 76676 8552 76678
rect 8576 76676 8632 76678
rect 8656 76676 8712 76678
rect 10016 86522 10072 86524
rect 10096 86522 10152 86524
rect 10176 86522 10232 86524
rect 10256 86522 10312 86524
rect 10016 86470 10062 86522
rect 10062 86470 10072 86522
rect 10096 86470 10126 86522
rect 10126 86470 10138 86522
rect 10138 86470 10152 86522
rect 10176 86470 10190 86522
rect 10190 86470 10202 86522
rect 10202 86470 10232 86522
rect 10256 86470 10266 86522
rect 10266 86470 10312 86522
rect 10016 86468 10072 86470
rect 10096 86468 10152 86470
rect 10176 86468 10232 86470
rect 10256 86468 10312 86470
rect 9356 85978 9412 85980
rect 9436 85978 9492 85980
rect 9516 85978 9572 85980
rect 9596 85978 9652 85980
rect 9356 85926 9402 85978
rect 9402 85926 9412 85978
rect 9436 85926 9466 85978
rect 9466 85926 9478 85978
rect 9478 85926 9492 85978
rect 9516 85926 9530 85978
rect 9530 85926 9542 85978
rect 9542 85926 9572 85978
rect 9596 85926 9606 85978
rect 9606 85926 9652 85978
rect 9356 85924 9412 85926
rect 9436 85924 9492 85926
rect 9516 85924 9572 85926
rect 9596 85924 9652 85926
rect 8416 75642 8472 75644
rect 8496 75642 8552 75644
rect 8576 75642 8632 75644
rect 8656 75642 8712 75644
rect 8416 75590 8462 75642
rect 8462 75590 8472 75642
rect 8496 75590 8526 75642
rect 8526 75590 8538 75642
rect 8538 75590 8552 75642
rect 8576 75590 8590 75642
rect 8590 75590 8602 75642
rect 8602 75590 8632 75642
rect 8656 75590 8666 75642
rect 8666 75590 8712 75642
rect 8416 75588 8472 75590
rect 8496 75588 8552 75590
rect 8576 75588 8632 75590
rect 8656 75588 8712 75590
rect 8416 74554 8472 74556
rect 8496 74554 8552 74556
rect 8576 74554 8632 74556
rect 8656 74554 8712 74556
rect 8416 74502 8462 74554
rect 8462 74502 8472 74554
rect 8496 74502 8526 74554
rect 8526 74502 8538 74554
rect 8538 74502 8552 74554
rect 8576 74502 8590 74554
rect 8590 74502 8602 74554
rect 8602 74502 8632 74554
rect 8656 74502 8666 74554
rect 8666 74502 8712 74554
rect 8416 74500 8472 74502
rect 8496 74500 8552 74502
rect 8576 74500 8632 74502
rect 8656 74500 8712 74502
rect 7746 73480 7802 73536
rect 8206 73480 8262 73536
rect 8114 73208 8170 73264
rect 7756 72922 7812 72924
rect 7836 72922 7892 72924
rect 7916 72922 7972 72924
rect 7996 72922 8052 72924
rect 7756 72870 7802 72922
rect 7802 72870 7812 72922
rect 7836 72870 7866 72922
rect 7866 72870 7878 72922
rect 7878 72870 7892 72922
rect 7916 72870 7930 72922
rect 7930 72870 7942 72922
rect 7942 72870 7972 72922
rect 7996 72870 8006 72922
rect 8006 72870 8052 72922
rect 7756 72868 7812 72870
rect 7836 72868 7892 72870
rect 7916 72868 7972 72870
rect 7996 72868 8052 72870
rect 7562 72800 7618 72856
rect 6826 71984 6882 72040
rect 7194 72140 7250 72176
rect 7194 72120 7196 72140
rect 7196 72120 7248 72140
rect 7248 72120 7250 72140
rect 6550 70932 6552 70952
rect 6552 70932 6604 70952
rect 6604 70932 6606 70952
rect 6550 70896 6606 70932
rect 6156 70746 6212 70748
rect 6236 70746 6292 70748
rect 6316 70746 6372 70748
rect 6396 70746 6452 70748
rect 6156 70694 6202 70746
rect 6202 70694 6212 70746
rect 6236 70694 6266 70746
rect 6266 70694 6278 70746
rect 6278 70694 6292 70746
rect 6316 70694 6330 70746
rect 6330 70694 6342 70746
rect 6342 70694 6372 70746
rect 6396 70694 6406 70746
rect 6406 70694 6452 70746
rect 6156 70692 6212 70694
rect 6236 70692 6292 70694
rect 6316 70692 6372 70694
rect 6396 70692 6452 70694
rect 5722 68720 5778 68776
rect 5216 68026 5272 68028
rect 5296 68026 5352 68028
rect 5376 68026 5432 68028
rect 5456 68026 5512 68028
rect 5216 67974 5262 68026
rect 5262 67974 5272 68026
rect 5296 67974 5326 68026
rect 5326 67974 5338 68026
rect 5338 67974 5352 68026
rect 5376 67974 5390 68026
rect 5390 67974 5402 68026
rect 5402 67974 5432 68026
rect 5456 67974 5466 68026
rect 5466 67974 5512 68026
rect 5216 67972 5272 67974
rect 5296 67972 5352 67974
rect 5376 67972 5432 67974
rect 5456 67972 5512 67974
rect 5354 67088 5410 67144
rect 5216 66938 5272 66940
rect 5296 66938 5352 66940
rect 5376 66938 5432 66940
rect 5456 66938 5512 66940
rect 5216 66886 5262 66938
rect 5262 66886 5272 66938
rect 5296 66886 5326 66938
rect 5326 66886 5338 66938
rect 5338 66886 5352 66938
rect 5376 66886 5390 66938
rect 5390 66886 5402 66938
rect 5402 66886 5432 66938
rect 5456 66886 5466 66938
rect 5466 66886 5512 66938
rect 5216 66884 5272 66886
rect 5296 66884 5352 66886
rect 5376 66884 5432 66886
rect 5456 66884 5512 66886
rect 5906 68720 5962 68776
rect 6156 69658 6212 69660
rect 6236 69658 6292 69660
rect 6316 69658 6372 69660
rect 6396 69658 6452 69660
rect 6156 69606 6202 69658
rect 6202 69606 6212 69658
rect 6236 69606 6266 69658
rect 6266 69606 6278 69658
rect 6278 69606 6292 69658
rect 6316 69606 6330 69658
rect 6330 69606 6342 69658
rect 6342 69606 6372 69658
rect 6396 69606 6406 69658
rect 6406 69606 6452 69658
rect 6156 69604 6212 69606
rect 6236 69604 6292 69606
rect 6316 69604 6372 69606
rect 6396 69604 6452 69606
rect 6816 71290 6872 71292
rect 6896 71290 6952 71292
rect 6976 71290 7032 71292
rect 7056 71290 7112 71292
rect 6816 71238 6862 71290
rect 6862 71238 6872 71290
rect 6896 71238 6926 71290
rect 6926 71238 6938 71290
rect 6938 71238 6952 71290
rect 6976 71238 6990 71290
rect 6990 71238 7002 71290
rect 7002 71238 7032 71290
rect 7056 71238 7066 71290
rect 7066 71238 7112 71290
rect 6816 71236 6872 71238
rect 6896 71236 6952 71238
rect 6976 71236 7032 71238
rect 7056 71236 7112 71238
rect 6918 70508 6974 70544
rect 6918 70488 6920 70508
rect 6920 70488 6972 70508
rect 6972 70488 6974 70508
rect 6816 70202 6872 70204
rect 6896 70202 6952 70204
rect 6976 70202 7032 70204
rect 7056 70202 7112 70204
rect 6816 70150 6862 70202
rect 6862 70150 6872 70202
rect 6896 70150 6926 70202
rect 6926 70150 6938 70202
rect 6938 70150 6952 70202
rect 6976 70150 6990 70202
rect 6990 70150 7002 70202
rect 7002 70150 7032 70202
rect 7056 70150 7066 70202
rect 7066 70150 7112 70202
rect 6816 70148 6872 70150
rect 6896 70148 6952 70150
rect 6976 70148 7032 70150
rect 7056 70148 7112 70150
rect 6816 69114 6872 69116
rect 6896 69114 6952 69116
rect 6976 69114 7032 69116
rect 7056 69114 7112 69116
rect 6816 69062 6862 69114
rect 6862 69062 6872 69114
rect 6896 69062 6926 69114
rect 6926 69062 6938 69114
rect 6938 69062 6952 69114
rect 6976 69062 6990 69114
rect 6990 69062 7002 69114
rect 7002 69062 7032 69114
rect 7056 69062 7066 69114
rect 7066 69062 7112 69114
rect 6816 69060 6872 69062
rect 6896 69060 6952 69062
rect 6976 69060 7032 69062
rect 7056 69060 7112 69062
rect 6156 68570 6212 68572
rect 6236 68570 6292 68572
rect 6316 68570 6372 68572
rect 6396 68570 6452 68572
rect 6156 68518 6202 68570
rect 6202 68518 6212 68570
rect 6236 68518 6266 68570
rect 6266 68518 6278 68570
rect 6278 68518 6292 68570
rect 6316 68518 6330 68570
rect 6330 68518 6342 68570
rect 6342 68518 6372 68570
rect 6396 68518 6406 68570
rect 6406 68518 6452 68570
rect 6156 68516 6212 68518
rect 6236 68516 6292 68518
rect 6316 68516 6372 68518
rect 6396 68516 6452 68518
rect 6090 68312 6146 68368
rect 6182 67632 6238 67688
rect 6918 68176 6974 68232
rect 6816 68026 6872 68028
rect 6896 68026 6952 68028
rect 6976 68026 7032 68028
rect 7056 68026 7112 68028
rect 6816 67974 6862 68026
rect 6862 67974 6872 68026
rect 6896 67974 6926 68026
rect 6926 67974 6938 68026
rect 6938 67974 6952 68026
rect 6976 67974 6990 68026
rect 6990 67974 7002 68026
rect 7002 67974 7032 68026
rect 7056 67974 7066 68026
rect 7066 67974 7112 68026
rect 6816 67972 6872 67974
rect 6896 67972 6952 67974
rect 6976 67972 7032 67974
rect 7056 67972 7112 67974
rect 6156 67482 6212 67484
rect 6236 67482 6292 67484
rect 6316 67482 6372 67484
rect 6396 67482 6452 67484
rect 6156 67430 6202 67482
rect 6202 67430 6212 67482
rect 6236 67430 6266 67482
rect 6266 67430 6278 67482
rect 6278 67430 6292 67482
rect 6316 67430 6330 67482
rect 6330 67430 6342 67482
rect 6342 67430 6372 67482
rect 6396 67430 6406 67482
rect 6406 67430 6452 67482
rect 6156 67428 6212 67430
rect 6236 67428 6292 67430
rect 6316 67428 6372 67430
rect 6396 67428 6452 67430
rect 5216 65850 5272 65852
rect 5296 65850 5352 65852
rect 5376 65850 5432 65852
rect 5456 65850 5512 65852
rect 5216 65798 5262 65850
rect 5262 65798 5272 65850
rect 5296 65798 5326 65850
rect 5326 65798 5338 65850
rect 5338 65798 5352 65850
rect 5376 65798 5390 65850
rect 5390 65798 5402 65850
rect 5402 65798 5432 65850
rect 5456 65798 5466 65850
rect 5466 65798 5512 65850
rect 5216 65796 5272 65798
rect 5296 65796 5352 65798
rect 5376 65796 5432 65798
rect 5456 65796 5512 65798
rect 5354 65592 5410 65648
rect 4556 65306 4612 65308
rect 4636 65306 4692 65308
rect 4716 65306 4772 65308
rect 4796 65306 4852 65308
rect 4556 65254 4602 65306
rect 4602 65254 4612 65306
rect 4636 65254 4666 65306
rect 4666 65254 4678 65306
rect 4678 65254 4692 65306
rect 4716 65254 4730 65306
rect 4730 65254 4742 65306
rect 4742 65254 4772 65306
rect 4796 65254 4806 65306
rect 4806 65254 4852 65306
rect 4556 65252 4612 65254
rect 4636 65252 4692 65254
rect 4716 65252 4772 65254
rect 4796 65252 4852 65254
rect 4556 64218 4612 64220
rect 4636 64218 4692 64220
rect 4716 64218 4772 64220
rect 4796 64218 4852 64220
rect 4556 64166 4602 64218
rect 4602 64166 4612 64218
rect 4636 64166 4666 64218
rect 4666 64166 4678 64218
rect 4678 64166 4692 64218
rect 4716 64166 4730 64218
rect 4730 64166 4742 64218
rect 4742 64166 4772 64218
rect 4796 64166 4806 64218
rect 4806 64166 4852 64218
rect 4556 64164 4612 64166
rect 4636 64164 4692 64166
rect 4716 64164 4772 64166
rect 4796 64164 4852 64166
rect 4556 63130 4612 63132
rect 4636 63130 4692 63132
rect 4716 63130 4772 63132
rect 4796 63130 4852 63132
rect 4556 63078 4602 63130
rect 4602 63078 4612 63130
rect 4636 63078 4666 63130
rect 4666 63078 4678 63130
rect 4678 63078 4692 63130
rect 4716 63078 4730 63130
rect 4730 63078 4742 63130
rect 4742 63078 4772 63130
rect 4796 63078 4806 63130
rect 4806 63078 4852 63130
rect 4556 63076 4612 63078
rect 4636 63076 4692 63078
rect 4716 63076 4772 63078
rect 4796 63076 4852 63078
rect 4556 62042 4612 62044
rect 4636 62042 4692 62044
rect 4716 62042 4772 62044
rect 4796 62042 4852 62044
rect 4556 61990 4602 62042
rect 4602 61990 4612 62042
rect 4636 61990 4666 62042
rect 4666 61990 4678 62042
rect 4678 61990 4692 62042
rect 4716 61990 4730 62042
rect 4730 61990 4742 62042
rect 4742 61990 4772 62042
rect 4796 61990 4806 62042
rect 4806 61990 4852 62042
rect 4556 61988 4612 61990
rect 4636 61988 4692 61990
rect 4716 61988 4772 61990
rect 4796 61988 4852 61990
rect 4556 60954 4612 60956
rect 4636 60954 4692 60956
rect 4716 60954 4772 60956
rect 4796 60954 4852 60956
rect 4556 60902 4602 60954
rect 4602 60902 4612 60954
rect 4636 60902 4666 60954
rect 4666 60902 4678 60954
rect 4678 60902 4692 60954
rect 4716 60902 4730 60954
rect 4730 60902 4742 60954
rect 4742 60902 4772 60954
rect 4796 60902 4806 60954
rect 4806 60902 4852 60954
rect 4556 60900 4612 60902
rect 4636 60900 4692 60902
rect 4716 60900 4772 60902
rect 4796 60900 4852 60902
rect 5216 64762 5272 64764
rect 5296 64762 5352 64764
rect 5376 64762 5432 64764
rect 5456 64762 5512 64764
rect 5216 64710 5262 64762
rect 5262 64710 5272 64762
rect 5296 64710 5326 64762
rect 5326 64710 5338 64762
rect 5338 64710 5352 64762
rect 5376 64710 5390 64762
rect 5390 64710 5402 64762
rect 5402 64710 5432 64762
rect 5456 64710 5466 64762
rect 5466 64710 5512 64762
rect 5216 64708 5272 64710
rect 5296 64708 5352 64710
rect 5376 64708 5432 64710
rect 5456 64708 5512 64710
rect 5216 63674 5272 63676
rect 5296 63674 5352 63676
rect 5376 63674 5432 63676
rect 5456 63674 5512 63676
rect 5216 63622 5262 63674
rect 5262 63622 5272 63674
rect 5296 63622 5326 63674
rect 5326 63622 5338 63674
rect 5338 63622 5352 63674
rect 5376 63622 5390 63674
rect 5390 63622 5402 63674
rect 5402 63622 5432 63674
rect 5456 63622 5466 63674
rect 5466 63622 5512 63674
rect 5216 63620 5272 63622
rect 5296 63620 5352 63622
rect 5376 63620 5432 63622
rect 5456 63620 5512 63622
rect 5216 62586 5272 62588
rect 5296 62586 5352 62588
rect 5376 62586 5432 62588
rect 5456 62586 5512 62588
rect 5216 62534 5262 62586
rect 5262 62534 5272 62586
rect 5296 62534 5326 62586
rect 5326 62534 5338 62586
rect 5338 62534 5352 62586
rect 5376 62534 5390 62586
rect 5390 62534 5402 62586
rect 5402 62534 5432 62586
rect 5456 62534 5466 62586
rect 5466 62534 5512 62586
rect 5216 62532 5272 62534
rect 5296 62532 5352 62534
rect 5376 62532 5432 62534
rect 5456 62532 5512 62534
rect 5216 61498 5272 61500
rect 5296 61498 5352 61500
rect 5376 61498 5432 61500
rect 5456 61498 5512 61500
rect 5216 61446 5262 61498
rect 5262 61446 5272 61498
rect 5296 61446 5326 61498
rect 5326 61446 5338 61498
rect 5338 61446 5352 61498
rect 5376 61446 5390 61498
rect 5390 61446 5402 61498
rect 5402 61446 5432 61498
rect 5456 61446 5466 61498
rect 5466 61446 5512 61498
rect 5216 61444 5272 61446
rect 5296 61444 5352 61446
rect 5376 61444 5432 61446
rect 5456 61444 5512 61446
rect 4556 59866 4612 59868
rect 4636 59866 4692 59868
rect 4716 59866 4772 59868
rect 4796 59866 4852 59868
rect 4556 59814 4602 59866
rect 4602 59814 4612 59866
rect 4636 59814 4666 59866
rect 4666 59814 4678 59866
rect 4678 59814 4692 59866
rect 4716 59814 4730 59866
rect 4730 59814 4742 59866
rect 4742 59814 4772 59866
rect 4796 59814 4806 59866
rect 4806 59814 4852 59866
rect 4556 59812 4612 59814
rect 4636 59812 4692 59814
rect 4716 59812 4772 59814
rect 4796 59812 4852 59814
rect 4556 58778 4612 58780
rect 4636 58778 4692 58780
rect 4716 58778 4772 58780
rect 4796 58778 4852 58780
rect 4556 58726 4602 58778
rect 4602 58726 4612 58778
rect 4636 58726 4666 58778
rect 4666 58726 4678 58778
rect 4678 58726 4692 58778
rect 4716 58726 4730 58778
rect 4730 58726 4742 58778
rect 4742 58726 4772 58778
rect 4796 58726 4806 58778
rect 4806 58726 4852 58778
rect 4556 58724 4612 58726
rect 4636 58724 4692 58726
rect 4716 58724 4772 58726
rect 4796 58724 4852 58726
rect 4556 57690 4612 57692
rect 4636 57690 4692 57692
rect 4716 57690 4772 57692
rect 4796 57690 4852 57692
rect 4556 57638 4602 57690
rect 4602 57638 4612 57690
rect 4636 57638 4666 57690
rect 4666 57638 4678 57690
rect 4678 57638 4692 57690
rect 4716 57638 4730 57690
rect 4730 57638 4742 57690
rect 4742 57638 4772 57690
rect 4796 57638 4806 57690
rect 4806 57638 4852 57690
rect 4556 57636 4612 57638
rect 4636 57636 4692 57638
rect 4716 57636 4772 57638
rect 4796 57636 4852 57638
rect 4158 54168 4214 54224
rect 4556 56602 4612 56604
rect 4636 56602 4692 56604
rect 4716 56602 4772 56604
rect 4796 56602 4852 56604
rect 4556 56550 4602 56602
rect 4602 56550 4612 56602
rect 4636 56550 4666 56602
rect 4666 56550 4678 56602
rect 4678 56550 4692 56602
rect 4716 56550 4730 56602
rect 4730 56550 4742 56602
rect 4742 56550 4772 56602
rect 4796 56550 4806 56602
rect 4806 56550 4852 56602
rect 4556 56548 4612 56550
rect 4636 56548 4692 56550
rect 4716 56548 4772 56550
rect 4796 56548 4852 56550
rect 4556 55514 4612 55516
rect 4636 55514 4692 55516
rect 4716 55514 4772 55516
rect 4796 55514 4852 55516
rect 4556 55462 4602 55514
rect 4602 55462 4612 55514
rect 4636 55462 4666 55514
rect 4666 55462 4678 55514
rect 4678 55462 4692 55514
rect 4716 55462 4730 55514
rect 4730 55462 4742 55514
rect 4742 55462 4772 55514
rect 4796 55462 4806 55514
rect 4806 55462 4852 55514
rect 4556 55460 4612 55462
rect 4636 55460 4692 55462
rect 4716 55460 4772 55462
rect 4796 55460 4852 55462
rect 4556 54426 4612 54428
rect 4636 54426 4692 54428
rect 4716 54426 4772 54428
rect 4796 54426 4852 54428
rect 4556 54374 4602 54426
rect 4602 54374 4612 54426
rect 4636 54374 4666 54426
rect 4666 54374 4678 54426
rect 4678 54374 4692 54426
rect 4716 54374 4730 54426
rect 4730 54374 4742 54426
rect 4742 54374 4772 54426
rect 4796 54374 4806 54426
rect 4806 54374 4852 54426
rect 4556 54372 4612 54374
rect 4636 54372 4692 54374
rect 4716 54372 4772 54374
rect 4796 54372 4852 54374
rect 5216 60410 5272 60412
rect 5296 60410 5352 60412
rect 5376 60410 5432 60412
rect 5456 60410 5512 60412
rect 5216 60358 5262 60410
rect 5262 60358 5272 60410
rect 5296 60358 5326 60410
rect 5326 60358 5338 60410
rect 5338 60358 5352 60410
rect 5376 60358 5390 60410
rect 5390 60358 5402 60410
rect 5402 60358 5432 60410
rect 5456 60358 5466 60410
rect 5466 60358 5512 60410
rect 5216 60356 5272 60358
rect 5296 60356 5352 60358
rect 5376 60356 5432 60358
rect 5456 60356 5512 60358
rect 5216 59322 5272 59324
rect 5296 59322 5352 59324
rect 5376 59322 5432 59324
rect 5456 59322 5512 59324
rect 5216 59270 5262 59322
rect 5262 59270 5272 59322
rect 5296 59270 5326 59322
rect 5326 59270 5338 59322
rect 5338 59270 5352 59322
rect 5376 59270 5390 59322
rect 5390 59270 5402 59322
rect 5402 59270 5432 59322
rect 5456 59270 5466 59322
rect 5466 59270 5512 59322
rect 5216 59268 5272 59270
rect 5296 59268 5352 59270
rect 5376 59268 5432 59270
rect 5456 59268 5512 59270
rect 5216 58234 5272 58236
rect 5296 58234 5352 58236
rect 5376 58234 5432 58236
rect 5456 58234 5512 58236
rect 5216 58182 5262 58234
rect 5262 58182 5272 58234
rect 5296 58182 5326 58234
rect 5326 58182 5338 58234
rect 5338 58182 5352 58234
rect 5376 58182 5390 58234
rect 5390 58182 5402 58234
rect 5402 58182 5432 58234
rect 5456 58182 5466 58234
rect 5466 58182 5512 58234
rect 5216 58180 5272 58182
rect 5296 58180 5352 58182
rect 5376 58180 5432 58182
rect 5456 58180 5512 58182
rect 6156 66394 6212 66396
rect 6236 66394 6292 66396
rect 6316 66394 6372 66396
rect 6396 66394 6452 66396
rect 6156 66342 6202 66394
rect 6202 66342 6212 66394
rect 6236 66342 6266 66394
rect 6266 66342 6278 66394
rect 6278 66342 6292 66394
rect 6316 66342 6330 66394
rect 6330 66342 6342 66394
rect 6342 66342 6372 66394
rect 6396 66342 6406 66394
rect 6406 66342 6452 66394
rect 6156 66340 6212 66342
rect 6236 66340 6292 66342
rect 6316 66340 6372 66342
rect 6396 66340 6452 66342
rect 6156 65306 6212 65308
rect 6236 65306 6292 65308
rect 6316 65306 6372 65308
rect 6396 65306 6452 65308
rect 6156 65254 6202 65306
rect 6202 65254 6212 65306
rect 6236 65254 6266 65306
rect 6266 65254 6278 65306
rect 6278 65254 6292 65306
rect 6316 65254 6330 65306
rect 6330 65254 6342 65306
rect 6342 65254 6372 65306
rect 6396 65254 6406 65306
rect 6406 65254 6452 65306
rect 6156 65252 6212 65254
rect 6236 65252 6292 65254
rect 6316 65252 6372 65254
rect 6396 65252 6452 65254
rect 6156 64218 6212 64220
rect 6236 64218 6292 64220
rect 6316 64218 6372 64220
rect 6396 64218 6452 64220
rect 6156 64166 6202 64218
rect 6202 64166 6212 64218
rect 6236 64166 6266 64218
rect 6266 64166 6278 64218
rect 6278 64166 6292 64218
rect 6316 64166 6330 64218
rect 6330 64166 6342 64218
rect 6342 64166 6372 64218
rect 6396 64166 6406 64218
rect 6406 64166 6452 64218
rect 6156 64164 6212 64166
rect 6236 64164 6292 64166
rect 6316 64164 6372 64166
rect 6396 64164 6452 64166
rect 5216 57146 5272 57148
rect 5296 57146 5352 57148
rect 5376 57146 5432 57148
rect 5456 57146 5512 57148
rect 5216 57094 5262 57146
rect 5262 57094 5272 57146
rect 5296 57094 5326 57146
rect 5326 57094 5338 57146
rect 5338 57094 5352 57146
rect 5376 57094 5390 57146
rect 5390 57094 5402 57146
rect 5402 57094 5432 57146
rect 5456 57094 5466 57146
rect 5466 57094 5512 57146
rect 5216 57092 5272 57094
rect 5296 57092 5352 57094
rect 5376 57092 5432 57094
rect 5456 57092 5512 57094
rect 4556 53338 4612 53340
rect 4636 53338 4692 53340
rect 4716 53338 4772 53340
rect 4796 53338 4852 53340
rect 4556 53286 4602 53338
rect 4602 53286 4612 53338
rect 4636 53286 4666 53338
rect 4666 53286 4678 53338
rect 4678 53286 4692 53338
rect 4716 53286 4730 53338
rect 4730 53286 4742 53338
rect 4742 53286 4772 53338
rect 4796 53286 4806 53338
rect 4806 53286 4852 53338
rect 4556 53284 4612 53286
rect 4636 53284 4692 53286
rect 4716 53284 4772 53286
rect 4796 53284 4852 53286
rect 4556 52250 4612 52252
rect 4636 52250 4692 52252
rect 4716 52250 4772 52252
rect 4796 52250 4852 52252
rect 4556 52198 4602 52250
rect 4602 52198 4612 52250
rect 4636 52198 4666 52250
rect 4666 52198 4678 52250
rect 4678 52198 4692 52250
rect 4716 52198 4730 52250
rect 4730 52198 4742 52250
rect 4742 52198 4772 52250
rect 4796 52198 4806 52250
rect 4806 52198 4852 52250
rect 4556 52196 4612 52198
rect 4636 52196 4692 52198
rect 4716 52196 4772 52198
rect 4796 52196 4852 52198
rect 5216 56058 5272 56060
rect 5296 56058 5352 56060
rect 5376 56058 5432 56060
rect 5456 56058 5512 56060
rect 5216 56006 5262 56058
rect 5262 56006 5272 56058
rect 5296 56006 5326 56058
rect 5326 56006 5338 56058
rect 5338 56006 5352 56058
rect 5376 56006 5390 56058
rect 5390 56006 5402 56058
rect 5402 56006 5432 56058
rect 5456 56006 5466 56058
rect 5466 56006 5512 56058
rect 5216 56004 5272 56006
rect 5296 56004 5352 56006
rect 5376 56004 5432 56006
rect 5456 56004 5512 56006
rect 5216 54970 5272 54972
rect 5296 54970 5352 54972
rect 5376 54970 5432 54972
rect 5456 54970 5512 54972
rect 5216 54918 5262 54970
rect 5262 54918 5272 54970
rect 5296 54918 5326 54970
rect 5326 54918 5338 54970
rect 5338 54918 5352 54970
rect 5376 54918 5390 54970
rect 5390 54918 5402 54970
rect 5402 54918 5432 54970
rect 5456 54918 5466 54970
rect 5466 54918 5512 54970
rect 5216 54916 5272 54918
rect 5296 54916 5352 54918
rect 5376 54916 5432 54918
rect 5456 54916 5512 54918
rect 5216 53882 5272 53884
rect 5296 53882 5352 53884
rect 5376 53882 5432 53884
rect 5456 53882 5512 53884
rect 5216 53830 5262 53882
rect 5262 53830 5272 53882
rect 5296 53830 5326 53882
rect 5326 53830 5338 53882
rect 5338 53830 5352 53882
rect 5376 53830 5390 53882
rect 5390 53830 5402 53882
rect 5402 53830 5432 53882
rect 5456 53830 5466 53882
rect 5466 53830 5512 53882
rect 5216 53828 5272 53830
rect 5296 53828 5352 53830
rect 5376 53828 5432 53830
rect 5456 53828 5512 53830
rect 4556 51162 4612 51164
rect 4636 51162 4692 51164
rect 4716 51162 4772 51164
rect 4796 51162 4852 51164
rect 4556 51110 4602 51162
rect 4602 51110 4612 51162
rect 4636 51110 4666 51162
rect 4666 51110 4678 51162
rect 4678 51110 4692 51162
rect 4716 51110 4730 51162
rect 4730 51110 4742 51162
rect 4742 51110 4772 51162
rect 4796 51110 4806 51162
rect 4806 51110 4852 51162
rect 4556 51108 4612 51110
rect 4636 51108 4692 51110
rect 4716 51108 4772 51110
rect 4796 51108 4852 51110
rect 4556 50074 4612 50076
rect 4636 50074 4692 50076
rect 4716 50074 4772 50076
rect 4796 50074 4852 50076
rect 4556 50022 4602 50074
rect 4602 50022 4612 50074
rect 4636 50022 4666 50074
rect 4666 50022 4678 50074
rect 4678 50022 4692 50074
rect 4716 50022 4730 50074
rect 4730 50022 4742 50074
rect 4742 50022 4772 50074
rect 4796 50022 4806 50074
rect 4806 50022 4852 50074
rect 4556 50020 4612 50022
rect 4636 50020 4692 50022
rect 4716 50020 4772 50022
rect 4796 50020 4852 50022
rect 5216 52794 5272 52796
rect 5296 52794 5352 52796
rect 5376 52794 5432 52796
rect 5456 52794 5512 52796
rect 5216 52742 5262 52794
rect 5262 52742 5272 52794
rect 5296 52742 5326 52794
rect 5326 52742 5338 52794
rect 5338 52742 5352 52794
rect 5376 52742 5390 52794
rect 5390 52742 5402 52794
rect 5402 52742 5432 52794
rect 5456 52742 5466 52794
rect 5466 52742 5512 52794
rect 5216 52740 5272 52742
rect 5296 52740 5352 52742
rect 5376 52740 5432 52742
rect 5456 52740 5512 52742
rect 5216 51706 5272 51708
rect 5296 51706 5352 51708
rect 5376 51706 5432 51708
rect 5456 51706 5512 51708
rect 5216 51654 5262 51706
rect 5262 51654 5272 51706
rect 5296 51654 5326 51706
rect 5326 51654 5338 51706
rect 5338 51654 5352 51706
rect 5376 51654 5390 51706
rect 5390 51654 5402 51706
rect 5402 51654 5432 51706
rect 5456 51654 5466 51706
rect 5466 51654 5512 51706
rect 5216 51652 5272 51654
rect 5296 51652 5352 51654
rect 5376 51652 5432 51654
rect 5456 51652 5512 51654
rect 6550 63280 6606 63336
rect 6156 63130 6212 63132
rect 6236 63130 6292 63132
rect 6316 63130 6372 63132
rect 6396 63130 6452 63132
rect 6156 63078 6202 63130
rect 6202 63078 6212 63130
rect 6236 63078 6266 63130
rect 6266 63078 6278 63130
rect 6278 63078 6292 63130
rect 6316 63078 6330 63130
rect 6330 63078 6342 63130
rect 6342 63078 6372 63130
rect 6396 63078 6406 63130
rect 6406 63078 6452 63130
rect 6156 63076 6212 63078
rect 6236 63076 6292 63078
rect 6316 63076 6372 63078
rect 6396 63076 6452 63078
rect 5216 50618 5272 50620
rect 5296 50618 5352 50620
rect 5376 50618 5432 50620
rect 5456 50618 5512 50620
rect 5216 50566 5262 50618
rect 5262 50566 5272 50618
rect 5296 50566 5326 50618
rect 5326 50566 5338 50618
rect 5338 50566 5352 50618
rect 5376 50566 5390 50618
rect 5390 50566 5402 50618
rect 5402 50566 5432 50618
rect 5456 50566 5466 50618
rect 5466 50566 5512 50618
rect 5216 50564 5272 50566
rect 5296 50564 5352 50566
rect 5376 50564 5432 50566
rect 5456 50564 5512 50566
rect 4556 48986 4612 48988
rect 4636 48986 4692 48988
rect 4716 48986 4772 48988
rect 4796 48986 4852 48988
rect 4556 48934 4602 48986
rect 4602 48934 4612 48986
rect 4636 48934 4666 48986
rect 4666 48934 4678 48986
rect 4678 48934 4692 48986
rect 4716 48934 4730 48986
rect 4730 48934 4742 48986
rect 4742 48934 4772 48986
rect 4796 48934 4806 48986
rect 4806 48934 4852 48986
rect 4556 48932 4612 48934
rect 4636 48932 4692 48934
rect 4716 48932 4772 48934
rect 4796 48932 4852 48934
rect 4556 47898 4612 47900
rect 4636 47898 4692 47900
rect 4716 47898 4772 47900
rect 4796 47898 4852 47900
rect 4556 47846 4602 47898
rect 4602 47846 4612 47898
rect 4636 47846 4666 47898
rect 4666 47846 4678 47898
rect 4678 47846 4692 47898
rect 4716 47846 4730 47898
rect 4730 47846 4742 47898
rect 4742 47846 4772 47898
rect 4796 47846 4806 47898
rect 4806 47846 4852 47898
rect 4556 47844 4612 47846
rect 4636 47844 4692 47846
rect 4716 47844 4772 47846
rect 4796 47844 4852 47846
rect 4434 46960 4490 47016
rect 4556 46810 4612 46812
rect 4636 46810 4692 46812
rect 4716 46810 4772 46812
rect 4796 46810 4852 46812
rect 4556 46758 4602 46810
rect 4602 46758 4612 46810
rect 4636 46758 4666 46810
rect 4666 46758 4678 46810
rect 4678 46758 4692 46810
rect 4716 46758 4730 46810
rect 4730 46758 4742 46810
rect 4742 46758 4772 46810
rect 4796 46758 4806 46810
rect 4806 46758 4852 46810
rect 4556 46756 4612 46758
rect 4636 46756 4692 46758
rect 4716 46756 4772 46758
rect 4796 46756 4852 46758
rect 4434 46552 4490 46608
rect 4066 45464 4122 45520
rect 3974 44920 4030 44976
rect 3616 44090 3672 44092
rect 3696 44090 3752 44092
rect 3776 44090 3832 44092
rect 3856 44090 3912 44092
rect 3616 44038 3662 44090
rect 3662 44038 3672 44090
rect 3696 44038 3726 44090
rect 3726 44038 3738 44090
rect 3738 44038 3752 44090
rect 3776 44038 3790 44090
rect 3790 44038 3802 44090
rect 3802 44038 3832 44090
rect 3856 44038 3866 44090
rect 3866 44038 3912 44090
rect 3616 44036 3672 44038
rect 3696 44036 3752 44038
rect 3776 44036 3832 44038
rect 3856 44036 3912 44038
rect 3616 43002 3672 43004
rect 3696 43002 3752 43004
rect 3776 43002 3832 43004
rect 3856 43002 3912 43004
rect 3616 42950 3662 43002
rect 3662 42950 3672 43002
rect 3696 42950 3726 43002
rect 3726 42950 3738 43002
rect 3738 42950 3752 43002
rect 3776 42950 3790 43002
rect 3790 42950 3802 43002
rect 3802 42950 3832 43002
rect 3856 42950 3866 43002
rect 3866 42950 3912 43002
rect 3616 42948 3672 42950
rect 3696 42948 3752 42950
rect 3776 42948 3832 42950
rect 3856 42948 3912 42950
rect 3616 41914 3672 41916
rect 3696 41914 3752 41916
rect 3776 41914 3832 41916
rect 3856 41914 3912 41916
rect 3616 41862 3662 41914
rect 3662 41862 3672 41914
rect 3696 41862 3726 41914
rect 3726 41862 3738 41914
rect 3738 41862 3752 41914
rect 3776 41862 3790 41914
rect 3790 41862 3802 41914
rect 3802 41862 3832 41914
rect 3856 41862 3866 41914
rect 3866 41862 3912 41914
rect 3616 41860 3672 41862
rect 3696 41860 3752 41862
rect 3776 41860 3832 41862
rect 3856 41860 3912 41862
rect 3616 40826 3672 40828
rect 3696 40826 3752 40828
rect 3776 40826 3832 40828
rect 3856 40826 3912 40828
rect 3616 40774 3662 40826
rect 3662 40774 3672 40826
rect 3696 40774 3726 40826
rect 3726 40774 3738 40826
rect 3738 40774 3752 40826
rect 3776 40774 3790 40826
rect 3790 40774 3802 40826
rect 3802 40774 3832 40826
rect 3856 40774 3866 40826
rect 3866 40774 3912 40826
rect 3616 40772 3672 40774
rect 3696 40772 3752 40774
rect 3776 40772 3832 40774
rect 3856 40772 3912 40774
rect 3616 39738 3672 39740
rect 3696 39738 3752 39740
rect 3776 39738 3832 39740
rect 3856 39738 3912 39740
rect 3616 39686 3662 39738
rect 3662 39686 3672 39738
rect 3696 39686 3726 39738
rect 3726 39686 3738 39738
rect 3738 39686 3752 39738
rect 3776 39686 3790 39738
rect 3790 39686 3802 39738
rect 3802 39686 3832 39738
rect 3856 39686 3866 39738
rect 3866 39686 3912 39738
rect 3616 39684 3672 39686
rect 3696 39684 3752 39686
rect 3776 39684 3832 39686
rect 3856 39684 3912 39686
rect 3616 38650 3672 38652
rect 3696 38650 3752 38652
rect 3776 38650 3832 38652
rect 3856 38650 3912 38652
rect 3616 38598 3662 38650
rect 3662 38598 3672 38650
rect 3696 38598 3726 38650
rect 3726 38598 3738 38650
rect 3738 38598 3752 38650
rect 3776 38598 3790 38650
rect 3790 38598 3802 38650
rect 3802 38598 3832 38650
rect 3856 38598 3866 38650
rect 3866 38598 3912 38650
rect 3616 38596 3672 38598
rect 3696 38596 3752 38598
rect 3776 38596 3832 38598
rect 3856 38596 3912 38598
rect 3616 37562 3672 37564
rect 3696 37562 3752 37564
rect 3776 37562 3832 37564
rect 3856 37562 3912 37564
rect 3616 37510 3662 37562
rect 3662 37510 3672 37562
rect 3696 37510 3726 37562
rect 3726 37510 3738 37562
rect 3738 37510 3752 37562
rect 3776 37510 3790 37562
rect 3790 37510 3802 37562
rect 3802 37510 3832 37562
rect 3856 37510 3866 37562
rect 3866 37510 3912 37562
rect 3616 37508 3672 37510
rect 3696 37508 3752 37510
rect 3776 37508 3832 37510
rect 3856 37508 3912 37510
rect 3616 36474 3672 36476
rect 3696 36474 3752 36476
rect 3776 36474 3832 36476
rect 3856 36474 3912 36476
rect 3616 36422 3662 36474
rect 3662 36422 3672 36474
rect 3696 36422 3726 36474
rect 3726 36422 3738 36474
rect 3738 36422 3752 36474
rect 3776 36422 3790 36474
rect 3790 36422 3802 36474
rect 3802 36422 3832 36474
rect 3856 36422 3866 36474
rect 3866 36422 3912 36474
rect 3616 36420 3672 36422
rect 3696 36420 3752 36422
rect 3776 36420 3832 36422
rect 3856 36420 3912 36422
rect 3616 35386 3672 35388
rect 3696 35386 3752 35388
rect 3776 35386 3832 35388
rect 3856 35386 3912 35388
rect 3616 35334 3662 35386
rect 3662 35334 3672 35386
rect 3696 35334 3726 35386
rect 3726 35334 3738 35386
rect 3738 35334 3752 35386
rect 3776 35334 3790 35386
rect 3790 35334 3802 35386
rect 3802 35334 3832 35386
rect 3856 35334 3866 35386
rect 3866 35334 3912 35386
rect 3616 35332 3672 35334
rect 3696 35332 3752 35334
rect 3776 35332 3832 35334
rect 3856 35332 3912 35334
rect 3616 34298 3672 34300
rect 3696 34298 3752 34300
rect 3776 34298 3832 34300
rect 3856 34298 3912 34300
rect 3616 34246 3662 34298
rect 3662 34246 3672 34298
rect 3696 34246 3726 34298
rect 3726 34246 3738 34298
rect 3738 34246 3752 34298
rect 3776 34246 3790 34298
rect 3790 34246 3802 34298
rect 3802 34246 3832 34298
rect 3856 34246 3866 34298
rect 3866 34246 3912 34298
rect 3616 34244 3672 34246
rect 3696 34244 3752 34246
rect 3776 34244 3832 34246
rect 3856 34244 3912 34246
rect 3616 33210 3672 33212
rect 3696 33210 3752 33212
rect 3776 33210 3832 33212
rect 3856 33210 3912 33212
rect 3616 33158 3662 33210
rect 3662 33158 3672 33210
rect 3696 33158 3726 33210
rect 3726 33158 3738 33210
rect 3738 33158 3752 33210
rect 3776 33158 3790 33210
rect 3790 33158 3802 33210
rect 3802 33158 3832 33210
rect 3856 33158 3866 33210
rect 3866 33158 3912 33210
rect 3616 33156 3672 33158
rect 3696 33156 3752 33158
rect 3776 33156 3832 33158
rect 3856 33156 3912 33158
rect 3616 32122 3672 32124
rect 3696 32122 3752 32124
rect 3776 32122 3832 32124
rect 3856 32122 3912 32124
rect 3616 32070 3662 32122
rect 3662 32070 3672 32122
rect 3696 32070 3726 32122
rect 3726 32070 3738 32122
rect 3738 32070 3752 32122
rect 3776 32070 3790 32122
rect 3790 32070 3802 32122
rect 3802 32070 3832 32122
rect 3856 32070 3866 32122
rect 3866 32070 3912 32122
rect 3616 32068 3672 32070
rect 3696 32068 3752 32070
rect 3776 32068 3832 32070
rect 3856 32068 3912 32070
rect 3616 31034 3672 31036
rect 3696 31034 3752 31036
rect 3776 31034 3832 31036
rect 3856 31034 3912 31036
rect 3616 30982 3662 31034
rect 3662 30982 3672 31034
rect 3696 30982 3726 31034
rect 3726 30982 3738 31034
rect 3738 30982 3752 31034
rect 3776 30982 3790 31034
rect 3790 30982 3802 31034
rect 3802 30982 3832 31034
rect 3856 30982 3866 31034
rect 3866 30982 3912 31034
rect 3616 30980 3672 30982
rect 3696 30980 3752 30982
rect 3776 30980 3832 30982
rect 3856 30980 3912 30982
rect 3616 29946 3672 29948
rect 3696 29946 3752 29948
rect 3776 29946 3832 29948
rect 3856 29946 3912 29948
rect 3616 29894 3662 29946
rect 3662 29894 3672 29946
rect 3696 29894 3726 29946
rect 3726 29894 3738 29946
rect 3738 29894 3752 29946
rect 3776 29894 3790 29946
rect 3790 29894 3802 29946
rect 3802 29894 3832 29946
rect 3856 29894 3866 29946
rect 3866 29894 3912 29946
rect 3616 29892 3672 29894
rect 3696 29892 3752 29894
rect 3776 29892 3832 29894
rect 3856 29892 3912 29894
rect 3616 28858 3672 28860
rect 3696 28858 3752 28860
rect 3776 28858 3832 28860
rect 3856 28858 3912 28860
rect 3616 28806 3662 28858
rect 3662 28806 3672 28858
rect 3696 28806 3726 28858
rect 3726 28806 3738 28858
rect 3738 28806 3752 28858
rect 3776 28806 3790 28858
rect 3790 28806 3802 28858
rect 3802 28806 3832 28858
rect 3856 28806 3866 28858
rect 3866 28806 3912 28858
rect 3616 28804 3672 28806
rect 3696 28804 3752 28806
rect 3776 28804 3832 28806
rect 3856 28804 3912 28806
rect 3616 27770 3672 27772
rect 3696 27770 3752 27772
rect 3776 27770 3832 27772
rect 3856 27770 3912 27772
rect 3616 27718 3662 27770
rect 3662 27718 3672 27770
rect 3696 27718 3726 27770
rect 3726 27718 3738 27770
rect 3738 27718 3752 27770
rect 3776 27718 3790 27770
rect 3790 27718 3802 27770
rect 3802 27718 3832 27770
rect 3856 27718 3866 27770
rect 3866 27718 3912 27770
rect 3616 27716 3672 27718
rect 3696 27716 3752 27718
rect 3776 27716 3832 27718
rect 3856 27716 3912 27718
rect 3616 26682 3672 26684
rect 3696 26682 3752 26684
rect 3776 26682 3832 26684
rect 3856 26682 3912 26684
rect 3616 26630 3662 26682
rect 3662 26630 3672 26682
rect 3696 26630 3726 26682
rect 3726 26630 3738 26682
rect 3738 26630 3752 26682
rect 3776 26630 3790 26682
rect 3790 26630 3802 26682
rect 3802 26630 3832 26682
rect 3856 26630 3866 26682
rect 3866 26630 3912 26682
rect 3616 26628 3672 26630
rect 3696 26628 3752 26630
rect 3776 26628 3832 26630
rect 3856 26628 3912 26630
rect 4066 42200 4122 42256
rect 3616 25594 3672 25596
rect 3696 25594 3752 25596
rect 3776 25594 3832 25596
rect 3856 25594 3912 25596
rect 3616 25542 3662 25594
rect 3662 25542 3672 25594
rect 3696 25542 3726 25594
rect 3726 25542 3738 25594
rect 3738 25542 3752 25594
rect 3776 25542 3790 25594
rect 3790 25542 3802 25594
rect 3802 25542 3832 25594
rect 3856 25542 3866 25594
rect 3866 25542 3912 25594
rect 3616 25540 3672 25542
rect 3696 25540 3752 25542
rect 3776 25540 3832 25542
rect 3856 25540 3912 25542
rect 3616 24506 3672 24508
rect 3696 24506 3752 24508
rect 3776 24506 3832 24508
rect 3856 24506 3912 24508
rect 3616 24454 3662 24506
rect 3662 24454 3672 24506
rect 3696 24454 3726 24506
rect 3726 24454 3738 24506
rect 3738 24454 3752 24506
rect 3776 24454 3790 24506
rect 3790 24454 3802 24506
rect 3802 24454 3832 24506
rect 3856 24454 3866 24506
rect 3866 24454 3912 24506
rect 3616 24452 3672 24454
rect 3696 24452 3752 24454
rect 3776 24452 3832 24454
rect 3856 24452 3912 24454
rect 3616 23418 3672 23420
rect 3696 23418 3752 23420
rect 3776 23418 3832 23420
rect 3856 23418 3912 23420
rect 3616 23366 3662 23418
rect 3662 23366 3672 23418
rect 3696 23366 3726 23418
rect 3726 23366 3738 23418
rect 3738 23366 3752 23418
rect 3776 23366 3790 23418
rect 3790 23366 3802 23418
rect 3802 23366 3832 23418
rect 3856 23366 3866 23418
rect 3866 23366 3912 23418
rect 3616 23364 3672 23366
rect 3696 23364 3752 23366
rect 3776 23364 3832 23366
rect 3856 23364 3912 23366
rect 3616 22330 3672 22332
rect 3696 22330 3752 22332
rect 3776 22330 3832 22332
rect 3856 22330 3912 22332
rect 3616 22278 3662 22330
rect 3662 22278 3672 22330
rect 3696 22278 3726 22330
rect 3726 22278 3738 22330
rect 3738 22278 3752 22330
rect 3776 22278 3790 22330
rect 3790 22278 3802 22330
rect 3802 22278 3832 22330
rect 3856 22278 3866 22330
rect 3866 22278 3912 22330
rect 3616 22276 3672 22278
rect 3696 22276 3752 22278
rect 3776 22276 3832 22278
rect 3856 22276 3912 22278
rect 3616 21242 3672 21244
rect 3696 21242 3752 21244
rect 3776 21242 3832 21244
rect 3856 21242 3912 21244
rect 3616 21190 3662 21242
rect 3662 21190 3672 21242
rect 3696 21190 3726 21242
rect 3726 21190 3738 21242
rect 3738 21190 3752 21242
rect 3776 21190 3790 21242
rect 3790 21190 3802 21242
rect 3802 21190 3832 21242
rect 3856 21190 3866 21242
rect 3866 21190 3912 21242
rect 3616 21188 3672 21190
rect 3696 21188 3752 21190
rect 3776 21188 3832 21190
rect 3856 21188 3912 21190
rect 3616 20154 3672 20156
rect 3696 20154 3752 20156
rect 3776 20154 3832 20156
rect 3856 20154 3912 20156
rect 3616 20102 3662 20154
rect 3662 20102 3672 20154
rect 3696 20102 3726 20154
rect 3726 20102 3738 20154
rect 3738 20102 3752 20154
rect 3776 20102 3790 20154
rect 3790 20102 3802 20154
rect 3802 20102 3832 20154
rect 3856 20102 3866 20154
rect 3866 20102 3912 20154
rect 3616 20100 3672 20102
rect 3696 20100 3752 20102
rect 3776 20100 3832 20102
rect 3856 20100 3912 20102
rect 3616 19066 3672 19068
rect 3696 19066 3752 19068
rect 3776 19066 3832 19068
rect 3856 19066 3912 19068
rect 3616 19014 3662 19066
rect 3662 19014 3672 19066
rect 3696 19014 3726 19066
rect 3726 19014 3738 19066
rect 3738 19014 3752 19066
rect 3776 19014 3790 19066
rect 3790 19014 3802 19066
rect 3802 19014 3832 19066
rect 3856 19014 3866 19066
rect 3866 19014 3912 19066
rect 3616 19012 3672 19014
rect 3696 19012 3752 19014
rect 3776 19012 3832 19014
rect 3856 19012 3912 19014
rect 3616 17978 3672 17980
rect 3696 17978 3752 17980
rect 3776 17978 3832 17980
rect 3856 17978 3912 17980
rect 3616 17926 3662 17978
rect 3662 17926 3672 17978
rect 3696 17926 3726 17978
rect 3726 17926 3738 17978
rect 3738 17926 3752 17978
rect 3776 17926 3790 17978
rect 3790 17926 3802 17978
rect 3802 17926 3832 17978
rect 3856 17926 3866 17978
rect 3866 17926 3912 17978
rect 3616 17924 3672 17926
rect 3696 17924 3752 17926
rect 3776 17924 3832 17926
rect 3856 17924 3912 17926
rect 3616 16890 3672 16892
rect 3696 16890 3752 16892
rect 3776 16890 3832 16892
rect 3856 16890 3912 16892
rect 3616 16838 3662 16890
rect 3662 16838 3672 16890
rect 3696 16838 3726 16890
rect 3726 16838 3738 16890
rect 3738 16838 3752 16890
rect 3776 16838 3790 16890
rect 3790 16838 3802 16890
rect 3802 16838 3832 16890
rect 3856 16838 3866 16890
rect 3866 16838 3912 16890
rect 3616 16836 3672 16838
rect 3696 16836 3752 16838
rect 3776 16836 3832 16838
rect 3856 16836 3912 16838
rect 3616 15802 3672 15804
rect 3696 15802 3752 15804
rect 3776 15802 3832 15804
rect 3856 15802 3912 15804
rect 3616 15750 3662 15802
rect 3662 15750 3672 15802
rect 3696 15750 3726 15802
rect 3726 15750 3738 15802
rect 3738 15750 3752 15802
rect 3776 15750 3790 15802
rect 3790 15750 3802 15802
rect 3802 15750 3832 15802
rect 3856 15750 3866 15802
rect 3866 15750 3912 15802
rect 3616 15748 3672 15750
rect 3696 15748 3752 15750
rect 3776 15748 3832 15750
rect 3856 15748 3912 15750
rect 3616 14714 3672 14716
rect 3696 14714 3752 14716
rect 3776 14714 3832 14716
rect 3856 14714 3912 14716
rect 3616 14662 3662 14714
rect 3662 14662 3672 14714
rect 3696 14662 3726 14714
rect 3726 14662 3738 14714
rect 3738 14662 3752 14714
rect 3776 14662 3790 14714
rect 3790 14662 3802 14714
rect 3802 14662 3832 14714
rect 3856 14662 3866 14714
rect 3866 14662 3912 14714
rect 3616 14660 3672 14662
rect 3696 14660 3752 14662
rect 3776 14660 3832 14662
rect 3856 14660 3912 14662
rect 3616 13626 3672 13628
rect 3696 13626 3752 13628
rect 3776 13626 3832 13628
rect 3856 13626 3912 13628
rect 3616 13574 3662 13626
rect 3662 13574 3672 13626
rect 3696 13574 3726 13626
rect 3726 13574 3738 13626
rect 3738 13574 3752 13626
rect 3776 13574 3790 13626
rect 3790 13574 3802 13626
rect 3802 13574 3832 13626
rect 3856 13574 3866 13626
rect 3866 13574 3912 13626
rect 3616 13572 3672 13574
rect 3696 13572 3752 13574
rect 3776 13572 3832 13574
rect 3856 13572 3912 13574
rect 3616 12538 3672 12540
rect 3696 12538 3752 12540
rect 3776 12538 3832 12540
rect 3856 12538 3912 12540
rect 3616 12486 3662 12538
rect 3662 12486 3672 12538
rect 3696 12486 3726 12538
rect 3726 12486 3738 12538
rect 3738 12486 3752 12538
rect 3776 12486 3790 12538
rect 3790 12486 3802 12538
rect 3802 12486 3832 12538
rect 3856 12486 3866 12538
rect 3866 12486 3912 12538
rect 3616 12484 3672 12486
rect 3696 12484 3752 12486
rect 3776 12484 3832 12486
rect 3856 12484 3912 12486
rect 3616 11450 3672 11452
rect 3696 11450 3752 11452
rect 3776 11450 3832 11452
rect 3856 11450 3912 11452
rect 3616 11398 3662 11450
rect 3662 11398 3672 11450
rect 3696 11398 3726 11450
rect 3726 11398 3738 11450
rect 3738 11398 3752 11450
rect 3776 11398 3790 11450
rect 3790 11398 3802 11450
rect 3802 11398 3832 11450
rect 3856 11398 3866 11450
rect 3866 11398 3912 11450
rect 3616 11396 3672 11398
rect 3696 11396 3752 11398
rect 3776 11396 3832 11398
rect 3856 11396 3912 11398
rect 3616 10362 3672 10364
rect 3696 10362 3752 10364
rect 3776 10362 3832 10364
rect 3856 10362 3912 10364
rect 3616 10310 3662 10362
rect 3662 10310 3672 10362
rect 3696 10310 3726 10362
rect 3726 10310 3738 10362
rect 3738 10310 3752 10362
rect 3776 10310 3790 10362
rect 3790 10310 3802 10362
rect 3802 10310 3832 10362
rect 3856 10310 3866 10362
rect 3866 10310 3912 10362
rect 3616 10308 3672 10310
rect 3696 10308 3752 10310
rect 3776 10308 3832 10310
rect 3856 10308 3912 10310
rect 3616 9274 3672 9276
rect 3696 9274 3752 9276
rect 3776 9274 3832 9276
rect 3856 9274 3912 9276
rect 3616 9222 3662 9274
rect 3662 9222 3672 9274
rect 3696 9222 3726 9274
rect 3726 9222 3738 9274
rect 3738 9222 3752 9274
rect 3776 9222 3790 9274
rect 3790 9222 3802 9274
rect 3802 9222 3832 9274
rect 3856 9222 3866 9274
rect 3866 9222 3912 9274
rect 3616 9220 3672 9222
rect 3696 9220 3752 9222
rect 3776 9220 3832 9222
rect 3856 9220 3912 9222
rect 3616 8186 3672 8188
rect 3696 8186 3752 8188
rect 3776 8186 3832 8188
rect 3856 8186 3912 8188
rect 3616 8134 3662 8186
rect 3662 8134 3672 8186
rect 3696 8134 3726 8186
rect 3726 8134 3738 8186
rect 3738 8134 3752 8186
rect 3776 8134 3790 8186
rect 3790 8134 3802 8186
rect 3802 8134 3832 8186
rect 3856 8134 3866 8186
rect 3866 8134 3912 8186
rect 3616 8132 3672 8134
rect 3696 8132 3752 8134
rect 3776 8132 3832 8134
rect 3856 8132 3912 8134
rect 3616 7098 3672 7100
rect 3696 7098 3752 7100
rect 3776 7098 3832 7100
rect 3856 7098 3912 7100
rect 3616 7046 3662 7098
rect 3662 7046 3672 7098
rect 3696 7046 3726 7098
rect 3726 7046 3738 7098
rect 3738 7046 3752 7098
rect 3776 7046 3790 7098
rect 3790 7046 3802 7098
rect 3802 7046 3832 7098
rect 3856 7046 3866 7098
rect 3866 7046 3912 7098
rect 3616 7044 3672 7046
rect 3696 7044 3752 7046
rect 3776 7044 3832 7046
rect 3856 7044 3912 7046
rect 2956 6554 3012 6556
rect 3036 6554 3092 6556
rect 3116 6554 3172 6556
rect 3196 6554 3252 6556
rect 2956 6502 3002 6554
rect 3002 6502 3012 6554
rect 3036 6502 3066 6554
rect 3066 6502 3078 6554
rect 3078 6502 3092 6554
rect 3116 6502 3130 6554
rect 3130 6502 3142 6554
rect 3142 6502 3172 6554
rect 3196 6502 3206 6554
rect 3206 6502 3252 6554
rect 2956 6500 3012 6502
rect 3036 6500 3092 6502
rect 3116 6500 3172 6502
rect 3196 6500 3252 6502
rect 3616 6010 3672 6012
rect 3696 6010 3752 6012
rect 3776 6010 3832 6012
rect 3856 6010 3912 6012
rect 3616 5958 3662 6010
rect 3662 5958 3672 6010
rect 3696 5958 3726 6010
rect 3726 5958 3738 6010
rect 3738 5958 3752 6010
rect 3776 5958 3790 6010
rect 3790 5958 3802 6010
rect 3802 5958 3832 6010
rect 3856 5958 3866 6010
rect 3866 5958 3912 6010
rect 3616 5956 3672 5958
rect 3696 5956 3752 5958
rect 3776 5956 3832 5958
rect 3856 5956 3912 5958
rect 4556 45722 4612 45724
rect 4636 45722 4692 45724
rect 4716 45722 4772 45724
rect 4796 45722 4852 45724
rect 4556 45670 4602 45722
rect 4602 45670 4612 45722
rect 4636 45670 4666 45722
rect 4666 45670 4678 45722
rect 4678 45670 4692 45722
rect 4716 45670 4730 45722
rect 4730 45670 4742 45722
rect 4742 45670 4772 45722
rect 4796 45670 4806 45722
rect 4806 45670 4852 45722
rect 4556 45668 4612 45670
rect 4636 45668 4692 45670
rect 4716 45668 4772 45670
rect 4796 45668 4852 45670
rect 4556 44634 4612 44636
rect 4636 44634 4692 44636
rect 4716 44634 4772 44636
rect 4796 44634 4852 44636
rect 4556 44582 4602 44634
rect 4602 44582 4612 44634
rect 4636 44582 4666 44634
rect 4666 44582 4678 44634
rect 4678 44582 4692 44634
rect 4716 44582 4730 44634
rect 4730 44582 4742 44634
rect 4742 44582 4772 44634
rect 4796 44582 4806 44634
rect 4806 44582 4852 44634
rect 4556 44580 4612 44582
rect 4636 44580 4692 44582
rect 4716 44580 4772 44582
rect 4796 44580 4852 44582
rect 5216 49530 5272 49532
rect 5296 49530 5352 49532
rect 5376 49530 5432 49532
rect 5456 49530 5512 49532
rect 5216 49478 5262 49530
rect 5262 49478 5272 49530
rect 5296 49478 5326 49530
rect 5326 49478 5338 49530
rect 5338 49478 5352 49530
rect 5376 49478 5390 49530
rect 5390 49478 5402 49530
rect 5402 49478 5432 49530
rect 5456 49478 5466 49530
rect 5466 49478 5512 49530
rect 5216 49476 5272 49478
rect 5296 49476 5352 49478
rect 5376 49476 5432 49478
rect 5456 49476 5512 49478
rect 5216 48442 5272 48444
rect 5296 48442 5352 48444
rect 5376 48442 5432 48444
rect 5456 48442 5512 48444
rect 5216 48390 5262 48442
rect 5262 48390 5272 48442
rect 5296 48390 5326 48442
rect 5326 48390 5338 48442
rect 5338 48390 5352 48442
rect 5376 48390 5390 48442
rect 5390 48390 5402 48442
rect 5402 48390 5432 48442
rect 5456 48390 5466 48442
rect 5466 48390 5512 48442
rect 5216 48388 5272 48390
rect 5296 48388 5352 48390
rect 5376 48388 5432 48390
rect 5456 48388 5512 48390
rect 5216 47354 5272 47356
rect 5296 47354 5352 47356
rect 5376 47354 5432 47356
rect 5456 47354 5512 47356
rect 5216 47302 5262 47354
rect 5262 47302 5272 47354
rect 5296 47302 5326 47354
rect 5326 47302 5338 47354
rect 5338 47302 5352 47354
rect 5376 47302 5390 47354
rect 5390 47302 5402 47354
rect 5402 47302 5432 47354
rect 5456 47302 5466 47354
rect 5466 47302 5512 47354
rect 5216 47300 5272 47302
rect 5296 47300 5352 47302
rect 5376 47300 5432 47302
rect 5456 47300 5512 47302
rect 5216 46266 5272 46268
rect 5296 46266 5352 46268
rect 5376 46266 5432 46268
rect 5456 46266 5512 46268
rect 5216 46214 5262 46266
rect 5262 46214 5272 46266
rect 5296 46214 5326 46266
rect 5326 46214 5338 46266
rect 5338 46214 5352 46266
rect 5376 46214 5390 46266
rect 5390 46214 5402 46266
rect 5402 46214 5432 46266
rect 5456 46214 5466 46266
rect 5466 46214 5512 46266
rect 5216 46212 5272 46214
rect 5296 46212 5352 46214
rect 5376 46212 5432 46214
rect 5456 46212 5512 46214
rect 5170 45328 5226 45384
rect 5216 45178 5272 45180
rect 5296 45178 5352 45180
rect 5376 45178 5432 45180
rect 5456 45178 5512 45180
rect 5216 45126 5262 45178
rect 5262 45126 5272 45178
rect 5296 45126 5326 45178
rect 5326 45126 5338 45178
rect 5338 45126 5352 45178
rect 5376 45126 5390 45178
rect 5390 45126 5402 45178
rect 5402 45126 5432 45178
rect 5456 45126 5466 45178
rect 5466 45126 5512 45178
rect 5216 45124 5272 45126
rect 5296 45124 5352 45126
rect 5376 45124 5432 45126
rect 5456 45124 5512 45126
rect 5170 44920 5226 44976
rect 5446 44820 5448 44840
rect 5448 44820 5500 44840
rect 5500 44820 5502 44840
rect 5446 44784 5502 44820
rect 4556 43546 4612 43548
rect 4636 43546 4692 43548
rect 4716 43546 4772 43548
rect 4796 43546 4852 43548
rect 4556 43494 4602 43546
rect 4602 43494 4612 43546
rect 4636 43494 4666 43546
rect 4666 43494 4678 43546
rect 4678 43494 4692 43546
rect 4716 43494 4730 43546
rect 4730 43494 4742 43546
rect 4742 43494 4772 43546
rect 4796 43494 4806 43546
rect 4806 43494 4852 43546
rect 4556 43492 4612 43494
rect 4636 43492 4692 43494
rect 4716 43492 4772 43494
rect 4796 43492 4852 43494
rect 4342 36624 4398 36680
rect 4250 36352 4306 36408
rect 4342 22888 4398 22944
rect 4250 22616 4306 22672
rect 2956 5466 3012 5468
rect 3036 5466 3092 5468
rect 3116 5466 3172 5468
rect 3196 5466 3252 5468
rect 2956 5414 3002 5466
rect 3002 5414 3012 5466
rect 3036 5414 3066 5466
rect 3066 5414 3078 5466
rect 3078 5414 3092 5466
rect 3116 5414 3130 5466
rect 3130 5414 3142 5466
rect 3142 5414 3172 5466
rect 3196 5414 3206 5466
rect 3206 5414 3252 5466
rect 2956 5412 3012 5414
rect 3036 5412 3092 5414
rect 3116 5412 3172 5414
rect 3196 5412 3252 5414
rect 3616 4922 3672 4924
rect 3696 4922 3752 4924
rect 3776 4922 3832 4924
rect 3856 4922 3912 4924
rect 3616 4870 3662 4922
rect 3662 4870 3672 4922
rect 3696 4870 3726 4922
rect 3726 4870 3738 4922
rect 3738 4870 3752 4922
rect 3776 4870 3790 4922
rect 3790 4870 3802 4922
rect 3802 4870 3832 4922
rect 3856 4870 3866 4922
rect 3866 4870 3912 4922
rect 3616 4868 3672 4870
rect 3696 4868 3752 4870
rect 3776 4868 3832 4870
rect 3856 4868 3912 4870
rect 4556 42458 4612 42460
rect 4636 42458 4692 42460
rect 4716 42458 4772 42460
rect 4796 42458 4852 42460
rect 4556 42406 4602 42458
rect 4602 42406 4612 42458
rect 4636 42406 4666 42458
rect 4666 42406 4678 42458
rect 4678 42406 4692 42458
rect 4716 42406 4730 42458
rect 4730 42406 4742 42458
rect 4742 42406 4772 42458
rect 4796 42406 4806 42458
rect 4806 42406 4852 42458
rect 4556 42404 4612 42406
rect 4636 42404 4692 42406
rect 4716 42404 4772 42406
rect 4796 42404 4852 42406
rect 4618 42200 4674 42256
rect 4556 41370 4612 41372
rect 4636 41370 4692 41372
rect 4716 41370 4772 41372
rect 4796 41370 4852 41372
rect 4556 41318 4602 41370
rect 4602 41318 4612 41370
rect 4636 41318 4666 41370
rect 4666 41318 4678 41370
rect 4678 41318 4692 41370
rect 4716 41318 4730 41370
rect 4730 41318 4742 41370
rect 4742 41318 4772 41370
rect 4796 41318 4806 41370
rect 4806 41318 4852 41370
rect 4556 41316 4612 41318
rect 4636 41316 4692 41318
rect 4716 41316 4772 41318
rect 4796 41316 4852 41318
rect 5216 44090 5272 44092
rect 5296 44090 5352 44092
rect 5376 44090 5432 44092
rect 5456 44090 5512 44092
rect 5216 44038 5262 44090
rect 5262 44038 5272 44090
rect 5296 44038 5326 44090
rect 5326 44038 5338 44090
rect 5338 44038 5352 44090
rect 5376 44038 5390 44090
rect 5390 44038 5402 44090
rect 5402 44038 5432 44090
rect 5456 44038 5466 44090
rect 5466 44038 5512 44090
rect 5216 44036 5272 44038
rect 5296 44036 5352 44038
rect 5376 44036 5432 44038
rect 5456 44036 5512 44038
rect 5216 43002 5272 43004
rect 5296 43002 5352 43004
rect 5376 43002 5432 43004
rect 5456 43002 5512 43004
rect 5216 42950 5262 43002
rect 5262 42950 5272 43002
rect 5296 42950 5326 43002
rect 5326 42950 5338 43002
rect 5338 42950 5352 43002
rect 5376 42950 5390 43002
rect 5390 42950 5402 43002
rect 5402 42950 5432 43002
rect 5456 42950 5466 43002
rect 5466 42950 5512 43002
rect 5216 42948 5272 42950
rect 5296 42948 5352 42950
rect 5376 42948 5432 42950
rect 5456 42948 5512 42950
rect 5262 42644 5264 42664
rect 5264 42644 5316 42664
rect 5316 42644 5318 42664
rect 5262 42608 5318 42644
rect 5630 44784 5686 44840
rect 5216 41914 5272 41916
rect 5296 41914 5352 41916
rect 5376 41914 5432 41916
rect 5456 41914 5512 41916
rect 5216 41862 5262 41914
rect 5262 41862 5272 41914
rect 5296 41862 5326 41914
rect 5326 41862 5338 41914
rect 5338 41862 5352 41914
rect 5376 41862 5390 41914
rect 5390 41862 5402 41914
rect 5402 41862 5432 41914
rect 5456 41862 5466 41914
rect 5466 41862 5512 41914
rect 5216 41860 5272 41862
rect 5296 41860 5352 41862
rect 5376 41860 5432 41862
rect 5456 41860 5512 41862
rect 5216 40826 5272 40828
rect 5296 40826 5352 40828
rect 5376 40826 5432 40828
rect 5456 40826 5512 40828
rect 5216 40774 5262 40826
rect 5262 40774 5272 40826
rect 5296 40774 5326 40826
rect 5326 40774 5338 40826
rect 5338 40774 5352 40826
rect 5376 40774 5390 40826
rect 5390 40774 5402 40826
rect 5402 40774 5432 40826
rect 5456 40774 5466 40826
rect 5466 40774 5512 40826
rect 5216 40772 5272 40774
rect 5296 40772 5352 40774
rect 5376 40772 5432 40774
rect 5456 40772 5512 40774
rect 4556 40282 4612 40284
rect 4636 40282 4692 40284
rect 4716 40282 4772 40284
rect 4796 40282 4852 40284
rect 4556 40230 4602 40282
rect 4602 40230 4612 40282
rect 4636 40230 4666 40282
rect 4666 40230 4678 40282
rect 4678 40230 4692 40282
rect 4716 40230 4730 40282
rect 4730 40230 4742 40282
rect 4742 40230 4772 40282
rect 4796 40230 4806 40282
rect 4806 40230 4852 40282
rect 4556 40228 4612 40230
rect 4636 40228 4692 40230
rect 4716 40228 4772 40230
rect 4796 40228 4852 40230
rect 4556 39194 4612 39196
rect 4636 39194 4692 39196
rect 4716 39194 4772 39196
rect 4796 39194 4852 39196
rect 4556 39142 4602 39194
rect 4602 39142 4612 39194
rect 4636 39142 4666 39194
rect 4666 39142 4678 39194
rect 4678 39142 4692 39194
rect 4716 39142 4730 39194
rect 4730 39142 4742 39194
rect 4742 39142 4772 39194
rect 4796 39142 4806 39194
rect 4806 39142 4852 39194
rect 4556 39140 4612 39142
rect 4636 39140 4692 39142
rect 4716 39140 4772 39142
rect 4796 39140 4852 39142
rect 4556 38106 4612 38108
rect 4636 38106 4692 38108
rect 4716 38106 4772 38108
rect 4796 38106 4852 38108
rect 4556 38054 4602 38106
rect 4602 38054 4612 38106
rect 4636 38054 4666 38106
rect 4666 38054 4678 38106
rect 4678 38054 4692 38106
rect 4716 38054 4730 38106
rect 4730 38054 4742 38106
rect 4742 38054 4772 38106
rect 4796 38054 4806 38106
rect 4806 38054 4852 38106
rect 4556 38052 4612 38054
rect 4636 38052 4692 38054
rect 4716 38052 4772 38054
rect 4796 38052 4852 38054
rect 4556 37018 4612 37020
rect 4636 37018 4692 37020
rect 4716 37018 4772 37020
rect 4796 37018 4852 37020
rect 4556 36966 4602 37018
rect 4602 36966 4612 37018
rect 4636 36966 4666 37018
rect 4666 36966 4678 37018
rect 4678 36966 4692 37018
rect 4716 36966 4730 37018
rect 4730 36966 4742 37018
rect 4742 36966 4772 37018
rect 4796 36966 4806 37018
rect 4806 36966 4852 37018
rect 4556 36964 4612 36966
rect 4636 36964 4692 36966
rect 4716 36964 4772 36966
rect 4796 36964 4852 36966
rect 4556 35930 4612 35932
rect 4636 35930 4692 35932
rect 4716 35930 4772 35932
rect 4796 35930 4852 35932
rect 4556 35878 4602 35930
rect 4602 35878 4612 35930
rect 4636 35878 4666 35930
rect 4666 35878 4678 35930
rect 4678 35878 4692 35930
rect 4716 35878 4730 35930
rect 4730 35878 4742 35930
rect 4742 35878 4772 35930
rect 4796 35878 4806 35930
rect 4806 35878 4852 35930
rect 4556 35876 4612 35878
rect 4636 35876 4692 35878
rect 4716 35876 4772 35878
rect 4796 35876 4852 35878
rect 4556 34842 4612 34844
rect 4636 34842 4692 34844
rect 4716 34842 4772 34844
rect 4796 34842 4852 34844
rect 4556 34790 4602 34842
rect 4602 34790 4612 34842
rect 4636 34790 4666 34842
rect 4666 34790 4678 34842
rect 4678 34790 4692 34842
rect 4716 34790 4730 34842
rect 4730 34790 4742 34842
rect 4742 34790 4772 34842
rect 4796 34790 4806 34842
rect 4806 34790 4852 34842
rect 4556 34788 4612 34790
rect 4636 34788 4692 34790
rect 4716 34788 4772 34790
rect 4796 34788 4852 34790
rect 4556 33754 4612 33756
rect 4636 33754 4692 33756
rect 4716 33754 4772 33756
rect 4796 33754 4852 33756
rect 4556 33702 4602 33754
rect 4602 33702 4612 33754
rect 4636 33702 4666 33754
rect 4666 33702 4678 33754
rect 4678 33702 4692 33754
rect 4716 33702 4730 33754
rect 4730 33702 4742 33754
rect 4742 33702 4772 33754
rect 4796 33702 4806 33754
rect 4806 33702 4852 33754
rect 4556 33700 4612 33702
rect 4636 33700 4692 33702
rect 4716 33700 4772 33702
rect 4796 33700 4852 33702
rect 4556 32666 4612 32668
rect 4636 32666 4692 32668
rect 4716 32666 4772 32668
rect 4796 32666 4852 32668
rect 4556 32614 4602 32666
rect 4602 32614 4612 32666
rect 4636 32614 4666 32666
rect 4666 32614 4678 32666
rect 4678 32614 4692 32666
rect 4716 32614 4730 32666
rect 4730 32614 4742 32666
rect 4742 32614 4772 32666
rect 4796 32614 4806 32666
rect 4806 32614 4852 32666
rect 4556 32612 4612 32614
rect 4636 32612 4692 32614
rect 4716 32612 4772 32614
rect 4796 32612 4852 32614
rect 4556 31578 4612 31580
rect 4636 31578 4692 31580
rect 4716 31578 4772 31580
rect 4796 31578 4852 31580
rect 4556 31526 4602 31578
rect 4602 31526 4612 31578
rect 4636 31526 4666 31578
rect 4666 31526 4678 31578
rect 4678 31526 4692 31578
rect 4716 31526 4730 31578
rect 4730 31526 4742 31578
rect 4742 31526 4772 31578
rect 4796 31526 4806 31578
rect 4806 31526 4852 31578
rect 4556 31524 4612 31526
rect 4636 31524 4692 31526
rect 4716 31524 4772 31526
rect 4796 31524 4852 31526
rect 4556 30490 4612 30492
rect 4636 30490 4692 30492
rect 4716 30490 4772 30492
rect 4796 30490 4852 30492
rect 4556 30438 4602 30490
rect 4602 30438 4612 30490
rect 4636 30438 4666 30490
rect 4666 30438 4678 30490
rect 4678 30438 4692 30490
rect 4716 30438 4730 30490
rect 4730 30438 4742 30490
rect 4742 30438 4772 30490
rect 4796 30438 4806 30490
rect 4806 30438 4852 30490
rect 4556 30436 4612 30438
rect 4636 30436 4692 30438
rect 4716 30436 4772 30438
rect 4796 30436 4852 30438
rect 4556 29402 4612 29404
rect 4636 29402 4692 29404
rect 4716 29402 4772 29404
rect 4796 29402 4852 29404
rect 4556 29350 4602 29402
rect 4602 29350 4612 29402
rect 4636 29350 4666 29402
rect 4666 29350 4678 29402
rect 4678 29350 4692 29402
rect 4716 29350 4730 29402
rect 4730 29350 4742 29402
rect 4742 29350 4772 29402
rect 4796 29350 4806 29402
rect 4806 29350 4852 29402
rect 4556 29348 4612 29350
rect 4636 29348 4692 29350
rect 4716 29348 4772 29350
rect 4796 29348 4852 29350
rect 4556 28314 4612 28316
rect 4636 28314 4692 28316
rect 4716 28314 4772 28316
rect 4796 28314 4852 28316
rect 4556 28262 4602 28314
rect 4602 28262 4612 28314
rect 4636 28262 4666 28314
rect 4666 28262 4678 28314
rect 4678 28262 4692 28314
rect 4716 28262 4730 28314
rect 4730 28262 4742 28314
rect 4742 28262 4772 28314
rect 4796 28262 4806 28314
rect 4806 28262 4852 28314
rect 4556 28260 4612 28262
rect 4636 28260 4692 28262
rect 4716 28260 4772 28262
rect 4796 28260 4852 28262
rect 4556 27226 4612 27228
rect 4636 27226 4692 27228
rect 4716 27226 4772 27228
rect 4796 27226 4852 27228
rect 4556 27174 4602 27226
rect 4602 27174 4612 27226
rect 4636 27174 4666 27226
rect 4666 27174 4678 27226
rect 4678 27174 4692 27226
rect 4716 27174 4730 27226
rect 4730 27174 4742 27226
rect 4742 27174 4772 27226
rect 4796 27174 4806 27226
rect 4806 27174 4852 27226
rect 4556 27172 4612 27174
rect 4636 27172 4692 27174
rect 4716 27172 4772 27174
rect 4796 27172 4852 27174
rect 4556 26138 4612 26140
rect 4636 26138 4692 26140
rect 4716 26138 4772 26140
rect 4796 26138 4852 26140
rect 4556 26086 4602 26138
rect 4602 26086 4612 26138
rect 4636 26086 4666 26138
rect 4666 26086 4678 26138
rect 4678 26086 4692 26138
rect 4716 26086 4730 26138
rect 4730 26086 4742 26138
rect 4742 26086 4772 26138
rect 4796 26086 4806 26138
rect 4806 26086 4852 26138
rect 4556 26084 4612 26086
rect 4636 26084 4692 26086
rect 4716 26084 4772 26086
rect 4796 26084 4852 26086
rect 4556 25050 4612 25052
rect 4636 25050 4692 25052
rect 4716 25050 4772 25052
rect 4796 25050 4852 25052
rect 4556 24998 4602 25050
rect 4602 24998 4612 25050
rect 4636 24998 4666 25050
rect 4666 24998 4678 25050
rect 4678 24998 4692 25050
rect 4716 24998 4730 25050
rect 4730 24998 4742 25050
rect 4742 24998 4772 25050
rect 4796 24998 4806 25050
rect 4806 24998 4852 25050
rect 4556 24996 4612 24998
rect 4636 24996 4692 24998
rect 4716 24996 4772 24998
rect 4796 24996 4852 24998
rect 4556 23962 4612 23964
rect 4636 23962 4692 23964
rect 4716 23962 4772 23964
rect 4796 23962 4852 23964
rect 4556 23910 4602 23962
rect 4602 23910 4612 23962
rect 4636 23910 4666 23962
rect 4666 23910 4678 23962
rect 4678 23910 4692 23962
rect 4716 23910 4730 23962
rect 4730 23910 4742 23962
rect 4742 23910 4772 23962
rect 4796 23910 4806 23962
rect 4806 23910 4852 23962
rect 4556 23908 4612 23910
rect 4636 23908 4692 23910
rect 4716 23908 4772 23910
rect 4796 23908 4852 23910
rect 4556 22874 4612 22876
rect 4636 22874 4692 22876
rect 4716 22874 4772 22876
rect 4796 22874 4852 22876
rect 4556 22822 4602 22874
rect 4602 22822 4612 22874
rect 4636 22822 4666 22874
rect 4666 22822 4678 22874
rect 4678 22822 4692 22874
rect 4716 22822 4730 22874
rect 4730 22822 4742 22874
rect 4742 22822 4772 22874
rect 4796 22822 4806 22874
rect 4806 22822 4852 22874
rect 4556 22820 4612 22822
rect 4636 22820 4692 22822
rect 4716 22820 4772 22822
rect 4796 22820 4852 22822
rect 4556 21786 4612 21788
rect 4636 21786 4692 21788
rect 4716 21786 4772 21788
rect 4796 21786 4852 21788
rect 4556 21734 4602 21786
rect 4602 21734 4612 21786
rect 4636 21734 4666 21786
rect 4666 21734 4678 21786
rect 4678 21734 4692 21786
rect 4716 21734 4730 21786
rect 4730 21734 4742 21786
rect 4742 21734 4772 21786
rect 4796 21734 4806 21786
rect 4806 21734 4852 21786
rect 4556 21732 4612 21734
rect 4636 21732 4692 21734
rect 4716 21732 4772 21734
rect 4796 21732 4852 21734
rect 4556 20698 4612 20700
rect 4636 20698 4692 20700
rect 4716 20698 4772 20700
rect 4796 20698 4852 20700
rect 4556 20646 4602 20698
rect 4602 20646 4612 20698
rect 4636 20646 4666 20698
rect 4666 20646 4678 20698
rect 4678 20646 4692 20698
rect 4716 20646 4730 20698
rect 4730 20646 4742 20698
rect 4742 20646 4772 20698
rect 4796 20646 4806 20698
rect 4806 20646 4852 20698
rect 4556 20644 4612 20646
rect 4636 20644 4692 20646
rect 4716 20644 4772 20646
rect 4796 20644 4852 20646
rect 4556 19610 4612 19612
rect 4636 19610 4692 19612
rect 4716 19610 4772 19612
rect 4796 19610 4852 19612
rect 4556 19558 4602 19610
rect 4602 19558 4612 19610
rect 4636 19558 4666 19610
rect 4666 19558 4678 19610
rect 4678 19558 4692 19610
rect 4716 19558 4730 19610
rect 4730 19558 4742 19610
rect 4742 19558 4772 19610
rect 4796 19558 4806 19610
rect 4806 19558 4852 19610
rect 4556 19556 4612 19558
rect 4636 19556 4692 19558
rect 4716 19556 4772 19558
rect 4796 19556 4852 19558
rect 5216 39738 5272 39740
rect 5296 39738 5352 39740
rect 5376 39738 5432 39740
rect 5456 39738 5512 39740
rect 5216 39686 5262 39738
rect 5262 39686 5272 39738
rect 5296 39686 5326 39738
rect 5326 39686 5338 39738
rect 5338 39686 5352 39738
rect 5376 39686 5390 39738
rect 5390 39686 5402 39738
rect 5402 39686 5432 39738
rect 5456 39686 5466 39738
rect 5466 39686 5512 39738
rect 5216 39684 5272 39686
rect 5296 39684 5352 39686
rect 5376 39684 5432 39686
rect 5456 39684 5512 39686
rect 6156 62042 6212 62044
rect 6236 62042 6292 62044
rect 6316 62042 6372 62044
rect 6396 62042 6452 62044
rect 6156 61990 6202 62042
rect 6202 61990 6212 62042
rect 6236 61990 6266 62042
rect 6266 61990 6278 62042
rect 6278 61990 6292 62042
rect 6316 61990 6330 62042
rect 6330 61990 6342 62042
rect 6342 61990 6372 62042
rect 6396 61990 6406 62042
rect 6406 61990 6452 62042
rect 6156 61988 6212 61990
rect 6236 61988 6292 61990
rect 6316 61988 6372 61990
rect 6396 61988 6452 61990
rect 6156 60954 6212 60956
rect 6236 60954 6292 60956
rect 6316 60954 6372 60956
rect 6396 60954 6452 60956
rect 6156 60902 6202 60954
rect 6202 60902 6212 60954
rect 6236 60902 6266 60954
rect 6266 60902 6278 60954
rect 6278 60902 6292 60954
rect 6316 60902 6330 60954
rect 6330 60902 6342 60954
rect 6342 60902 6372 60954
rect 6396 60902 6406 60954
rect 6406 60902 6452 60954
rect 6156 60900 6212 60902
rect 6236 60900 6292 60902
rect 6316 60900 6372 60902
rect 6396 60900 6452 60902
rect 6156 59866 6212 59868
rect 6236 59866 6292 59868
rect 6316 59866 6372 59868
rect 6396 59866 6452 59868
rect 6156 59814 6202 59866
rect 6202 59814 6212 59866
rect 6236 59814 6266 59866
rect 6266 59814 6278 59866
rect 6278 59814 6292 59866
rect 6316 59814 6330 59866
rect 6330 59814 6342 59866
rect 6342 59814 6372 59866
rect 6396 59814 6406 59866
rect 6406 59814 6452 59866
rect 6156 59812 6212 59814
rect 6236 59812 6292 59814
rect 6316 59812 6372 59814
rect 6396 59812 6452 59814
rect 6156 58778 6212 58780
rect 6236 58778 6292 58780
rect 6316 58778 6372 58780
rect 6396 58778 6452 58780
rect 6156 58726 6202 58778
rect 6202 58726 6212 58778
rect 6236 58726 6266 58778
rect 6266 58726 6278 58778
rect 6278 58726 6292 58778
rect 6316 58726 6330 58778
rect 6330 58726 6342 58778
rect 6342 58726 6372 58778
rect 6396 58726 6406 58778
rect 6406 58726 6452 58778
rect 6156 58724 6212 58726
rect 6236 58724 6292 58726
rect 6316 58724 6372 58726
rect 6396 58724 6452 58726
rect 6458 57840 6514 57896
rect 6156 57690 6212 57692
rect 6236 57690 6292 57692
rect 6316 57690 6372 57692
rect 6396 57690 6452 57692
rect 6156 57638 6202 57690
rect 6202 57638 6212 57690
rect 6236 57638 6266 57690
rect 6266 57638 6278 57690
rect 6278 57638 6292 57690
rect 6316 57638 6330 57690
rect 6330 57638 6342 57690
rect 6342 57638 6372 57690
rect 6396 57638 6406 57690
rect 6406 57638 6452 57690
rect 6156 57636 6212 57638
rect 6236 57636 6292 57638
rect 6316 57636 6372 57638
rect 6396 57636 6452 57638
rect 6550 57432 6606 57488
rect 6156 56602 6212 56604
rect 6236 56602 6292 56604
rect 6316 56602 6372 56604
rect 6396 56602 6452 56604
rect 6156 56550 6202 56602
rect 6202 56550 6212 56602
rect 6236 56550 6266 56602
rect 6266 56550 6278 56602
rect 6278 56550 6292 56602
rect 6316 56550 6330 56602
rect 6330 56550 6342 56602
rect 6342 56550 6372 56602
rect 6396 56550 6406 56602
rect 6406 56550 6452 56602
rect 6156 56548 6212 56550
rect 6236 56548 6292 56550
rect 6316 56548 6372 56550
rect 6396 56548 6452 56550
rect 6156 55514 6212 55516
rect 6236 55514 6292 55516
rect 6316 55514 6372 55516
rect 6396 55514 6452 55516
rect 6156 55462 6202 55514
rect 6202 55462 6212 55514
rect 6236 55462 6266 55514
rect 6266 55462 6278 55514
rect 6278 55462 6292 55514
rect 6316 55462 6330 55514
rect 6330 55462 6342 55514
rect 6342 55462 6372 55514
rect 6396 55462 6406 55514
rect 6406 55462 6452 55514
rect 6156 55460 6212 55462
rect 6236 55460 6292 55462
rect 6316 55460 6372 55462
rect 6396 55460 6452 55462
rect 6156 54426 6212 54428
rect 6236 54426 6292 54428
rect 6316 54426 6372 54428
rect 6396 54426 6452 54428
rect 6156 54374 6202 54426
rect 6202 54374 6212 54426
rect 6236 54374 6266 54426
rect 6266 54374 6278 54426
rect 6278 54374 6292 54426
rect 6316 54374 6330 54426
rect 6330 54374 6342 54426
rect 6342 54374 6372 54426
rect 6396 54374 6406 54426
rect 6406 54374 6452 54426
rect 6156 54372 6212 54374
rect 6236 54372 6292 54374
rect 6316 54372 6372 54374
rect 6396 54372 6452 54374
rect 5998 53488 6054 53544
rect 6156 53338 6212 53340
rect 6236 53338 6292 53340
rect 6316 53338 6372 53340
rect 6396 53338 6452 53340
rect 6156 53286 6202 53338
rect 6202 53286 6212 53338
rect 6236 53286 6266 53338
rect 6266 53286 6278 53338
rect 6278 53286 6292 53338
rect 6316 53286 6330 53338
rect 6330 53286 6342 53338
rect 6342 53286 6372 53338
rect 6396 53286 6406 53338
rect 6406 53286 6452 53338
rect 6156 53284 6212 53286
rect 6236 53284 6292 53286
rect 6316 53284 6372 53286
rect 6396 53284 6452 53286
rect 6156 52250 6212 52252
rect 6236 52250 6292 52252
rect 6316 52250 6372 52252
rect 6396 52250 6452 52252
rect 6156 52198 6202 52250
rect 6202 52198 6212 52250
rect 6236 52198 6266 52250
rect 6266 52198 6278 52250
rect 6278 52198 6292 52250
rect 6316 52198 6330 52250
rect 6330 52198 6342 52250
rect 6342 52198 6372 52250
rect 6396 52198 6406 52250
rect 6406 52198 6452 52250
rect 6156 52196 6212 52198
rect 6236 52196 6292 52198
rect 6316 52196 6372 52198
rect 6396 52196 6452 52198
rect 6918 67224 6974 67280
rect 7378 68720 7434 68776
rect 7930 72156 7932 72176
rect 7932 72156 7984 72176
rect 7984 72156 7986 72176
rect 7930 72120 7986 72156
rect 7756 71834 7812 71836
rect 7836 71834 7892 71836
rect 7916 71834 7972 71836
rect 7996 71834 8052 71836
rect 7756 71782 7802 71834
rect 7802 71782 7812 71834
rect 7836 71782 7866 71834
rect 7866 71782 7878 71834
rect 7878 71782 7892 71834
rect 7916 71782 7930 71834
rect 7930 71782 7942 71834
rect 7942 71782 7972 71834
rect 7996 71782 8006 71834
rect 8006 71782 8052 71834
rect 7756 71780 7812 71782
rect 7836 71780 7892 71782
rect 7916 71780 7972 71782
rect 7996 71780 8052 71782
rect 7838 71576 7894 71632
rect 7756 70746 7812 70748
rect 7836 70746 7892 70748
rect 7916 70746 7972 70748
rect 7996 70746 8052 70748
rect 7756 70694 7802 70746
rect 7802 70694 7812 70746
rect 7836 70694 7866 70746
rect 7866 70694 7878 70746
rect 7878 70694 7892 70746
rect 7916 70694 7930 70746
rect 7930 70694 7942 70746
rect 7942 70694 7972 70746
rect 7996 70694 8006 70746
rect 8006 70694 8052 70746
rect 7756 70692 7812 70694
rect 7836 70692 7892 70694
rect 7916 70692 7972 70694
rect 7996 70692 8052 70694
rect 7746 70488 7802 70544
rect 8022 70488 8078 70544
rect 7756 69658 7812 69660
rect 7836 69658 7892 69660
rect 7916 69658 7972 69660
rect 7996 69658 8052 69660
rect 7756 69606 7802 69658
rect 7802 69606 7812 69658
rect 7836 69606 7866 69658
rect 7866 69606 7878 69658
rect 7878 69606 7892 69658
rect 7916 69606 7930 69658
rect 7930 69606 7942 69658
rect 7942 69606 7972 69658
rect 7996 69606 8006 69658
rect 8006 69606 8052 69658
rect 7756 69604 7812 69606
rect 7836 69604 7892 69606
rect 7916 69604 7972 69606
rect 7996 69604 8052 69606
rect 7756 68570 7812 68572
rect 7836 68570 7892 68572
rect 7916 68570 7972 68572
rect 7996 68570 8052 68572
rect 7756 68518 7802 68570
rect 7802 68518 7812 68570
rect 7836 68518 7866 68570
rect 7866 68518 7878 68570
rect 7878 68518 7892 68570
rect 7916 68518 7930 68570
rect 7930 68518 7942 68570
rect 7942 68518 7972 68570
rect 7996 68518 8006 68570
rect 8006 68518 8052 68570
rect 7756 68516 7812 68518
rect 7836 68516 7892 68518
rect 7916 68516 7972 68518
rect 7996 68516 8052 68518
rect 8206 70896 8262 70952
rect 7930 68176 7986 68232
rect 6816 66938 6872 66940
rect 6896 66938 6952 66940
rect 6976 66938 7032 66940
rect 7056 66938 7112 66940
rect 6816 66886 6862 66938
rect 6862 66886 6872 66938
rect 6896 66886 6926 66938
rect 6926 66886 6938 66938
rect 6938 66886 6952 66938
rect 6976 66886 6990 66938
rect 6990 66886 7002 66938
rect 7002 66886 7032 66938
rect 7056 66886 7066 66938
rect 7066 66886 7112 66938
rect 6816 66884 6872 66886
rect 6896 66884 6952 66886
rect 6976 66884 7032 66886
rect 7056 66884 7112 66886
rect 6816 65850 6872 65852
rect 6896 65850 6952 65852
rect 6976 65850 7032 65852
rect 7056 65850 7112 65852
rect 6816 65798 6862 65850
rect 6862 65798 6872 65850
rect 6896 65798 6926 65850
rect 6926 65798 6938 65850
rect 6938 65798 6952 65850
rect 6976 65798 6990 65850
rect 6990 65798 7002 65850
rect 7002 65798 7032 65850
rect 7056 65798 7066 65850
rect 7066 65798 7112 65850
rect 6816 65796 6872 65798
rect 6896 65796 6952 65798
rect 6976 65796 7032 65798
rect 7056 65796 7112 65798
rect 7010 64912 7066 64968
rect 6816 64762 6872 64764
rect 6896 64762 6952 64764
rect 6976 64762 7032 64764
rect 7056 64762 7112 64764
rect 6816 64710 6862 64762
rect 6862 64710 6872 64762
rect 6896 64710 6926 64762
rect 6926 64710 6938 64762
rect 6938 64710 6952 64762
rect 6976 64710 6990 64762
rect 6990 64710 7002 64762
rect 7002 64710 7032 64762
rect 7056 64710 7066 64762
rect 7066 64710 7112 64762
rect 6816 64708 6872 64710
rect 6896 64708 6952 64710
rect 6976 64708 7032 64710
rect 7056 64708 7112 64710
rect 6826 64504 6882 64560
rect 8416 73466 8472 73468
rect 8496 73466 8552 73468
rect 8576 73466 8632 73468
rect 8656 73466 8712 73468
rect 8416 73414 8462 73466
rect 8462 73414 8472 73466
rect 8496 73414 8526 73466
rect 8526 73414 8538 73466
rect 8538 73414 8552 73466
rect 8576 73414 8590 73466
rect 8590 73414 8602 73466
rect 8602 73414 8632 73466
rect 8656 73414 8666 73466
rect 8666 73414 8712 73466
rect 8416 73412 8472 73414
rect 8496 73412 8552 73414
rect 8576 73412 8632 73414
rect 8656 73412 8712 73414
rect 8666 73208 8722 73264
rect 8482 73072 8538 73128
rect 8390 72684 8446 72720
rect 8390 72664 8392 72684
rect 8392 72664 8444 72684
rect 8444 72664 8446 72684
rect 9356 84890 9412 84892
rect 9436 84890 9492 84892
rect 9516 84890 9572 84892
rect 9596 84890 9652 84892
rect 9356 84838 9402 84890
rect 9402 84838 9412 84890
rect 9436 84838 9466 84890
rect 9466 84838 9478 84890
rect 9478 84838 9492 84890
rect 9516 84838 9530 84890
rect 9530 84838 9542 84890
rect 9542 84838 9572 84890
rect 9596 84838 9606 84890
rect 9606 84838 9652 84890
rect 9356 84836 9412 84838
rect 9436 84836 9492 84838
rect 9516 84836 9572 84838
rect 9596 84836 9652 84838
rect 9356 83802 9412 83804
rect 9436 83802 9492 83804
rect 9516 83802 9572 83804
rect 9596 83802 9652 83804
rect 9356 83750 9402 83802
rect 9402 83750 9412 83802
rect 9436 83750 9466 83802
rect 9466 83750 9478 83802
rect 9478 83750 9492 83802
rect 9516 83750 9530 83802
rect 9530 83750 9542 83802
rect 9542 83750 9572 83802
rect 9596 83750 9606 83802
rect 9606 83750 9652 83802
rect 9356 83748 9412 83750
rect 9436 83748 9492 83750
rect 9516 83748 9572 83750
rect 9596 83748 9652 83750
rect 9356 82714 9412 82716
rect 9436 82714 9492 82716
rect 9516 82714 9572 82716
rect 9596 82714 9652 82716
rect 9356 82662 9402 82714
rect 9402 82662 9412 82714
rect 9436 82662 9466 82714
rect 9466 82662 9478 82714
rect 9478 82662 9492 82714
rect 9516 82662 9530 82714
rect 9530 82662 9542 82714
rect 9542 82662 9572 82714
rect 9596 82662 9606 82714
rect 9606 82662 9652 82714
rect 9356 82660 9412 82662
rect 9436 82660 9492 82662
rect 9516 82660 9572 82662
rect 9596 82660 9652 82662
rect 9356 81626 9412 81628
rect 9436 81626 9492 81628
rect 9516 81626 9572 81628
rect 9596 81626 9652 81628
rect 9356 81574 9402 81626
rect 9402 81574 9412 81626
rect 9436 81574 9466 81626
rect 9466 81574 9478 81626
rect 9478 81574 9492 81626
rect 9516 81574 9530 81626
rect 9530 81574 9542 81626
rect 9542 81574 9572 81626
rect 9596 81574 9606 81626
rect 9606 81574 9652 81626
rect 9356 81572 9412 81574
rect 9436 81572 9492 81574
rect 9516 81572 9572 81574
rect 9596 81572 9652 81574
rect 9356 80538 9412 80540
rect 9436 80538 9492 80540
rect 9516 80538 9572 80540
rect 9596 80538 9652 80540
rect 9356 80486 9402 80538
rect 9402 80486 9412 80538
rect 9436 80486 9466 80538
rect 9466 80486 9478 80538
rect 9478 80486 9492 80538
rect 9516 80486 9530 80538
rect 9530 80486 9542 80538
rect 9542 80486 9572 80538
rect 9596 80486 9606 80538
rect 9606 80486 9652 80538
rect 9356 80484 9412 80486
rect 9436 80484 9492 80486
rect 9516 80484 9572 80486
rect 9596 80484 9652 80486
rect 9356 79450 9412 79452
rect 9436 79450 9492 79452
rect 9516 79450 9572 79452
rect 9596 79450 9652 79452
rect 9356 79398 9402 79450
rect 9402 79398 9412 79450
rect 9436 79398 9466 79450
rect 9466 79398 9478 79450
rect 9478 79398 9492 79450
rect 9516 79398 9530 79450
rect 9530 79398 9542 79450
rect 9542 79398 9572 79450
rect 9596 79398 9606 79450
rect 9606 79398 9652 79450
rect 9356 79396 9412 79398
rect 9436 79396 9492 79398
rect 9516 79396 9572 79398
rect 9596 79396 9652 79398
rect 9356 78362 9412 78364
rect 9436 78362 9492 78364
rect 9516 78362 9572 78364
rect 9596 78362 9652 78364
rect 9356 78310 9402 78362
rect 9402 78310 9412 78362
rect 9436 78310 9466 78362
rect 9466 78310 9478 78362
rect 9478 78310 9492 78362
rect 9516 78310 9530 78362
rect 9530 78310 9542 78362
rect 9542 78310 9572 78362
rect 9596 78310 9606 78362
rect 9606 78310 9652 78362
rect 9356 78308 9412 78310
rect 9436 78308 9492 78310
rect 9516 78308 9572 78310
rect 9596 78308 9652 78310
rect 9356 77274 9412 77276
rect 9436 77274 9492 77276
rect 9516 77274 9572 77276
rect 9596 77274 9652 77276
rect 9356 77222 9402 77274
rect 9402 77222 9412 77274
rect 9436 77222 9466 77274
rect 9466 77222 9478 77274
rect 9478 77222 9492 77274
rect 9516 77222 9530 77274
rect 9530 77222 9542 77274
rect 9542 77222 9572 77274
rect 9596 77222 9606 77274
rect 9606 77222 9652 77274
rect 9356 77220 9412 77222
rect 9436 77220 9492 77222
rect 9516 77220 9572 77222
rect 9596 77220 9652 77222
rect 9356 76186 9412 76188
rect 9436 76186 9492 76188
rect 9516 76186 9572 76188
rect 9596 76186 9652 76188
rect 9356 76134 9402 76186
rect 9402 76134 9412 76186
rect 9436 76134 9466 76186
rect 9466 76134 9478 76186
rect 9478 76134 9492 76186
rect 9516 76134 9530 76186
rect 9530 76134 9542 76186
rect 9542 76134 9572 76186
rect 9596 76134 9606 76186
rect 9606 76134 9652 76186
rect 9356 76132 9412 76134
rect 9436 76132 9492 76134
rect 9516 76132 9572 76134
rect 9596 76132 9652 76134
rect 9356 75098 9412 75100
rect 9436 75098 9492 75100
rect 9516 75098 9572 75100
rect 9596 75098 9652 75100
rect 9356 75046 9402 75098
rect 9402 75046 9412 75098
rect 9436 75046 9466 75098
rect 9466 75046 9478 75098
rect 9478 75046 9492 75098
rect 9516 75046 9530 75098
rect 9530 75046 9542 75098
rect 9542 75046 9572 75098
rect 9596 75046 9606 75098
rect 9606 75046 9652 75098
rect 9356 75044 9412 75046
rect 9436 75044 9492 75046
rect 9516 75044 9572 75046
rect 9596 75044 9652 75046
rect 8416 72378 8472 72380
rect 8496 72378 8552 72380
rect 8576 72378 8632 72380
rect 8656 72378 8712 72380
rect 8416 72326 8462 72378
rect 8462 72326 8472 72378
rect 8496 72326 8526 72378
rect 8526 72326 8538 72378
rect 8538 72326 8552 72378
rect 8576 72326 8590 72378
rect 8590 72326 8602 72378
rect 8602 72326 8632 72378
rect 8656 72326 8666 72378
rect 8666 72326 8712 72378
rect 8416 72324 8472 72326
rect 8496 72324 8552 72326
rect 8576 72324 8632 72326
rect 8656 72324 8712 72326
rect 8390 71440 8446 71496
rect 8416 71290 8472 71292
rect 8496 71290 8552 71292
rect 8576 71290 8632 71292
rect 8656 71290 8712 71292
rect 8416 71238 8462 71290
rect 8462 71238 8472 71290
rect 8496 71238 8526 71290
rect 8526 71238 8538 71290
rect 8538 71238 8552 71290
rect 8576 71238 8590 71290
rect 8590 71238 8602 71290
rect 8602 71238 8632 71290
rect 8656 71238 8666 71290
rect 8666 71238 8712 71290
rect 8416 71236 8472 71238
rect 8496 71236 8552 71238
rect 8576 71236 8632 71238
rect 8656 71236 8712 71238
rect 8482 71052 8538 71088
rect 8482 71032 8484 71052
rect 8484 71032 8536 71052
rect 8536 71032 8538 71052
rect 8482 70488 8538 70544
rect 8574 70352 8630 70408
rect 8416 70202 8472 70204
rect 8496 70202 8552 70204
rect 8576 70202 8632 70204
rect 8656 70202 8712 70204
rect 8416 70150 8462 70202
rect 8462 70150 8472 70202
rect 8496 70150 8526 70202
rect 8526 70150 8538 70202
rect 8538 70150 8552 70202
rect 8576 70150 8590 70202
rect 8590 70150 8602 70202
rect 8602 70150 8632 70202
rect 8656 70150 8666 70202
rect 8666 70150 8712 70202
rect 8416 70148 8472 70150
rect 8496 70148 8552 70150
rect 8576 70148 8632 70150
rect 8656 70148 8712 70150
rect 8416 69114 8472 69116
rect 8496 69114 8552 69116
rect 8576 69114 8632 69116
rect 8656 69114 8712 69116
rect 8416 69062 8462 69114
rect 8462 69062 8472 69114
rect 8496 69062 8526 69114
rect 8526 69062 8538 69114
rect 8538 69062 8552 69114
rect 8576 69062 8590 69114
rect 8590 69062 8602 69114
rect 8602 69062 8632 69114
rect 8656 69062 8666 69114
rect 8666 69062 8712 69114
rect 8416 69060 8472 69062
rect 8496 69060 8552 69062
rect 8576 69060 8632 69062
rect 8656 69060 8712 69062
rect 8390 68856 8446 68912
rect 8574 68892 8576 68912
rect 8576 68892 8628 68912
rect 8628 68892 8630 68912
rect 8574 68856 8630 68892
rect 8482 68176 8538 68232
rect 8416 68026 8472 68028
rect 8496 68026 8552 68028
rect 8576 68026 8632 68028
rect 8656 68026 8712 68028
rect 8416 67974 8462 68026
rect 8462 67974 8472 68026
rect 8496 67974 8526 68026
rect 8526 67974 8538 68026
rect 8538 67974 8552 68026
rect 8576 67974 8590 68026
rect 8590 67974 8602 68026
rect 8602 67974 8632 68026
rect 8656 67974 8666 68026
rect 8666 67974 8712 68026
rect 8416 67972 8472 67974
rect 8496 67972 8552 67974
rect 8576 67972 8632 67974
rect 8656 67972 8712 67974
rect 7756 67482 7812 67484
rect 7836 67482 7892 67484
rect 7916 67482 7972 67484
rect 7996 67482 8052 67484
rect 7756 67430 7802 67482
rect 7802 67430 7812 67482
rect 7836 67430 7866 67482
rect 7866 67430 7878 67482
rect 7878 67430 7892 67482
rect 7916 67430 7930 67482
rect 7930 67430 7942 67482
rect 7942 67430 7972 67482
rect 7996 67430 8006 67482
rect 8006 67430 8052 67482
rect 7756 67428 7812 67430
rect 7836 67428 7892 67430
rect 7916 67428 7972 67430
rect 7996 67428 8052 67430
rect 7756 66394 7812 66396
rect 7836 66394 7892 66396
rect 7916 66394 7972 66396
rect 7996 66394 8052 66396
rect 7756 66342 7802 66394
rect 7802 66342 7812 66394
rect 7836 66342 7866 66394
rect 7866 66342 7878 66394
rect 7878 66342 7892 66394
rect 7916 66342 7930 66394
rect 7930 66342 7942 66394
rect 7942 66342 7972 66394
rect 7996 66342 8006 66394
rect 8006 66342 8052 66394
rect 7756 66340 7812 66342
rect 7836 66340 7892 66342
rect 7916 66340 7972 66342
rect 7996 66340 8052 66342
rect 7378 66000 7434 66056
rect 6816 63674 6872 63676
rect 6896 63674 6952 63676
rect 6976 63674 7032 63676
rect 7056 63674 7112 63676
rect 6816 63622 6862 63674
rect 6862 63622 6872 63674
rect 6896 63622 6926 63674
rect 6926 63622 6938 63674
rect 6938 63622 6952 63674
rect 6976 63622 6990 63674
rect 6990 63622 7002 63674
rect 7002 63622 7032 63674
rect 7056 63622 7066 63674
rect 7066 63622 7112 63674
rect 6816 63620 6872 63622
rect 6896 63620 6952 63622
rect 6976 63620 7032 63622
rect 7056 63620 7112 63622
rect 6826 62736 6882 62792
rect 6816 62586 6872 62588
rect 6896 62586 6952 62588
rect 6976 62586 7032 62588
rect 7056 62586 7112 62588
rect 6816 62534 6862 62586
rect 6862 62534 6872 62586
rect 6896 62534 6926 62586
rect 6926 62534 6938 62586
rect 6938 62534 6952 62586
rect 6976 62534 6990 62586
rect 6990 62534 7002 62586
rect 7002 62534 7032 62586
rect 7056 62534 7066 62586
rect 7066 62534 7112 62586
rect 6816 62532 6872 62534
rect 6896 62532 6952 62534
rect 6976 62532 7032 62534
rect 7056 62532 7112 62534
rect 6816 61498 6872 61500
rect 6896 61498 6952 61500
rect 6976 61498 7032 61500
rect 7056 61498 7112 61500
rect 6816 61446 6862 61498
rect 6862 61446 6872 61498
rect 6896 61446 6926 61498
rect 6926 61446 6938 61498
rect 6938 61446 6952 61498
rect 6976 61446 6990 61498
rect 6990 61446 7002 61498
rect 7002 61446 7032 61498
rect 7056 61446 7066 61498
rect 7066 61446 7112 61498
rect 6816 61444 6872 61446
rect 6896 61444 6952 61446
rect 6976 61444 7032 61446
rect 7056 61444 7112 61446
rect 7286 62192 7342 62248
rect 7756 65306 7812 65308
rect 7836 65306 7892 65308
rect 7916 65306 7972 65308
rect 7996 65306 8052 65308
rect 7756 65254 7802 65306
rect 7802 65254 7812 65306
rect 7836 65254 7866 65306
rect 7866 65254 7878 65306
rect 7878 65254 7892 65306
rect 7916 65254 7930 65306
rect 7930 65254 7942 65306
rect 7942 65254 7972 65306
rect 7996 65254 8006 65306
rect 8006 65254 8052 65306
rect 7756 65252 7812 65254
rect 7836 65252 7892 65254
rect 7916 65252 7972 65254
rect 7996 65252 8052 65254
rect 8482 67360 8538 67416
rect 8574 67224 8630 67280
rect 8416 66938 8472 66940
rect 8496 66938 8552 66940
rect 8576 66938 8632 66940
rect 8656 66938 8712 66940
rect 8416 66886 8462 66938
rect 8462 66886 8472 66938
rect 8496 66886 8526 66938
rect 8526 66886 8538 66938
rect 8538 66886 8552 66938
rect 8576 66886 8590 66938
rect 8590 66886 8602 66938
rect 8602 66886 8632 66938
rect 8656 66886 8666 66938
rect 8666 66886 8712 66938
rect 8416 66884 8472 66886
rect 8496 66884 8552 66886
rect 8576 66884 8632 66886
rect 8656 66884 8712 66886
rect 8482 66000 8538 66056
rect 8416 65850 8472 65852
rect 8496 65850 8552 65852
rect 8576 65850 8632 65852
rect 8656 65850 8712 65852
rect 8416 65798 8462 65850
rect 8462 65798 8472 65850
rect 8496 65798 8526 65850
rect 8526 65798 8538 65850
rect 8538 65798 8552 65850
rect 8576 65798 8590 65850
rect 8590 65798 8602 65850
rect 8602 65798 8632 65850
rect 8656 65798 8666 65850
rect 8666 65798 8712 65850
rect 8416 65796 8472 65798
rect 8496 65796 8552 65798
rect 8576 65796 8632 65798
rect 8656 65796 8712 65798
rect 9126 73616 9182 73672
rect 9356 74010 9412 74012
rect 9436 74010 9492 74012
rect 9516 74010 9572 74012
rect 9596 74010 9652 74012
rect 9356 73958 9402 74010
rect 9402 73958 9412 74010
rect 9436 73958 9466 74010
rect 9466 73958 9478 74010
rect 9478 73958 9492 74010
rect 9516 73958 9530 74010
rect 9530 73958 9542 74010
rect 9542 73958 9572 74010
rect 9596 73958 9606 74010
rect 9606 73958 9652 74010
rect 9356 73956 9412 73958
rect 9436 73956 9492 73958
rect 9516 73956 9572 73958
rect 9596 73956 9652 73958
rect 9356 72922 9412 72924
rect 9436 72922 9492 72924
rect 9516 72922 9572 72924
rect 9596 72922 9652 72924
rect 9356 72870 9402 72922
rect 9402 72870 9412 72922
rect 9436 72870 9466 72922
rect 9466 72870 9478 72922
rect 9478 72870 9492 72922
rect 9516 72870 9530 72922
rect 9530 72870 9542 72922
rect 9542 72870 9572 72922
rect 9596 72870 9606 72922
rect 9606 72870 9652 72922
rect 9356 72868 9412 72870
rect 9436 72868 9492 72870
rect 9516 72868 9572 72870
rect 9596 72868 9652 72870
rect 9402 72564 9404 72584
rect 9404 72564 9456 72584
rect 9456 72564 9458 72584
rect 9402 72528 9458 72564
rect 9402 71984 9458 72040
rect 9356 71834 9412 71836
rect 9436 71834 9492 71836
rect 9516 71834 9572 71836
rect 9596 71834 9652 71836
rect 9356 71782 9402 71834
rect 9402 71782 9412 71834
rect 9436 71782 9466 71834
rect 9466 71782 9478 71834
rect 9478 71782 9492 71834
rect 9516 71782 9530 71834
rect 9530 71782 9542 71834
rect 9542 71782 9572 71834
rect 9596 71782 9606 71834
rect 9606 71782 9652 71834
rect 9356 71780 9412 71782
rect 9436 71780 9492 71782
rect 9516 71780 9572 71782
rect 9596 71780 9652 71782
rect 9218 70896 9274 70952
rect 9356 70746 9412 70748
rect 9436 70746 9492 70748
rect 9516 70746 9572 70748
rect 9596 70746 9652 70748
rect 9356 70694 9402 70746
rect 9402 70694 9412 70746
rect 9436 70694 9466 70746
rect 9466 70694 9478 70746
rect 9478 70694 9492 70746
rect 9516 70694 9530 70746
rect 9530 70694 9542 70746
rect 9542 70694 9572 70746
rect 9596 70694 9606 70746
rect 9606 70694 9652 70746
rect 9356 70692 9412 70694
rect 9436 70692 9492 70694
rect 9516 70692 9572 70694
rect 9596 70692 9652 70694
rect 9126 70216 9182 70272
rect 9310 70100 9366 70136
rect 9310 70080 9312 70100
rect 9312 70080 9364 70100
rect 9364 70080 9366 70100
rect 9586 69944 9642 70000
rect 9954 74296 10010 74352
rect 9356 69658 9412 69660
rect 9436 69658 9492 69660
rect 9516 69658 9572 69660
rect 9596 69658 9652 69660
rect 9356 69606 9402 69658
rect 9402 69606 9412 69658
rect 9436 69606 9466 69658
rect 9466 69606 9478 69658
rect 9478 69606 9492 69658
rect 9516 69606 9530 69658
rect 9530 69606 9542 69658
rect 9542 69606 9572 69658
rect 9596 69606 9606 69658
rect 9606 69606 9652 69658
rect 9356 69604 9412 69606
rect 9436 69604 9492 69606
rect 9516 69604 9572 69606
rect 9596 69604 9652 69606
rect 9126 68312 9182 68368
rect 9356 68570 9412 68572
rect 9436 68570 9492 68572
rect 9516 68570 9572 68572
rect 9596 68570 9652 68572
rect 9356 68518 9402 68570
rect 9402 68518 9412 68570
rect 9436 68518 9466 68570
rect 9466 68518 9478 68570
rect 9478 68518 9492 68570
rect 9516 68518 9530 68570
rect 9530 68518 9542 68570
rect 9542 68518 9572 68570
rect 9596 68518 9606 68570
rect 9606 68518 9652 68570
rect 9356 68516 9412 68518
rect 9436 68516 9492 68518
rect 9516 68516 9572 68518
rect 9596 68516 9652 68518
rect 9310 67632 9366 67688
rect 9356 67482 9412 67484
rect 9436 67482 9492 67484
rect 9516 67482 9572 67484
rect 9596 67482 9652 67484
rect 9356 67430 9402 67482
rect 9402 67430 9412 67482
rect 9436 67430 9466 67482
rect 9466 67430 9478 67482
rect 9478 67430 9492 67482
rect 9516 67430 9530 67482
rect 9530 67430 9542 67482
rect 9542 67430 9572 67482
rect 9596 67430 9606 67482
rect 9606 67430 9652 67482
rect 9356 67428 9412 67430
rect 9436 67428 9492 67430
rect 9516 67428 9572 67430
rect 9596 67428 9652 67430
rect 9310 67224 9366 67280
rect 9126 67124 9128 67144
rect 9128 67124 9180 67144
rect 9180 67124 9182 67144
rect 9126 67088 9182 67124
rect 7756 64218 7812 64220
rect 7836 64218 7892 64220
rect 7916 64218 7972 64220
rect 7996 64218 8052 64220
rect 7756 64166 7802 64218
rect 7802 64166 7812 64218
rect 7836 64166 7866 64218
rect 7866 64166 7878 64218
rect 7878 64166 7892 64218
rect 7916 64166 7930 64218
rect 7930 64166 7942 64218
rect 7942 64166 7972 64218
rect 7996 64166 8006 64218
rect 8006 64166 8052 64218
rect 7756 64164 7812 64166
rect 7836 64164 7892 64166
rect 7916 64164 7972 64166
rect 7996 64164 8052 64166
rect 8416 64762 8472 64764
rect 8496 64762 8552 64764
rect 8576 64762 8632 64764
rect 8656 64762 8712 64764
rect 8416 64710 8462 64762
rect 8462 64710 8472 64762
rect 8496 64710 8526 64762
rect 8526 64710 8538 64762
rect 8538 64710 8552 64762
rect 8576 64710 8590 64762
rect 8590 64710 8602 64762
rect 8602 64710 8632 64762
rect 8656 64710 8666 64762
rect 8666 64710 8712 64762
rect 8416 64708 8472 64710
rect 8496 64708 8552 64710
rect 8576 64708 8632 64710
rect 8656 64708 8712 64710
rect 8206 63416 8262 63472
rect 7756 63130 7812 63132
rect 7836 63130 7892 63132
rect 7916 63130 7972 63132
rect 7996 63130 8052 63132
rect 7756 63078 7802 63130
rect 7802 63078 7812 63130
rect 7836 63078 7866 63130
rect 7866 63078 7878 63130
rect 7878 63078 7892 63130
rect 7916 63078 7930 63130
rect 7930 63078 7942 63130
rect 7942 63078 7972 63130
rect 7996 63078 8006 63130
rect 8006 63078 8052 63130
rect 7756 63076 7812 63078
rect 7836 63076 7892 63078
rect 7916 63076 7972 63078
rect 7996 63076 8052 63078
rect 6816 60410 6872 60412
rect 6896 60410 6952 60412
rect 6976 60410 7032 60412
rect 7056 60410 7112 60412
rect 6816 60358 6862 60410
rect 6862 60358 6872 60410
rect 6896 60358 6926 60410
rect 6926 60358 6938 60410
rect 6938 60358 6952 60410
rect 6976 60358 6990 60410
rect 6990 60358 7002 60410
rect 7002 60358 7032 60410
rect 7056 60358 7066 60410
rect 7066 60358 7112 60410
rect 6816 60356 6872 60358
rect 6896 60356 6952 60358
rect 6976 60356 7032 60358
rect 7056 60356 7112 60358
rect 6816 59322 6872 59324
rect 6896 59322 6952 59324
rect 6976 59322 7032 59324
rect 7056 59322 7112 59324
rect 6816 59270 6862 59322
rect 6862 59270 6872 59322
rect 6896 59270 6926 59322
rect 6926 59270 6938 59322
rect 6938 59270 6952 59322
rect 6976 59270 6990 59322
rect 6990 59270 7002 59322
rect 7002 59270 7032 59322
rect 7056 59270 7066 59322
rect 7066 59270 7112 59322
rect 6816 59268 6872 59270
rect 6896 59268 6952 59270
rect 6976 59268 7032 59270
rect 7056 59268 7112 59270
rect 6816 58234 6872 58236
rect 6896 58234 6952 58236
rect 6976 58234 7032 58236
rect 7056 58234 7112 58236
rect 6816 58182 6862 58234
rect 6862 58182 6872 58234
rect 6896 58182 6926 58234
rect 6926 58182 6938 58234
rect 6938 58182 6952 58234
rect 6976 58182 6990 58234
rect 6990 58182 7002 58234
rect 7002 58182 7032 58234
rect 7056 58182 7066 58234
rect 7066 58182 7112 58234
rect 6816 58180 6872 58182
rect 6896 58180 6952 58182
rect 6976 58180 7032 58182
rect 7056 58180 7112 58182
rect 6816 57146 6872 57148
rect 6896 57146 6952 57148
rect 6976 57146 7032 57148
rect 7056 57146 7112 57148
rect 6816 57094 6862 57146
rect 6862 57094 6872 57146
rect 6896 57094 6926 57146
rect 6926 57094 6938 57146
rect 6938 57094 6952 57146
rect 6976 57094 6990 57146
rect 6990 57094 7002 57146
rect 7002 57094 7032 57146
rect 7056 57094 7066 57146
rect 7066 57094 7112 57146
rect 6816 57092 6872 57094
rect 6896 57092 6952 57094
rect 6976 57092 7032 57094
rect 7056 57092 7112 57094
rect 6090 51312 6146 51368
rect 6156 51162 6212 51164
rect 6236 51162 6292 51164
rect 6316 51162 6372 51164
rect 6396 51162 6452 51164
rect 6156 51110 6202 51162
rect 6202 51110 6212 51162
rect 6236 51110 6266 51162
rect 6266 51110 6278 51162
rect 6278 51110 6292 51162
rect 6316 51110 6330 51162
rect 6330 51110 6342 51162
rect 6342 51110 6372 51162
rect 6396 51110 6406 51162
rect 6406 51110 6452 51162
rect 6156 51108 6212 51110
rect 6236 51108 6292 51110
rect 6316 51108 6372 51110
rect 6396 51108 6452 51110
rect 6090 50904 6146 50960
rect 6156 50074 6212 50076
rect 6236 50074 6292 50076
rect 6316 50074 6372 50076
rect 6396 50074 6452 50076
rect 6156 50022 6202 50074
rect 6202 50022 6212 50074
rect 6236 50022 6266 50074
rect 6266 50022 6278 50074
rect 6278 50022 6292 50074
rect 6316 50022 6330 50074
rect 6330 50022 6342 50074
rect 6342 50022 6372 50074
rect 6396 50022 6406 50074
rect 6406 50022 6452 50074
rect 6156 50020 6212 50022
rect 6236 50020 6292 50022
rect 6316 50020 6372 50022
rect 6396 50020 6452 50022
rect 6156 48986 6212 48988
rect 6236 48986 6292 48988
rect 6316 48986 6372 48988
rect 6396 48986 6452 48988
rect 6156 48934 6202 48986
rect 6202 48934 6212 48986
rect 6236 48934 6266 48986
rect 6266 48934 6278 48986
rect 6278 48934 6292 48986
rect 6316 48934 6330 48986
rect 6330 48934 6342 48986
rect 6342 48934 6372 48986
rect 6396 48934 6406 48986
rect 6406 48934 6452 48986
rect 6156 48932 6212 48934
rect 6236 48932 6292 48934
rect 6316 48932 6372 48934
rect 6396 48932 6452 48934
rect 6156 47898 6212 47900
rect 6236 47898 6292 47900
rect 6316 47898 6372 47900
rect 6396 47898 6452 47900
rect 6156 47846 6202 47898
rect 6202 47846 6212 47898
rect 6236 47846 6266 47898
rect 6266 47846 6278 47898
rect 6278 47846 6292 47898
rect 6316 47846 6330 47898
rect 6330 47846 6342 47898
rect 6342 47846 6372 47898
rect 6396 47846 6406 47898
rect 6406 47846 6452 47898
rect 6156 47844 6212 47846
rect 6236 47844 6292 47846
rect 6316 47844 6372 47846
rect 6396 47844 6452 47846
rect 6156 46810 6212 46812
rect 6236 46810 6292 46812
rect 6316 46810 6372 46812
rect 6396 46810 6452 46812
rect 6156 46758 6202 46810
rect 6202 46758 6212 46810
rect 6236 46758 6266 46810
rect 6266 46758 6278 46810
rect 6278 46758 6292 46810
rect 6316 46758 6330 46810
rect 6330 46758 6342 46810
rect 6342 46758 6372 46810
rect 6396 46758 6406 46810
rect 6406 46758 6452 46810
rect 6156 46756 6212 46758
rect 6236 46756 6292 46758
rect 6316 46756 6372 46758
rect 6396 46756 6452 46758
rect 5998 45872 6054 45928
rect 5216 38650 5272 38652
rect 5296 38650 5352 38652
rect 5376 38650 5432 38652
rect 5456 38650 5512 38652
rect 5216 38598 5262 38650
rect 5262 38598 5272 38650
rect 5296 38598 5326 38650
rect 5326 38598 5338 38650
rect 5338 38598 5352 38650
rect 5376 38598 5390 38650
rect 5390 38598 5402 38650
rect 5402 38598 5432 38650
rect 5456 38598 5466 38650
rect 5466 38598 5512 38650
rect 5216 38596 5272 38598
rect 5296 38596 5352 38598
rect 5376 38596 5432 38598
rect 5456 38596 5512 38598
rect 5216 37562 5272 37564
rect 5296 37562 5352 37564
rect 5376 37562 5432 37564
rect 5456 37562 5512 37564
rect 5216 37510 5262 37562
rect 5262 37510 5272 37562
rect 5296 37510 5326 37562
rect 5326 37510 5338 37562
rect 5338 37510 5352 37562
rect 5376 37510 5390 37562
rect 5390 37510 5402 37562
rect 5402 37510 5432 37562
rect 5456 37510 5466 37562
rect 5466 37510 5512 37562
rect 5216 37508 5272 37510
rect 5296 37508 5352 37510
rect 5376 37508 5432 37510
rect 5456 37508 5512 37510
rect 5216 36474 5272 36476
rect 5296 36474 5352 36476
rect 5376 36474 5432 36476
rect 5456 36474 5512 36476
rect 5216 36422 5262 36474
rect 5262 36422 5272 36474
rect 5296 36422 5326 36474
rect 5326 36422 5338 36474
rect 5338 36422 5352 36474
rect 5376 36422 5390 36474
rect 5390 36422 5402 36474
rect 5402 36422 5432 36474
rect 5456 36422 5466 36474
rect 5466 36422 5512 36474
rect 5216 36420 5272 36422
rect 5296 36420 5352 36422
rect 5376 36420 5432 36422
rect 5456 36420 5512 36422
rect 5216 35386 5272 35388
rect 5296 35386 5352 35388
rect 5376 35386 5432 35388
rect 5456 35386 5512 35388
rect 5216 35334 5262 35386
rect 5262 35334 5272 35386
rect 5296 35334 5326 35386
rect 5326 35334 5338 35386
rect 5338 35334 5352 35386
rect 5376 35334 5390 35386
rect 5390 35334 5402 35386
rect 5402 35334 5432 35386
rect 5456 35334 5466 35386
rect 5466 35334 5512 35386
rect 5216 35332 5272 35334
rect 5296 35332 5352 35334
rect 5376 35332 5432 35334
rect 5456 35332 5512 35334
rect 5216 34298 5272 34300
rect 5296 34298 5352 34300
rect 5376 34298 5432 34300
rect 5456 34298 5512 34300
rect 5216 34246 5262 34298
rect 5262 34246 5272 34298
rect 5296 34246 5326 34298
rect 5326 34246 5338 34298
rect 5338 34246 5352 34298
rect 5376 34246 5390 34298
rect 5390 34246 5402 34298
rect 5402 34246 5432 34298
rect 5456 34246 5466 34298
rect 5466 34246 5512 34298
rect 5216 34244 5272 34246
rect 5296 34244 5352 34246
rect 5376 34244 5432 34246
rect 5456 34244 5512 34246
rect 5216 33210 5272 33212
rect 5296 33210 5352 33212
rect 5376 33210 5432 33212
rect 5456 33210 5512 33212
rect 5216 33158 5262 33210
rect 5262 33158 5272 33210
rect 5296 33158 5326 33210
rect 5326 33158 5338 33210
rect 5338 33158 5352 33210
rect 5376 33158 5390 33210
rect 5390 33158 5402 33210
rect 5402 33158 5432 33210
rect 5456 33158 5466 33210
rect 5466 33158 5512 33210
rect 5216 33156 5272 33158
rect 5296 33156 5352 33158
rect 5376 33156 5432 33158
rect 5456 33156 5512 33158
rect 5216 32122 5272 32124
rect 5296 32122 5352 32124
rect 5376 32122 5432 32124
rect 5456 32122 5512 32124
rect 5216 32070 5262 32122
rect 5262 32070 5272 32122
rect 5296 32070 5326 32122
rect 5326 32070 5338 32122
rect 5338 32070 5352 32122
rect 5376 32070 5390 32122
rect 5390 32070 5402 32122
rect 5402 32070 5432 32122
rect 5456 32070 5466 32122
rect 5466 32070 5512 32122
rect 5216 32068 5272 32070
rect 5296 32068 5352 32070
rect 5376 32068 5432 32070
rect 5456 32068 5512 32070
rect 5216 31034 5272 31036
rect 5296 31034 5352 31036
rect 5376 31034 5432 31036
rect 5456 31034 5512 31036
rect 5216 30982 5262 31034
rect 5262 30982 5272 31034
rect 5296 30982 5326 31034
rect 5326 30982 5338 31034
rect 5338 30982 5352 31034
rect 5376 30982 5390 31034
rect 5390 30982 5402 31034
rect 5402 30982 5432 31034
rect 5456 30982 5466 31034
rect 5466 30982 5512 31034
rect 5216 30980 5272 30982
rect 5296 30980 5352 30982
rect 5376 30980 5432 30982
rect 5456 30980 5512 30982
rect 5216 29946 5272 29948
rect 5296 29946 5352 29948
rect 5376 29946 5432 29948
rect 5456 29946 5512 29948
rect 5216 29894 5262 29946
rect 5262 29894 5272 29946
rect 5296 29894 5326 29946
rect 5326 29894 5338 29946
rect 5338 29894 5352 29946
rect 5376 29894 5390 29946
rect 5390 29894 5402 29946
rect 5402 29894 5432 29946
rect 5456 29894 5466 29946
rect 5466 29894 5512 29946
rect 5216 29892 5272 29894
rect 5296 29892 5352 29894
rect 5376 29892 5432 29894
rect 5456 29892 5512 29894
rect 6156 45722 6212 45724
rect 6236 45722 6292 45724
rect 6316 45722 6372 45724
rect 6396 45722 6452 45724
rect 6156 45670 6202 45722
rect 6202 45670 6212 45722
rect 6236 45670 6266 45722
rect 6266 45670 6278 45722
rect 6278 45670 6292 45722
rect 6316 45670 6330 45722
rect 6330 45670 6342 45722
rect 6342 45670 6372 45722
rect 6396 45670 6406 45722
rect 6406 45670 6452 45722
rect 6156 45668 6212 45670
rect 6236 45668 6292 45670
rect 6316 45668 6372 45670
rect 6396 45668 6452 45670
rect 6090 45464 6146 45520
rect 6156 44634 6212 44636
rect 6236 44634 6292 44636
rect 6316 44634 6372 44636
rect 6396 44634 6452 44636
rect 6156 44582 6202 44634
rect 6202 44582 6212 44634
rect 6236 44582 6266 44634
rect 6266 44582 6278 44634
rect 6278 44582 6292 44634
rect 6316 44582 6330 44634
rect 6330 44582 6342 44634
rect 6342 44582 6372 44634
rect 6396 44582 6406 44634
rect 6406 44582 6452 44634
rect 6156 44580 6212 44582
rect 6236 44580 6292 44582
rect 6316 44580 6372 44582
rect 6396 44580 6452 44582
rect 6156 43546 6212 43548
rect 6236 43546 6292 43548
rect 6316 43546 6372 43548
rect 6396 43546 6452 43548
rect 6156 43494 6202 43546
rect 6202 43494 6212 43546
rect 6236 43494 6266 43546
rect 6266 43494 6278 43546
rect 6278 43494 6292 43546
rect 6316 43494 6330 43546
rect 6330 43494 6342 43546
rect 6342 43494 6372 43546
rect 6396 43494 6406 43546
rect 6406 43494 6452 43546
rect 6156 43492 6212 43494
rect 6236 43492 6292 43494
rect 6316 43492 6372 43494
rect 6396 43492 6452 43494
rect 6156 42458 6212 42460
rect 6236 42458 6292 42460
rect 6316 42458 6372 42460
rect 6396 42458 6452 42460
rect 6156 42406 6202 42458
rect 6202 42406 6212 42458
rect 6236 42406 6266 42458
rect 6266 42406 6278 42458
rect 6278 42406 6292 42458
rect 6316 42406 6330 42458
rect 6330 42406 6342 42458
rect 6342 42406 6372 42458
rect 6396 42406 6406 42458
rect 6406 42406 6452 42458
rect 6156 42404 6212 42406
rect 6236 42404 6292 42406
rect 6316 42404 6372 42406
rect 6396 42404 6452 42406
rect 6156 41370 6212 41372
rect 6236 41370 6292 41372
rect 6316 41370 6372 41372
rect 6396 41370 6452 41372
rect 6156 41318 6202 41370
rect 6202 41318 6212 41370
rect 6236 41318 6266 41370
rect 6266 41318 6278 41370
rect 6278 41318 6292 41370
rect 6316 41318 6330 41370
rect 6330 41318 6342 41370
rect 6342 41318 6372 41370
rect 6396 41318 6406 41370
rect 6406 41318 6452 41370
rect 6156 41316 6212 41318
rect 6236 41316 6292 41318
rect 6316 41316 6372 41318
rect 6396 41316 6452 41318
rect 5216 28858 5272 28860
rect 5296 28858 5352 28860
rect 5376 28858 5432 28860
rect 5456 28858 5512 28860
rect 5216 28806 5262 28858
rect 5262 28806 5272 28858
rect 5296 28806 5326 28858
rect 5326 28806 5338 28858
rect 5338 28806 5352 28858
rect 5376 28806 5390 28858
rect 5390 28806 5402 28858
rect 5402 28806 5432 28858
rect 5456 28806 5466 28858
rect 5466 28806 5512 28858
rect 5216 28804 5272 28806
rect 5296 28804 5352 28806
rect 5376 28804 5432 28806
rect 5456 28804 5512 28806
rect 5446 27920 5502 27976
rect 5216 27770 5272 27772
rect 5296 27770 5352 27772
rect 5376 27770 5432 27772
rect 5456 27770 5512 27772
rect 5216 27718 5262 27770
rect 5262 27718 5272 27770
rect 5296 27718 5326 27770
rect 5326 27718 5338 27770
rect 5338 27718 5352 27770
rect 5376 27718 5390 27770
rect 5390 27718 5402 27770
rect 5402 27718 5432 27770
rect 5456 27718 5466 27770
rect 5466 27718 5512 27770
rect 5216 27716 5272 27718
rect 5296 27716 5352 27718
rect 5376 27716 5432 27718
rect 5456 27716 5512 27718
rect 5446 27512 5502 27568
rect 5216 26682 5272 26684
rect 5296 26682 5352 26684
rect 5376 26682 5432 26684
rect 5456 26682 5512 26684
rect 5216 26630 5262 26682
rect 5262 26630 5272 26682
rect 5296 26630 5326 26682
rect 5326 26630 5338 26682
rect 5338 26630 5352 26682
rect 5376 26630 5390 26682
rect 5390 26630 5402 26682
rect 5402 26630 5432 26682
rect 5456 26630 5466 26682
rect 5466 26630 5512 26682
rect 5216 26628 5272 26630
rect 5296 26628 5352 26630
rect 5376 26628 5432 26630
rect 5456 26628 5512 26630
rect 5216 25594 5272 25596
rect 5296 25594 5352 25596
rect 5376 25594 5432 25596
rect 5456 25594 5512 25596
rect 5216 25542 5262 25594
rect 5262 25542 5272 25594
rect 5296 25542 5326 25594
rect 5326 25542 5338 25594
rect 5338 25542 5352 25594
rect 5376 25542 5390 25594
rect 5390 25542 5402 25594
rect 5402 25542 5432 25594
rect 5456 25542 5466 25594
rect 5466 25542 5512 25594
rect 5216 25540 5272 25542
rect 5296 25540 5352 25542
rect 5376 25540 5432 25542
rect 5456 25540 5512 25542
rect 4556 18522 4612 18524
rect 4636 18522 4692 18524
rect 4716 18522 4772 18524
rect 4796 18522 4852 18524
rect 4556 18470 4602 18522
rect 4602 18470 4612 18522
rect 4636 18470 4666 18522
rect 4666 18470 4678 18522
rect 4678 18470 4692 18522
rect 4716 18470 4730 18522
rect 4730 18470 4742 18522
rect 4742 18470 4772 18522
rect 4796 18470 4806 18522
rect 4806 18470 4852 18522
rect 4556 18468 4612 18470
rect 4636 18468 4692 18470
rect 4716 18468 4772 18470
rect 4796 18468 4852 18470
rect 4556 17434 4612 17436
rect 4636 17434 4692 17436
rect 4716 17434 4772 17436
rect 4796 17434 4852 17436
rect 4556 17382 4602 17434
rect 4602 17382 4612 17434
rect 4636 17382 4666 17434
rect 4666 17382 4678 17434
rect 4678 17382 4692 17434
rect 4716 17382 4730 17434
rect 4730 17382 4742 17434
rect 4742 17382 4772 17434
rect 4796 17382 4806 17434
rect 4806 17382 4852 17434
rect 4556 17380 4612 17382
rect 4636 17380 4692 17382
rect 4716 17380 4772 17382
rect 4796 17380 4852 17382
rect 4556 16346 4612 16348
rect 4636 16346 4692 16348
rect 4716 16346 4772 16348
rect 4796 16346 4852 16348
rect 4556 16294 4602 16346
rect 4602 16294 4612 16346
rect 4636 16294 4666 16346
rect 4666 16294 4678 16346
rect 4678 16294 4692 16346
rect 4716 16294 4730 16346
rect 4730 16294 4742 16346
rect 4742 16294 4772 16346
rect 4796 16294 4806 16346
rect 4806 16294 4852 16346
rect 4556 16292 4612 16294
rect 4636 16292 4692 16294
rect 4716 16292 4772 16294
rect 4796 16292 4852 16294
rect 4556 15258 4612 15260
rect 4636 15258 4692 15260
rect 4716 15258 4772 15260
rect 4796 15258 4852 15260
rect 4556 15206 4602 15258
rect 4602 15206 4612 15258
rect 4636 15206 4666 15258
rect 4666 15206 4678 15258
rect 4678 15206 4692 15258
rect 4716 15206 4730 15258
rect 4730 15206 4742 15258
rect 4742 15206 4772 15258
rect 4796 15206 4806 15258
rect 4806 15206 4852 15258
rect 4556 15204 4612 15206
rect 4636 15204 4692 15206
rect 4716 15204 4772 15206
rect 4796 15204 4852 15206
rect 4556 14170 4612 14172
rect 4636 14170 4692 14172
rect 4716 14170 4772 14172
rect 4796 14170 4852 14172
rect 4556 14118 4602 14170
rect 4602 14118 4612 14170
rect 4636 14118 4666 14170
rect 4666 14118 4678 14170
rect 4678 14118 4692 14170
rect 4716 14118 4730 14170
rect 4730 14118 4742 14170
rect 4742 14118 4772 14170
rect 4796 14118 4806 14170
rect 4806 14118 4852 14170
rect 4556 14116 4612 14118
rect 4636 14116 4692 14118
rect 4716 14116 4772 14118
rect 4796 14116 4852 14118
rect 4556 13082 4612 13084
rect 4636 13082 4692 13084
rect 4716 13082 4772 13084
rect 4796 13082 4852 13084
rect 4556 13030 4602 13082
rect 4602 13030 4612 13082
rect 4636 13030 4666 13082
rect 4666 13030 4678 13082
rect 4678 13030 4692 13082
rect 4716 13030 4730 13082
rect 4730 13030 4742 13082
rect 4742 13030 4772 13082
rect 4796 13030 4806 13082
rect 4806 13030 4852 13082
rect 4556 13028 4612 13030
rect 4636 13028 4692 13030
rect 4716 13028 4772 13030
rect 4796 13028 4852 13030
rect 4556 11994 4612 11996
rect 4636 11994 4692 11996
rect 4716 11994 4772 11996
rect 4796 11994 4852 11996
rect 4556 11942 4602 11994
rect 4602 11942 4612 11994
rect 4636 11942 4666 11994
rect 4666 11942 4678 11994
rect 4678 11942 4692 11994
rect 4716 11942 4730 11994
rect 4730 11942 4742 11994
rect 4742 11942 4772 11994
rect 4796 11942 4806 11994
rect 4806 11942 4852 11994
rect 4556 11940 4612 11942
rect 4636 11940 4692 11942
rect 4716 11940 4772 11942
rect 4796 11940 4852 11942
rect 4556 10906 4612 10908
rect 4636 10906 4692 10908
rect 4716 10906 4772 10908
rect 4796 10906 4852 10908
rect 4556 10854 4602 10906
rect 4602 10854 4612 10906
rect 4636 10854 4666 10906
rect 4666 10854 4678 10906
rect 4678 10854 4692 10906
rect 4716 10854 4730 10906
rect 4730 10854 4742 10906
rect 4742 10854 4772 10906
rect 4796 10854 4806 10906
rect 4806 10854 4852 10906
rect 4556 10852 4612 10854
rect 4636 10852 4692 10854
rect 4716 10852 4772 10854
rect 4796 10852 4852 10854
rect 4556 9818 4612 9820
rect 4636 9818 4692 9820
rect 4716 9818 4772 9820
rect 4796 9818 4852 9820
rect 4556 9766 4602 9818
rect 4602 9766 4612 9818
rect 4636 9766 4666 9818
rect 4666 9766 4678 9818
rect 4678 9766 4692 9818
rect 4716 9766 4730 9818
rect 4730 9766 4742 9818
rect 4742 9766 4772 9818
rect 4796 9766 4806 9818
rect 4806 9766 4852 9818
rect 4556 9764 4612 9766
rect 4636 9764 4692 9766
rect 4716 9764 4772 9766
rect 4796 9764 4852 9766
rect 4556 8730 4612 8732
rect 4636 8730 4692 8732
rect 4716 8730 4772 8732
rect 4796 8730 4852 8732
rect 4556 8678 4602 8730
rect 4602 8678 4612 8730
rect 4636 8678 4666 8730
rect 4666 8678 4678 8730
rect 4678 8678 4692 8730
rect 4716 8678 4730 8730
rect 4730 8678 4742 8730
rect 4742 8678 4772 8730
rect 4796 8678 4806 8730
rect 4806 8678 4852 8730
rect 4556 8676 4612 8678
rect 4636 8676 4692 8678
rect 4716 8676 4772 8678
rect 4796 8676 4852 8678
rect 4556 7642 4612 7644
rect 4636 7642 4692 7644
rect 4716 7642 4772 7644
rect 4796 7642 4852 7644
rect 4556 7590 4602 7642
rect 4602 7590 4612 7642
rect 4636 7590 4666 7642
rect 4666 7590 4678 7642
rect 4678 7590 4692 7642
rect 4716 7590 4730 7642
rect 4730 7590 4742 7642
rect 4742 7590 4772 7642
rect 4796 7590 4806 7642
rect 4806 7590 4852 7642
rect 4556 7588 4612 7590
rect 4636 7588 4692 7590
rect 4716 7588 4772 7590
rect 4796 7588 4852 7590
rect 4556 6554 4612 6556
rect 4636 6554 4692 6556
rect 4716 6554 4772 6556
rect 4796 6554 4852 6556
rect 4556 6502 4602 6554
rect 4602 6502 4612 6554
rect 4636 6502 4666 6554
rect 4666 6502 4678 6554
rect 4678 6502 4692 6554
rect 4716 6502 4730 6554
rect 4730 6502 4742 6554
rect 4742 6502 4772 6554
rect 4796 6502 4806 6554
rect 4806 6502 4852 6554
rect 4556 6500 4612 6502
rect 4636 6500 4692 6502
rect 4716 6500 4772 6502
rect 4796 6500 4852 6502
rect 4556 5466 4612 5468
rect 4636 5466 4692 5468
rect 4716 5466 4772 5468
rect 4796 5466 4852 5468
rect 4556 5414 4602 5466
rect 4602 5414 4612 5466
rect 4636 5414 4666 5466
rect 4666 5414 4678 5466
rect 4678 5414 4692 5466
rect 4716 5414 4730 5466
rect 4730 5414 4742 5466
rect 4742 5414 4772 5466
rect 4796 5414 4806 5466
rect 4806 5414 4852 5466
rect 4556 5412 4612 5414
rect 4636 5412 4692 5414
rect 4716 5412 4772 5414
rect 4796 5412 4852 5414
rect 2956 4378 3012 4380
rect 3036 4378 3092 4380
rect 3116 4378 3172 4380
rect 3196 4378 3252 4380
rect 2956 4326 3002 4378
rect 3002 4326 3012 4378
rect 3036 4326 3066 4378
rect 3066 4326 3078 4378
rect 3078 4326 3092 4378
rect 3116 4326 3130 4378
rect 3130 4326 3142 4378
rect 3142 4326 3172 4378
rect 3196 4326 3206 4378
rect 3206 4326 3252 4378
rect 2956 4324 3012 4326
rect 3036 4324 3092 4326
rect 3116 4324 3172 4326
rect 3196 4324 3252 4326
rect 4556 4378 4612 4380
rect 4636 4378 4692 4380
rect 4716 4378 4772 4380
rect 4796 4378 4852 4380
rect 4556 4326 4602 4378
rect 4602 4326 4612 4378
rect 4636 4326 4666 4378
rect 4666 4326 4678 4378
rect 4678 4326 4692 4378
rect 4716 4326 4730 4378
rect 4730 4326 4742 4378
rect 4742 4326 4772 4378
rect 4796 4326 4806 4378
rect 4806 4326 4852 4378
rect 4556 4324 4612 4326
rect 4636 4324 4692 4326
rect 4716 4324 4772 4326
rect 4796 4324 4852 4326
rect 3616 3834 3672 3836
rect 3696 3834 3752 3836
rect 3776 3834 3832 3836
rect 3856 3834 3912 3836
rect 3616 3782 3662 3834
rect 3662 3782 3672 3834
rect 3696 3782 3726 3834
rect 3726 3782 3738 3834
rect 3738 3782 3752 3834
rect 3776 3782 3790 3834
rect 3790 3782 3802 3834
rect 3802 3782 3832 3834
rect 3856 3782 3866 3834
rect 3866 3782 3912 3834
rect 3616 3780 3672 3782
rect 3696 3780 3752 3782
rect 3776 3780 3832 3782
rect 3856 3780 3912 3782
rect 2956 3290 3012 3292
rect 3036 3290 3092 3292
rect 3116 3290 3172 3292
rect 3196 3290 3252 3292
rect 2956 3238 3002 3290
rect 3002 3238 3012 3290
rect 3036 3238 3066 3290
rect 3066 3238 3078 3290
rect 3078 3238 3092 3290
rect 3116 3238 3130 3290
rect 3130 3238 3142 3290
rect 3142 3238 3172 3290
rect 3196 3238 3206 3290
rect 3206 3238 3252 3290
rect 2956 3236 3012 3238
rect 3036 3236 3092 3238
rect 3116 3236 3172 3238
rect 3196 3236 3252 3238
rect 4556 3290 4612 3292
rect 4636 3290 4692 3292
rect 4716 3290 4772 3292
rect 4796 3290 4852 3292
rect 4556 3238 4602 3290
rect 4602 3238 4612 3290
rect 4636 3238 4666 3290
rect 4666 3238 4678 3290
rect 4678 3238 4692 3290
rect 4716 3238 4730 3290
rect 4730 3238 4742 3290
rect 4742 3238 4772 3290
rect 4796 3238 4806 3290
rect 4806 3238 4852 3290
rect 4556 3236 4612 3238
rect 4636 3236 4692 3238
rect 4716 3236 4772 3238
rect 4796 3236 4852 3238
rect 3616 2746 3672 2748
rect 3696 2746 3752 2748
rect 3776 2746 3832 2748
rect 3856 2746 3912 2748
rect 3616 2694 3662 2746
rect 3662 2694 3672 2746
rect 3696 2694 3726 2746
rect 3726 2694 3738 2746
rect 3738 2694 3752 2746
rect 3776 2694 3790 2746
rect 3790 2694 3802 2746
rect 3802 2694 3832 2746
rect 3856 2694 3866 2746
rect 3866 2694 3912 2746
rect 3616 2692 3672 2694
rect 3696 2692 3752 2694
rect 3776 2692 3832 2694
rect 3856 2692 3912 2694
rect 2956 2202 3012 2204
rect 3036 2202 3092 2204
rect 3116 2202 3172 2204
rect 3196 2202 3252 2204
rect 2956 2150 3002 2202
rect 3002 2150 3012 2202
rect 3036 2150 3066 2202
rect 3066 2150 3078 2202
rect 3078 2150 3092 2202
rect 3116 2150 3130 2202
rect 3130 2150 3142 2202
rect 3142 2150 3172 2202
rect 3196 2150 3206 2202
rect 3206 2150 3252 2202
rect 2956 2148 3012 2150
rect 3036 2148 3092 2150
rect 3116 2148 3172 2150
rect 3196 2148 3252 2150
rect 4556 2202 4612 2204
rect 4636 2202 4692 2204
rect 4716 2202 4772 2204
rect 4796 2202 4852 2204
rect 4556 2150 4602 2202
rect 4602 2150 4612 2202
rect 4636 2150 4666 2202
rect 4666 2150 4678 2202
rect 4678 2150 4692 2202
rect 4716 2150 4730 2202
rect 4730 2150 4742 2202
rect 4742 2150 4772 2202
rect 4796 2150 4806 2202
rect 4806 2150 4852 2202
rect 4556 2148 4612 2150
rect 4636 2148 4692 2150
rect 4716 2148 4772 2150
rect 4796 2148 4852 2150
rect 1674 1944 1730 2000
rect 3616 1658 3672 1660
rect 3696 1658 3752 1660
rect 3776 1658 3832 1660
rect 3856 1658 3912 1660
rect 3616 1606 3662 1658
rect 3662 1606 3672 1658
rect 3696 1606 3726 1658
rect 3726 1606 3738 1658
rect 3738 1606 3752 1658
rect 3776 1606 3790 1658
rect 3790 1606 3802 1658
rect 3802 1606 3832 1658
rect 3856 1606 3866 1658
rect 3866 1606 3912 1658
rect 3616 1604 3672 1606
rect 3696 1604 3752 1606
rect 3776 1604 3832 1606
rect 3856 1604 3912 1606
rect 2956 1114 3012 1116
rect 3036 1114 3092 1116
rect 3116 1114 3172 1116
rect 3196 1114 3252 1116
rect 2956 1062 3002 1114
rect 3002 1062 3012 1114
rect 3036 1062 3066 1114
rect 3066 1062 3078 1114
rect 3078 1062 3092 1114
rect 3116 1062 3130 1114
rect 3130 1062 3142 1114
rect 3142 1062 3172 1114
rect 3196 1062 3206 1114
rect 3206 1062 3252 1114
rect 2956 1060 3012 1062
rect 3036 1060 3092 1062
rect 3116 1060 3172 1062
rect 3196 1060 3252 1062
rect 4556 1114 4612 1116
rect 4636 1114 4692 1116
rect 4716 1114 4772 1116
rect 4796 1114 4852 1116
rect 4556 1062 4602 1114
rect 4602 1062 4612 1114
rect 4636 1062 4666 1114
rect 4666 1062 4678 1114
rect 4678 1062 4692 1114
rect 4716 1062 4730 1114
rect 4730 1062 4742 1114
rect 4742 1062 4772 1114
rect 4796 1062 4806 1114
rect 4806 1062 4852 1114
rect 4556 1060 4612 1062
rect 4636 1060 4692 1062
rect 4716 1060 4772 1062
rect 4796 1060 4852 1062
rect 5216 24506 5272 24508
rect 5296 24506 5352 24508
rect 5376 24506 5432 24508
rect 5456 24506 5512 24508
rect 5216 24454 5262 24506
rect 5262 24454 5272 24506
rect 5296 24454 5326 24506
rect 5326 24454 5338 24506
rect 5338 24454 5352 24506
rect 5376 24454 5390 24506
rect 5390 24454 5402 24506
rect 5402 24454 5432 24506
rect 5456 24454 5466 24506
rect 5466 24454 5512 24506
rect 5216 24452 5272 24454
rect 5296 24452 5352 24454
rect 5376 24452 5432 24454
rect 5456 24452 5512 24454
rect 5216 23418 5272 23420
rect 5296 23418 5352 23420
rect 5376 23418 5432 23420
rect 5456 23418 5512 23420
rect 5216 23366 5262 23418
rect 5262 23366 5272 23418
rect 5296 23366 5326 23418
rect 5326 23366 5338 23418
rect 5338 23366 5352 23418
rect 5376 23366 5390 23418
rect 5390 23366 5402 23418
rect 5402 23366 5432 23418
rect 5456 23366 5466 23418
rect 5466 23366 5512 23418
rect 5216 23364 5272 23366
rect 5296 23364 5352 23366
rect 5376 23364 5432 23366
rect 5456 23364 5512 23366
rect 5216 22330 5272 22332
rect 5296 22330 5352 22332
rect 5376 22330 5432 22332
rect 5456 22330 5512 22332
rect 5216 22278 5262 22330
rect 5262 22278 5272 22330
rect 5296 22278 5326 22330
rect 5326 22278 5338 22330
rect 5338 22278 5352 22330
rect 5376 22278 5390 22330
rect 5390 22278 5402 22330
rect 5402 22278 5432 22330
rect 5456 22278 5466 22330
rect 5466 22278 5512 22330
rect 5216 22276 5272 22278
rect 5296 22276 5352 22278
rect 5376 22276 5432 22278
rect 5456 22276 5512 22278
rect 5216 21242 5272 21244
rect 5296 21242 5352 21244
rect 5376 21242 5432 21244
rect 5456 21242 5512 21244
rect 5216 21190 5262 21242
rect 5262 21190 5272 21242
rect 5296 21190 5326 21242
rect 5326 21190 5338 21242
rect 5338 21190 5352 21242
rect 5376 21190 5390 21242
rect 5390 21190 5402 21242
rect 5402 21190 5432 21242
rect 5456 21190 5466 21242
rect 5466 21190 5512 21242
rect 5216 21188 5272 21190
rect 5296 21188 5352 21190
rect 5376 21188 5432 21190
rect 5456 21188 5512 21190
rect 5216 20154 5272 20156
rect 5296 20154 5352 20156
rect 5376 20154 5432 20156
rect 5456 20154 5512 20156
rect 5216 20102 5262 20154
rect 5262 20102 5272 20154
rect 5296 20102 5326 20154
rect 5326 20102 5338 20154
rect 5338 20102 5352 20154
rect 5376 20102 5390 20154
rect 5390 20102 5402 20154
rect 5402 20102 5432 20154
rect 5456 20102 5466 20154
rect 5466 20102 5512 20154
rect 5216 20100 5272 20102
rect 5296 20100 5352 20102
rect 5376 20100 5432 20102
rect 5456 20100 5512 20102
rect 5216 19066 5272 19068
rect 5296 19066 5352 19068
rect 5376 19066 5432 19068
rect 5456 19066 5512 19068
rect 5216 19014 5262 19066
rect 5262 19014 5272 19066
rect 5296 19014 5326 19066
rect 5326 19014 5338 19066
rect 5338 19014 5352 19066
rect 5376 19014 5390 19066
rect 5390 19014 5402 19066
rect 5402 19014 5432 19066
rect 5456 19014 5466 19066
rect 5466 19014 5512 19066
rect 5216 19012 5272 19014
rect 5296 19012 5352 19014
rect 5376 19012 5432 19014
rect 5456 19012 5512 19014
rect 5216 17978 5272 17980
rect 5296 17978 5352 17980
rect 5376 17978 5432 17980
rect 5456 17978 5512 17980
rect 5216 17926 5262 17978
rect 5262 17926 5272 17978
rect 5296 17926 5326 17978
rect 5326 17926 5338 17978
rect 5338 17926 5352 17978
rect 5376 17926 5390 17978
rect 5390 17926 5402 17978
rect 5402 17926 5432 17978
rect 5456 17926 5466 17978
rect 5466 17926 5512 17978
rect 5216 17924 5272 17926
rect 5296 17924 5352 17926
rect 5376 17924 5432 17926
rect 5456 17924 5512 17926
rect 5216 16890 5272 16892
rect 5296 16890 5352 16892
rect 5376 16890 5432 16892
rect 5456 16890 5512 16892
rect 5216 16838 5262 16890
rect 5262 16838 5272 16890
rect 5296 16838 5326 16890
rect 5326 16838 5338 16890
rect 5338 16838 5352 16890
rect 5376 16838 5390 16890
rect 5390 16838 5402 16890
rect 5402 16838 5432 16890
rect 5456 16838 5466 16890
rect 5466 16838 5512 16890
rect 5216 16836 5272 16838
rect 5296 16836 5352 16838
rect 5376 16836 5432 16838
rect 5456 16836 5512 16838
rect 5216 15802 5272 15804
rect 5296 15802 5352 15804
rect 5376 15802 5432 15804
rect 5456 15802 5512 15804
rect 5216 15750 5262 15802
rect 5262 15750 5272 15802
rect 5296 15750 5326 15802
rect 5326 15750 5338 15802
rect 5338 15750 5352 15802
rect 5376 15750 5390 15802
rect 5390 15750 5402 15802
rect 5402 15750 5432 15802
rect 5456 15750 5466 15802
rect 5466 15750 5512 15802
rect 5216 15748 5272 15750
rect 5296 15748 5352 15750
rect 5376 15748 5432 15750
rect 5456 15748 5512 15750
rect 5216 14714 5272 14716
rect 5296 14714 5352 14716
rect 5376 14714 5432 14716
rect 5456 14714 5512 14716
rect 5216 14662 5262 14714
rect 5262 14662 5272 14714
rect 5296 14662 5326 14714
rect 5326 14662 5338 14714
rect 5338 14662 5352 14714
rect 5376 14662 5390 14714
rect 5390 14662 5402 14714
rect 5402 14662 5432 14714
rect 5456 14662 5466 14714
rect 5466 14662 5512 14714
rect 5216 14660 5272 14662
rect 5296 14660 5352 14662
rect 5376 14660 5432 14662
rect 5456 14660 5512 14662
rect 5216 13626 5272 13628
rect 5296 13626 5352 13628
rect 5376 13626 5432 13628
rect 5456 13626 5512 13628
rect 5216 13574 5262 13626
rect 5262 13574 5272 13626
rect 5296 13574 5326 13626
rect 5326 13574 5338 13626
rect 5338 13574 5352 13626
rect 5376 13574 5390 13626
rect 5390 13574 5402 13626
rect 5402 13574 5432 13626
rect 5456 13574 5466 13626
rect 5466 13574 5512 13626
rect 5216 13572 5272 13574
rect 5296 13572 5352 13574
rect 5376 13572 5432 13574
rect 5456 13572 5512 13574
rect 5216 12538 5272 12540
rect 5296 12538 5352 12540
rect 5376 12538 5432 12540
rect 5456 12538 5512 12540
rect 5216 12486 5262 12538
rect 5262 12486 5272 12538
rect 5296 12486 5326 12538
rect 5326 12486 5338 12538
rect 5338 12486 5352 12538
rect 5376 12486 5390 12538
rect 5390 12486 5402 12538
rect 5402 12486 5432 12538
rect 5456 12486 5466 12538
rect 5466 12486 5512 12538
rect 5216 12484 5272 12486
rect 5296 12484 5352 12486
rect 5376 12484 5432 12486
rect 5456 12484 5512 12486
rect 5216 11450 5272 11452
rect 5296 11450 5352 11452
rect 5376 11450 5432 11452
rect 5456 11450 5512 11452
rect 5216 11398 5262 11450
rect 5262 11398 5272 11450
rect 5296 11398 5326 11450
rect 5326 11398 5338 11450
rect 5338 11398 5352 11450
rect 5376 11398 5390 11450
rect 5390 11398 5402 11450
rect 5402 11398 5432 11450
rect 5456 11398 5466 11450
rect 5466 11398 5512 11450
rect 5216 11396 5272 11398
rect 5296 11396 5352 11398
rect 5376 11396 5432 11398
rect 5456 11396 5512 11398
rect 6156 40282 6212 40284
rect 6236 40282 6292 40284
rect 6316 40282 6372 40284
rect 6396 40282 6452 40284
rect 6156 40230 6202 40282
rect 6202 40230 6212 40282
rect 6236 40230 6266 40282
rect 6266 40230 6278 40282
rect 6278 40230 6292 40282
rect 6316 40230 6330 40282
rect 6330 40230 6342 40282
rect 6342 40230 6372 40282
rect 6396 40230 6406 40282
rect 6406 40230 6452 40282
rect 6156 40228 6212 40230
rect 6236 40228 6292 40230
rect 6316 40228 6372 40230
rect 6396 40228 6452 40230
rect 6156 39194 6212 39196
rect 6236 39194 6292 39196
rect 6316 39194 6372 39196
rect 6396 39194 6452 39196
rect 6156 39142 6202 39194
rect 6202 39142 6212 39194
rect 6236 39142 6266 39194
rect 6266 39142 6278 39194
rect 6278 39142 6292 39194
rect 6316 39142 6330 39194
rect 6330 39142 6342 39194
rect 6342 39142 6372 39194
rect 6396 39142 6406 39194
rect 6406 39142 6452 39194
rect 6156 39140 6212 39142
rect 6236 39140 6292 39142
rect 6316 39140 6372 39142
rect 6396 39140 6452 39142
rect 6156 38106 6212 38108
rect 6236 38106 6292 38108
rect 6316 38106 6372 38108
rect 6396 38106 6452 38108
rect 6156 38054 6202 38106
rect 6202 38054 6212 38106
rect 6236 38054 6266 38106
rect 6266 38054 6278 38106
rect 6278 38054 6292 38106
rect 6316 38054 6330 38106
rect 6330 38054 6342 38106
rect 6342 38054 6372 38106
rect 6396 38054 6406 38106
rect 6406 38054 6452 38106
rect 6156 38052 6212 38054
rect 6236 38052 6292 38054
rect 6316 38052 6372 38054
rect 6396 38052 6452 38054
rect 6156 37018 6212 37020
rect 6236 37018 6292 37020
rect 6316 37018 6372 37020
rect 6396 37018 6452 37020
rect 6156 36966 6202 37018
rect 6202 36966 6212 37018
rect 6236 36966 6266 37018
rect 6266 36966 6278 37018
rect 6278 36966 6292 37018
rect 6316 36966 6330 37018
rect 6330 36966 6342 37018
rect 6342 36966 6372 37018
rect 6396 36966 6406 37018
rect 6406 36966 6452 37018
rect 6156 36964 6212 36966
rect 6236 36964 6292 36966
rect 6316 36964 6372 36966
rect 6396 36964 6452 36966
rect 6816 56058 6872 56060
rect 6896 56058 6952 56060
rect 6976 56058 7032 56060
rect 7056 56058 7112 56060
rect 6816 56006 6862 56058
rect 6862 56006 6872 56058
rect 6896 56006 6926 56058
rect 6926 56006 6938 56058
rect 6938 56006 6952 56058
rect 6976 56006 6990 56058
rect 6990 56006 7002 56058
rect 7002 56006 7032 56058
rect 7056 56006 7066 56058
rect 7066 56006 7112 56058
rect 6816 56004 6872 56006
rect 6896 56004 6952 56006
rect 6976 56004 7032 56006
rect 7056 56004 7112 56006
rect 6816 54970 6872 54972
rect 6896 54970 6952 54972
rect 6976 54970 7032 54972
rect 7056 54970 7112 54972
rect 6816 54918 6862 54970
rect 6862 54918 6872 54970
rect 6896 54918 6926 54970
rect 6926 54918 6938 54970
rect 6938 54918 6952 54970
rect 6976 54918 6990 54970
rect 6990 54918 7002 54970
rect 7002 54918 7032 54970
rect 7056 54918 7066 54970
rect 7066 54918 7112 54970
rect 6816 54916 6872 54918
rect 6896 54916 6952 54918
rect 6976 54916 7032 54918
rect 7056 54916 7112 54918
rect 6816 53882 6872 53884
rect 6896 53882 6952 53884
rect 6976 53882 7032 53884
rect 7056 53882 7112 53884
rect 6816 53830 6862 53882
rect 6862 53830 6872 53882
rect 6896 53830 6926 53882
rect 6926 53830 6938 53882
rect 6938 53830 6952 53882
rect 6976 53830 6990 53882
rect 6990 53830 7002 53882
rect 7002 53830 7032 53882
rect 7056 53830 7066 53882
rect 7066 53830 7112 53882
rect 6816 53828 6872 53830
rect 6896 53828 6952 53830
rect 6976 53828 7032 53830
rect 7056 53828 7112 53830
rect 7102 53524 7104 53544
rect 7104 53524 7156 53544
rect 7156 53524 7158 53544
rect 7102 53488 7158 53524
rect 7756 62042 7812 62044
rect 7836 62042 7892 62044
rect 7916 62042 7972 62044
rect 7996 62042 8052 62044
rect 7756 61990 7802 62042
rect 7802 61990 7812 62042
rect 7836 61990 7866 62042
rect 7866 61990 7878 62042
rect 7878 61990 7892 62042
rect 7916 61990 7930 62042
rect 7930 61990 7942 62042
rect 7942 61990 7972 62042
rect 7996 61990 8006 62042
rect 8006 61990 8052 62042
rect 7756 61988 7812 61990
rect 7836 61988 7892 61990
rect 7916 61988 7972 61990
rect 7996 61988 8052 61990
rect 8416 63674 8472 63676
rect 8496 63674 8552 63676
rect 8576 63674 8632 63676
rect 8656 63674 8712 63676
rect 8416 63622 8462 63674
rect 8462 63622 8472 63674
rect 8496 63622 8526 63674
rect 8526 63622 8538 63674
rect 8538 63622 8552 63674
rect 8576 63622 8590 63674
rect 8590 63622 8602 63674
rect 8602 63622 8632 63674
rect 8656 63622 8666 63674
rect 8666 63622 8712 63674
rect 8416 63620 8472 63622
rect 8496 63620 8552 63622
rect 8576 63620 8632 63622
rect 8656 63620 8712 63622
rect 9402 67124 9404 67144
rect 9404 67124 9456 67144
rect 9456 67124 9458 67144
rect 9402 67088 9458 67124
rect 9356 66394 9412 66396
rect 9436 66394 9492 66396
rect 9516 66394 9572 66396
rect 9596 66394 9652 66396
rect 9356 66342 9402 66394
rect 9402 66342 9412 66394
rect 9436 66342 9466 66394
rect 9466 66342 9478 66394
rect 9478 66342 9492 66394
rect 9516 66342 9530 66394
rect 9530 66342 9542 66394
rect 9542 66342 9572 66394
rect 9596 66342 9606 66394
rect 9606 66342 9652 66394
rect 9356 66340 9412 66342
rect 9436 66340 9492 66342
rect 9516 66340 9572 66342
rect 9596 66340 9652 66342
rect 9356 65306 9412 65308
rect 9436 65306 9492 65308
rect 9516 65306 9572 65308
rect 9596 65306 9652 65308
rect 9356 65254 9402 65306
rect 9402 65254 9412 65306
rect 9436 65254 9466 65306
rect 9466 65254 9478 65306
rect 9478 65254 9492 65306
rect 9516 65254 9530 65306
rect 9530 65254 9542 65306
rect 9542 65254 9572 65306
rect 9596 65254 9606 65306
rect 9606 65254 9652 65306
rect 9356 65252 9412 65254
rect 9436 65252 9492 65254
rect 9516 65252 9572 65254
rect 9596 65252 9652 65254
rect 9356 64218 9412 64220
rect 9436 64218 9492 64220
rect 9516 64218 9572 64220
rect 9596 64218 9652 64220
rect 9356 64166 9402 64218
rect 9402 64166 9412 64218
rect 9436 64166 9466 64218
rect 9466 64166 9478 64218
rect 9478 64166 9492 64218
rect 9516 64166 9530 64218
rect 9530 64166 9542 64218
rect 9542 64166 9572 64218
rect 9596 64166 9606 64218
rect 9606 64166 9652 64218
rect 9356 64164 9412 64166
rect 9436 64164 9492 64166
rect 9516 64164 9572 64166
rect 9596 64164 9652 64166
rect 8390 63280 8446 63336
rect 8942 63280 8998 63336
rect 8666 62892 8722 62928
rect 8666 62872 8668 62892
rect 8668 62872 8720 62892
rect 8720 62872 8722 62892
rect 8416 62586 8472 62588
rect 8496 62586 8552 62588
rect 8576 62586 8632 62588
rect 8656 62586 8712 62588
rect 8416 62534 8462 62586
rect 8462 62534 8472 62586
rect 8496 62534 8526 62586
rect 8526 62534 8538 62586
rect 8538 62534 8552 62586
rect 8576 62534 8590 62586
rect 8590 62534 8602 62586
rect 8602 62534 8632 62586
rect 8656 62534 8666 62586
rect 8666 62534 8712 62586
rect 8416 62532 8472 62534
rect 8496 62532 8552 62534
rect 8576 62532 8632 62534
rect 8656 62532 8712 62534
rect 7756 60954 7812 60956
rect 7836 60954 7892 60956
rect 7916 60954 7972 60956
rect 7996 60954 8052 60956
rect 7756 60902 7802 60954
rect 7802 60902 7812 60954
rect 7836 60902 7866 60954
rect 7866 60902 7878 60954
rect 7878 60902 7892 60954
rect 7916 60902 7930 60954
rect 7930 60902 7942 60954
rect 7942 60902 7972 60954
rect 7996 60902 8006 60954
rect 8006 60902 8052 60954
rect 7756 60900 7812 60902
rect 7836 60900 7892 60902
rect 7916 60900 7972 60902
rect 7996 60900 8052 60902
rect 7756 59866 7812 59868
rect 7836 59866 7892 59868
rect 7916 59866 7972 59868
rect 7996 59866 8052 59868
rect 7756 59814 7802 59866
rect 7802 59814 7812 59866
rect 7836 59814 7866 59866
rect 7866 59814 7878 59866
rect 7878 59814 7892 59866
rect 7916 59814 7930 59866
rect 7930 59814 7942 59866
rect 7942 59814 7972 59866
rect 7996 59814 8006 59866
rect 8006 59814 8052 59866
rect 7756 59812 7812 59814
rect 7836 59812 7892 59814
rect 7916 59812 7972 59814
rect 7996 59812 8052 59814
rect 7756 58778 7812 58780
rect 7836 58778 7892 58780
rect 7916 58778 7972 58780
rect 7996 58778 8052 58780
rect 7756 58726 7802 58778
rect 7802 58726 7812 58778
rect 7836 58726 7866 58778
rect 7866 58726 7878 58778
rect 7878 58726 7892 58778
rect 7916 58726 7930 58778
rect 7930 58726 7942 58778
rect 7942 58726 7972 58778
rect 7996 58726 8006 58778
rect 8006 58726 8052 58778
rect 7756 58724 7812 58726
rect 7836 58724 7892 58726
rect 7916 58724 7972 58726
rect 7996 58724 8052 58726
rect 7756 57690 7812 57692
rect 7836 57690 7892 57692
rect 7916 57690 7972 57692
rect 7996 57690 8052 57692
rect 7756 57638 7802 57690
rect 7802 57638 7812 57690
rect 7836 57638 7866 57690
rect 7866 57638 7878 57690
rect 7878 57638 7892 57690
rect 7916 57638 7930 57690
rect 7930 57638 7942 57690
rect 7942 57638 7972 57690
rect 7996 57638 8006 57690
rect 8006 57638 8052 57690
rect 7756 57636 7812 57638
rect 7836 57636 7892 57638
rect 7916 57636 7972 57638
rect 7996 57636 8052 57638
rect 7756 56602 7812 56604
rect 7836 56602 7892 56604
rect 7916 56602 7972 56604
rect 7996 56602 8052 56604
rect 7756 56550 7802 56602
rect 7802 56550 7812 56602
rect 7836 56550 7866 56602
rect 7866 56550 7878 56602
rect 7878 56550 7892 56602
rect 7916 56550 7930 56602
rect 7930 56550 7942 56602
rect 7942 56550 7972 56602
rect 7996 56550 8006 56602
rect 8006 56550 8052 56602
rect 7756 56548 7812 56550
rect 7836 56548 7892 56550
rect 7916 56548 7972 56550
rect 7996 56548 8052 56550
rect 8416 61498 8472 61500
rect 8496 61498 8552 61500
rect 8576 61498 8632 61500
rect 8656 61498 8712 61500
rect 8416 61446 8462 61498
rect 8462 61446 8472 61498
rect 8496 61446 8526 61498
rect 8526 61446 8538 61498
rect 8538 61446 8552 61498
rect 8576 61446 8590 61498
rect 8590 61446 8602 61498
rect 8602 61446 8632 61498
rect 8656 61446 8666 61498
rect 8666 61446 8712 61498
rect 8416 61444 8472 61446
rect 8496 61444 8552 61446
rect 8576 61444 8632 61446
rect 8656 61444 8712 61446
rect 8416 60410 8472 60412
rect 8496 60410 8552 60412
rect 8576 60410 8632 60412
rect 8656 60410 8712 60412
rect 8416 60358 8462 60410
rect 8462 60358 8472 60410
rect 8496 60358 8526 60410
rect 8526 60358 8538 60410
rect 8538 60358 8552 60410
rect 8576 60358 8590 60410
rect 8590 60358 8602 60410
rect 8602 60358 8632 60410
rect 8656 60358 8666 60410
rect 8666 60358 8712 60410
rect 8416 60356 8472 60358
rect 8496 60356 8552 60358
rect 8576 60356 8632 60358
rect 8656 60356 8712 60358
rect 8416 59322 8472 59324
rect 8496 59322 8552 59324
rect 8576 59322 8632 59324
rect 8656 59322 8712 59324
rect 8416 59270 8462 59322
rect 8462 59270 8472 59322
rect 8496 59270 8526 59322
rect 8526 59270 8538 59322
rect 8538 59270 8552 59322
rect 8576 59270 8590 59322
rect 8590 59270 8602 59322
rect 8602 59270 8632 59322
rect 8656 59270 8666 59322
rect 8666 59270 8712 59322
rect 8416 59268 8472 59270
rect 8496 59268 8552 59270
rect 8576 59268 8632 59270
rect 8656 59268 8712 59270
rect 9034 60424 9090 60480
rect 8416 58234 8472 58236
rect 8496 58234 8552 58236
rect 8576 58234 8632 58236
rect 8656 58234 8712 58236
rect 8416 58182 8462 58234
rect 8462 58182 8472 58234
rect 8496 58182 8526 58234
rect 8526 58182 8538 58234
rect 8538 58182 8552 58234
rect 8576 58182 8590 58234
rect 8590 58182 8602 58234
rect 8602 58182 8632 58234
rect 8656 58182 8666 58234
rect 8666 58182 8712 58234
rect 8416 58180 8472 58182
rect 8496 58180 8552 58182
rect 8576 58180 8632 58182
rect 8656 58180 8712 58182
rect 8298 57840 8354 57896
rect 8206 57704 8262 57760
rect 8942 60152 8998 60208
rect 8850 57840 8906 57896
rect 8416 57146 8472 57148
rect 8496 57146 8552 57148
rect 8576 57146 8632 57148
rect 8656 57146 8712 57148
rect 8416 57094 8462 57146
rect 8462 57094 8472 57146
rect 8496 57094 8526 57146
rect 8526 57094 8538 57146
rect 8538 57094 8552 57146
rect 8576 57094 8590 57146
rect 8590 57094 8602 57146
rect 8602 57094 8632 57146
rect 8656 57094 8666 57146
rect 8666 57094 8712 57146
rect 8416 57092 8472 57094
rect 8496 57092 8552 57094
rect 8576 57092 8632 57094
rect 8656 57092 8712 57094
rect 8416 56058 8472 56060
rect 8496 56058 8552 56060
rect 8576 56058 8632 56060
rect 8656 56058 8712 56060
rect 8416 56006 8462 56058
rect 8462 56006 8472 56058
rect 8496 56006 8526 56058
rect 8526 56006 8538 56058
rect 8538 56006 8552 56058
rect 8576 56006 8590 56058
rect 8590 56006 8602 56058
rect 8602 56006 8632 56058
rect 8656 56006 8666 56058
rect 8666 56006 8712 56058
rect 8416 56004 8472 56006
rect 8496 56004 8552 56006
rect 8576 56004 8632 56006
rect 8656 56004 8712 56006
rect 7756 55514 7812 55516
rect 7836 55514 7892 55516
rect 7916 55514 7972 55516
rect 7996 55514 8052 55516
rect 7756 55462 7802 55514
rect 7802 55462 7812 55514
rect 7836 55462 7866 55514
rect 7866 55462 7878 55514
rect 7878 55462 7892 55514
rect 7916 55462 7930 55514
rect 7930 55462 7942 55514
rect 7942 55462 7972 55514
rect 7996 55462 8006 55514
rect 8006 55462 8052 55514
rect 7756 55460 7812 55462
rect 7836 55460 7892 55462
rect 7916 55460 7972 55462
rect 7996 55460 8052 55462
rect 7756 54426 7812 54428
rect 7836 54426 7892 54428
rect 7916 54426 7972 54428
rect 7996 54426 8052 54428
rect 7756 54374 7802 54426
rect 7802 54374 7812 54426
rect 7836 54374 7866 54426
rect 7866 54374 7878 54426
rect 7878 54374 7892 54426
rect 7916 54374 7930 54426
rect 7930 54374 7942 54426
rect 7942 54374 7972 54426
rect 7996 54374 8006 54426
rect 8006 54374 8052 54426
rect 7756 54372 7812 54374
rect 7836 54372 7892 54374
rect 7916 54372 7972 54374
rect 7996 54372 8052 54374
rect 7838 54188 7894 54224
rect 7838 54168 7840 54188
rect 7840 54168 7892 54188
rect 7892 54168 7894 54188
rect 7756 53338 7812 53340
rect 7836 53338 7892 53340
rect 7916 53338 7972 53340
rect 7996 53338 8052 53340
rect 7756 53286 7802 53338
rect 7802 53286 7812 53338
rect 7836 53286 7866 53338
rect 7866 53286 7878 53338
rect 7878 53286 7892 53338
rect 7916 53286 7930 53338
rect 7930 53286 7942 53338
rect 7942 53286 7972 53338
rect 7996 53286 8006 53338
rect 8006 53286 8052 53338
rect 7756 53284 7812 53286
rect 7836 53284 7892 53286
rect 7916 53284 7972 53286
rect 7996 53284 8052 53286
rect 7194 52944 7250 53000
rect 6816 52794 6872 52796
rect 6896 52794 6952 52796
rect 6976 52794 7032 52796
rect 7056 52794 7112 52796
rect 6816 52742 6862 52794
rect 6862 52742 6872 52794
rect 6896 52742 6926 52794
rect 6926 52742 6938 52794
rect 6938 52742 6952 52794
rect 6976 52742 6990 52794
rect 6990 52742 7002 52794
rect 7002 52742 7032 52794
rect 7056 52742 7066 52794
rect 7066 52742 7112 52794
rect 6816 52740 6872 52742
rect 6896 52740 6952 52742
rect 6976 52740 7032 52742
rect 7056 52740 7112 52742
rect 6816 51706 6872 51708
rect 6896 51706 6952 51708
rect 6976 51706 7032 51708
rect 7056 51706 7112 51708
rect 6816 51654 6862 51706
rect 6862 51654 6872 51706
rect 6896 51654 6926 51706
rect 6926 51654 6938 51706
rect 6938 51654 6952 51706
rect 6976 51654 6990 51706
rect 6990 51654 7002 51706
rect 7002 51654 7032 51706
rect 7056 51654 7066 51706
rect 7066 51654 7112 51706
rect 6816 51652 6872 51654
rect 6896 51652 6952 51654
rect 6976 51652 7032 51654
rect 7056 51652 7112 51654
rect 7470 52944 7526 53000
rect 7378 52128 7434 52184
rect 7562 51856 7618 51912
rect 6816 50618 6872 50620
rect 6896 50618 6952 50620
rect 6976 50618 7032 50620
rect 7056 50618 7112 50620
rect 6816 50566 6862 50618
rect 6862 50566 6872 50618
rect 6896 50566 6926 50618
rect 6926 50566 6938 50618
rect 6938 50566 6952 50618
rect 6976 50566 6990 50618
rect 6990 50566 7002 50618
rect 7002 50566 7032 50618
rect 7056 50566 7066 50618
rect 7066 50566 7112 50618
rect 6816 50564 6872 50566
rect 6896 50564 6952 50566
rect 6976 50564 7032 50566
rect 7056 50564 7112 50566
rect 6816 49530 6872 49532
rect 6896 49530 6952 49532
rect 6976 49530 7032 49532
rect 7056 49530 7112 49532
rect 6816 49478 6862 49530
rect 6862 49478 6872 49530
rect 6896 49478 6926 49530
rect 6926 49478 6938 49530
rect 6938 49478 6952 49530
rect 6976 49478 6990 49530
rect 6990 49478 7002 49530
rect 7002 49478 7032 49530
rect 7056 49478 7066 49530
rect 7066 49478 7112 49530
rect 6816 49476 6872 49478
rect 6896 49476 6952 49478
rect 6976 49476 7032 49478
rect 7056 49476 7112 49478
rect 6816 48442 6872 48444
rect 6896 48442 6952 48444
rect 6976 48442 7032 48444
rect 7056 48442 7112 48444
rect 6816 48390 6862 48442
rect 6862 48390 6872 48442
rect 6896 48390 6926 48442
rect 6926 48390 6938 48442
rect 6938 48390 6952 48442
rect 6976 48390 6990 48442
rect 6990 48390 7002 48442
rect 7002 48390 7032 48442
rect 7056 48390 7066 48442
rect 7066 48390 7112 48442
rect 6816 48388 6872 48390
rect 6896 48388 6952 48390
rect 6976 48388 7032 48390
rect 7056 48388 7112 48390
rect 6816 47354 6872 47356
rect 6896 47354 6952 47356
rect 6976 47354 7032 47356
rect 7056 47354 7112 47356
rect 6816 47302 6862 47354
rect 6862 47302 6872 47354
rect 6896 47302 6926 47354
rect 6926 47302 6938 47354
rect 6938 47302 6952 47354
rect 6976 47302 6990 47354
rect 6990 47302 7002 47354
rect 7002 47302 7032 47354
rect 7056 47302 7066 47354
rect 7066 47302 7112 47354
rect 6816 47300 6872 47302
rect 6896 47300 6952 47302
rect 6976 47300 7032 47302
rect 7056 47300 7112 47302
rect 7102 46416 7158 46472
rect 6816 46266 6872 46268
rect 6896 46266 6952 46268
rect 6976 46266 7032 46268
rect 7056 46266 7112 46268
rect 6816 46214 6862 46266
rect 6862 46214 6872 46266
rect 6896 46214 6926 46266
rect 6926 46214 6938 46266
rect 6938 46214 6952 46266
rect 6976 46214 6990 46266
rect 6990 46214 7002 46266
rect 7002 46214 7032 46266
rect 7056 46214 7066 46266
rect 7066 46214 7112 46266
rect 6816 46212 6872 46214
rect 6896 46212 6952 46214
rect 6976 46212 7032 46214
rect 7056 46212 7112 46214
rect 6816 45178 6872 45180
rect 6896 45178 6952 45180
rect 6976 45178 7032 45180
rect 7056 45178 7112 45180
rect 6816 45126 6862 45178
rect 6862 45126 6872 45178
rect 6896 45126 6926 45178
rect 6926 45126 6938 45178
rect 6938 45126 6952 45178
rect 6976 45126 6990 45178
rect 6990 45126 7002 45178
rect 7002 45126 7032 45178
rect 7056 45126 7066 45178
rect 7066 45126 7112 45178
rect 6816 45124 6872 45126
rect 6896 45124 6952 45126
rect 6976 45124 7032 45126
rect 7056 45124 7112 45126
rect 6816 44090 6872 44092
rect 6896 44090 6952 44092
rect 6976 44090 7032 44092
rect 7056 44090 7112 44092
rect 6816 44038 6862 44090
rect 6862 44038 6872 44090
rect 6896 44038 6926 44090
rect 6926 44038 6938 44090
rect 6938 44038 6952 44090
rect 6976 44038 6990 44090
rect 6990 44038 7002 44090
rect 7002 44038 7032 44090
rect 7056 44038 7066 44090
rect 7066 44038 7112 44090
rect 6816 44036 6872 44038
rect 6896 44036 6952 44038
rect 6976 44036 7032 44038
rect 7056 44036 7112 44038
rect 6734 43832 6790 43888
rect 7194 43832 7250 43888
rect 6816 43002 6872 43004
rect 6896 43002 6952 43004
rect 6976 43002 7032 43004
rect 7056 43002 7112 43004
rect 6816 42950 6862 43002
rect 6862 42950 6872 43002
rect 6896 42950 6926 43002
rect 6926 42950 6938 43002
rect 6938 42950 6952 43002
rect 6976 42950 6990 43002
rect 6990 42950 7002 43002
rect 7002 42950 7032 43002
rect 7056 42950 7066 43002
rect 7066 42950 7112 43002
rect 6816 42948 6872 42950
rect 6896 42948 6952 42950
rect 6976 42948 7032 42950
rect 7056 42948 7112 42950
rect 7756 52250 7812 52252
rect 7836 52250 7892 52252
rect 7916 52250 7972 52252
rect 7996 52250 8052 52252
rect 7756 52198 7802 52250
rect 7802 52198 7812 52250
rect 7836 52198 7866 52250
rect 7866 52198 7878 52250
rect 7878 52198 7892 52250
rect 7916 52198 7930 52250
rect 7930 52198 7942 52250
rect 7942 52198 7972 52250
rect 7996 52198 8006 52250
rect 8006 52198 8052 52250
rect 7756 52196 7812 52198
rect 7836 52196 7892 52198
rect 7916 52196 7972 52198
rect 7996 52196 8052 52198
rect 7756 51162 7812 51164
rect 7836 51162 7892 51164
rect 7916 51162 7972 51164
rect 7996 51162 8052 51164
rect 7756 51110 7802 51162
rect 7802 51110 7812 51162
rect 7836 51110 7866 51162
rect 7866 51110 7878 51162
rect 7878 51110 7892 51162
rect 7916 51110 7930 51162
rect 7930 51110 7942 51162
rect 7942 51110 7972 51162
rect 7996 51110 8006 51162
rect 8006 51110 8052 51162
rect 7756 51108 7812 51110
rect 7836 51108 7892 51110
rect 7916 51108 7972 51110
rect 7996 51108 8052 51110
rect 7756 50074 7812 50076
rect 7836 50074 7892 50076
rect 7916 50074 7972 50076
rect 7996 50074 8052 50076
rect 7756 50022 7802 50074
rect 7802 50022 7812 50074
rect 7836 50022 7866 50074
rect 7866 50022 7878 50074
rect 7878 50022 7892 50074
rect 7916 50022 7930 50074
rect 7930 50022 7942 50074
rect 7942 50022 7972 50074
rect 7996 50022 8006 50074
rect 8006 50022 8052 50074
rect 7756 50020 7812 50022
rect 7836 50020 7892 50022
rect 7916 50020 7972 50022
rect 7996 50020 8052 50022
rect 8416 54970 8472 54972
rect 8496 54970 8552 54972
rect 8576 54970 8632 54972
rect 8656 54970 8712 54972
rect 8416 54918 8462 54970
rect 8462 54918 8472 54970
rect 8496 54918 8526 54970
rect 8526 54918 8538 54970
rect 8538 54918 8552 54970
rect 8576 54918 8590 54970
rect 8590 54918 8602 54970
rect 8602 54918 8632 54970
rect 8656 54918 8666 54970
rect 8666 54918 8712 54970
rect 8416 54916 8472 54918
rect 8496 54916 8552 54918
rect 8576 54916 8632 54918
rect 8656 54916 8712 54918
rect 8416 53882 8472 53884
rect 8496 53882 8552 53884
rect 8576 53882 8632 53884
rect 8656 53882 8712 53884
rect 8416 53830 8462 53882
rect 8462 53830 8472 53882
rect 8496 53830 8526 53882
rect 8526 53830 8538 53882
rect 8538 53830 8552 53882
rect 8576 53830 8590 53882
rect 8590 53830 8602 53882
rect 8602 53830 8632 53882
rect 8656 53830 8666 53882
rect 8666 53830 8712 53882
rect 8416 53828 8472 53830
rect 8496 53828 8552 53830
rect 8576 53828 8632 53830
rect 8656 53828 8712 53830
rect 8416 52794 8472 52796
rect 8496 52794 8552 52796
rect 8576 52794 8632 52796
rect 8656 52794 8712 52796
rect 8416 52742 8462 52794
rect 8462 52742 8472 52794
rect 8496 52742 8526 52794
rect 8526 52742 8538 52794
rect 8538 52742 8552 52794
rect 8576 52742 8590 52794
rect 8590 52742 8602 52794
rect 8602 52742 8632 52794
rect 8656 52742 8666 52794
rect 8666 52742 8712 52794
rect 8416 52740 8472 52742
rect 8496 52740 8552 52742
rect 8576 52740 8632 52742
rect 8656 52740 8712 52742
rect 8416 51706 8472 51708
rect 8496 51706 8552 51708
rect 8576 51706 8632 51708
rect 8656 51706 8712 51708
rect 8416 51654 8462 51706
rect 8462 51654 8472 51706
rect 8496 51654 8526 51706
rect 8526 51654 8538 51706
rect 8538 51654 8552 51706
rect 8576 51654 8590 51706
rect 8590 51654 8602 51706
rect 8602 51654 8632 51706
rect 8656 51654 8666 51706
rect 8666 51654 8712 51706
rect 8416 51652 8472 51654
rect 8496 51652 8552 51654
rect 8576 51652 8632 51654
rect 8656 51652 8712 51654
rect 7756 48986 7812 48988
rect 7836 48986 7892 48988
rect 7916 48986 7972 48988
rect 7996 48986 8052 48988
rect 7756 48934 7802 48986
rect 7802 48934 7812 48986
rect 7836 48934 7866 48986
rect 7866 48934 7878 48986
rect 7878 48934 7892 48986
rect 7916 48934 7930 48986
rect 7930 48934 7942 48986
rect 7942 48934 7972 48986
rect 7996 48934 8006 48986
rect 8006 48934 8052 48986
rect 7756 48932 7812 48934
rect 7836 48932 7892 48934
rect 7916 48932 7972 48934
rect 7996 48932 8052 48934
rect 7756 47898 7812 47900
rect 7836 47898 7892 47900
rect 7916 47898 7972 47900
rect 7996 47898 8052 47900
rect 7756 47846 7802 47898
rect 7802 47846 7812 47898
rect 7836 47846 7866 47898
rect 7866 47846 7878 47898
rect 7878 47846 7892 47898
rect 7916 47846 7930 47898
rect 7930 47846 7942 47898
rect 7942 47846 7972 47898
rect 7996 47846 8006 47898
rect 8006 47846 8052 47898
rect 7756 47844 7812 47846
rect 7836 47844 7892 47846
rect 7916 47844 7972 47846
rect 7996 47844 8052 47846
rect 7756 46810 7812 46812
rect 7836 46810 7892 46812
rect 7916 46810 7972 46812
rect 7996 46810 8052 46812
rect 7756 46758 7802 46810
rect 7802 46758 7812 46810
rect 7836 46758 7866 46810
rect 7866 46758 7878 46810
rect 7878 46758 7892 46810
rect 7916 46758 7930 46810
rect 7930 46758 7942 46810
rect 7942 46758 7972 46810
rect 7996 46758 8006 46810
rect 8006 46758 8052 46810
rect 7756 46756 7812 46758
rect 7836 46756 7892 46758
rect 7916 46756 7972 46758
rect 7996 46756 8052 46758
rect 9356 63130 9412 63132
rect 9436 63130 9492 63132
rect 9516 63130 9572 63132
rect 9596 63130 9652 63132
rect 9356 63078 9402 63130
rect 9402 63078 9412 63130
rect 9436 63078 9466 63130
rect 9466 63078 9478 63130
rect 9478 63078 9492 63130
rect 9516 63078 9530 63130
rect 9530 63078 9542 63130
rect 9542 63078 9572 63130
rect 9596 63078 9606 63130
rect 9606 63078 9652 63130
rect 9356 63076 9412 63078
rect 9436 63076 9492 63078
rect 9516 63076 9572 63078
rect 9596 63076 9652 63078
rect 10230 71032 10286 71088
rect 9356 62042 9412 62044
rect 9436 62042 9492 62044
rect 9516 62042 9572 62044
rect 9596 62042 9652 62044
rect 9356 61990 9402 62042
rect 9402 61990 9412 62042
rect 9436 61990 9466 62042
rect 9466 61990 9478 62042
rect 9478 61990 9492 62042
rect 9516 61990 9530 62042
rect 9530 61990 9542 62042
rect 9542 61990 9572 62042
rect 9596 61990 9606 62042
rect 9606 61990 9652 62042
rect 9356 61988 9412 61990
rect 9436 61988 9492 61990
rect 9516 61988 9572 61990
rect 9596 61988 9652 61990
rect 9356 60954 9412 60956
rect 9436 60954 9492 60956
rect 9516 60954 9572 60956
rect 9596 60954 9652 60956
rect 9356 60902 9402 60954
rect 9402 60902 9412 60954
rect 9436 60902 9466 60954
rect 9466 60902 9478 60954
rect 9478 60902 9492 60954
rect 9516 60902 9530 60954
rect 9530 60902 9542 60954
rect 9542 60902 9572 60954
rect 9596 60902 9606 60954
rect 9606 60902 9652 60954
rect 9356 60900 9412 60902
rect 9436 60900 9492 60902
rect 9516 60900 9572 60902
rect 9596 60900 9652 60902
rect 8416 50618 8472 50620
rect 8496 50618 8552 50620
rect 8576 50618 8632 50620
rect 8656 50618 8712 50620
rect 8416 50566 8462 50618
rect 8462 50566 8472 50618
rect 8496 50566 8526 50618
rect 8526 50566 8538 50618
rect 8538 50566 8552 50618
rect 8576 50566 8590 50618
rect 8590 50566 8602 50618
rect 8602 50566 8632 50618
rect 8656 50566 8666 50618
rect 8666 50566 8712 50618
rect 8416 50564 8472 50566
rect 8496 50564 8552 50566
rect 8576 50564 8632 50566
rect 8656 50564 8712 50566
rect 8416 49530 8472 49532
rect 8496 49530 8552 49532
rect 8576 49530 8632 49532
rect 8656 49530 8712 49532
rect 8416 49478 8462 49530
rect 8462 49478 8472 49530
rect 8496 49478 8526 49530
rect 8526 49478 8538 49530
rect 8538 49478 8552 49530
rect 8576 49478 8590 49530
rect 8590 49478 8602 49530
rect 8602 49478 8632 49530
rect 8656 49478 8666 49530
rect 8666 49478 8712 49530
rect 8416 49476 8472 49478
rect 8496 49476 8552 49478
rect 8576 49476 8632 49478
rect 8656 49476 8712 49478
rect 8416 48442 8472 48444
rect 8496 48442 8552 48444
rect 8576 48442 8632 48444
rect 8656 48442 8712 48444
rect 8416 48390 8462 48442
rect 8462 48390 8472 48442
rect 8496 48390 8526 48442
rect 8526 48390 8538 48442
rect 8538 48390 8552 48442
rect 8576 48390 8590 48442
rect 8590 48390 8602 48442
rect 8602 48390 8632 48442
rect 8656 48390 8666 48442
rect 8666 48390 8712 48442
rect 8416 48388 8472 48390
rect 8496 48388 8552 48390
rect 8576 48388 8632 48390
rect 8656 48388 8712 48390
rect 8416 47354 8472 47356
rect 8496 47354 8552 47356
rect 8576 47354 8632 47356
rect 8656 47354 8712 47356
rect 8416 47302 8462 47354
rect 8462 47302 8472 47354
rect 8496 47302 8526 47354
rect 8526 47302 8538 47354
rect 8538 47302 8552 47354
rect 8576 47302 8590 47354
rect 8590 47302 8602 47354
rect 8602 47302 8632 47354
rect 8656 47302 8666 47354
rect 8666 47302 8712 47354
rect 8416 47300 8472 47302
rect 8496 47300 8552 47302
rect 8576 47300 8632 47302
rect 8656 47300 8712 47302
rect 8416 46266 8472 46268
rect 8496 46266 8552 46268
rect 8576 46266 8632 46268
rect 8656 46266 8712 46268
rect 8416 46214 8462 46266
rect 8462 46214 8472 46266
rect 8496 46214 8526 46266
rect 8526 46214 8538 46266
rect 8538 46214 8552 46266
rect 8576 46214 8590 46266
rect 8590 46214 8602 46266
rect 8602 46214 8632 46266
rect 8656 46214 8666 46266
rect 8666 46214 8712 46266
rect 8416 46212 8472 46214
rect 8496 46212 8552 46214
rect 8576 46212 8632 46214
rect 8656 46212 8712 46214
rect 7756 45722 7812 45724
rect 7836 45722 7892 45724
rect 7916 45722 7972 45724
rect 7996 45722 8052 45724
rect 7756 45670 7802 45722
rect 7802 45670 7812 45722
rect 7836 45670 7866 45722
rect 7866 45670 7878 45722
rect 7878 45670 7892 45722
rect 7916 45670 7930 45722
rect 7930 45670 7942 45722
rect 7942 45670 7972 45722
rect 7996 45670 8006 45722
rect 8006 45670 8052 45722
rect 7756 45668 7812 45670
rect 7836 45668 7892 45670
rect 7916 45668 7972 45670
rect 7996 45668 8052 45670
rect 8206 45600 8262 45656
rect 7756 44634 7812 44636
rect 7836 44634 7892 44636
rect 7916 44634 7972 44636
rect 7996 44634 8052 44636
rect 7756 44582 7802 44634
rect 7802 44582 7812 44634
rect 7836 44582 7866 44634
rect 7866 44582 7878 44634
rect 7878 44582 7892 44634
rect 7916 44582 7930 44634
rect 7930 44582 7942 44634
rect 7942 44582 7972 44634
rect 7996 44582 8006 44634
rect 8006 44582 8052 44634
rect 7756 44580 7812 44582
rect 7836 44580 7892 44582
rect 7916 44580 7972 44582
rect 7996 44580 8052 44582
rect 6816 41914 6872 41916
rect 6896 41914 6952 41916
rect 6976 41914 7032 41916
rect 7056 41914 7112 41916
rect 6816 41862 6862 41914
rect 6862 41862 6872 41914
rect 6896 41862 6926 41914
rect 6926 41862 6938 41914
rect 6938 41862 6952 41914
rect 6976 41862 6990 41914
rect 6990 41862 7002 41914
rect 7002 41862 7032 41914
rect 7056 41862 7066 41914
rect 7066 41862 7112 41914
rect 6816 41860 6872 41862
rect 6896 41860 6952 41862
rect 6976 41860 7032 41862
rect 7056 41860 7112 41862
rect 6816 40826 6872 40828
rect 6896 40826 6952 40828
rect 6976 40826 7032 40828
rect 7056 40826 7112 40828
rect 6816 40774 6862 40826
rect 6862 40774 6872 40826
rect 6896 40774 6926 40826
rect 6926 40774 6938 40826
rect 6938 40774 6952 40826
rect 6976 40774 6990 40826
rect 6990 40774 7002 40826
rect 7002 40774 7032 40826
rect 7056 40774 7066 40826
rect 7066 40774 7112 40826
rect 6816 40772 6872 40774
rect 6896 40772 6952 40774
rect 6976 40772 7032 40774
rect 7056 40772 7112 40774
rect 6816 39738 6872 39740
rect 6896 39738 6952 39740
rect 6976 39738 7032 39740
rect 7056 39738 7112 39740
rect 6816 39686 6862 39738
rect 6862 39686 6872 39738
rect 6896 39686 6926 39738
rect 6926 39686 6938 39738
rect 6938 39686 6952 39738
rect 6976 39686 6990 39738
rect 6990 39686 7002 39738
rect 7002 39686 7032 39738
rect 7056 39686 7066 39738
rect 7066 39686 7112 39738
rect 6816 39684 6872 39686
rect 6896 39684 6952 39686
rect 6976 39684 7032 39686
rect 7056 39684 7112 39686
rect 6816 38650 6872 38652
rect 6896 38650 6952 38652
rect 6976 38650 7032 38652
rect 7056 38650 7112 38652
rect 6816 38598 6862 38650
rect 6862 38598 6872 38650
rect 6896 38598 6926 38650
rect 6926 38598 6938 38650
rect 6938 38598 6952 38650
rect 6976 38598 6990 38650
rect 6990 38598 7002 38650
rect 7002 38598 7032 38650
rect 7056 38598 7066 38650
rect 7066 38598 7112 38650
rect 6816 38596 6872 38598
rect 6896 38596 6952 38598
rect 6976 38596 7032 38598
rect 7056 38596 7112 38598
rect 6816 37562 6872 37564
rect 6896 37562 6952 37564
rect 6976 37562 7032 37564
rect 7056 37562 7112 37564
rect 6816 37510 6862 37562
rect 6862 37510 6872 37562
rect 6896 37510 6926 37562
rect 6926 37510 6938 37562
rect 6938 37510 6952 37562
rect 6976 37510 6990 37562
rect 6990 37510 7002 37562
rect 7002 37510 7032 37562
rect 7056 37510 7066 37562
rect 7066 37510 7112 37562
rect 6816 37508 6872 37510
rect 6896 37508 6952 37510
rect 6976 37508 7032 37510
rect 7056 37508 7112 37510
rect 6918 37324 6974 37360
rect 6918 37304 6920 37324
rect 6920 37304 6972 37324
rect 6972 37304 6974 37324
rect 6816 36474 6872 36476
rect 6896 36474 6952 36476
rect 6976 36474 7032 36476
rect 7056 36474 7112 36476
rect 6816 36422 6862 36474
rect 6862 36422 6872 36474
rect 6896 36422 6926 36474
rect 6926 36422 6938 36474
rect 6938 36422 6952 36474
rect 6976 36422 6990 36474
rect 6990 36422 7002 36474
rect 7002 36422 7032 36474
rect 7056 36422 7066 36474
rect 7066 36422 7112 36474
rect 6816 36420 6872 36422
rect 6896 36420 6952 36422
rect 6976 36420 7032 36422
rect 7056 36420 7112 36422
rect 6156 35930 6212 35932
rect 6236 35930 6292 35932
rect 6316 35930 6372 35932
rect 6396 35930 6452 35932
rect 6156 35878 6202 35930
rect 6202 35878 6212 35930
rect 6236 35878 6266 35930
rect 6266 35878 6278 35930
rect 6278 35878 6292 35930
rect 6316 35878 6330 35930
rect 6330 35878 6342 35930
rect 6342 35878 6372 35930
rect 6396 35878 6406 35930
rect 6406 35878 6452 35930
rect 6156 35876 6212 35878
rect 6236 35876 6292 35878
rect 6316 35876 6372 35878
rect 6396 35876 6452 35878
rect 6156 34842 6212 34844
rect 6236 34842 6292 34844
rect 6316 34842 6372 34844
rect 6396 34842 6452 34844
rect 6156 34790 6202 34842
rect 6202 34790 6212 34842
rect 6236 34790 6266 34842
rect 6266 34790 6278 34842
rect 6278 34790 6292 34842
rect 6316 34790 6330 34842
rect 6330 34790 6342 34842
rect 6342 34790 6372 34842
rect 6396 34790 6406 34842
rect 6406 34790 6452 34842
rect 6156 34788 6212 34790
rect 6236 34788 6292 34790
rect 6316 34788 6372 34790
rect 6396 34788 6452 34790
rect 6156 33754 6212 33756
rect 6236 33754 6292 33756
rect 6316 33754 6372 33756
rect 6396 33754 6452 33756
rect 6156 33702 6202 33754
rect 6202 33702 6212 33754
rect 6236 33702 6266 33754
rect 6266 33702 6278 33754
rect 6278 33702 6292 33754
rect 6316 33702 6330 33754
rect 6330 33702 6342 33754
rect 6342 33702 6372 33754
rect 6396 33702 6406 33754
rect 6406 33702 6452 33754
rect 6156 33700 6212 33702
rect 6236 33700 6292 33702
rect 6316 33700 6372 33702
rect 6396 33700 6452 33702
rect 6156 32666 6212 32668
rect 6236 32666 6292 32668
rect 6316 32666 6372 32668
rect 6396 32666 6452 32668
rect 6156 32614 6202 32666
rect 6202 32614 6212 32666
rect 6236 32614 6266 32666
rect 6266 32614 6278 32666
rect 6278 32614 6292 32666
rect 6316 32614 6330 32666
rect 6330 32614 6342 32666
rect 6342 32614 6372 32666
rect 6396 32614 6406 32666
rect 6406 32614 6452 32666
rect 6156 32612 6212 32614
rect 6236 32612 6292 32614
rect 6316 32612 6372 32614
rect 6396 32612 6452 32614
rect 5998 31864 6054 31920
rect 6156 31578 6212 31580
rect 6236 31578 6292 31580
rect 6316 31578 6372 31580
rect 6396 31578 6452 31580
rect 6156 31526 6202 31578
rect 6202 31526 6212 31578
rect 6236 31526 6266 31578
rect 6266 31526 6278 31578
rect 6278 31526 6292 31578
rect 6316 31526 6330 31578
rect 6330 31526 6342 31578
rect 6342 31526 6372 31578
rect 6396 31526 6406 31578
rect 6406 31526 6452 31578
rect 6156 31524 6212 31526
rect 6236 31524 6292 31526
rect 6316 31524 6372 31526
rect 6396 31524 6452 31526
rect 5998 31320 6054 31376
rect 6090 30640 6146 30696
rect 6156 30490 6212 30492
rect 6236 30490 6292 30492
rect 6316 30490 6372 30492
rect 6396 30490 6452 30492
rect 6156 30438 6202 30490
rect 6202 30438 6212 30490
rect 6236 30438 6266 30490
rect 6266 30438 6278 30490
rect 6278 30438 6292 30490
rect 6316 30438 6330 30490
rect 6330 30438 6342 30490
rect 6342 30438 6372 30490
rect 6396 30438 6406 30490
rect 6406 30438 6452 30490
rect 6156 30436 6212 30438
rect 6236 30436 6292 30438
rect 6316 30436 6372 30438
rect 6396 30436 6452 30438
rect 6156 29402 6212 29404
rect 6236 29402 6292 29404
rect 6316 29402 6372 29404
rect 6396 29402 6452 29404
rect 6156 29350 6202 29402
rect 6202 29350 6212 29402
rect 6236 29350 6266 29402
rect 6266 29350 6278 29402
rect 6278 29350 6292 29402
rect 6316 29350 6330 29402
rect 6330 29350 6342 29402
rect 6342 29350 6372 29402
rect 6396 29350 6406 29402
rect 6406 29350 6452 29402
rect 6156 29348 6212 29350
rect 6236 29348 6292 29350
rect 6316 29348 6372 29350
rect 6396 29348 6452 29350
rect 6090 29144 6146 29200
rect 5906 28464 5962 28520
rect 5906 28192 5962 28248
rect 6156 28314 6212 28316
rect 6236 28314 6292 28316
rect 6316 28314 6372 28316
rect 6396 28314 6452 28316
rect 6156 28262 6202 28314
rect 6202 28262 6212 28314
rect 6236 28262 6266 28314
rect 6266 28262 6278 28314
rect 6278 28262 6292 28314
rect 6316 28262 6330 28314
rect 6330 28262 6342 28314
rect 6342 28262 6372 28314
rect 6396 28262 6406 28314
rect 6406 28262 6452 28314
rect 6156 28260 6212 28262
rect 6236 28260 6292 28262
rect 6316 28260 6372 28262
rect 6396 28260 6452 28262
rect 6156 27226 6212 27228
rect 6236 27226 6292 27228
rect 6316 27226 6372 27228
rect 6396 27226 6452 27228
rect 6156 27174 6202 27226
rect 6202 27174 6212 27226
rect 6236 27174 6266 27226
rect 6266 27174 6278 27226
rect 6278 27174 6292 27226
rect 6316 27174 6330 27226
rect 6330 27174 6342 27226
rect 6342 27174 6372 27226
rect 6396 27174 6406 27226
rect 6406 27174 6452 27226
rect 6156 27172 6212 27174
rect 6236 27172 6292 27174
rect 6316 27172 6372 27174
rect 6396 27172 6452 27174
rect 6816 35386 6872 35388
rect 6896 35386 6952 35388
rect 6976 35386 7032 35388
rect 7056 35386 7112 35388
rect 6816 35334 6862 35386
rect 6862 35334 6872 35386
rect 6896 35334 6926 35386
rect 6926 35334 6938 35386
rect 6938 35334 6952 35386
rect 6976 35334 6990 35386
rect 6990 35334 7002 35386
rect 7002 35334 7032 35386
rect 7056 35334 7066 35386
rect 7066 35334 7112 35386
rect 6816 35332 6872 35334
rect 6896 35332 6952 35334
rect 6976 35332 7032 35334
rect 7056 35332 7112 35334
rect 6816 34298 6872 34300
rect 6896 34298 6952 34300
rect 6976 34298 7032 34300
rect 7056 34298 7112 34300
rect 6816 34246 6862 34298
rect 6862 34246 6872 34298
rect 6896 34246 6926 34298
rect 6926 34246 6938 34298
rect 6938 34246 6952 34298
rect 6976 34246 6990 34298
rect 6990 34246 7002 34298
rect 7002 34246 7032 34298
rect 7056 34246 7066 34298
rect 7066 34246 7112 34298
rect 6816 34244 6872 34246
rect 6896 34244 6952 34246
rect 6976 34244 7032 34246
rect 7056 34244 7112 34246
rect 7756 43546 7812 43548
rect 7836 43546 7892 43548
rect 7916 43546 7972 43548
rect 7996 43546 8052 43548
rect 7756 43494 7802 43546
rect 7802 43494 7812 43546
rect 7836 43494 7866 43546
rect 7866 43494 7878 43546
rect 7878 43494 7892 43546
rect 7916 43494 7930 43546
rect 7930 43494 7942 43546
rect 7942 43494 7972 43546
rect 7996 43494 8006 43546
rect 8006 43494 8052 43546
rect 7756 43492 7812 43494
rect 7836 43492 7892 43494
rect 7916 43492 7972 43494
rect 7996 43492 8052 43494
rect 7756 42458 7812 42460
rect 7836 42458 7892 42460
rect 7916 42458 7972 42460
rect 7996 42458 8052 42460
rect 7756 42406 7802 42458
rect 7802 42406 7812 42458
rect 7836 42406 7866 42458
rect 7866 42406 7878 42458
rect 7878 42406 7892 42458
rect 7916 42406 7930 42458
rect 7930 42406 7942 42458
rect 7942 42406 7972 42458
rect 7996 42406 8006 42458
rect 8006 42406 8052 42458
rect 7756 42404 7812 42406
rect 7836 42404 7892 42406
rect 7916 42404 7972 42406
rect 7996 42404 8052 42406
rect 7756 41370 7812 41372
rect 7836 41370 7892 41372
rect 7916 41370 7972 41372
rect 7996 41370 8052 41372
rect 7756 41318 7802 41370
rect 7802 41318 7812 41370
rect 7836 41318 7866 41370
rect 7866 41318 7878 41370
rect 7878 41318 7892 41370
rect 7916 41318 7930 41370
rect 7930 41318 7942 41370
rect 7942 41318 7972 41370
rect 7996 41318 8006 41370
rect 8006 41318 8052 41370
rect 7756 41316 7812 41318
rect 7836 41316 7892 41318
rect 7916 41316 7972 41318
rect 7996 41316 8052 41318
rect 9356 59866 9412 59868
rect 9436 59866 9492 59868
rect 9516 59866 9572 59868
rect 9596 59866 9652 59868
rect 9356 59814 9402 59866
rect 9402 59814 9412 59866
rect 9436 59814 9466 59866
rect 9466 59814 9478 59866
rect 9478 59814 9492 59866
rect 9516 59814 9530 59866
rect 9530 59814 9542 59866
rect 9542 59814 9572 59866
rect 9596 59814 9606 59866
rect 9606 59814 9652 59866
rect 9356 59812 9412 59814
rect 9436 59812 9492 59814
rect 9516 59812 9572 59814
rect 9596 59812 9652 59814
rect 9356 58778 9412 58780
rect 9436 58778 9492 58780
rect 9516 58778 9572 58780
rect 9596 58778 9652 58780
rect 9356 58726 9402 58778
rect 9402 58726 9412 58778
rect 9436 58726 9466 58778
rect 9466 58726 9478 58778
rect 9478 58726 9492 58778
rect 9516 58726 9530 58778
rect 9530 58726 9542 58778
rect 9542 58726 9572 58778
rect 9596 58726 9606 58778
rect 9606 58726 9652 58778
rect 9356 58724 9412 58726
rect 9436 58724 9492 58726
rect 9516 58724 9572 58726
rect 9596 58724 9652 58726
rect 9310 57840 9366 57896
rect 9356 57690 9412 57692
rect 9436 57690 9492 57692
rect 9516 57690 9572 57692
rect 9596 57690 9652 57692
rect 9356 57638 9402 57690
rect 9402 57638 9412 57690
rect 9436 57638 9466 57690
rect 9466 57638 9478 57690
rect 9478 57638 9492 57690
rect 9516 57638 9530 57690
rect 9530 57638 9542 57690
rect 9542 57638 9572 57690
rect 9596 57638 9606 57690
rect 9606 57638 9652 57690
rect 9356 57636 9412 57638
rect 9436 57636 9492 57638
rect 9516 57636 9572 57638
rect 9596 57636 9652 57638
rect 9356 56602 9412 56604
rect 9436 56602 9492 56604
rect 9516 56602 9572 56604
rect 9596 56602 9652 56604
rect 9356 56550 9402 56602
rect 9402 56550 9412 56602
rect 9436 56550 9466 56602
rect 9466 56550 9478 56602
rect 9478 56550 9492 56602
rect 9516 56550 9530 56602
rect 9530 56550 9542 56602
rect 9542 56550 9572 56602
rect 9596 56550 9606 56602
rect 9606 56550 9652 56602
rect 9356 56548 9412 56550
rect 9436 56548 9492 56550
rect 9516 56548 9572 56550
rect 9596 56548 9652 56550
rect 9356 55514 9412 55516
rect 9436 55514 9492 55516
rect 9516 55514 9572 55516
rect 9596 55514 9652 55516
rect 9356 55462 9402 55514
rect 9402 55462 9412 55514
rect 9436 55462 9466 55514
rect 9466 55462 9478 55514
rect 9478 55462 9492 55514
rect 9516 55462 9530 55514
rect 9530 55462 9542 55514
rect 9542 55462 9572 55514
rect 9596 55462 9606 55514
rect 9606 55462 9652 55514
rect 9356 55460 9412 55462
rect 9436 55460 9492 55462
rect 9516 55460 9572 55462
rect 9596 55460 9652 55462
rect 9356 54426 9412 54428
rect 9436 54426 9492 54428
rect 9516 54426 9572 54428
rect 9596 54426 9652 54428
rect 9356 54374 9402 54426
rect 9402 54374 9412 54426
rect 9436 54374 9466 54426
rect 9466 54374 9478 54426
rect 9478 54374 9492 54426
rect 9516 54374 9530 54426
rect 9530 54374 9542 54426
rect 9542 54374 9572 54426
rect 9596 54374 9606 54426
rect 9606 54374 9652 54426
rect 9356 54372 9412 54374
rect 9436 54372 9492 54374
rect 9516 54372 9572 54374
rect 9596 54372 9652 54374
rect 9356 53338 9412 53340
rect 9436 53338 9492 53340
rect 9516 53338 9572 53340
rect 9596 53338 9652 53340
rect 9356 53286 9402 53338
rect 9402 53286 9412 53338
rect 9436 53286 9466 53338
rect 9466 53286 9478 53338
rect 9478 53286 9492 53338
rect 9516 53286 9530 53338
rect 9530 53286 9542 53338
rect 9542 53286 9572 53338
rect 9596 53286 9606 53338
rect 9606 53286 9652 53338
rect 9356 53284 9412 53286
rect 9436 53284 9492 53286
rect 9516 53284 9572 53286
rect 9596 53284 9652 53286
rect 9356 52250 9412 52252
rect 9436 52250 9492 52252
rect 9516 52250 9572 52252
rect 9596 52250 9652 52252
rect 9356 52198 9402 52250
rect 9402 52198 9412 52250
rect 9436 52198 9466 52250
rect 9466 52198 9478 52250
rect 9478 52198 9492 52250
rect 9516 52198 9530 52250
rect 9530 52198 9542 52250
rect 9542 52198 9572 52250
rect 9596 52198 9606 52250
rect 9606 52198 9652 52250
rect 9356 52196 9412 52198
rect 9436 52196 9492 52198
rect 9516 52196 9572 52198
rect 9596 52196 9652 52198
rect 9356 51162 9412 51164
rect 9436 51162 9492 51164
rect 9516 51162 9572 51164
rect 9596 51162 9652 51164
rect 9356 51110 9402 51162
rect 9402 51110 9412 51162
rect 9436 51110 9466 51162
rect 9466 51110 9478 51162
rect 9478 51110 9492 51162
rect 9516 51110 9530 51162
rect 9530 51110 9542 51162
rect 9542 51110 9572 51162
rect 9596 51110 9606 51162
rect 9606 51110 9652 51162
rect 9356 51108 9412 51110
rect 9436 51108 9492 51110
rect 9516 51108 9572 51110
rect 9596 51108 9652 51110
rect 9494 50224 9550 50280
rect 9356 50074 9412 50076
rect 9436 50074 9492 50076
rect 9516 50074 9572 50076
rect 9596 50074 9652 50076
rect 9356 50022 9402 50074
rect 9402 50022 9412 50074
rect 9436 50022 9466 50074
rect 9466 50022 9478 50074
rect 9478 50022 9492 50074
rect 9516 50022 9530 50074
rect 9530 50022 9542 50074
rect 9542 50022 9572 50074
rect 9596 50022 9606 50074
rect 9606 50022 9652 50074
rect 9356 50020 9412 50022
rect 9436 50020 9492 50022
rect 9516 50020 9572 50022
rect 9596 50020 9652 50022
rect 8416 45178 8472 45180
rect 8496 45178 8552 45180
rect 8576 45178 8632 45180
rect 8656 45178 8712 45180
rect 8416 45126 8462 45178
rect 8462 45126 8472 45178
rect 8496 45126 8526 45178
rect 8526 45126 8538 45178
rect 8538 45126 8552 45178
rect 8576 45126 8590 45178
rect 8590 45126 8602 45178
rect 8602 45126 8632 45178
rect 8656 45126 8666 45178
rect 8666 45126 8712 45178
rect 8416 45124 8472 45126
rect 8496 45124 8552 45126
rect 8576 45124 8632 45126
rect 8656 45124 8712 45126
rect 8416 44090 8472 44092
rect 8496 44090 8552 44092
rect 8576 44090 8632 44092
rect 8656 44090 8712 44092
rect 8416 44038 8462 44090
rect 8462 44038 8472 44090
rect 8496 44038 8526 44090
rect 8526 44038 8538 44090
rect 8538 44038 8552 44090
rect 8576 44038 8590 44090
rect 8590 44038 8602 44090
rect 8602 44038 8632 44090
rect 8656 44038 8666 44090
rect 8666 44038 8712 44090
rect 8416 44036 8472 44038
rect 8496 44036 8552 44038
rect 8576 44036 8632 44038
rect 8656 44036 8712 44038
rect 8416 43002 8472 43004
rect 8496 43002 8552 43004
rect 8576 43002 8632 43004
rect 8656 43002 8712 43004
rect 8416 42950 8462 43002
rect 8462 42950 8472 43002
rect 8496 42950 8526 43002
rect 8526 42950 8538 43002
rect 8538 42950 8552 43002
rect 8576 42950 8590 43002
rect 8590 42950 8602 43002
rect 8602 42950 8632 43002
rect 8656 42950 8666 43002
rect 8666 42950 8712 43002
rect 8416 42948 8472 42950
rect 8496 42948 8552 42950
rect 8576 42948 8632 42950
rect 8656 42948 8712 42950
rect 7756 40282 7812 40284
rect 7836 40282 7892 40284
rect 7916 40282 7972 40284
rect 7996 40282 8052 40284
rect 7756 40230 7802 40282
rect 7802 40230 7812 40282
rect 7836 40230 7866 40282
rect 7866 40230 7878 40282
rect 7878 40230 7892 40282
rect 7916 40230 7930 40282
rect 7930 40230 7942 40282
rect 7942 40230 7972 40282
rect 7996 40230 8006 40282
rect 8006 40230 8052 40282
rect 7756 40228 7812 40230
rect 7836 40228 7892 40230
rect 7916 40228 7972 40230
rect 7996 40228 8052 40230
rect 9356 48986 9412 48988
rect 9436 48986 9492 48988
rect 9516 48986 9572 48988
rect 9596 48986 9652 48988
rect 9356 48934 9402 48986
rect 9402 48934 9412 48986
rect 9436 48934 9466 48986
rect 9466 48934 9478 48986
rect 9478 48934 9492 48986
rect 9516 48934 9530 48986
rect 9530 48934 9542 48986
rect 9542 48934 9572 48986
rect 9596 48934 9606 48986
rect 9606 48934 9652 48986
rect 9356 48932 9412 48934
rect 9436 48932 9492 48934
rect 9516 48932 9572 48934
rect 9596 48932 9652 48934
rect 9310 48728 9366 48784
rect 9310 48048 9366 48104
rect 9356 47898 9412 47900
rect 9436 47898 9492 47900
rect 9516 47898 9572 47900
rect 9596 47898 9652 47900
rect 9356 47846 9402 47898
rect 9402 47846 9412 47898
rect 9436 47846 9466 47898
rect 9466 47846 9478 47898
rect 9478 47846 9492 47898
rect 9516 47846 9530 47898
rect 9530 47846 9542 47898
rect 9542 47846 9572 47898
rect 9596 47846 9606 47898
rect 9606 47846 9652 47898
rect 9356 47844 9412 47846
rect 9436 47844 9492 47846
rect 9516 47844 9572 47846
rect 9596 47844 9652 47846
rect 8942 42608 8998 42664
rect 8416 41914 8472 41916
rect 8496 41914 8552 41916
rect 8576 41914 8632 41916
rect 8656 41914 8712 41916
rect 8416 41862 8462 41914
rect 8462 41862 8472 41914
rect 8496 41862 8526 41914
rect 8526 41862 8538 41914
rect 8538 41862 8552 41914
rect 8576 41862 8590 41914
rect 8590 41862 8602 41914
rect 8602 41862 8632 41914
rect 8656 41862 8666 41914
rect 8666 41862 8712 41914
rect 8416 41860 8472 41862
rect 8496 41860 8552 41862
rect 8576 41860 8632 41862
rect 8656 41860 8712 41862
rect 8416 40826 8472 40828
rect 8496 40826 8552 40828
rect 8576 40826 8632 40828
rect 8656 40826 8712 40828
rect 8416 40774 8462 40826
rect 8462 40774 8472 40826
rect 8496 40774 8526 40826
rect 8526 40774 8538 40826
rect 8538 40774 8552 40826
rect 8576 40774 8590 40826
rect 8590 40774 8602 40826
rect 8602 40774 8632 40826
rect 8656 40774 8666 40826
rect 8666 40774 8712 40826
rect 8416 40772 8472 40774
rect 8496 40772 8552 40774
rect 8576 40772 8632 40774
rect 8656 40772 8712 40774
rect 7838 39888 7894 39944
rect 6816 33210 6872 33212
rect 6896 33210 6952 33212
rect 6976 33210 7032 33212
rect 7056 33210 7112 33212
rect 6816 33158 6862 33210
rect 6862 33158 6872 33210
rect 6896 33158 6926 33210
rect 6926 33158 6938 33210
rect 6938 33158 6952 33210
rect 6976 33158 6990 33210
rect 6990 33158 7002 33210
rect 7002 33158 7032 33210
rect 7056 33158 7066 33210
rect 7066 33158 7112 33210
rect 6816 33156 6872 33158
rect 6896 33156 6952 33158
rect 6976 33156 7032 33158
rect 7056 33156 7112 33158
rect 6816 32122 6872 32124
rect 6896 32122 6952 32124
rect 6976 32122 7032 32124
rect 7056 32122 7112 32124
rect 6816 32070 6862 32122
rect 6862 32070 6872 32122
rect 6896 32070 6926 32122
rect 6926 32070 6938 32122
rect 6938 32070 6952 32122
rect 6976 32070 6990 32122
rect 6990 32070 7002 32122
rect 7002 32070 7032 32122
rect 7056 32070 7066 32122
rect 7066 32070 7112 32122
rect 6816 32068 6872 32070
rect 6896 32068 6952 32070
rect 6976 32068 7032 32070
rect 7056 32068 7112 32070
rect 7010 31864 7066 31920
rect 7286 32272 7342 32328
rect 7756 39194 7812 39196
rect 7836 39194 7892 39196
rect 7916 39194 7972 39196
rect 7996 39194 8052 39196
rect 7756 39142 7802 39194
rect 7802 39142 7812 39194
rect 7836 39142 7866 39194
rect 7866 39142 7878 39194
rect 7878 39142 7892 39194
rect 7916 39142 7930 39194
rect 7930 39142 7942 39194
rect 7942 39142 7972 39194
rect 7996 39142 8006 39194
rect 8006 39142 8052 39194
rect 7756 39140 7812 39142
rect 7836 39140 7892 39142
rect 7916 39140 7972 39142
rect 7996 39140 8052 39142
rect 8206 38392 8262 38448
rect 7756 38106 7812 38108
rect 7836 38106 7892 38108
rect 7916 38106 7972 38108
rect 7996 38106 8052 38108
rect 7756 38054 7802 38106
rect 7802 38054 7812 38106
rect 7836 38054 7866 38106
rect 7866 38054 7878 38106
rect 7878 38054 7892 38106
rect 7916 38054 7930 38106
rect 7930 38054 7942 38106
rect 7942 38054 7972 38106
rect 7996 38054 8006 38106
rect 8006 38054 8052 38106
rect 7756 38052 7812 38054
rect 7836 38052 7892 38054
rect 7916 38052 7972 38054
rect 7996 38052 8052 38054
rect 7756 37018 7812 37020
rect 7836 37018 7892 37020
rect 7916 37018 7972 37020
rect 7996 37018 8052 37020
rect 7756 36966 7802 37018
rect 7802 36966 7812 37018
rect 7836 36966 7866 37018
rect 7866 36966 7878 37018
rect 7878 36966 7892 37018
rect 7916 36966 7930 37018
rect 7930 36966 7942 37018
rect 7942 36966 7972 37018
rect 7996 36966 8006 37018
rect 8006 36966 8052 37018
rect 7756 36964 7812 36966
rect 7836 36964 7892 36966
rect 7916 36964 7972 36966
rect 7996 36964 8052 36966
rect 7756 35930 7812 35932
rect 7836 35930 7892 35932
rect 7916 35930 7972 35932
rect 7996 35930 8052 35932
rect 7756 35878 7802 35930
rect 7802 35878 7812 35930
rect 7836 35878 7866 35930
rect 7866 35878 7878 35930
rect 7878 35878 7892 35930
rect 7916 35878 7930 35930
rect 7930 35878 7942 35930
rect 7942 35878 7972 35930
rect 7996 35878 8006 35930
rect 8006 35878 8052 35930
rect 7756 35876 7812 35878
rect 7836 35876 7892 35878
rect 7916 35876 7972 35878
rect 7996 35876 8052 35878
rect 7756 34842 7812 34844
rect 7836 34842 7892 34844
rect 7916 34842 7972 34844
rect 7996 34842 8052 34844
rect 7756 34790 7802 34842
rect 7802 34790 7812 34842
rect 7836 34790 7866 34842
rect 7866 34790 7878 34842
rect 7878 34790 7892 34842
rect 7916 34790 7930 34842
rect 7930 34790 7942 34842
rect 7942 34790 7972 34842
rect 7996 34790 8006 34842
rect 8006 34790 8052 34842
rect 7756 34788 7812 34790
rect 7836 34788 7892 34790
rect 7916 34788 7972 34790
rect 7996 34788 8052 34790
rect 7756 33754 7812 33756
rect 7836 33754 7892 33756
rect 7916 33754 7972 33756
rect 7996 33754 8052 33756
rect 7756 33702 7802 33754
rect 7802 33702 7812 33754
rect 7836 33702 7866 33754
rect 7866 33702 7878 33754
rect 7878 33702 7892 33754
rect 7916 33702 7930 33754
rect 7930 33702 7942 33754
rect 7942 33702 7972 33754
rect 7996 33702 8006 33754
rect 8006 33702 8052 33754
rect 7756 33700 7812 33702
rect 7836 33700 7892 33702
rect 7916 33700 7972 33702
rect 7996 33700 8052 33702
rect 8416 39738 8472 39740
rect 8496 39738 8552 39740
rect 8576 39738 8632 39740
rect 8656 39738 8712 39740
rect 8416 39686 8462 39738
rect 8462 39686 8472 39738
rect 8496 39686 8526 39738
rect 8526 39686 8538 39738
rect 8538 39686 8552 39738
rect 8576 39686 8590 39738
rect 8590 39686 8602 39738
rect 8602 39686 8632 39738
rect 8656 39686 8666 39738
rect 8666 39686 8712 39738
rect 8416 39684 8472 39686
rect 8496 39684 8552 39686
rect 8576 39684 8632 39686
rect 8656 39684 8712 39686
rect 8416 38650 8472 38652
rect 8496 38650 8552 38652
rect 8576 38650 8632 38652
rect 8656 38650 8712 38652
rect 8416 38598 8462 38650
rect 8462 38598 8472 38650
rect 8496 38598 8526 38650
rect 8526 38598 8538 38650
rect 8538 38598 8552 38650
rect 8576 38598 8590 38650
rect 8590 38598 8602 38650
rect 8602 38598 8632 38650
rect 8656 38598 8666 38650
rect 8666 38598 8712 38650
rect 8416 38596 8472 38598
rect 8496 38596 8552 38598
rect 8576 38596 8632 38598
rect 8656 38596 8712 38598
rect 8416 37562 8472 37564
rect 8496 37562 8552 37564
rect 8576 37562 8632 37564
rect 8656 37562 8712 37564
rect 8416 37510 8462 37562
rect 8462 37510 8472 37562
rect 8496 37510 8526 37562
rect 8526 37510 8538 37562
rect 8538 37510 8552 37562
rect 8576 37510 8590 37562
rect 8590 37510 8602 37562
rect 8602 37510 8632 37562
rect 8656 37510 8666 37562
rect 8666 37510 8712 37562
rect 8416 37508 8472 37510
rect 8496 37508 8552 37510
rect 8576 37508 8632 37510
rect 8656 37508 8712 37510
rect 8298 36760 8354 36816
rect 8416 36474 8472 36476
rect 8496 36474 8552 36476
rect 8576 36474 8632 36476
rect 8656 36474 8712 36476
rect 8416 36422 8462 36474
rect 8462 36422 8472 36474
rect 8496 36422 8526 36474
rect 8526 36422 8538 36474
rect 8538 36422 8552 36474
rect 8576 36422 8590 36474
rect 8590 36422 8602 36474
rect 8602 36422 8632 36474
rect 8656 36422 8666 36474
rect 8666 36422 8712 36474
rect 8416 36420 8472 36422
rect 8496 36420 8552 36422
rect 8576 36420 8632 36422
rect 8656 36420 8712 36422
rect 8416 35386 8472 35388
rect 8496 35386 8552 35388
rect 8576 35386 8632 35388
rect 8656 35386 8712 35388
rect 8416 35334 8462 35386
rect 8462 35334 8472 35386
rect 8496 35334 8526 35386
rect 8526 35334 8538 35386
rect 8538 35334 8552 35386
rect 8576 35334 8590 35386
rect 8590 35334 8602 35386
rect 8602 35334 8632 35386
rect 8656 35334 8666 35386
rect 8666 35334 8712 35386
rect 8416 35332 8472 35334
rect 8496 35332 8552 35334
rect 8576 35332 8632 35334
rect 8656 35332 8712 35334
rect 8298 35128 8354 35184
rect 8416 34298 8472 34300
rect 8496 34298 8552 34300
rect 8576 34298 8632 34300
rect 8656 34298 8712 34300
rect 8416 34246 8462 34298
rect 8462 34246 8472 34298
rect 8496 34246 8526 34298
rect 8526 34246 8538 34298
rect 8538 34246 8552 34298
rect 8576 34246 8590 34298
rect 8590 34246 8602 34298
rect 8602 34246 8632 34298
rect 8656 34246 8666 34298
rect 8666 34246 8712 34298
rect 8416 34244 8472 34246
rect 8496 34244 8552 34246
rect 8576 34244 8632 34246
rect 8656 34244 8712 34246
rect 7756 32666 7812 32668
rect 7836 32666 7892 32668
rect 7916 32666 7972 32668
rect 7996 32666 8052 32668
rect 7756 32614 7802 32666
rect 7802 32614 7812 32666
rect 7836 32614 7866 32666
rect 7866 32614 7878 32666
rect 7878 32614 7892 32666
rect 7916 32614 7930 32666
rect 7930 32614 7942 32666
rect 7942 32614 7972 32666
rect 7996 32614 8006 32666
rect 8006 32614 8052 32666
rect 7756 32612 7812 32614
rect 7836 32612 7892 32614
rect 7916 32612 7972 32614
rect 7996 32612 8052 32614
rect 6816 31034 6872 31036
rect 6896 31034 6952 31036
rect 6976 31034 7032 31036
rect 7056 31034 7112 31036
rect 6816 30982 6862 31034
rect 6862 30982 6872 31034
rect 6896 30982 6926 31034
rect 6926 30982 6938 31034
rect 6938 30982 6952 31034
rect 6976 30982 6990 31034
rect 6990 30982 7002 31034
rect 7002 30982 7032 31034
rect 7056 30982 7066 31034
rect 7066 30982 7112 31034
rect 6816 30980 6872 30982
rect 6896 30980 6952 30982
rect 6976 30980 7032 30982
rect 7056 30980 7112 30982
rect 6816 29946 6872 29948
rect 6896 29946 6952 29948
rect 6976 29946 7032 29948
rect 7056 29946 7112 29948
rect 6816 29894 6862 29946
rect 6862 29894 6872 29946
rect 6896 29894 6926 29946
rect 6926 29894 6938 29946
rect 6938 29894 6952 29946
rect 6976 29894 6990 29946
rect 6990 29894 7002 29946
rect 7002 29894 7032 29946
rect 7056 29894 7066 29946
rect 7066 29894 7112 29946
rect 6816 29892 6872 29894
rect 6896 29892 6952 29894
rect 6976 29892 7032 29894
rect 7056 29892 7112 29894
rect 6816 28858 6872 28860
rect 6896 28858 6952 28860
rect 6976 28858 7032 28860
rect 7056 28858 7112 28860
rect 6816 28806 6862 28858
rect 6862 28806 6872 28858
rect 6896 28806 6926 28858
rect 6926 28806 6938 28858
rect 6938 28806 6952 28858
rect 6976 28806 6990 28858
rect 6990 28806 7002 28858
rect 7002 28806 7032 28858
rect 7056 28806 7066 28858
rect 7066 28806 7112 28858
rect 6816 28804 6872 28806
rect 6896 28804 6952 28806
rect 6976 28804 7032 28806
rect 7056 28804 7112 28806
rect 7010 27920 7066 27976
rect 6816 27770 6872 27772
rect 6896 27770 6952 27772
rect 6976 27770 7032 27772
rect 7056 27770 7112 27772
rect 6816 27718 6862 27770
rect 6862 27718 6872 27770
rect 6896 27718 6926 27770
rect 6926 27718 6938 27770
rect 6938 27718 6952 27770
rect 6976 27718 6990 27770
rect 6990 27718 7002 27770
rect 7002 27718 7032 27770
rect 7056 27718 7066 27770
rect 7066 27718 7112 27770
rect 6816 27716 6872 27718
rect 6896 27716 6952 27718
rect 6976 27716 7032 27718
rect 7056 27716 7112 27718
rect 6090 26288 6146 26344
rect 6156 26138 6212 26140
rect 6236 26138 6292 26140
rect 6316 26138 6372 26140
rect 6396 26138 6452 26140
rect 6156 26086 6202 26138
rect 6202 26086 6212 26138
rect 6236 26086 6266 26138
rect 6266 26086 6278 26138
rect 6278 26086 6292 26138
rect 6316 26086 6330 26138
rect 6330 26086 6342 26138
rect 6342 26086 6372 26138
rect 6396 26086 6406 26138
rect 6406 26086 6452 26138
rect 6156 26084 6212 26086
rect 6236 26084 6292 26086
rect 6316 26084 6372 26086
rect 6396 26084 6452 26086
rect 5814 25900 5870 25936
rect 5814 25880 5816 25900
rect 5816 25880 5868 25900
rect 5868 25880 5870 25900
rect 5216 10362 5272 10364
rect 5296 10362 5352 10364
rect 5376 10362 5432 10364
rect 5456 10362 5512 10364
rect 5216 10310 5262 10362
rect 5262 10310 5272 10362
rect 5296 10310 5326 10362
rect 5326 10310 5338 10362
rect 5338 10310 5352 10362
rect 5376 10310 5390 10362
rect 5390 10310 5402 10362
rect 5402 10310 5432 10362
rect 5456 10310 5466 10362
rect 5466 10310 5512 10362
rect 5216 10308 5272 10310
rect 5296 10308 5352 10310
rect 5376 10308 5432 10310
rect 5456 10308 5512 10310
rect 5216 9274 5272 9276
rect 5296 9274 5352 9276
rect 5376 9274 5432 9276
rect 5456 9274 5512 9276
rect 5216 9222 5262 9274
rect 5262 9222 5272 9274
rect 5296 9222 5326 9274
rect 5326 9222 5338 9274
rect 5338 9222 5352 9274
rect 5376 9222 5390 9274
rect 5390 9222 5402 9274
rect 5402 9222 5432 9274
rect 5456 9222 5466 9274
rect 5466 9222 5512 9274
rect 5216 9220 5272 9222
rect 5296 9220 5352 9222
rect 5376 9220 5432 9222
rect 5456 9220 5512 9222
rect 5216 8186 5272 8188
rect 5296 8186 5352 8188
rect 5376 8186 5432 8188
rect 5456 8186 5512 8188
rect 5216 8134 5262 8186
rect 5262 8134 5272 8186
rect 5296 8134 5326 8186
rect 5326 8134 5338 8186
rect 5338 8134 5352 8186
rect 5376 8134 5390 8186
rect 5390 8134 5402 8186
rect 5402 8134 5432 8186
rect 5456 8134 5466 8186
rect 5466 8134 5512 8186
rect 5216 8132 5272 8134
rect 5296 8132 5352 8134
rect 5376 8132 5432 8134
rect 5456 8132 5512 8134
rect 5216 7098 5272 7100
rect 5296 7098 5352 7100
rect 5376 7098 5432 7100
rect 5456 7098 5512 7100
rect 5216 7046 5262 7098
rect 5262 7046 5272 7098
rect 5296 7046 5326 7098
rect 5326 7046 5338 7098
rect 5338 7046 5352 7098
rect 5376 7046 5390 7098
rect 5390 7046 5402 7098
rect 5402 7046 5432 7098
rect 5456 7046 5466 7098
rect 5466 7046 5512 7098
rect 5216 7044 5272 7046
rect 5296 7044 5352 7046
rect 5376 7044 5432 7046
rect 5456 7044 5512 7046
rect 5216 6010 5272 6012
rect 5296 6010 5352 6012
rect 5376 6010 5432 6012
rect 5456 6010 5512 6012
rect 5216 5958 5262 6010
rect 5262 5958 5272 6010
rect 5296 5958 5326 6010
rect 5326 5958 5338 6010
rect 5338 5958 5352 6010
rect 5376 5958 5390 6010
rect 5390 5958 5402 6010
rect 5402 5958 5432 6010
rect 5456 5958 5466 6010
rect 5466 5958 5512 6010
rect 5216 5956 5272 5958
rect 5296 5956 5352 5958
rect 5376 5956 5432 5958
rect 5456 5956 5512 5958
rect 5216 4922 5272 4924
rect 5296 4922 5352 4924
rect 5376 4922 5432 4924
rect 5456 4922 5512 4924
rect 5216 4870 5262 4922
rect 5262 4870 5272 4922
rect 5296 4870 5326 4922
rect 5326 4870 5338 4922
rect 5338 4870 5352 4922
rect 5376 4870 5390 4922
rect 5390 4870 5402 4922
rect 5402 4870 5432 4922
rect 5456 4870 5466 4922
rect 5466 4870 5512 4922
rect 5216 4868 5272 4870
rect 5296 4868 5352 4870
rect 5376 4868 5432 4870
rect 5456 4868 5512 4870
rect 5216 3834 5272 3836
rect 5296 3834 5352 3836
rect 5376 3834 5432 3836
rect 5456 3834 5512 3836
rect 5216 3782 5262 3834
rect 5262 3782 5272 3834
rect 5296 3782 5326 3834
rect 5326 3782 5338 3834
rect 5338 3782 5352 3834
rect 5376 3782 5390 3834
rect 5390 3782 5402 3834
rect 5402 3782 5432 3834
rect 5456 3782 5466 3834
rect 5466 3782 5512 3834
rect 5216 3780 5272 3782
rect 5296 3780 5352 3782
rect 5376 3780 5432 3782
rect 5456 3780 5512 3782
rect 5216 2746 5272 2748
rect 5296 2746 5352 2748
rect 5376 2746 5432 2748
rect 5456 2746 5512 2748
rect 5216 2694 5262 2746
rect 5262 2694 5272 2746
rect 5296 2694 5326 2746
rect 5326 2694 5338 2746
rect 5338 2694 5352 2746
rect 5376 2694 5390 2746
rect 5390 2694 5402 2746
rect 5402 2694 5432 2746
rect 5456 2694 5466 2746
rect 5466 2694 5512 2746
rect 5216 2692 5272 2694
rect 5296 2692 5352 2694
rect 5376 2692 5432 2694
rect 5456 2692 5512 2694
rect 5216 1658 5272 1660
rect 5296 1658 5352 1660
rect 5376 1658 5432 1660
rect 5456 1658 5512 1660
rect 5216 1606 5262 1658
rect 5262 1606 5272 1658
rect 5296 1606 5326 1658
rect 5326 1606 5338 1658
rect 5338 1606 5352 1658
rect 5376 1606 5390 1658
rect 5390 1606 5402 1658
rect 5402 1606 5432 1658
rect 5456 1606 5466 1658
rect 5466 1606 5512 1658
rect 5216 1604 5272 1606
rect 5296 1604 5352 1606
rect 5376 1604 5432 1606
rect 5456 1604 5512 1606
rect 5722 3440 5778 3496
rect 6156 25050 6212 25052
rect 6236 25050 6292 25052
rect 6316 25050 6372 25052
rect 6396 25050 6452 25052
rect 6156 24998 6202 25050
rect 6202 24998 6212 25050
rect 6236 24998 6266 25050
rect 6266 24998 6278 25050
rect 6278 24998 6292 25050
rect 6316 24998 6330 25050
rect 6330 24998 6342 25050
rect 6342 24998 6372 25050
rect 6396 24998 6406 25050
rect 6406 24998 6452 25050
rect 6156 24996 6212 24998
rect 6236 24996 6292 24998
rect 6316 24996 6372 24998
rect 6396 24996 6452 24998
rect 6156 23962 6212 23964
rect 6236 23962 6292 23964
rect 6316 23962 6372 23964
rect 6396 23962 6452 23964
rect 6156 23910 6202 23962
rect 6202 23910 6212 23962
rect 6236 23910 6266 23962
rect 6266 23910 6278 23962
rect 6278 23910 6292 23962
rect 6316 23910 6330 23962
rect 6330 23910 6342 23962
rect 6342 23910 6372 23962
rect 6396 23910 6406 23962
rect 6406 23910 6452 23962
rect 6156 23908 6212 23910
rect 6236 23908 6292 23910
rect 6316 23908 6372 23910
rect 6396 23908 6452 23910
rect 6156 22874 6212 22876
rect 6236 22874 6292 22876
rect 6316 22874 6372 22876
rect 6396 22874 6452 22876
rect 6156 22822 6202 22874
rect 6202 22822 6212 22874
rect 6236 22822 6266 22874
rect 6266 22822 6278 22874
rect 6278 22822 6292 22874
rect 6316 22822 6330 22874
rect 6330 22822 6342 22874
rect 6342 22822 6372 22874
rect 6396 22822 6406 22874
rect 6406 22822 6452 22874
rect 6156 22820 6212 22822
rect 6236 22820 6292 22822
rect 6316 22820 6372 22822
rect 6396 22820 6452 22822
rect 6156 21786 6212 21788
rect 6236 21786 6292 21788
rect 6316 21786 6372 21788
rect 6396 21786 6452 21788
rect 6156 21734 6202 21786
rect 6202 21734 6212 21786
rect 6236 21734 6266 21786
rect 6266 21734 6278 21786
rect 6278 21734 6292 21786
rect 6316 21734 6330 21786
rect 6330 21734 6342 21786
rect 6342 21734 6372 21786
rect 6396 21734 6406 21786
rect 6406 21734 6452 21786
rect 6156 21732 6212 21734
rect 6236 21732 6292 21734
rect 6316 21732 6372 21734
rect 6396 21732 6452 21734
rect 5906 3576 5962 3632
rect 6156 20698 6212 20700
rect 6236 20698 6292 20700
rect 6316 20698 6372 20700
rect 6396 20698 6452 20700
rect 6156 20646 6202 20698
rect 6202 20646 6212 20698
rect 6236 20646 6266 20698
rect 6266 20646 6278 20698
rect 6278 20646 6292 20698
rect 6316 20646 6330 20698
rect 6330 20646 6342 20698
rect 6342 20646 6372 20698
rect 6396 20646 6406 20698
rect 6406 20646 6452 20698
rect 6156 20644 6212 20646
rect 6236 20644 6292 20646
rect 6316 20644 6372 20646
rect 6396 20644 6452 20646
rect 6156 19610 6212 19612
rect 6236 19610 6292 19612
rect 6316 19610 6372 19612
rect 6396 19610 6452 19612
rect 6156 19558 6202 19610
rect 6202 19558 6212 19610
rect 6236 19558 6266 19610
rect 6266 19558 6278 19610
rect 6278 19558 6292 19610
rect 6316 19558 6330 19610
rect 6330 19558 6342 19610
rect 6342 19558 6372 19610
rect 6396 19558 6406 19610
rect 6406 19558 6452 19610
rect 6156 19556 6212 19558
rect 6236 19556 6292 19558
rect 6316 19556 6372 19558
rect 6396 19556 6452 19558
rect 6156 18522 6212 18524
rect 6236 18522 6292 18524
rect 6316 18522 6372 18524
rect 6396 18522 6452 18524
rect 6156 18470 6202 18522
rect 6202 18470 6212 18522
rect 6236 18470 6266 18522
rect 6266 18470 6278 18522
rect 6278 18470 6292 18522
rect 6316 18470 6330 18522
rect 6330 18470 6342 18522
rect 6342 18470 6372 18522
rect 6396 18470 6406 18522
rect 6406 18470 6452 18522
rect 6156 18468 6212 18470
rect 6236 18468 6292 18470
rect 6316 18468 6372 18470
rect 6396 18468 6452 18470
rect 6156 17434 6212 17436
rect 6236 17434 6292 17436
rect 6316 17434 6372 17436
rect 6396 17434 6452 17436
rect 6156 17382 6202 17434
rect 6202 17382 6212 17434
rect 6236 17382 6266 17434
rect 6266 17382 6278 17434
rect 6278 17382 6292 17434
rect 6316 17382 6330 17434
rect 6330 17382 6342 17434
rect 6342 17382 6372 17434
rect 6396 17382 6406 17434
rect 6406 17382 6452 17434
rect 6156 17380 6212 17382
rect 6236 17380 6292 17382
rect 6316 17380 6372 17382
rect 6396 17380 6452 17382
rect 6156 16346 6212 16348
rect 6236 16346 6292 16348
rect 6316 16346 6372 16348
rect 6396 16346 6452 16348
rect 6156 16294 6202 16346
rect 6202 16294 6212 16346
rect 6236 16294 6266 16346
rect 6266 16294 6278 16346
rect 6278 16294 6292 16346
rect 6316 16294 6330 16346
rect 6330 16294 6342 16346
rect 6342 16294 6372 16346
rect 6396 16294 6406 16346
rect 6406 16294 6452 16346
rect 6156 16292 6212 16294
rect 6236 16292 6292 16294
rect 6316 16292 6372 16294
rect 6396 16292 6452 16294
rect 6156 15258 6212 15260
rect 6236 15258 6292 15260
rect 6316 15258 6372 15260
rect 6396 15258 6452 15260
rect 6156 15206 6202 15258
rect 6202 15206 6212 15258
rect 6236 15206 6266 15258
rect 6266 15206 6278 15258
rect 6278 15206 6292 15258
rect 6316 15206 6330 15258
rect 6330 15206 6342 15258
rect 6342 15206 6372 15258
rect 6396 15206 6406 15258
rect 6406 15206 6452 15258
rect 6156 15204 6212 15206
rect 6236 15204 6292 15206
rect 6316 15204 6372 15206
rect 6396 15204 6452 15206
rect 6156 14170 6212 14172
rect 6236 14170 6292 14172
rect 6316 14170 6372 14172
rect 6396 14170 6452 14172
rect 6156 14118 6202 14170
rect 6202 14118 6212 14170
rect 6236 14118 6266 14170
rect 6266 14118 6278 14170
rect 6278 14118 6292 14170
rect 6316 14118 6330 14170
rect 6330 14118 6342 14170
rect 6342 14118 6372 14170
rect 6396 14118 6406 14170
rect 6406 14118 6452 14170
rect 6156 14116 6212 14118
rect 6236 14116 6292 14118
rect 6316 14116 6372 14118
rect 6396 14116 6452 14118
rect 6156 13082 6212 13084
rect 6236 13082 6292 13084
rect 6316 13082 6372 13084
rect 6396 13082 6452 13084
rect 6156 13030 6202 13082
rect 6202 13030 6212 13082
rect 6236 13030 6266 13082
rect 6266 13030 6278 13082
rect 6278 13030 6292 13082
rect 6316 13030 6330 13082
rect 6330 13030 6342 13082
rect 6342 13030 6372 13082
rect 6396 13030 6406 13082
rect 6406 13030 6452 13082
rect 6156 13028 6212 13030
rect 6236 13028 6292 13030
rect 6316 13028 6372 13030
rect 6396 13028 6452 13030
rect 6156 11994 6212 11996
rect 6236 11994 6292 11996
rect 6316 11994 6372 11996
rect 6396 11994 6452 11996
rect 6156 11942 6202 11994
rect 6202 11942 6212 11994
rect 6236 11942 6266 11994
rect 6266 11942 6278 11994
rect 6278 11942 6292 11994
rect 6316 11942 6330 11994
rect 6330 11942 6342 11994
rect 6342 11942 6372 11994
rect 6396 11942 6406 11994
rect 6406 11942 6452 11994
rect 6156 11940 6212 11942
rect 6236 11940 6292 11942
rect 6316 11940 6372 11942
rect 6396 11940 6452 11942
rect 6156 10906 6212 10908
rect 6236 10906 6292 10908
rect 6316 10906 6372 10908
rect 6396 10906 6452 10908
rect 6156 10854 6202 10906
rect 6202 10854 6212 10906
rect 6236 10854 6266 10906
rect 6266 10854 6278 10906
rect 6278 10854 6292 10906
rect 6316 10854 6330 10906
rect 6330 10854 6342 10906
rect 6342 10854 6372 10906
rect 6396 10854 6406 10906
rect 6406 10854 6452 10906
rect 6156 10852 6212 10854
rect 6236 10852 6292 10854
rect 6316 10852 6372 10854
rect 6396 10852 6452 10854
rect 6156 9818 6212 9820
rect 6236 9818 6292 9820
rect 6316 9818 6372 9820
rect 6396 9818 6452 9820
rect 6156 9766 6202 9818
rect 6202 9766 6212 9818
rect 6236 9766 6266 9818
rect 6266 9766 6278 9818
rect 6278 9766 6292 9818
rect 6316 9766 6330 9818
rect 6330 9766 6342 9818
rect 6342 9766 6372 9818
rect 6396 9766 6406 9818
rect 6406 9766 6452 9818
rect 6156 9764 6212 9766
rect 6236 9764 6292 9766
rect 6316 9764 6372 9766
rect 6396 9764 6452 9766
rect 6156 8730 6212 8732
rect 6236 8730 6292 8732
rect 6316 8730 6372 8732
rect 6396 8730 6452 8732
rect 6156 8678 6202 8730
rect 6202 8678 6212 8730
rect 6236 8678 6266 8730
rect 6266 8678 6278 8730
rect 6278 8678 6292 8730
rect 6316 8678 6330 8730
rect 6330 8678 6342 8730
rect 6342 8678 6372 8730
rect 6396 8678 6406 8730
rect 6406 8678 6452 8730
rect 6156 8676 6212 8678
rect 6236 8676 6292 8678
rect 6316 8676 6372 8678
rect 6396 8676 6452 8678
rect 6156 7642 6212 7644
rect 6236 7642 6292 7644
rect 6316 7642 6372 7644
rect 6396 7642 6452 7644
rect 6156 7590 6202 7642
rect 6202 7590 6212 7642
rect 6236 7590 6266 7642
rect 6266 7590 6278 7642
rect 6278 7590 6292 7642
rect 6316 7590 6330 7642
rect 6330 7590 6342 7642
rect 6342 7590 6372 7642
rect 6396 7590 6406 7642
rect 6406 7590 6452 7642
rect 6156 7588 6212 7590
rect 6236 7588 6292 7590
rect 6316 7588 6372 7590
rect 6396 7588 6452 7590
rect 6156 6554 6212 6556
rect 6236 6554 6292 6556
rect 6316 6554 6372 6556
rect 6396 6554 6452 6556
rect 6156 6502 6202 6554
rect 6202 6502 6212 6554
rect 6236 6502 6266 6554
rect 6266 6502 6278 6554
rect 6278 6502 6292 6554
rect 6316 6502 6330 6554
rect 6330 6502 6342 6554
rect 6342 6502 6372 6554
rect 6396 6502 6406 6554
rect 6406 6502 6452 6554
rect 6156 6500 6212 6502
rect 6236 6500 6292 6502
rect 6316 6500 6372 6502
rect 6396 6500 6452 6502
rect 6156 5466 6212 5468
rect 6236 5466 6292 5468
rect 6316 5466 6372 5468
rect 6396 5466 6452 5468
rect 6156 5414 6202 5466
rect 6202 5414 6212 5466
rect 6236 5414 6266 5466
rect 6266 5414 6278 5466
rect 6278 5414 6292 5466
rect 6316 5414 6330 5466
rect 6330 5414 6342 5466
rect 6342 5414 6372 5466
rect 6396 5414 6406 5466
rect 6406 5414 6452 5466
rect 6156 5412 6212 5414
rect 6236 5412 6292 5414
rect 6316 5412 6372 5414
rect 6396 5412 6452 5414
rect 6156 4378 6212 4380
rect 6236 4378 6292 4380
rect 6316 4378 6372 4380
rect 6396 4378 6452 4380
rect 6156 4326 6202 4378
rect 6202 4326 6212 4378
rect 6236 4326 6266 4378
rect 6266 4326 6278 4378
rect 6278 4326 6292 4378
rect 6316 4326 6330 4378
rect 6330 4326 6342 4378
rect 6342 4326 6372 4378
rect 6396 4326 6406 4378
rect 6406 4326 6452 4378
rect 6156 4324 6212 4326
rect 6236 4324 6292 4326
rect 6316 4324 6372 4326
rect 6396 4324 6452 4326
rect 6156 3290 6212 3292
rect 6236 3290 6292 3292
rect 6316 3290 6372 3292
rect 6396 3290 6452 3292
rect 6156 3238 6202 3290
rect 6202 3238 6212 3290
rect 6236 3238 6266 3290
rect 6266 3238 6278 3290
rect 6278 3238 6292 3290
rect 6316 3238 6330 3290
rect 6330 3238 6342 3290
rect 6342 3238 6372 3290
rect 6396 3238 6406 3290
rect 6406 3238 6452 3290
rect 6156 3236 6212 3238
rect 6236 3236 6292 3238
rect 6316 3236 6372 3238
rect 6396 3236 6452 3238
rect 6156 2202 6212 2204
rect 6236 2202 6292 2204
rect 6316 2202 6372 2204
rect 6396 2202 6452 2204
rect 6156 2150 6202 2202
rect 6202 2150 6212 2202
rect 6236 2150 6266 2202
rect 6266 2150 6278 2202
rect 6278 2150 6292 2202
rect 6316 2150 6330 2202
rect 6330 2150 6342 2202
rect 6342 2150 6372 2202
rect 6396 2150 6406 2202
rect 6406 2150 6452 2202
rect 6156 2148 6212 2150
rect 6236 2148 6292 2150
rect 6316 2148 6372 2150
rect 6396 2148 6452 2150
rect 7194 27512 7250 27568
rect 6816 26682 6872 26684
rect 6896 26682 6952 26684
rect 6976 26682 7032 26684
rect 7056 26682 7112 26684
rect 6816 26630 6862 26682
rect 6862 26630 6872 26682
rect 6896 26630 6926 26682
rect 6926 26630 6938 26682
rect 6938 26630 6952 26682
rect 6976 26630 6990 26682
rect 6990 26630 7002 26682
rect 7002 26630 7032 26682
rect 7056 26630 7066 26682
rect 7066 26630 7112 26682
rect 6816 26628 6872 26630
rect 6896 26628 6952 26630
rect 6976 26628 7032 26630
rect 7056 26628 7112 26630
rect 6816 25594 6872 25596
rect 6896 25594 6952 25596
rect 6976 25594 7032 25596
rect 7056 25594 7112 25596
rect 6816 25542 6862 25594
rect 6862 25542 6872 25594
rect 6896 25542 6926 25594
rect 6926 25542 6938 25594
rect 6938 25542 6952 25594
rect 6976 25542 6990 25594
rect 6990 25542 7002 25594
rect 7002 25542 7032 25594
rect 7056 25542 7066 25594
rect 7066 25542 7112 25594
rect 6816 25540 6872 25542
rect 6896 25540 6952 25542
rect 6976 25540 7032 25542
rect 7056 25540 7112 25542
rect 7470 28328 7526 28384
rect 6816 24506 6872 24508
rect 6896 24506 6952 24508
rect 6976 24506 7032 24508
rect 7056 24506 7112 24508
rect 6816 24454 6862 24506
rect 6862 24454 6872 24506
rect 6896 24454 6926 24506
rect 6926 24454 6938 24506
rect 6938 24454 6952 24506
rect 6976 24454 6990 24506
rect 6990 24454 7002 24506
rect 7002 24454 7032 24506
rect 7056 24454 7066 24506
rect 7066 24454 7112 24506
rect 6816 24452 6872 24454
rect 6896 24452 6952 24454
rect 6976 24452 7032 24454
rect 7056 24452 7112 24454
rect 6816 23418 6872 23420
rect 6896 23418 6952 23420
rect 6976 23418 7032 23420
rect 7056 23418 7112 23420
rect 6816 23366 6862 23418
rect 6862 23366 6872 23418
rect 6896 23366 6926 23418
rect 6926 23366 6938 23418
rect 6938 23366 6952 23418
rect 6976 23366 6990 23418
rect 6990 23366 7002 23418
rect 7002 23366 7032 23418
rect 7056 23366 7066 23418
rect 7066 23366 7112 23418
rect 6816 23364 6872 23366
rect 6896 23364 6952 23366
rect 6976 23364 7032 23366
rect 7056 23364 7112 23366
rect 9356 46810 9412 46812
rect 9436 46810 9492 46812
rect 9516 46810 9572 46812
rect 9596 46810 9652 46812
rect 9356 46758 9402 46810
rect 9402 46758 9412 46810
rect 9436 46758 9466 46810
rect 9466 46758 9478 46810
rect 9478 46758 9492 46810
rect 9516 46758 9530 46810
rect 9530 46758 9542 46810
rect 9542 46758 9572 46810
rect 9596 46758 9606 46810
rect 9606 46758 9652 46810
rect 9356 46756 9412 46758
rect 9436 46756 9492 46758
rect 9516 46756 9572 46758
rect 9596 46756 9652 46758
rect 9310 46552 9366 46608
rect 9356 45722 9412 45724
rect 9436 45722 9492 45724
rect 9516 45722 9572 45724
rect 9596 45722 9652 45724
rect 9356 45670 9402 45722
rect 9402 45670 9412 45722
rect 9436 45670 9466 45722
rect 9466 45670 9478 45722
rect 9478 45670 9492 45722
rect 9516 45670 9530 45722
rect 9530 45670 9542 45722
rect 9542 45670 9572 45722
rect 9596 45670 9606 45722
rect 9606 45670 9652 45722
rect 9356 45668 9412 45670
rect 9436 45668 9492 45670
rect 9516 45668 9572 45670
rect 9596 45668 9652 45670
rect 9356 44634 9412 44636
rect 9436 44634 9492 44636
rect 9516 44634 9572 44636
rect 9596 44634 9652 44636
rect 9356 44582 9402 44634
rect 9402 44582 9412 44634
rect 9436 44582 9466 44634
rect 9466 44582 9478 44634
rect 9478 44582 9492 44634
rect 9516 44582 9530 44634
rect 9530 44582 9542 44634
rect 9542 44582 9572 44634
rect 9596 44582 9606 44634
rect 9606 44582 9652 44634
rect 9356 44580 9412 44582
rect 9436 44580 9492 44582
rect 9516 44580 9572 44582
rect 9596 44580 9652 44582
rect 9356 43546 9412 43548
rect 9436 43546 9492 43548
rect 9516 43546 9572 43548
rect 9596 43546 9652 43548
rect 9356 43494 9402 43546
rect 9402 43494 9412 43546
rect 9436 43494 9466 43546
rect 9466 43494 9478 43546
rect 9478 43494 9492 43546
rect 9516 43494 9530 43546
rect 9530 43494 9542 43546
rect 9542 43494 9572 43546
rect 9596 43494 9606 43546
rect 9606 43494 9652 43546
rect 9356 43492 9412 43494
rect 9436 43492 9492 43494
rect 9516 43492 9572 43494
rect 9596 43492 9652 43494
rect 9356 42458 9412 42460
rect 9436 42458 9492 42460
rect 9516 42458 9572 42460
rect 9596 42458 9652 42460
rect 9356 42406 9402 42458
rect 9402 42406 9412 42458
rect 9436 42406 9466 42458
rect 9466 42406 9478 42458
rect 9478 42406 9492 42458
rect 9516 42406 9530 42458
rect 9530 42406 9542 42458
rect 9542 42406 9572 42458
rect 9596 42406 9606 42458
rect 9606 42406 9652 42458
rect 9356 42404 9412 42406
rect 9436 42404 9492 42406
rect 9516 42404 9572 42406
rect 9596 42404 9652 42406
rect 9356 41370 9412 41372
rect 9436 41370 9492 41372
rect 9516 41370 9572 41372
rect 9596 41370 9652 41372
rect 9356 41318 9402 41370
rect 9402 41318 9412 41370
rect 9436 41318 9466 41370
rect 9466 41318 9478 41370
rect 9478 41318 9492 41370
rect 9516 41318 9530 41370
rect 9530 41318 9542 41370
rect 9542 41318 9572 41370
rect 9596 41318 9606 41370
rect 9606 41318 9652 41370
rect 9356 41316 9412 41318
rect 9436 41316 9492 41318
rect 9516 41316 9572 41318
rect 9596 41316 9652 41318
rect 9356 40282 9412 40284
rect 9436 40282 9492 40284
rect 9516 40282 9572 40284
rect 9596 40282 9652 40284
rect 9356 40230 9402 40282
rect 9402 40230 9412 40282
rect 9436 40230 9466 40282
rect 9466 40230 9478 40282
rect 9478 40230 9492 40282
rect 9516 40230 9530 40282
rect 9530 40230 9542 40282
rect 9542 40230 9572 40282
rect 9596 40230 9606 40282
rect 9606 40230 9652 40282
rect 9356 40228 9412 40230
rect 9436 40228 9492 40230
rect 9516 40228 9572 40230
rect 9596 40228 9652 40230
rect 9356 39194 9412 39196
rect 9436 39194 9492 39196
rect 9516 39194 9572 39196
rect 9596 39194 9652 39196
rect 9356 39142 9402 39194
rect 9402 39142 9412 39194
rect 9436 39142 9466 39194
rect 9466 39142 9478 39194
rect 9478 39142 9492 39194
rect 9516 39142 9530 39194
rect 9530 39142 9542 39194
rect 9542 39142 9572 39194
rect 9596 39142 9606 39194
rect 9606 39142 9652 39194
rect 9356 39140 9412 39142
rect 9436 39140 9492 39142
rect 9516 39140 9572 39142
rect 9596 39140 9652 39142
rect 8850 36352 8906 36408
rect 9356 38106 9412 38108
rect 9436 38106 9492 38108
rect 9516 38106 9572 38108
rect 9596 38106 9652 38108
rect 9356 38054 9402 38106
rect 9402 38054 9412 38106
rect 9436 38054 9466 38106
rect 9466 38054 9478 38106
rect 9478 38054 9492 38106
rect 9516 38054 9530 38106
rect 9530 38054 9542 38106
rect 9542 38054 9572 38106
rect 9596 38054 9606 38106
rect 9606 38054 9652 38106
rect 9356 38052 9412 38054
rect 9436 38052 9492 38054
rect 9516 38052 9572 38054
rect 9596 38052 9652 38054
rect 9770 37304 9826 37360
rect 9356 37018 9412 37020
rect 9436 37018 9492 37020
rect 9516 37018 9572 37020
rect 9596 37018 9652 37020
rect 9356 36966 9402 37018
rect 9402 36966 9412 37018
rect 9436 36966 9466 37018
rect 9466 36966 9478 37018
rect 9478 36966 9492 37018
rect 9516 36966 9530 37018
rect 9530 36966 9542 37018
rect 9542 36966 9572 37018
rect 9596 36966 9606 37018
rect 9606 36966 9652 37018
rect 9356 36964 9412 36966
rect 9436 36964 9492 36966
rect 9516 36964 9572 36966
rect 9596 36964 9652 36966
rect 7756 31578 7812 31580
rect 7836 31578 7892 31580
rect 7916 31578 7972 31580
rect 7996 31578 8052 31580
rect 7756 31526 7802 31578
rect 7802 31526 7812 31578
rect 7836 31526 7866 31578
rect 7866 31526 7878 31578
rect 7878 31526 7892 31578
rect 7916 31526 7930 31578
rect 7930 31526 7942 31578
rect 7942 31526 7972 31578
rect 7996 31526 8006 31578
rect 8006 31526 8052 31578
rect 7756 31524 7812 31526
rect 7836 31524 7892 31526
rect 7916 31524 7972 31526
rect 7996 31524 8052 31526
rect 7756 30490 7812 30492
rect 7836 30490 7892 30492
rect 7916 30490 7972 30492
rect 7996 30490 8052 30492
rect 7756 30438 7802 30490
rect 7802 30438 7812 30490
rect 7836 30438 7866 30490
rect 7866 30438 7878 30490
rect 7878 30438 7892 30490
rect 7916 30438 7930 30490
rect 7930 30438 7942 30490
rect 7942 30438 7972 30490
rect 7996 30438 8006 30490
rect 8006 30438 8052 30490
rect 7756 30436 7812 30438
rect 7836 30436 7892 30438
rect 7916 30436 7972 30438
rect 7996 30436 8052 30438
rect 7756 29402 7812 29404
rect 7836 29402 7892 29404
rect 7916 29402 7972 29404
rect 7996 29402 8052 29404
rect 7756 29350 7802 29402
rect 7802 29350 7812 29402
rect 7836 29350 7866 29402
rect 7866 29350 7878 29402
rect 7878 29350 7892 29402
rect 7916 29350 7930 29402
rect 7930 29350 7942 29402
rect 7942 29350 7972 29402
rect 7996 29350 8006 29402
rect 8006 29350 8052 29402
rect 7756 29348 7812 29350
rect 7836 29348 7892 29350
rect 7916 29348 7972 29350
rect 7996 29348 8052 29350
rect 7930 28464 7986 28520
rect 8416 33210 8472 33212
rect 8496 33210 8552 33212
rect 8576 33210 8632 33212
rect 8656 33210 8712 33212
rect 8416 33158 8462 33210
rect 8462 33158 8472 33210
rect 8496 33158 8526 33210
rect 8526 33158 8538 33210
rect 8538 33158 8552 33210
rect 8576 33158 8590 33210
rect 8590 33158 8602 33210
rect 8602 33158 8632 33210
rect 8656 33158 8666 33210
rect 8666 33158 8712 33210
rect 8416 33156 8472 33158
rect 8496 33156 8552 33158
rect 8576 33156 8632 33158
rect 8656 33156 8712 33158
rect 8416 32122 8472 32124
rect 8496 32122 8552 32124
rect 8576 32122 8632 32124
rect 8656 32122 8712 32124
rect 8416 32070 8462 32122
rect 8462 32070 8472 32122
rect 8496 32070 8526 32122
rect 8526 32070 8538 32122
rect 8538 32070 8552 32122
rect 8576 32070 8590 32122
rect 8590 32070 8602 32122
rect 8602 32070 8632 32122
rect 8656 32070 8666 32122
rect 8666 32070 8712 32122
rect 8416 32068 8472 32070
rect 8496 32068 8552 32070
rect 8576 32068 8632 32070
rect 8656 32068 8712 32070
rect 8416 31034 8472 31036
rect 8496 31034 8552 31036
rect 8576 31034 8632 31036
rect 8656 31034 8712 31036
rect 8416 30982 8462 31034
rect 8462 30982 8472 31034
rect 8496 30982 8526 31034
rect 8526 30982 8538 31034
rect 8538 30982 8552 31034
rect 8576 30982 8590 31034
rect 8590 30982 8602 31034
rect 8602 30982 8632 31034
rect 8656 30982 8666 31034
rect 8666 30982 8712 31034
rect 8416 30980 8472 30982
rect 8496 30980 8552 30982
rect 8576 30980 8632 30982
rect 8656 30980 8712 30982
rect 8416 29946 8472 29948
rect 8496 29946 8552 29948
rect 8576 29946 8632 29948
rect 8656 29946 8712 29948
rect 8416 29894 8462 29946
rect 8462 29894 8472 29946
rect 8496 29894 8526 29946
rect 8526 29894 8538 29946
rect 8538 29894 8552 29946
rect 8576 29894 8590 29946
rect 8590 29894 8602 29946
rect 8602 29894 8632 29946
rect 8656 29894 8666 29946
rect 8666 29894 8712 29946
rect 8416 29892 8472 29894
rect 8496 29892 8552 29894
rect 8576 29892 8632 29894
rect 8656 29892 8712 29894
rect 8942 31728 8998 31784
rect 7756 28314 7812 28316
rect 7836 28314 7892 28316
rect 7916 28314 7972 28316
rect 7996 28314 8052 28316
rect 7756 28262 7802 28314
rect 7802 28262 7812 28314
rect 7836 28262 7866 28314
rect 7866 28262 7878 28314
rect 7878 28262 7892 28314
rect 7916 28262 7930 28314
rect 7930 28262 7942 28314
rect 7942 28262 7972 28314
rect 7996 28262 8006 28314
rect 8006 28262 8052 28314
rect 7756 28260 7812 28262
rect 7836 28260 7892 28262
rect 7916 28260 7972 28262
rect 7996 28260 8052 28262
rect 7756 27226 7812 27228
rect 7836 27226 7892 27228
rect 7916 27226 7972 27228
rect 7996 27226 8052 27228
rect 7756 27174 7802 27226
rect 7802 27174 7812 27226
rect 7836 27174 7866 27226
rect 7866 27174 7878 27226
rect 7878 27174 7892 27226
rect 7916 27174 7930 27226
rect 7930 27174 7942 27226
rect 7942 27174 7972 27226
rect 7996 27174 8006 27226
rect 8006 27174 8052 27226
rect 7756 27172 7812 27174
rect 7836 27172 7892 27174
rect 7916 27172 7972 27174
rect 7996 27172 8052 27174
rect 7756 26138 7812 26140
rect 7836 26138 7892 26140
rect 7916 26138 7972 26140
rect 7996 26138 8052 26140
rect 7756 26086 7802 26138
rect 7802 26086 7812 26138
rect 7836 26086 7866 26138
rect 7866 26086 7878 26138
rect 7878 26086 7892 26138
rect 7916 26086 7930 26138
rect 7930 26086 7942 26138
rect 7942 26086 7972 26138
rect 7996 26086 8006 26138
rect 8006 26086 8052 26138
rect 7756 26084 7812 26086
rect 7836 26084 7892 26086
rect 7916 26084 7972 26086
rect 7996 26084 8052 26086
rect 6816 22330 6872 22332
rect 6896 22330 6952 22332
rect 6976 22330 7032 22332
rect 7056 22330 7112 22332
rect 6816 22278 6862 22330
rect 6862 22278 6872 22330
rect 6896 22278 6926 22330
rect 6926 22278 6938 22330
rect 6938 22278 6952 22330
rect 6976 22278 6990 22330
rect 6990 22278 7002 22330
rect 7002 22278 7032 22330
rect 7056 22278 7066 22330
rect 7066 22278 7112 22330
rect 6816 22276 6872 22278
rect 6896 22276 6952 22278
rect 6976 22276 7032 22278
rect 7056 22276 7112 22278
rect 7654 25780 7656 25800
rect 7656 25780 7708 25800
rect 7708 25780 7710 25800
rect 7654 25744 7710 25780
rect 7756 25050 7812 25052
rect 7836 25050 7892 25052
rect 7916 25050 7972 25052
rect 7996 25050 8052 25052
rect 7756 24998 7802 25050
rect 7802 24998 7812 25050
rect 7836 24998 7866 25050
rect 7866 24998 7878 25050
rect 7878 24998 7892 25050
rect 7916 24998 7930 25050
rect 7930 24998 7942 25050
rect 7942 24998 7972 25050
rect 7996 24998 8006 25050
rect 8006 24998 8052 25050
rect 7756 24996 7812 24998
rect 7836 24996 7892 24998
rect 7916 24996 7972 24998
rect 7996 24996 8052 24998
rect 7756 23962 7812 23964
rect 7836 23962 7892 23964
rect 7916 23962 7972 23964
rect 7996 23962 8052 23964
rect 7756 23910 7802 23962
rect 7802 23910 7812 23962
rect 7836 23910 7866 23962
rect 7866 23910 7878 23962
rect 7878 23910 7892 23962
rect 7916 23910 7930 23962
rect 7930 23910 7942 23962
rect 7942 23910 7972 23962
rect 7996 23910 8006 23962
rect 8006 23910 8052 23962
rect 7756 23908 7812 23910
rect 7836 23908 7892 23910
rect 7916 23908 7972 23910
rect 7996 23908 8052 23910
rect 7756 22874 7812 22876
rect 7836 22874 7892 22876
rect 7916 22874 7972 22876
rect 7996 22874 8052 22876
rect 7756 22822 7802 22874
rect 7802 22822 7812 22874
rect 7836 22822 7866 22874
rect 7866 22822 7878 22874
rect 7878 22822 7892 22874
rect 7916 22822 7930 22874
rect 7930 22822 7942 22874
rect 7942 22822 7972 22874
rect 7996 22822 8006 22874
rect 8006 22822 8052 22874
rect 7756 22820 7812 22822
rect 7836 22820 7892 22822
rect 7916 22820 7972 22822
rect 7996 22820 8052 22822
rect 6816 21242 6872 21244
rect 6896 21242 6952 21244
rect 6976 21242 7032 21244
rect 7056 21242 7112 21244
rect 6816 21190 6862 21242
rect 6862 21190 6872 21242
rect 6896 21190 6926 21242
rect 6926 21190 6938 21242
rect 6938 21190 6952 21242
rect 6976 21190 6990 21242
rect 6990 21190 7002 21242
rect 7002 21190 7032 21242
rect 7056 21190 7066 21242
rect 7066 21190 7112 21242
rect 6816 21188 6872 21190
rect 6896 21188 6952 21190
rect 6976 21188 7032 21190
rect 7056 21188 7112 21190
rect 6816 20154 6872 20156
rect 6896 20154 6952 20156
rect 6976 20154 7032 20156
rect 7056 20154 7112 20156
rect 6816 20102 6862 20154
rect 6862 20102 6872 20154
rect 6896 20102 6926 20154
rect 6926 20102 6938 20154
rect 6938 20102 6952 20154
rect 6976 20102 6990 20154
rect 6990 20102 7002 20154
rect 7002 20102 7032 20154
rect 7056 20102 7066 20154
rect 7066 20102 7112 20154
rect 6816 20100 6872 20102
rect 6896 20100 6952 20102
rect 6976 20100 7032 20102
rect 7056 20100 7112 20102
rect 6816 19066 6872 19068
rect 6896 19066 6952 19068
rect 6976 19066 7032 19068
rect 7056 19066 7112 19068
rect 6816 19014 6862 19066
rect 6862 19014 6872 19066
rect 6896 19014 6926 19066
rect 6926 19014 6938 19066
rect 6938 19014 6952 19066
rect 6976 19014 6990 19066
rect 6990 19014 7002 19066
rect 7002 19014 7032 19066
rect 7056 19014 7066 19066
rect 7066 19014 7112 19066
rect 6816 19012 6872 19014
rect 6896 19012 6952 19014
rect 6976 19012 7032 19014
rect 7056 19012 7112 19014
rect 6816 17978 6872 17980
rect 6896 17978 6952 17980
rect 6976 17978 7032 17980
rect 7056 17978 7112 17980
rect 6816 17926 6862 17978
rect 6862 17926 6872 17978
rect 6896 17926 6926 17978
rect 6926 17926 6938 17978
rect 6938 17926 6952 17978
rect 6976 17926 6990 17978
rect 6990 17926 7002 17978
rect 7002 17926 7032 17978
rect 7056 17926 7066 17978
rect 7066 17926 7112 17978
rect 6816 17924 6872 17926
rect 6896 17924 6952 17926
rect 6976 17924 7032 17926
rect 7056 17924 7112 17926
rect 6816 16890 6872 16892
rect 6896 16890 6952 16892
rect 6976 16890 7032 16892
rect 7056 16890 7112 16892
rect 6816 16838 6862 16890
rect 6862 16838 6872 16890
rect 6896 16838 6926 16890
rect 6926 16838 6938 16890
rect 6938 16838 6952 16890
rect 6976 16838 6990 16890
rect 6990 16838 7002 16890
rect 7002 16838 7032 16890
rect 7056 16838 7066 16890
rect 7066 16838 7112 16890
rect 6816 16836 6872 16838
rect 6896 16836 6952 16838
rect 6976 16836 7032 16838
rect 7056 16836 7112 16838
rect 6816 15802 6872 15804
rect 6896 15802 6952 15804
rect 6976 15802 7032 15804
rect 7056 15802 7112 15804
rect 6816 15750 6862 15802
rect 6862 15750 6872 15802
rect 6896 15750 6926 15802
rect 6926 15750 6938 15802
rect 6938 15750 6952 15802
rect 6976 15750 6990 15802
rect 6990 15750 7002 15802
rect 7002 15750 7032 15802
rect 7056 15750 7066 15802
rect 7066 15750 7112 15802
rect 6816 15748 6872 15750
rect 6896 15748 6952 15750
rect 6976 15748 7032 15750
rect 7056 15748 7112 15750
rect 6816 14714 6872 14716
rect 6896 14714 6952 14716
rect 6976 14714 7032 14716
rect 7056 14714 7112 14716
rect 6816 14662 6862 14714
rect 6862 14662 6872 14714
rect 6896 14662 6926 14714
rect 6926 14662 6938 14714
rect 6938 14662 6952 14714
rect 6976 14662 6990 14714
rect 6990 14662 7002 14714
rect 7002 14662 7032 14714
rect 7056 14662 7066 14714
rect 7066 14662 7112 14714
rect 6816 14660 6872 14662
rect 6896 14660 6952 14662
rect 6976 14660 7032 14662
rect 7056 14660 7112 14662
rect 7756 21786 7812 21788
rect 7836 21786 7892 21788
rect 7916 21786 7972 21788
rect 7996 21786 8052 21788
rect 7756 21734 7802 21786
rect 7802 21734 7812 21786
rect 7836 21734 7866 21786
rect 7866 21734 7878 21786
rect 7878 21734 7892 21786
rect 7916 21734 7930 21786
rect 7930 21734 7942 21786
rect 7942 21734 7972 21786
rect 7996 21734 8006 21786
rect 8006 21734 8052 21786
rect 7756 21732 7812 21734
rect 7836 21732 7892 21734
rect 7916 21732 7972 21734
rect 7996 21732 8052 21734
rect 7756 20698 7812 20700
rect 7836 20698 7892 20700
rect 7916 20698 7972 20700
rect 7996 20698 8052 20700
rect 7756 20646 7802 20698
rect 7802 20646 7812 20698
rect 7836 20646 7866 20698
rect 7866 20646 7878 20698
rect 7878 20646 7892 20698
rect 7916 20646 7930 20698
rect 7930 20646 7942 20698
rect 7942 20646 7972 20698
rect 7996 20646 8006 20698
rect 8006 20646 8052 20698
rect 7756 20644 7812 20646
rect 7836 20644 7892 20646
rect 7916 20644 7972 20646
rect 7996 20644 8052 20646
rect 7756 19610 7812 19612
rect 7836 19610 7892 19612
rect 7916 19610 7972 19612
rect 7996 19610 8052 19612
rect 7756 19558 7802 19610
rect 7802 19558 7812 19610
rect 7836 19558 7866 19610
rect 7866 19558 7878 19610
rect 7878 19558 7892 19610
rect 7916 19558 7930 19610
rect 7930 19558 7942 19610
rect 7942 19558 7972 19610
rect 7996 19558 8006 19610
rect 8006 19558 8052 19610
rect 7756 19556 7812 19558
rect 7836 19556 7892 19558
rect 7916 19556 7972 19558
rect 7996 19556 8052 19558
rect 6816 13626 6872 13628
rect 6896 13626 6952 13628
rect 6976 13626 7032 13628
rect 7056 13626 7112 13628
rect 6816 13574 6862 13626
rect 6862 13574 6872 13626
rect 6896 13574 6926 13626
rect 6926 13574 6938 13626
rect 6938 13574 6952 13626
rect 6976 13574 6990 13626
rect 6990 13574 7002 13626
rect 7002 13574 7032 13626
rect 7056 13574 7066 13626
rect 7066 13574 7112 13626
rect 6816 13572 6872 13574
rect 6896 13572 6952 13574
rect 6976 13572 7032 13574
rect 7056 13572 7112 13574
rect 6816 12538 6872 12540
rect 6896 12538 6952 12540
rect 6976 12538 7032 12540
rect 7056 12538 7112 12540
rect 6816 12486 6862 12538
rect 6862 12486 6872 12538
rect 6896 12486 6926 12538
rect 6926 12486 6938 12538
rect 6938 12486 6952 12538
rect 6976 12486 6990 12538
rect 6990 12486 7002 12538
rect 7002 12486 7032 12538
rect 7056 12486 7066 12538
rect 7066 12486 7112 12538
rect 6816 12484 6872 12486
rect 6896 12484 6952 12486
rect 6976 12484 7032 12486
rect 7056 12484 7112 12486
rect 6816 11450 6872 11452
rect 6896 11450 6952 11452
rect 6976 11450 7032 11452
rect 7056 11450 7112 11452
rect 6816 11398 6862 11450
rect 6862 11398 6872 11450
rect 6896 11398 6926 11450
rect 6926 11398 6938 11450
rect 6938 11398 6952 11450
rect 6976 11398 6990 11450
rect 6990 11398 7002 11450
rect 7002 11398 7032 11450
rect 7056 11398 7066 11450
rect 7066 11398 7112 11450
rect 6816 11396 6872 11398
rect 6896 11396 6952 11398
rect 6976 11396 7032 11398
rect 7056 11396 7112 11398
rect 6816 10362 6872 10364
rect 6896 10362 6952 10364
rect 6976 10362 7032 10364
rect 7056 10362 7112 10364
rect 6816 10310 6862 10362
rect 6862 10310 6872 10362
rect 6896 10310 6926 10362
rect 6926 10310 6938 10362
rect 6938 10310 6952 10362
rect 6976 10310 6990 10362
rect 6990 10310 7002 10362
rect 7002 10310 7032 10362
rect 7056 10310 7066 10362
rect 7066 10310 7112 10362
rect 6816 10308 6872 10310
rect 6896 10308 6952 10310
rect 6976 10308 7032 10310
rect 7056 10308 7112 10310
rect 7756 18522 7812 18524
rect 7836 18522 7892 18524
rect 7916 18522 7972 18524
rect 7996 18522 8052 18524
rect 7756 18470 7802 18522
rect 7802 18470 7812 18522
rect 7836 18470 7866 18522
rect 7866 18470 7878 18522
rect 7878 18470 7892 18522
rect 7916 18470 7930 18522
rect 7930 18470 7942 18522
rect 7942 18470 7972 18522
rect 7996 18470 8006 18522
rect 8006 18470 8052 18522
rect 7756 18468 7812 18470
rect 7836 18468 7892 18470
rect 7916 18468 7972 18470
rect 7996 18468 8052 18470
rect 7756 17434 7812 17436
rect 7836 17434 7892 17436
rect 7916 17434 7972 17436
rect 7996 17434 8052 17436
rect 7756 17382 7802 17434
rect 7802 17382 7812 17434
rect 7836 17382 7866 17434
rect 7866 17382 7878 17434
rect 7878 17382 7892 17434
rect 7916 17382 7930 17434
rect 7930 17382 7942 17434
rect 7942 17382 7972 17434
rect 7996 17382 8006 17434
rect 8006 17382 8052 17434
rect 7756 17380 7812 17382
rect 7836 17380 7892 17382
rect 7916 17380 7972 17382
rect 7996 17380 8052 17382
rect 7756 16346 7812 16348
rect 7836 16346 7892 16348
rect 7916 16346 7972 16348
rect 7996 16346 8052 16348
rect 7756 16294 7802 16346
rect 7802 16294 7812 16346
rect 7836 16294 7866 16346
rect 7866 16294 7878 16346
rect 7878 16294 7892 16346
rect 7916 16294 7930 16346
rect 7930 16294 7942 16346
rect 7942 16294 7972 16346
rect 7996 16294 8006 16346
rect 8006 16294 8052 16346
rect 7756 16292 7812 16294
rect 7836 16292 7892 16294
rect 7916 16292 7972 16294
rect 7996 16292 8052 16294
rect 7756 15258 7812 15260
rect 7836 15258 7892 15260
rect 7916 15258 7972 15260
rect 7996 15258 8052 15260
rect 7756 15206 7802 15258
rect 7802 15206 7812 15258
rect 7836 15206 7866 15258
rect 7866 15206 7878 15258
rect 7878 15206 7892 15258
rect 7916 15206 7930 15258
rect 7930 15206 7942 15258
rect 7942 15206 7972 15258
rect 7996 15206 8006 15258
rect 8006 15206 8052 15258
rect 7756 15204 7812 15206
rect 7836 15204 7892 15206
rect 7916 15204 7972 15206
rect 7996 15204 8052 15206
rect 6816 9274 6872 9276
rect 6896 9274 6952 9276
rect 6976 9274 7032 9276
rect 7056 9274 7112 9276
rect 6816 9222 6862 9274
rect 6862 9222 6872 9274
rect 6896 9222 6926 9274
rect 6926 9222 6938 9274
rect 6938 9222 6952 9274
rect 6976 9222 6990 9274
rect 6990 9222 7002 9274
rect 7002 9222 7032 9274
rect 7056 9222 7066 9274
rect 7066 9222 7112 9274
rect 6816 9220 6872 9222
rect 6896 9220 6952 9222
rect 6976 9220 7032 9222
rect 7056 9220 7112 9222
rect 6816 8186 6872 8188
rect 6896 8186 6952 8188
rect 6976 8186 7032 8188
rect 7056 8186 7112 8188
rect 6816 8134 6862 8186
rect 6862 8134 6872 8186
rect 6896 8134 6926 8186
rect 6926 8134 6938 8186
rect 6938 8134 6952 8186
rect 6976 8134 6990 8186
rect 6990 8134 7002 8186
rect 7002 8134 7032 8186
rect 7056 8134 7066 8186
rect 7066 8134 7112 8186
rect 6816 8132 6872 8134
rect 6896 8132 6952 8134
rect 6976 8132 7032 8134
rect 7056 8132 7112 8134
rect 6816 7098 6872 7100
rect 6896 7098 6952 7100
rect 6976 7098 7032 7100
rect 7056 7098 7112 7100
rect 6816 7046 6862 7098
rect 6862 7046 6872 7098
rect 6896 7046 6926 7098
rect 6926 7046 6938 7098
rect 6938 7046 6952 7098
rect 6976 7046 6990 7098
rect 6990 7046 7002 7098
rect 7002 7046 7032 7098
rect 7056 7046 7066 7098
rect 7066 7046 7112 7098
rect 6816 7044 6872 7046
rect 6896 7044 6952 7046
rect 6976 7044 7032 7046
rect 7056 7044 7112 7046
rect 6816 6010 6872 6012
rect 6896 6010 6952 6012
rect 6976 6010 7032 6012
rect 7056 6010 7112 6012
rect 6816 5958 6862 6010
rect 6862 5958 6872 6010
rect 6896 5958 6926 6010
rect 6926 5958 6938 6010
rect 6938 5958 6952 6010
rect 6976 5958 6990 6010
rect 6990 5958 7002 6010
rect 7002 5958 7032 6010
rect 7056 5958 7066 6010
rect 7066 5958 7112 6010
rect 6816 5956 6872 5958
rect 6896 5956 6952 5958
rect 6976 5956 7032 5958
rect 7056 5956 7112 5958
rect 6816 4922 6872 4924
rect 6896 4922 6952 4924
rect 6976 4922 7032 4924
rect 7056 4922 7112 4924
rect 6816 4870 6862 4922
rect 6862 4870 6872 4922
rect 6896 4870 6926 4922
rect 6926 4870 6938 4922
rect 6938 4870 6952 4922
rect 6976 4870 6990 4922
rect 6990 4870 7002 4922
rect 7002 4870 7032 4922
rect 7056 4870 7066 4922
rect 7066 4870 7112 4922
rect 6816 4868 6872 4870
rect 6896 4868 6952 4870
rect 6976 4868 7032 4870
rect 7056 4868 7112 4870
rect 6816 3834 6872 3836
rect 6896 3834 6952 3836
rect 6976 3834 7032 3836
rect 7056 3834 7112 3836
rect 6816 3782 6862 3834
rect 6862 3782 6872 3834
rect 6896 3782 6926 3834
rect 6926 3782 6938 3834
rect 6938 3782 6952 3834
rect 6976 3782 6990 3834
rect 6990 3782 7002 3834
rect 7002 3782 7032 3834
rect 7056 3782 7066 3834
rect 7066 3782 7112 3834
rect 6816 3780 6872 3782
rect 6896 3780 6952 3782
rect 6976 3780 7032 3782
rect 7056 3780 7112 3782
rect 6816 2746 6872 2748
rect 6896 2746 6952 2748
rect 6976 2746 7032 2748
rect 7056 2746 7112 2748
rect 6816 2694 6862 2746
rect 6862 2694 6872 2746
rect 6896 2694 6926 2746
rect 6926 2694 6938 2746
rect 6938 2694 6952 2746
rect 6976 2694 6990 2746
rect 6990 2694 7002 2746
rect 7002 2694 7032 2746
rect 7056 2694 7066 2746
rect 7066 2694 7112 2746
rect 6816 2692 6872 2694
rect 6896 2692 6952 2694
rect 6976 2692 7032 2694
rect 7056 2692 7112 2694
rect 6816 1658 6872 1660
rect 6896 1658 6952 1660
rect 6976 1658 7032 1660
rect 7056 1658 7112 1660
rect 6816 1606 6862 1658
rect 6862 1606 6872 1658
rect 6896 1606 6926 1658
rect 6926 1606 6938 1658
rect 6938 1606 6952 1658
rect 6976 1606 6990 1658
rect 6990 1606 7002 1658
rect 7002 1606 7032 1658
rect 7056 1606 7066 1658
rect 7066 1606 7112 1658
rect 6816 1604 6872 1606
rect 6896 1604 6952 1606
rect 6976 1604 7032 1606
rect 7056 1604 7112 1606
rect 6156 1114 6212 1116
rect 6236 1114 6292 1116
rect 6316 1114 6372 1116
rect 6396 1114 6452 1116
rect 6156 1062 6202 1114
rect 6202 1062 6212 1114
rect 6236 1062 6266 1114
rect 6266 1062 6278 1114
rect 6278 1062 6292 1114
rect 6316 1062 6330 1114
rect 6330 1062 6342 1114
rect 6342 1062 6372 1114
rect 6396 1062 6406 1114
rect 6406 1062 6452 1114
rect 6156 1060 6212 1062
rect 6236 1060 6292 1062
rect 6316 1060 6372 1062
rect 6396 1060 6452 1062
rect 4986 720 5042 776
rect 7756 14170 7812 14172
rect 7836 14170 7892 14172
rect 7916 14170 7972 14172
rect 7996 14170 8052 14172
rect 7756 14118 7802 14170
rect 7802 14118 7812 14170
rect 7836 14118 7866 14170
rect 7866 14118 7878 14170
rect 7878 14118 7892 14170
rect 7916 14118 7930 14170
rect 7930 14118 7942 14170
rect 7942 14118 7972 14170
rect 7996 14118 8006 14170
rect 8006 14118 8052 14170
rect 7756 14116 7812 14118
rect 7836 14116 7892 14118
rect 7916 14116 7972 14118
rect 7996 14116 8052 14118
rect 8416 28858 8472 28860
rect 8496 28858 8552 28860
rect 8576 28858 8632 28860
rect 8656 28858 8712 28860
rect 8416 28806 8462 28858
rect 8462 28806 8472 28858
rect 8496 28806 8526 28858
rect 8526 28806 8538 28858
rect 8538 28806 8552 28858
rect 8576 28806 8590 28858
rect 8590 28806 8602 28858
rect 8602 28806 8632 28858
rect 8656 28806 8666 28858
rect 8666 28806 8712 28858
rect 8416 28804 8472 28806
rect 8496 28804 8552 28806
rect 8576 28804 8632 28806
rect 8656 28804 8712 28806
rect 8416 27770 8472 27772
rect 8496 27770 8552 27772
rect 8576 27770 8632 27772
rect 8656 27770 8712 27772
rect 8416 27718 8462 27770
rect 8462 27718 8472 27770
rect 8496 27718 8526 27770
rect 8526 27718 8538 27770
rect 8538 27718 8552 27770
rect 8576 27718 8590 27770
rect 8590 27718 8602 27770
rect 8602 27718 8632 27770
rect 8656 27718 8666 27770
rect 8666 27718 8712 27770
rect 8416 27716 8472 27718
rect 8496 27716 8552 27718
rect 8576 27716 8632 27718
rect 8656 27716 8712 27718
rect 8416 26682 8472 26684
rect 8496 26682 8552 26684
rect 8576 26682 8632 26684
rect 8656 26682 8712 26684
rect 8416 26630 8462 26682
rect 8462 26630 8472 26682
rect 8496 26630 8526 26682
rect 8526 26630 8538 26682
rect 8538 26630 8552 26682
rect 8576 26630 8590 26682
rect 8590 26630 8602 26682
rect 8602 26630 8632 26682
rect 8656 26630 8666 26682
rect 8666 26630 8712 26682
rect 8416 26628 8472 26630
rect 8496 26628 8552 26630
rect 8576 26628 8632 26630
rect 8656 26628 8712 26630
rect 8416 25594 8472 25596
rect 8496 25594 8552 25596
rect 8576 25594 8632 25596
rect 8656 25594 8712 25596
rect 8416 25542 8462 25594
rect 8462 25542 8472 25594
rect 8496 25542 8526 25594
rect 8526 25542 8538 25594
rect 8538 25542 8552 25594
rect 8576 25542 8590 25594
rect 8590 25542 8602 25594
rect 8602 25542 8632 25594
rect 8656 25542 8666 25594
rect 8666 25542 8712 25594
rect 8416 25540 8472 25542
rect 8496 25540 8552 25542
rect 8576 25540 8632 25542
rect 8656 25540 8712 25542
rect 8416 24506 8472 24508
rect 8496 24506 8552 24508
rect 8576 24506 8632 24508
rect 8656 24506 8712 24508
rect 8416 24454 8462 24506
rect 8462 24454 8472 24506
rect 8496 24454 8526 24506
rect 8526 24454 8538 24506
rect 8538 24454 8552 24506
rect 8576 24454 8590 24506
rect 8590 24454 8602 24506
rect 8602 24454 8632 24506
rect 8656 24454 8666 24506
rect 8666 24454 8712 24506
rect 8416 24452 8472 24454
rect 8496 24452 8552 24454
rect 8576 24452 8632 24454
rect 8656 24452 8712 24454
rect 8416 23418 8472 23420
rect 8496 23418 8552 23420
rect 8576 23418 8632 23420
rect 8656 23418 8712 23420
rect 8416 23366 8462 23418
rect 8462 23366 8472 23418
rect 8496 23366 8526 23418
rect 8526 23366 8538 23418
rect 8538 23366 8552 23418
rect 8576 23366 8590 23418
rect 8590 23366 8602 23418
rect 8602 23366 8632 23418
rect 8656 23366 8666 23418
rect 8666 23366 8712 23418
rect 8416 23364 8472 23366
rect 8496 23364 8552 23366
rect 8576 23364 8632 23366
rect 8656 23364 8712 23366
rect 8416 22330 8472 22332
rect 8496 22330 8552 22332
rect 8576 22330 8632 22332
rect 8656 22330 8712 22332
rect 8416 22278 8462 22330
rect 8462 22278 8472 22330
rect 8496 22278 8526 22330
rect 8526 22278 8538 22330
rect 8538 22278 8552 22330
rect 8576 22278 8590 22330
rect 8590 22278 8602 22330
rect 8602 22278 8632 22330
rect 8656 22278 8666 22330
rect 8666 22278 8712 22330
rect 8416 22276 8472 22278
rect 8496 22276 8552 22278
rect 8576 22276 8632 22278
rect 8656 22276 8712 22278
rect 8416 21242 8472 21244
rect 8496 21242 8552 21244
rect 8576 21242 8632 21244
rect 8656 21242 8712 21244
rect 8416 21190 8462 21242
rect 8462 21190 8472 21242
rect 8496 21190 8526 21242
rect 8526 21190 8538 21242
rect 8538 21190 8552 21242
rect 8576 21190 8590 21242
rect 8590 21190 8602 21242
rect 8602 21190 8632 21242
rect 8656 21190 8666 21242
rect 8666 21190 8712 21242
rect 8416 21188 8472 21190
rect 8496 21188 8552 21190
rect 8576 21188 8632 21190
rect 8656 21188 8712 21190
rect 8416 20154 8472 20156
rect 8496 20154 8552 20156
rect 8576 20154 8632 20156
rect 8656 20154 8712 20156
rect 8416 20102 8462 20154
rect 8462 20102 8472 20154
rect 8496 20102 8526 20154
rect 8526 20102 8538 20154
rect 8538 20102 8552 20154
rect 8576 20102 8590 20154
rect 8590 20102 8602 20154
rect 8602 20102 8632 20154
rect 8656 20102 8666 20154
rect 8666 20102 8712 20154
rect 8416 20100 8472 20102
rect 8496 20100 8552 20102
rect 8576 20100 8632 20102
rect 8656 20100 8712 20102
rect 8416 19066 8472 19068
rect 8496 19066 8552 19068
rect 8576 19066 8632 19068
rect 8656 19066 8712 19068
rect 8416 19014 8462 19066
rect 8462 19014 8472 19066
rect 8496 19014 8526 19066
rect 8526 19014 8538 19066
rect 8538 19014 8552 19066
rect 8576 19014 8590 19066
rect 8590 19014 8602 19066
rect 8602 19014 8632 19066
rect 8656 19014 8666 19066
rect 8666 19014 8712 19066
rect 8416 19012 8472 19014
rect 8496 19012 8552 19014
rect 8576 19012 8632 19014
rect 8656 19012 8712 19014
rect 8416 17978 8472 17980
rect 8496 17978 8552 17980
rect 8576 17978 8632 17980
rect 8656 17978 8712 17980
rect 8416 17926 8462 17978
rect 8462 17926 8472 17978
rect 8496 17926 8526 17978
rect 8526 17926 8538 17978
rect 8538 17926 8552 17978
rect 8576 17926 8590 17978
rect 8590 17926 8602 17978
rect 8602 17926 8632 17978
rect 8656 17926 8666 17978
rect 8666 17926 8712 17978
rect 8416 17924 8472 17926
rect 8496 17924 8552 17926
rect 8576 17924 8632 17926
rect 8656 17924 8712 17926
rect 8416 16890 8472 16892
rect 8496 16890 8552 16892
rect 8576 16890 8632 16892
rect 8656 16890 8712 16892
rect 8416 16838 8462 16890
rect 8462 16838 8472 16890
rect 8496 16838 8526 16890
rect 8526 16838 8538 16890
rect 8538 16838 8552 16890
rect 8576 16838 8590 16890
rect 8590 16838 8602 16890
rect 8602 16838 8632 16890
rect 8656 16838 8666 16890
rect 8666 16838 8712 16890
rect 8416 16836 8472 16838
rect 8496 16836 8552 16838
rect 8576 16836 8632 16838
rect 8656 16836 8712 16838
rect 9356 35930 9412 35932
rect 9436 35930 9492 35932
rect 9516 35930 9572 35932
rect 9596 35930 9652 35932
rect 9356 35878 9402 35930
rect 9402 35878 9412 35930
rect 9436 35878 9466 35930
rect 9466 35878 9478 35930
rect 9478 35878 9492 35930
rect 9516 35878 9530 35930
rect 9530 35878 9542 35930
rect 9542 35878 9572 35930
rect 9596 35878 9606 35930
rect 9606 35878 9652 35930
rect 9356 35876 9412 35878
rect 9436 35876 9492 35878
rect 9516 35876 9572 35878
rect 9596 35876 9652 35878
rect 9356 34842 9412 34844
rect 9436 34842 9492 34844
rect 9516 34842 9572 34844
rect 9596 34842 9652 34844
rect 9356 34790 9402 34842
rect 9402 34790 9412 34842
rect 9436 34790 9466 34842
rect 9466 34790 9478 34842
rect 9478 34790 9492 34842
rect 9516 34790 9530 34842
rect 9530 34790 9542 34842
rect 9542 34790 9572 34842
rect 9596 34790 9606 34842
rect 9606 34790 9652 34842
rect 9356 34788 9412 34790
rect 9436 34788 9492 34790
rect 9516 34788 9572 34790
rect 9596 34788 9652 34790
rect 9356 33754 9412 33756
rect 9436 33754 9492 33756
rect 9516 33754 9572 33756
rect 9596 33754 9652 33756
rect 9356 33702 9402 33754
rect 9402 33702 9412 33754
rect 9436 33702 9466 33754
rect 9466 33702 9478 33754
rect 9478 33702 9492 33754
rect 9516 33702 9530 33754
rect 9530 33702 9542 33754
rect 9542 33702 9572 33754
rect 9596 33702 9606 33754
rect 9606 33702 9652 33754
rect 9356 33700 9412 33702
rect 9436 33700 9492 33702
rect 9516 33700 9572 33702
rect 9596 33700 9652 33702
rect 9356 32666 9412 32668
rect 9436 32666 9492 32668
rect 9516 32666 9572 32668
rect 9596 32666 9652 32668
rect 9356 32614 9402 32666
rect 9402 32614 9412 32666
rect 9436 32614 9466 32666
rect 9466 32614 9478 32666
rect 9478 32614 9492 32666
rect 9516 32614 9530 32666
rect 9530 32614 9542 32666
rect 9542 32614 9572 32666
rect 9596 32614 9606 32666
rect 9606 32614 9652 32666
rect 9356 32612 9412 32614
rect 9436 32612 9492 32614
rect 9516 32612 9572 32614
rect 9596 32612 9652 32614
rect 9494 31728 9550 31784
rect 9356 31578 9412 31580
rect 9436 31578 9492 31580
rect 9516 31578 9572 31580
rect 9596 31578 9652 31580
rect 9356 31526 9402 31578
rect 9402 31526 9412 31578
rect 9436 31526 9466 31578
rect 9466 31526 9478 31578
rect 9478 31526 9492 31578
rect 9516 31526 9530 31578
rect 9530 31526 9542 31578
rect 9542 31526 9572 31578
rect 9596 31526 9606 31578
rect 9606 31526 9652 31578
rect 9356 31524 9412 31526
rect 9436 31524 9492 31526
rect 9516 31524 9572 31526
rect 9596 31524 9652 31526
rect 9356 30490 9412 30492
rect 9436 30490 9492 30492
rect 9516 30490 9572 30492
rect 9596 30490 9652 30492
rect 9356 30438 9402 30490
rect 9402 30438 9412 30490
rect 9436 30438 9466 30490
rect 9466 30438 9478 30490
rect 9478 30438 9492 30490
rect 9516 30438 9530 30490
rect 9530 30438 9542 30490
rect 9542 30438 9572 30490
rect 9596 30438 9606 30490
rect 9606 30438 9652 30490
rect 9356 30436 9412 30438
rect 9436 30436 9492 30438
rect 9516 30436 9572 30438
rect 9596 30436 9652 30438
rect 9356 29402 9412 29404
rect 9436 29402 9492 29404
rect 9516 29402 9572 29404
rect 9596 29402 9652 29404
rect 9356 29350 9402 29402
rect 9402 29350 9412 29402
rect 9436 29350 9466 29402
rect 9466 29350 9478 29402
rect 9478 29350 9492 29402
rect 9516 29350 9530 29402
rect 9530 29350 9542 29402
rect 9542 29350 9572 29402
rect 9596 29350 9606 29402
rect 9606 29350 9652 29402
rect 9356 29348 9412 29350
rect 9436 29348 9492 29350
rect 9516 29348 9572 29350
rect 9596 29348 9652 29350
rect 7756 13082 7812 13084
rect 7836 13082 7892 13084
rect 7916 13082 7972 13084
rect 7996 13082 8052 13084
rect 7756 13030 7802 13082
rect 7802 13030 7812 13082
rect 7836 13030 7866 13082
rect 7866 13030 7878 13082
rect 7878 13030 7892 13082
rect 7916 13030 7930 13082
rect 7930 13030 7942 13082
rect 7942 13030 7972 13082
rect 7996 13030 8006 13082
rect 8006 13030 8052 13082
rect 7756 13028 7812 13030
rect 7836 13028 7892 13030
rect 7916 13028 7972 13030
rect 7996 13028 8052 13030
rect 7756 11994 7812 11996
rect 7836 11994 7892 11996
rect 7916 11994 7972 11996
rect 7996 11994 8052 11996
rect 7756 11942 7802 11994
rect 7802 11942 7812 11994
rect 7836 11942 7866 11994
rect 7866 11942 7878 11994
rect 7878 11942 7892 11994
rect 7916 11942 7930 11994
rect 7930 11942 7942 11994
rect 7942 11942 7972 11994
rect 7996 11942 8006 11994
rect 8006 11942 8052 11994
rect 7756 11940 7812 11942
rect 7836 11940 7892 11942
rect 7916 11940 7972 11942
rect 7996 11940 8052 11942
rect 7756 10906 7812 10908
rect 7836 10906 7892 10908
rect 7916 10906 7972 10908
rect 7996 10906 8052 10908
rect 7756 10854 7802 10906
rect 7802 10854 7812 10906
rect 7836 10854 7866 10906
rect 7866 10854 7878 10906
rect 7878 10854 7892 10906
rect 7916 10854 7930 10906
rect 7930 10854 7942 10906
rect 7942 10854 7972 10906
rect 7996 10854 8006 10906
rect 8006 10854 8052 10906
rect 7756 10852 7812 10854
rect 7836 10852 7892 10854
rect 7916 10852 7972 10854
rect 7996 10852 8052 10854
rect 7756 9818 7812 9820
rect 7836 9818 7892 9820
rect 7916 9818 7972 9820
rect 7996 9818 8052 9820
rect 7756 9766 7802 9818
rect 7802 9766 7812 9818
rect 7836 9766 7866 9818
rect 7866 9766 7878 9818
rect 7878 9766 7892 9818
rect 7916 9766 7930 9818
rect 7930 9766 7942 9818
rect 7942 9766 7972 9818
rect 7996 9766 8006 9818
rect 8006 9766 8052 9818
rect 7756 9764 7812 9766
rect 7836 9764 7892 9766
rect 7916 9764 7972 9766
rect 7996 9764 8052 9766
rect 7756 8730 7812 8732
rect 7836 8730 7892 8732
rect 7916 8730 7972 8732
rect 7996 8730 8052 8732
rect 7756 8678 7802 8730
rect 7802 8678 7812 8730
rect 7836 8678 7866 8730
rect 7866 8678 7878 8730
rect 7878 8678 7892 8730
rect 7916 8678 7930 8730
rect 7930 8678 7942 8730
rect 7942 8678 7972 8730
rect 7996 8678 8006 8730
rect 8006 8678 8052 8730
rect 7756 8676 7812 8678
rect 7836 8676 7892 8678
rect 7916 8676 7972 8678
rect 7996 8676 8052 8678
rect 7756 7642 7812 7644
rect 7836 7642 7892 7644
rect 7916 7642 7972 7644
rect 7996 7642 8052 7644
rect 7756 7590 7802 7642
rect 7802 7590 7812 7642
rect 7836 7590 7866 7642
rect 7866 7590 7878 7642
rect 7878 7590 7892 7642
rect 7916 7590 7930 7642
rect 7930 7590 7942 7642
rect 7942 7590 7972 7642
rect 7996 7590 8006 7642
rect 8006 7590 8052 7642
rect 7756 7588 7812 7590
rect 7836 7588 7892 7590
rect 7916 7588 7972 7590
rect 7996 7588 8052 7590
rect 7756 6554 7812 6556
rect 7836 6554 7892 6556
rect 7916 6554 7972 6556
rect 7996 6554 8052 6556
rect 7756 6502 7802 6554
rect 7802 6502 7812 6554
rect 7836 6502 7866 6554
rect 7866 6502 7878 6554
rect 7878 6502 7892 6554
rect 7916 6502 7930 6554
rect 7930 6502 7942 6554
rect 7942 6502 7972 6554
rect 7996 6502 8006 6554
rect 8006 6502 8052 6554
rect 7756 6500 7812 6502
rect 7836 6500 7892 6502
rect 7916 6500 7972 6502
rect 7996 6500 8052 6502
rect 7756 5466 7812 5468
rect 7836 5466 7892 5468
rect 7916 5466 7972 5468
rect 7996 5466 8052 5468
rect 7756 5414 7802 5466
rect 7802 5414 7812 5466
rect 7836 5414 7866 5466
rect 7866 5414 7878 5466
rect 7878 5414 7892 5466
rect 7916 5414 7930 5466
rect 7930 5414 7942 5466
rect 7942 5414 7972 5466
rect 7996 5414 8006 5466
rect 8006 5414 8052 5466
rect 7756 5412 7812 5414
rect 7836 5412 7892 5414
rect 7916 5412 7972 5414
rect 7996 5412 8052 5414
rect 7756 4378 7812 4380
rect 7836 4378 7892 4380
rect 7916 4378 7972 4380
rect 7996 4378 8052 4380
rect 7756 4326 7802 4378
rect 7802 4326 7812 4378
rect 7836 4326 7866 4378
rect 7866 4326 7878 4378
rect 7878 4326 7892 4378
rect 7916 4326 7930 4378
rect 7930 4326 7942 4378
rect 7942 4326 7972 4378
rect 7996 4326 8006 4378
rect 8006 4326 8052 4378
rect 7756 4324 7812 4326
rect 7836 4324 7892 4326
rect 7916 4324 7972 4326
rect 7996 4324 8052 4326
rect 7756 3290 7812 3292
rect 7836 3290 7892 3292
rect 7916 3290 7972 3292
rect 7996 3290 8052 3292
rect 7756 3238 7802 3290
rect 7802 3238 7812 3290
rect 7836 3238 7866 3290
rect 7866 3238 7878 3290
rect 7878 3238 7892 3290
rect 7916 3238 7930 3290
rect 7930 3238 7942 3290
rect 7942 3238 7972 3290
rect 7996 3238 8006 3290
rect 8006 3238 8052 3290
rect 7756 3236 7812 3238
rect 7836 3236 7892 3238
rect 7916 3236 7972 3238
rect 7996 3236 8052 3238
rect 7756 2202 7812 2204
rect 7836 2202 7892 2204
rect 7916 2202 7972 2204
rect 7996 2202 8052 2204
rect 7756 2150 7802 2202
rect 7802 2150 7812 2202
rect 7836 2150 7866 2202
rect 7866 2150 7878 2202
rect 7878 2150 7892 2202
rect 7916 2150 7930 2202
rect 7930 2150 7942 2202
rect 7942 2150 7972 2202
rect 7996 2150 8006 2202
rect 8006 2150 8052 2202
rect 7756 2148 7812 2150
rect 7836 2148 7892 2150
rect 7916 2148 7972 2150
rect 7996 2148 8052 2150
rect 7756 1114 7812 1116
rect 7836 1114 7892 1116
rect 7916 1114 7972 1116
rect 7996 1114 8052 1116
rect 7756 1062 7802 1114
rect 7802 1062 7812 1114
rect 7836 1062 7866 1114
rect 7866 1062 7878 1114
rect 7878 1062 7892 1114
rect 7916 1062 7930 1114
rect 7930 1062 7942 1114
rect 7942 1062 7972 1114
rect 7996 1062 8006 1114
rect 8006 1062 8052 1114
rect 7756 1060 7812 1062
rect 7836 1060 7892 1062
rect 7916 1060 7972 1062
rect 7996 1060 8052 1062
rect 8416 15802 8472 15804
rect 8496 15802 8552 15804
rect 8576 15802 8632 15804
rect 8656 15802 8712 15804
rect 8416 15750 8462 15802
rect 8462 15750 8472 15802
rect 8496 15750 8526 15802
rect 8526 15750 8538 15802
rect 8538 15750 8552 15802
rect 8576 15750 8590 15802
rect 8590 15750 8602 15802
rect 8602 15750 8632 15802
rect 8656 15750 8666 15802
rect 8666 15750 8712 15802
rect 8416 15748 8472 15750
rect 8496 15748 8552 15750
rect 8576 15748 8632 15750
rect 8656 15748 8712 15750
rect 8416 14714 8472 14716
rect 8496 14714 8552 14716
rect 8576 14714 8632 14716
rect 8656 14714 8712 14716
rect 8416 14662 8462 14714
rect 8462 14662 8472 14714
rect 8496 14662 8526 14714
rect 8526 14662 8538 14714
rect 8538 14662 8552 14714
rect 8576 14662 8590 14714
rect 8590 14662 8602 14714
rect 8602 14662 8632 14714
rect 8656 14662 8666 14714
rect 8666 14662 8712 14714
rect 8416 14660 8472 14662
rect 8496 14660 8552 14662
rect 8576 14660 8632 14662
rect 8656 14660 8712 14662
rect 8416 13626 8472 13628
rect 8496 13626 8552 13628
rect 8576 13626 8632 13628
rect 8656 13626 8712 13628
rect 8416 13574 8462 13626
rect 8462 13574 8472 13626
rect 8496 13574 8526 13626
rect 8526 13574 8538 13626
rect 8538 13574 8552 13626
rect 8576 13574 8590 13626
rect 8590 13574 8602 13626
rect 8602 13574 8632 13626
rect 8656 13574 8666 13626
rect 8666 13574 8712 13626
rect 8416 13572 8472 13574
rect 8496 13572 8552 13574
rect 8576 13572 8632 13574
rect 8656 13572 8712 13574
rect 8416 12538 8472 12540
rect 8496 12538 8552 12540
rect 8576 12538 8632 12540
rect 8656 12538 8712 12540
rect 8416 12486 8462 12538
rect 8462 12486 8472 12538
rect 8496 12486 8526 12538
rect 8526 12486 8538 12538
rect 8538 12486 8552 12538
rect 8576 12486 8590 12538
rect 8590 12486 8602 12538
rect 8602 12486 8632 12538
rect 8656 12486 8666 12538
rect 8666 12486 8712 12538
rect 8416 12484 8472 12486
rect 8496 12484 8552 12486
rect 8576 12484 8632 12486
rect 8656 12484 8712 12486
rect 8416 11450 8472 11452
rect 8496 11450 8552 11452
rect 8576 11450 8632 11452
rect 8656 11450 8712 11452
rect 8416 11398 8462 11450
rect 8462 11398 8472 11450
rect 8496 11398 8526 11450
rect 8526 11398 8538 11450
rect 8538 11398 8552 11450
rect 8576 11398 8590 11450
rect 8590 11398 8602 11450
rect 8602 11398 8632 11450
rect 8656 11398 8666 11450
rect 8666 11398 8712 11450
rect 8416 11396 8472 11398
rect 8496 11396 8552 11398
rect 8576 11396 8632 11398
rect 8656 11396 8712 11398
rect 8416 10362 8472 10364
rect 8496 10362 8552 10364
rect 8576 10362 8632 10364
rect 8656 10362 8712 10364
rect 8416 10310 8462 10362
rect 8462 10310 8472 10362
rect 8496 10310 8526 10362
rect 8526 10310 8538 10362
rect 8538 10310 8552 10362
rect 8576 10310 8590 10362
rect 8590 10310 8602 10362
rect 8602 10310 8632 10362
rect 8656 10310 8666 10362
rect 8666 10310 8712 10362
rect 8416 10308 8472 10310
rect 8496 10308 8552 10310
rect 8576 10308 8632 10310
rect 8656 10308 8712 10310
rect 8416 9274 8472 9276
rect 8496 9274 8552 9276
rect 8576 9274 8632 9276
rect 8656 9274 8712 9276
rect 8416 9222 8462 9274
rect 8462 9222 8472 9274
rect 8496 9222 8526 9274
rect 8526 9222 8538 9274
rect 8538 9222 8552 9274
rect 8576 9222 8590 9274
rect 8590 9222 8602 9274
rect 8602 9222 8632 9274
rect 8656 9222 8666 9274
rect 8666 9222 8712 9274
rect 8416 9220 8472 9222
rect 8496 9220 8552 9222
rect 8576 9220 8632 9222
rect 8656 9220 8712 9222
rect 8416 8186 8472 8188
rect 8496 8186 8552 8188
rect 8576 8186 8632 8188
rect 8656 8186 8712 8188
rect 8416 8134 8462 8186
rect 8462 8134 8472 8186
rect 8496 8134 8526 8186
rect 8526 8134 8538 8186
rect 8538 8134 8552 8186
rect 8576 8134 8590 8186
rect 8590 8134 8602 8186
rect 8602 8134 8632 8186
rect 8656 8134 8666 8186
rect 8666 8134 8712 8186
rect 8416 8132 8472 8134
rect 8496 8132 8552 8134
rect 8576 8132 8632 8134
rect 8656 8132 8712 8134
rect 8416 7098 8472 7100
rect 8496 7098 8552 7100
rect 8576 7098 8632 7100
rect 8656 7098 8712 7100
rect 8416 7046 8462 7098
rect 8462 7046 8472 7098
rect 8496 7046 8526 7098
rect 8526 7046 8538 7098
rect 8538 7046 8552 7098
rect 8576 7046 8590 7098
rect 8590 7046 8602 7098
rect 8602 7046 8632 7098
rect 8656 7046 8666 7098
rect 8666 7046 8712 7098
rect 8416 7044 8472 7046
rect 8496 7044 8552 7046
rect 8576 7044 8632 7046
rect 8656 7044 8712 7046
rect 8416 6010 8472 6012
rect 8496 6010 8552 6012
rect 8576 6010 8632 6012
rect 8656 6010 8712 6012
rect 8416 5958 8462 6010
rect 8462 5958 8472 6010
rect 8496 5958 8526 6010
rect 8526 5958 8538 6010
rect 8538 5958 8552 6010
rect 8576 5958 8590 6010
rect 8590 5958 8602 6010
rect 8602 5958 8632 6010
rect 8656 5958 8666 6010
rect 8666 5958 8712 6010
rect 8416 5956 8472 5958
rect 8496 5956 8552 5958
rect 8576 5956 8632 5958
rect 8656 5956 8712 5958
rect 8416 4922 8472 4924
rect 8496 4922 8552 4924
rect 8576 4922 8632 4924
rect 8656 4922 8712 4924
rect 8416 4870 8462 4922
rect 8462 4870 8472 4922
rect 8496 4870 8526 4922
rect 8526 4870 8538 4922
rect 8538 4870 8552 4922
rect 8576 4870 8590 4922
rect 8590 4870 8602 4922
rect 8602 4870 8632 4922
rect 8656 4870 8666 4922
rect 8666 4870 8712 4922
rect 8416 4868 8472 4870
rect 8496 4868 8552 4870
rect 8576 4868 8632 4870
rect 8656 4868 8712 4870
rect 8416 3834 8472 3836
rect 8496 3834 8552 3836
rect 8576 3834 8632 3836
rect 8656 3834 8712 3836
rect 8416 3782 8462 3834
rect 8462 3782 8472 3834
rect 8496 3782 8526 3834
rect 8526 3782 8538 3834
rect 8538 3782 8552 3834
rect 8576 3782 8590 3834
rect 8590 3782 8602 3834
rect 8602 3782 8632 3834
rect 8656 3782 8666 3834
rect 8666 3782 8712 3834
rect 8416 3780 8472 3782
rect 8496 3780 8552 3782
rect 8576 3780 8632 3782
rect 8656 3780 8712 3782
rect 8416 2746 8472 2748
rect 8496 2746 8552 2748
rect 8576 2746 8632 2748
rect 8656 2746 8712 2748
rect 8416 2694 8462 2746
rect 8462 2694 8472 2746
rect 8496 2694 8526 2746
rect 8526 2694 8538 2746
rect 8538 2694 8552 2746
rect 8576 2694 8590 2746
rect 8590 2694 8602 2746
rect 8602 2694 8632 2746
rect 8656 2694 8666 2746
rect 8666 2694 8712 2746
rect 8416 2692 8472 2694
rect 8496 2692 8552 2694
rect 8576 2692 8632 2694
rect 8656 2692 8712 2694
rect 8416 1658 8472 1660
rect 8496 1658 8552 1660
rect 8576 1658 8632 1660
rect 8656 1658 8712 1660
rect 8416 1606 8462 1658
rect 8462 1606 8472 1658
rect 8496 1606 8526 1658
rect 8526 1606 8538 1658
rect 8538 1606 8552 1658
rect 8576 1606 8590 1658
rect 8590 1606 8602 1658
rect 8602 1606 8632 1658
rect 8656 1606 8666 1658
rect 8666 1606 8712 1658
rect 8416 1604 8472 1606
rect 8496 1604 8552 1606
rect 8576 1604 8632 1606
rect 8656 1604 8712 1606
rect 9356 28314 9412 28316
rect 9436 28314 9492 28316
rect 9516 28314 9572 28316
rect 9596 28314 9652 28316
rect 9356 28262 9402 28314
rect 9402 28262 9412 28314
rect 9436 28262 9466 28314
rect 9466 28262 9478 28314
rect 9478 28262 9492 28314
rect 9516 28262 9530 28314
rect 9530 28262 9542 28314
rect 9542 28262 9572 28314
rect 9596 28262 9606 28314
rect 9606 28262 9652 28314
rect 9356 28260 9412 28262
rect 9436 28260 9492 28262
rect 9516 28260 9572 28262
rect 9596 28260 9652 28262
rect 9356 27226 9412 27228
rect 9436 27226 9492 27228
rect 9516 27226 9572 27228
rect 9596 27226 9652 27228
rect 9356 27174 9402 27226
rect 9402 27174 9412 27226
rect 9436 27174 9466 27226
rect 9466 27174 9478 27226
rect 9478 27174 9492 27226
rect 9516 27174 9530 27226
rect 9530 27174 9542 27226
rect 9542 27174 9572 27226
rect 9596 27174 9606 27226
rect 9606 27174 9652 27226
rect 9356 27172 9412 27174
rect 9436 27172 9492 27174
rect 9516 27172 9572 27174
rect 9596 27172 9652 27174
rect 9356 26138 9412 26140
rect 9436 26138 9492 26140
rect 9516 26138 9572 26140
rect 9596 26138 9652 26140
rect 9356 26086 9402 26138
rect 9402 26086 9412 26138
rect 9436 26086 9466 26138
rect 9466 26086 9478 26138
rect 9478 26086 9492 26138
rect 9516 26086 9530 26138
rect 9530 26086 9542 26138
rect 9542 26086 9572 26138
rect 9596 26086 9606 26138
rect 9606 26086 9652 26138
rect 9356 26084 9412 26086
rect 9436 26084 9492 26086
rect 9516 26084 9572 26086
rect 9596 26084 9652 26086
rect 9356 25050 9412 25052
rect 9436 25050 9492 25052
rect 9516 25050 9572 25052
rect 9596 25050 9652 25052
rect 9356 24998 9402 25050
rect 9402 24998 9412 25050
rect 9436 24998 9466 25050
rect 9466 24998 9478 25050
rect 9478 24998 9492 25050
rect 9516 24998 9530 25050
rect 9530 24998 9542 25050
rect 9542 24998 9572 25050
rect 9596 24998 9606 25050
rect 9606 24998 9652 25050
rect 9356 24996 9412 24998
rect 9436 24996 9492 24998
rect 9516 24996 9572 24998
rect 9596 24996 9652 24998
rect 9356 23962 9412 23964
rect 9436 23962 9492 23964
rect 9516 23962 9572 23964
rect 9596 23962 9652 23964
rect 9356 23910 9402 23962
rect 9402 23910 9412 23962
rect 9436 23910 9466 23962
rect 9466 23910 9478 23962
rect 9478 23910 9492 23962
rect 9516 23910 9530 23962
rect 9530 23910 9542 23962
rect 9542 23910 9572 23962
rect 9596 23910 9606 23962
rect 9606 23910 9652 23962
rect 9356 23908 9412 23910
rect 9436 23908 9492 23910
rect 9516 23908 9572 23910
rect 9596 23908 9652 23910
rect 9356 22874 9412 22876
rect 9436 22874 9492 22876
rect 9516 22874 9572 22876
rect 9596 22874 9652 22876
rect 9356 22822 9402 22874
rect 9402 22822 9412 22874
rect 9436 22822 9466 22874
rect 9466 22822 9478 22874
rect 9478 22822 9492 22874
rect 9516 22822 9530 22874
rect 9530 22822 9542 22874
rect 9542 22822 9572 22874
rect 9596 22822 9606 22874
rect 9606 22822 9652 22874
rect 9356 22820 9412 22822
rect 9436 22820 9492 22822
rect 9516 22820 9572 22822
rect 9596 22820 9652 22822
rect 9356 21786 9412 21788
rect 9436 21786 9492 21788
rect 9516 21786 9572 21788
rect 9596 21786 9652 21788
rect 9356 21734 9402 21786
rect 9402 21734 9412 21786
rect 9436 21734 9466 21786
rect 9466 21734 9478 21786
rect 9478 21734 9492 21786
rect 9516 21734 9530 21786
rect 9530 21734 9542 21786
rect 9542 21734 9572 21786
rect 9596 21734 9606 21786
rect 9606 21734 9652 21786
rect 9356 21732 9412 21734
rect 9436 21732 9492 21734
rect 9516 21732 9572 21734
rect 9596 21732 9652 21734
rect 9356 20698 9412 20700
rect 9436 20698 9492 20700
rect 9516 20698 9572 20700
rect 9596 20698 9652 20700
rect 9356 20646 9402 20698
rect 9402 20646 9412 20698
rect 9436 20646 9466 20698
rect 9466 20646 9478 20698
rect 9478 20646 9492 20698
rect 9516 20646 9530 20698
rect 9530 20646 9542 20698
rect 9542 20646 9572 20698
rect 9596 20646 9606 20698
rect 9606 20646 9652 20698
rect 9356 20644 9412 20646
rect 9436 20644 9492 20646
rect 9516 20644 9572 20646
rect 9596 20644 9652 20646
rect 9356 19610 9412 19612
rect 9436 19610 9492 19612
rect 9516 19610 9572 19612
rect 9596 19610 9652 19612
rect 9356 19558 9402 19610
rect 9402 19558 9412 19610
rect 9436 19558 9466 19610
rect 9466 19558 9478 19610
rect 9478 19558 9492 19610
rect 9516 19558 9530 19610
rect 9530 19558 9542 19610
rect 9542 19558 9572 19610
rect 9596 19558 9606 19610
rect 9606 19558 9652 19610
rect 9356 19556 9412 19558
rect 9436 19556 9492 19558
rect 9516 19556 9572 19558
rect 9596 19556 9652 19558
rect 9356 18522 9412 18524
rect 9436 18522 9492 18524
rect 9516 18522 9572 18524
rect 9596 18522 9652 18524
rect 9356 18470 9402 18522
rect 9402 18470 9412 18522
rect 9436 18470 9466 18522
rect 9466 18470 9478 18522
rect 9478 18470 9492 18522
rect 9516 18470 9530 18522
rect 9530 18470 9542 18522
rect 9542 18470 9572 18522
rect 9596 18470 9606 18522
rect 9606 18470 9652 18522
rect 9356 18468 9412 18470
rect 9436 18468 9492 18470
rect 9516 18468 9572 18470
rect 9596 18468 9652 18470
rect 9356 17434 9412 17436
rect 9436 17434 9492 17436
rect 9516 17434 9572 17436
rect 9596 17434 9652 17436
rect 9356 17382 9402 17434
rect 9402 17382 9412 17434
rect 9436 17382 9466 17434
rect 9466 17382 9478 17434
rect 9478 17382 9492 17434
rect 9516 17382 9530 17434
rect 9530 17382 9542 17434
rect 9542 17382 9572 17434
rect 9596 17382 9606 17434
rect 9606 17382 9652 17434
rect 9356 17380 9412 17382
rect 9436 17380 9492 17382
rect 9516 17380 9572 17382
rect 9596 17380 9652 17382
rect 9356 16346 9412 16348
rect 9436 16346 9492 16348
rect 9516 16346 9572 16348
rect 9596 16346 9652 16348
rect 9356 16294 9402 16346
rect 9402 16294 9412 16346
rect 9436 16294 9466 16346
rect 9466 16294 9478 16346
rect 9478 16294 9492 16346
rect 9516 16294 9530 16346
rect 9530 16294 9542 16346
rect 9542 16294 9572 16346
rect 9596 16294 9606 16346
rect 9606 16294 9652 16346
rect 9356 16292 9412 16294
rect 9436 16292 9492 16294
rect 9516 16292 9572 16294
rect 9596 16292 9652 16294
rect 9356 15258 9412 15260
rect 9436 15258 9492 15260
rect 9516 15258 9572 15260
rect 9596 15258 9652 15260
rect 9356 15206 9402 15258
rect 9402 15206 9412 15258
rect 9436 15206 9466 15258
rect 9466 15206 9478 15258
rect 9478 15206 9492 15258
rect 9516 15206 9530 15258
rect 9530 15206 9542 15258
rect 9542 15206 9572 15258
rect 9596 15206 9606 15258
rect 9606 15206 9652 15258
rect 9356 15204 9412 15206
rect 9436 15204 9492 15206
rect 9516 15204 9572 15206
rect 9596 15204 9652 15206
rect 10506 69264 10562 69320
rect 10956 85978 11012 85980
rect 11036 85978 11092 85980
rect 11116 85978 11172 85980
rect 11196 85978 11252 85980
rect 10956 85926 11002 85978
rect 11002 85926 11012 85978
rect 11036 85926 11066 85978
rect 11066 85926 11078 85978
rect 11078 85926 11092 85978
rect 11116 85926 11130 85978
rect 11130 85926 11142 85978
rect 11142 85926 11172 85978
rect 11196 85926 11206 85978
rect 11206 85926 11252 85978
rect 10956 85924 11012 85926
rect 11036 85924 11092 85926
rect 11116 85924 11172 85926
rect 11196 85924 11252 85926
rect 10506 38120 10562 38176
rect 10414 31456 10470 31512
rect 10322 29688 10378 29744
rect 9356 14170 9412 14172
rect 9436 14170 9492 14172
rect 9516 14170 9572 14172
rect 9596 14170 9652 14172
rect 9356 14118 9402 14170
rect 9402 14118 9412 14170
rect 9436 14118 9466 14170
rect 9466 14118 9478 14170
rect 9478 14118 9492 14170
rect 9516 14118 9530 14170
rect 9530 14118 9542 14170
rect 9542 14118 9572 14170
rect 9596 14118 9606 14170
rect 9606 14118 9652 14170
rect 9356 14116 9412 14118
rect 9436 14116 9492 14118
rect 9516 14116 9572 14118
rect 9596 14116 9652 14118
rect 9356 13082 9412 13084
rect 9436 13082 9492 13084
rect 9516 13082 9572 13084
rect 9596 13082 9652 13084
rect 9356 13030 9402 13082
rect 9402 13030 9412 13082
rect 9436 13030 9466 13082
rect 9466 13030 9478 13082
rect 9478 13030 9492 13082
rect 9516 13030 9530 13082
rect 9530 13030 9542 13082
rect 9542 13030 9572 13082
rect 9596 13030 9606 13082
rect 9606 13030 9652 13082
rect 9356 13028 9412 13030
rect 9436 13028 9492 13030
rect 9516 13028 9572 13030
rect 9596 13028 9652 13030
rect 9356 11994 9412 11996
rect 9436 11994 9492 11996
rect 9516 11994 9572 11996
rect 9596 11994 9652 11996
rect 9356 11942 9402 11994
rect 9402 11942 9412 11994
rect 9436 11942 9466 11994
rect 9466 11942 9478 11994
rect 9478 11942 9492 11994
rect 9516 11942 9530 11994
rect 9530 11942 9542 11994
rect 9542 11942 9572 11994
rect 9596 11942 9606 11994
rect 9606 11942 9652 11994
rect 9356 11940 9412 11942
rect 9436 11940 9492 11942
rect 9516 11940 9572 11942
rect 9596 11940 9652 11942
rect 9586 11192 9642 11248
rect 9356 10906 9412 10908
rect 9436 10906 9492 10908
rect 9516 10906 9572 10908
rect 9596 10906 9652 10908
rect 9356 10854 9402 10906
rect 9402 10854 9412 10906
rect 9436 10854 9466 10906
rect 9466 10854 9478 10906
rect 9478 10854 9492 10906
rect 9516 10854 9530 10906
rect 9530 10854 9542 10906
rect 9542 10854 9572 10906
rect 9596 10854 9606 10906
rect 9606 10854 9652 10906
rect 9356 10852 9412 10854
rect 9436 10852 9492 10854
rect 9516 10852 9572 10854
rect 9596 10852 9652 10854
rect 9356 9818 9412 9820
rect 9436 9818 9492 9820
rect 9516 9818 9572 9820
rect 9596 9818 9652 9820
rect 9356 9766 9402 9818
rect 9402 9766 9412 9818
rect 9436 9766 9466 9818
rect 9466 9766 9478 9818
rect 9478 9766 9492 9818
rect 9516 9766 9530 9818
rect 9530 9766 9542 9818
rect 9542 9766 9572 9818
rect 9596 9766 9606 9818
rect 9606 9766 9652 9818
rect 9356 9764 9412 9766
rect 9436 9764 9492 9766
rect 9516 9764 9572 9766
rect 9596 9764 9652 9766
rect 9356 8730 9412 8732
rect 9436 8730 9492 8732
rect 9516 8730 9572 8732
rect 9596 8730 9652 8732
rect 9356 8678 9402 8730
rect 9402 8678 9412 8730
rect 9436 8678 9466 8730
rect 9466 8678 9478 8730
rect 9478 8678 9492 8730
rect 9516 8678 9530 8730
rect 9530 8678 9542 8730
rect 9542 8678 9572 8730
rect 9596 8678 9606 8730
rect 9606 8678 9652 8730
rect 9356 8676 9412 8678
rect 9436 8676 9492 8678
rect 9516 8676 9572 8678
rect 9596 8676 9652 8678
rect 9356 7642 9412 7644
rect 9436 7642 9492 7644
rect 9516 7642 9572 7644
rect 9596 7642 9652 7644
rect 9356 7590 9402 7642
rect 9402 7590 9412 7642
rect 9436 7590 9466 7642
rect 9466 7590 9478 7642
rect 9478 7590 9492 7642
rect 9516 7590 9530 7642
rect 9530 7590 9542 7642
rect 9542 7590 9572 7642
rect 9596 7590 9606 7642
rect 9606 7590 9652 7642
rect 9356 7588 9412 7590
rect 9436 7588 9492 7590
rect 9516 7588 9572 7590
rect 9596 7588 9652 7590
rect 9356 6554 9412 6556
rect 9436 6554 9492 6556
rect 9516 6554 9572 6556
rect 9596 6554 9652 6556
rect 9356 6502 9402 6554
rect 9402 6502 9412 6554
rect 9436 6502 9466 6554
rect 9466 6502 9478 6554
rect 9478 6502 9492 6554
rect 9516 6502 9530 6554
rect 9530 6502 9542 6554
rect 9542 6502 9572 6554
rect 9596 6502 9606 6554
rect 9606 6502 9652 6554
rect 9356 6500 9412 6502
rect 9436 6500 9492 6502
rect 9516 6500 9572 6502
rect 9596 6500 9652 6502
rect 9356 5466 9412 5468
rect 9436 5466 9492 5468
rect 9516 5466 9572 5468
rect 9596 5466 9652 5468
rect 9356 5414 9402 5466
rect 9402 5414 9412 5466
rect 9436 5414 9466 5466
rect 9466 5414 9478 5466
rect 9478 5414 9492 5466
rect 9516 5414 9530 5466
rect 9530 5414 9542 5466
rect 9542 5414 9572 5466
rect 9596 5414 9606 5466
rect 9606 5414 9652 5466
rect 9356 5412 9412 5414
rect 9436 5412 9492 5414
rect 9516 5412 9572 5414
rect 9596 5412 9652 5414
rect 9356 4378 9412 4380
rect 9436 4378 9492 4380
rect 9516 4378 9572 4380
rect 9596 4378 9652 4380
rect 9356 4326 9402 4378
rect 9402 4326 9412 4378
rect 9436 4326 9466 4378
rect 9466 4326 9478 4378
rect 9478 4326 9492 4378
rect 9516 4326 9530 4378
rect 9530 4326 9542 4378
rect 9542 4326 9572 4378
rect 9596 4326 9606 4378
rect 9606 4326 9652 4378
rect 9356 4324 9412 4326
rect 9436 4324 9492 4326
rect 9516 4324 9572 4326
rect 9596 4324 9652 4326
rect 9356 3290 9412 3292
rect 9436 3290 9492 3292
rect 9516 3290 9572 3292
rect 9596 3290 9652 3292
rect 9356 3238 9402 3290
rect 9402 3238 9412 3290
rect 9436 3238 9466 3290
rect 9466 3238 9478 3290
rect 9478 3238 9492 3290
rect 9516 3238 9530 3290
rect 9530 3238 9542 3290
rect 9542 3238 9572 3290
rect 9596 3238 9606 3290
rect 9606 3238 9652 3290
rect 9356 3236 9412 3238
rect 9436 3236 9492 3238
rect 9516 3236 9572 3238
rect 9596 3236 9652 3238
rect 9356 2202 9412 2204
rect 9436 2202 9492 2204
rect 9516 2202 9572 2204
rect 9596 2202 9652 2204
rect 9356 2150 9402 2202
rect 9402 2150 9412 2202
rect 9436 2150 9466 2202
rect 9466 2150 9478 2202
rect 9478 2150 9492 2202
rect 9516 2150 9530 2202
rect 9530 2150 9542 2202
rect 9542 2150 9572 2202
rect 9596 2150 9606 2202
rect 9606 2150 9652 2202
rect 9356 2148 9412 2150
rect 9436 2148 9492 2150
rect 9516 2148 9572 2150
rect 9596 2148 9652 2150
rect 9356 1114 9412 1116
rect 9436 1114 9492 1116
rect 9516 1114 9572 1116
rect 9596 1114 9652 1116
rect 9356 1062 9402 1114
rect 9402 1062 9412 1114
rect 9436 1062 9466 1114
rect 9466 1062 9478 1114
rect 9478 1062 9492 1114
rect 9516 1062 9530 1114
rect 9530 1062 9542 1114
rect 9542 1062 9572 1114
rect 9596 1062 9606 1114
rect 9606 1062 9652 1114
rect 9356 1060 9412 1062
rect 9436 1060 9492 1062
rect 9516 1060 9572 1062
rect 9596 1060 9652 1062
rect 1306 312 1362 368
rect 10016 1658 10072 1660
rect 10096 1658 10152 1660
rect 10176 1658 10232 1660
rect 10256 1658 10312 1660
rect 10016 1606 10062 1658
rect 10062 1606 10072 1658
rect 10096 1606 10126 1658
rect 10126 1606 10138 1658
rect 10138 1606 10152 1658
rect 10176 1606 10190 1658
rect 10190 1606 10202 1658
rect 10202 1606 10232 1658
rect 10256 1606 10266 1658
rect 10266 1606 10312 1658
rect 10016 1604 10072 1606
rect 10096 1604 10152 1606
rect 10176 1604 10232 1606
rect 10256 1604 10312 1606
rect 11616 86522 11672 86524
rect 11696 86522 11752 86524
rect 11776 86522 11832 86524
rect 11856 86522 11912 86524
rect 11616 86470 11662 86522
rect 11662 86470 11672 86522
rect 11696 86470 11726 86522
rect 11726 86470 11738 86522
rect 11738 86470 11752 86522
rect 11776 86470 11790 86522
rect 11790 86470 11802 86522
rect 11802 86470 11832 86522
rect 11856 86470 11866 86522
rect 11866 86470 11912 86522
rect 11616 86468 11672 86470
rect 11696 86468 11752 86470
rect 11776 86468 11832 86470
rect 11856 86468 11912 86470
rect 13216 86522 13272 86524
rect 13296 86522 13352 86524
rect 13376 86522 13432 86524
rect 13456 86522 13512 86524
rect 13216 86470 13262 86522
rect 13262 86470 13272 86522
rect 13296 86470 13326 86522
rect 13326 86470 13338 86522
rect 13338 86470 13352 86522
rect 13376 86470 13390 86522
rect 13390 86470 13402 86522
rect 13402 86470 13432 86522
rect 13456 86470 13466 86522
rect 13466 86470 13512 86522
rect 13216 86468 13272 86470
rect 13296 86468 13352 86470
rect 13376 86468 13432 86470
rect 13456 86468 13512 86470
rect 14816 86522 14872 86524
rect 14896 86522 14952 86524
rect 14976 86522 15032 86524
rect 15056 86522 15112 86524
rect 14816 86470 14862 86522
rect 14862 86470 14872 86522
rect 14896 86470 14926 86522
rect 14926 86470 14938 86522
rect 14938 86470 14952 86522
rect 14976 86470 14990 86522
rect 14990 86470 15002 86522
rect 15002 86470 15032 86522
rect 15056 86470 15066 86522
rect 15066 86470 15112 86522
rect 14816 86468 14872 86470
rect 14896 86468 14952 86470
rect 14976 86468 15032 86470
rect 15056 86468 15112 86470
rect 16416 86522 16472 86524
rect 16496 86522 16552 86524
rect 16576 86522 16632 86524
rect 16656 86522 16712 86524
rect 16416 86470 16462 86522
rect 16462 86470 16472 86522
rect 16496 86470 16526 86522
rect 16526 86470 16538 86522
rect 16538 86470 16552 86522
rect 16576 86470 16590 86522
rect 16590 86470 16602 86522
rect 16602 86470 16632 86522
rect 16656 86470 16666 86522
rect 16666 86470 16712 86522
rect 16416 86468 16472 86470
rect 16496 86468 16552 86470
rect 16576 86468 16632 86470
rect 16656 86468 16712 86470
rect 11886 65048 11942 65104
rect 10690 3304 10746 3360
rect 11334 11192 11390 11248
rect 11334 9560 11390 9616
rect 12556 85978 12612 85980
rect 12636 85978 12692 85980
rect 12716 85978 12772 85980
rect 12796 85978 12852 85980
rect 12556 85926 12602 85978
rect 12602 85926 12612 85978
rect 12636 85926 12666 85978
rect 12666 85926 12678 85978
rect 12678 85926 12692 85978
rect 12716 85926 12730 85978
rect 12730 85926 12742 85978
rect 12742 85926 12772 85978
rect 12796 85926 12806 85978
rect 12806 85926 12852 85978
rect 12556 85924 12612 85926
rect 12636 85924 12692 85926
rect 12716 85924 12772 85926
rect 12796 85924 12852 85926
rect 18016 86522 18072 86524
rect 18096 86522 18152 86524
rect 18176 86522 18232 86524
rect 18256 86522 18312 86524
rect 18016 86470 18062 86522
rect 18062 86470 18072 86522
rect 18096 86470 18126 86522
rect 18126 86470 18138 86522
rect 18138 86470 18152 86522
rect 18176 86470 18190 86522
rect 18190 86470 18202 86522
rect 18202 86470 18232 86522
rect 18256 86470 18266 86522
rect 18266 86470 18312 86522
rect 18016 86468 18072 86470
rect 18096 86468 18152 86470
rect 18176 86468 18232 86470
rect 18256 86468 18312 86470
rect 19616 86522 19672 86524
rect 19696 86522 19752 86524
rect 19776 86522 19832 86524
rect 19856 86522 19912 86524
rect 19616 86470 19662 86522
rect 19662 86470 19672 86522
rect 19696 86470 19726 86522
rect 19726 86470 19738 86522
rect 19738 86470 19752 86522
rect 19776 86470 19790 86522
rect 19790 86470 19802 86522
rect 19802 86470 19832 86522
rect 19856 86470 19866 86522
rect 19866 86470 19912 86522
rect 19616 86468 19672 86470
rect 19696 86468 19752 86470
rect 19776 86468 19832 86470
rect 19856 86468 19912 86470
rect 21216 86522 21272 86524
rect 21296 86522 21352 86524
rect 21376 86522 21432 86524
rect 21456 86522 21512 86524
rect 21216 86470 21262 86522
rect 21262 86470 21272 86522
rect 21296 86470 21326 86522
rect 21326 86470 21338 86522
rect 21338 86470 21352 86522
rect 21376 86470 21390 86522
rect 21390 86470 21402 86522
rect 21402 86470 21432 86522
rect 21456 86470 21466 86522
rect 21466 86470 21512 86522
rect 21216 86468 21272 86470
rect 21296 86468 21352 86470
rect 21376 86468 21432 86470
rect 21456 86468 21512 86470
rect 22816 86522 22872 86524
rect 22896 86522 22952 86524
rect 22976 86522 23032 86524
rect 23056 86522 23112 86524
rect 22816 86470 22862 86522
rect 22862 86470 22872 86522
rect 22896 86470 22926 86522
rect 22926 86470 22938 86522
rect 22938 86470 22952 86522
rect 22976 86470 22990 86522
rect 22990 86470 23002 86522
rect 23002 86470 23032 86522
rect 23056 86470 23066 86522
rect 23066 86470 23112 86522
rect 22816 86468 22872 86470
rect 22896 86468 22952 86470
rect 22976 86468 23032 86470
rect 23056 86468 23112 86470
rect 24416 86522 24472 86524
rect 24496 86522 24552 86524
rect 24576 86522 24632 86524
rect 24656 86522 24712 86524
rect 24416 86470 24462 86522
rect 24462 86470 24472 86522
rect 24496 86470 24526 86522
rect 24526 86470 24538 86522
rect 24538 86470 24552 86522
rect 24576 86470 24590 86522
rect 24590 86470 24602 86522
rect 24602 86470 24632 86522
rect 24656 86470 24666 86522
rect 24666 86470 24712 86522
rect 24416 86468 24472 86470
rect 24496 86468 24552 86470
rect 24576 86468 24632 86470
rect 24656 86468 24712 86470
rect 26016 86522 26072 86524
rect 26096 86522 26152 86524
rect 26176 86522 26232 86524
rect 26256 86522 26312 86524
rect 26016 86470 26062 86522
rect 26062 86470 26072 86522
rect 26096 86470 26126 86522
rect 26126 86470 26138 86522
rect 26138 86470 26152 86522
rect 26176 86470 26190 86522
rect 26190 86470 26202 86522
rect 26202 86470 26232 86522
rect 26256 86470 26266 86522
rect 26266 86470 26312 86522
rect 26016 86468 26072 86470
rect 26096 86468 26152 86470
rect 26176 86468 26232 86470
rect 26256 86468 26312 86470
rect 14156 85978 14212 85980
rect 14236 85978 14292 85980
rect 14316 85978 14372 85980
rect 14396 85978 14452 85980
rect 14156 85926 14202 85978
rect 14202 85926 14212 85978
rect 14236 85926 14266 85978
rect 14266 85926 14278 85978
rect 14278 85926 14292 85978
rect 14316 85926 14330 85978
rect 14330 85926 14342 85978
rect 14342 85926 14372 85978
rect 14396 85926 14406 85978
rect 14406 85926 14452 85978
rect 14156 85924 14212 85926
rect 14236 85924 14292 85926
rect 14316 85924 14372 85926
rect 14396 85924 14452 85926
rect 15756 85978 15812 85980
rect 15836 85978 15892 85980
rect 15916 85978 15972 85980
rect 15996 85978 16052 85980
rect 15756 85926 15802 85978
rect 15802 85926 15812 85978
rect 15836 85926 15866 85978
rect 15866 85926 15878 85978
rect 15878 85926 15892 85978
rect 15916 85926 15930 85978
rect 15930 85926 15942 85978
rect 15942 85926 15972 85978
rect 15996 85926 16006 85978
rect 16006 85926 16052 85978
rect 15756 85924 15812 85926
rect 15836 85924 15892 85926
rect 15916 85924 15972 85926
rect 15996 85924 16052 85926
rect 17356 85978 17412 85980
rect 17436 85978 17492 85980
rect 17516 85978 17572 85980
rect 17596 85978 17652 85980
rect 17356 85926 17402 85978
rect 17402 85926 17412 85978
rect 17436 85926 17466 85978
rect 17466 85926 17478 85978
rect 17478 85926 17492 85978
rect 17516 85926 17530 85978
rect 17530 85926 17542 85978
rect 17542 85926 17572 85978
rect 17596 85926 17606 85978
rect 17606 85926 17652 85978
rect 17356 85924 17412 85926
rect 17436 85924 17492 85926
rect 17516 85924 17572 85926
rect 17596 85924 17652 85926
rect 18956 85978 19012 85980
rect 19036 85978 19092 85980
rect 19116 85978 19172 85980
rect 19196 85978 19252 85980
rect 18956 85926 19002 85978
rect 19002 85926 19012 85978
rect 19036 85926 19066 85978
rect 19066 85926 19078 85978
rect 19078 85926 19092 85978
rect 19116 85926 19130 85978
rect 19130 85926 19142 85978
rect 19142 85926 19172 85978
rect 19196 85926 19206 85978
rect 19206 85926 19252 85978
rect 18956 85924 19012 85926
rect 19036 85924 19092 85926
rect 19116 85924 19172 85926
rect 19196 85924 19252 85926
rect 20556 85978 20612 85980
rect 20636 85978 20692 85980
rect 20716 85978 20772 85980
rect 20796 85978 20852 85980
rect 20556 85926 20602 85978
rect 20602 85926 20612 85978
rect 20636 85926 20666 85978
rect 20666 85926 20678 85978
rect 20678 85926 20692 85978
rect 20716 85926 20730 85978
rect 20730 85926 20742 85978
rect 20742 85926 20772 85978
rect 20796 85926 20806 85978
rect 20806 85926 20852 85978
rect 20556 85924 20612 85926
rect 20636 85924 20692 85926
rect 20716 85924 20772 85926
rect 20796 85924 20852 85926
rect 22156 85978 22212 85980
rect 22236 85978 22292 85980
rect 22316 85978 22372 85980
rect 22396 85978 22452 85980
rect 22156 85926 22202 85978
rect 22202 85926 22212 85978
rect 22236 85926 22266 85978
rect 22266 85926 22278 85978
rect 22278 85926 22292 85978
rect 22316 85926 22330 85978
rect 22330 85926 22342 85978
rect 22342 85926 22372 85978
rect 22396 85926 22406 85978
rect 22406 85926 22452 85978
rect 22156 85924 22212 85926
rect 22236 85924 22292 85926
rect 22316 85924 22372 85926
rect 22396 85924 22452 85926
rect 23756 85978 23812 85980
rect 23836 85978 23892 85980
rect 23916 85978 23972 85980
rect 23996 85978 24052 85980
rect 23756 85926 23802 85978
rect 23802 85926 23812 85978
rect 23836 85926 23866 85978
rect 23866 85926 23878 85978
rect 23878 85926 23892 85978
rect 23916 85926 23930 85978
rect 23930 85926 23942 85978
rect 23942 85926 23972 85978
rect 23996 85926 24006 85978
rect 24006 85926 24052 85978
rect 23756 85924 23812 85926
rect 23836 85924 23892 85926
rect 23916 85924 23972 85926
rect 23996 85924 24052 85926
rect 25356 85978 25412 85980
rect 25436 85978 25492 85980
rect 25516 85978 25572 85980
rect 25596 85978 25652 85980
rect 25356 85926 25402 85978
rect 25402 85926 25412 85978
rect 25436 85926 25466 85978
rect 25466 85926 25478 85978
rect 25478 85926 25492 85978
rect 25516 85926 25530 85978
rect 25530 85926 25542 85978
rect 25542 85926 25572 85978
rect 25596 85926 25606 85978
rect 25606 85926 25652 85978
rect 25356 85924 25412 85926
rect 25436 85924 25492 85926
rect 25516 85924 25572 85926
rect 25596 85924 25652 85926
rect 26956 85978 27012 85980
rect 27036 85978 27092 85980
rect 27116 85978 27172 85980
rect 27196 85978 27252 85980
rect 26956 85926 27002 85978
rect 27002 85926 27012 85978
rect 27036 85926 27066 85978
rect 27066 85926 27078 85978
rect 27078 85926 27092 85978
rect 27116 85926 27130 85978
rect 27130 85926 27142 85978
rect 27142 85926 27172 85978
rect 27196 85926 27206 85978
rect 27206 85926 27252 85978
rect 26956 85924 27012 85926
rect 27036 85924 27092 85926
rect 27116 85924 27172 85926
rect 27196 85924 27252 85926
rect 27616 86522 27672 86524
rect 27696 86522 27752 86524
rect 27776 86522 27832 86524
rect 27856 86522 27912 86524
rect 27616 86470 27662 86522
rect 27662 86470 27672 86522
rect 27696 86470 27726 86522
rect 27726 86470 27738 86522
rect 27738 86470 27752 86522
rect 27776 86470 27790 86522
rect 27790 86470 27802 86522
rect 27802 86470 27832 86522
rect 27856 86470 27866 86522
rect 27866 86470 27912 86522
rect 27616 86468 27672 86470
rect 27696 86468 27752 86470
rect 27776 86468 27832 86470
rect 27856 86468 27912 86470
rect 29216 86522 29272 86524
rect 29296 86522 29352 86524
rect 29376 86522 29432 86524
rect 29456 86522 29512 86524
rect 29216 86470 29262 86522
rect 29262 86470 29272 86522
rect 29296 86470 29326 86522
rect 29326 86470 29338 86522
rect 29338 86470 29352 86522
rect 29376 86470 29390 86522
rect 29390 86470 29402 86522
rect 29402 86470 29432 86522
rect 29456 86470 29466 86522
rect 29466 86470 29512 86522
rect 29216 86468 29272 86470
rect 29296 86468 29352 86470
rect 29376 86468 29432 86470
rect 29456 86468 29512 86470
rect 28556 85978 28612 85980
rect 28636 85978 28692 85980
rect 28716 85978 28772 85980
rect 28796 85978 28852 85980
rect 28556 85926 28602 85978
rect 28602 85926 28612 85978
rect 28636 85926 28666 85978
rect 28666 85926 28678 85978
rect 28678 85926 28692 85978
rect 28716 85926 28730 85978
rect 28730 85926 28742 85978
rect 28742 85926 28772 85978
rect 28796 85926 28806 85978
rect 28806 85926 28852 85978
rect 28556 85924 28612 85926
rect 28636 85924 28692 85926
rect 28716 85924 28772 85926
rect 28796 85924 28852 85926
rect 30816 86522 30872 86524
rect 30896 86522 30952 86524
rect 30976 86522 31032 86524
rect 31056 86522 31112 86524
rect 30816 86470 30862 86522
rect 30862 86470 30872 86522
rect 30896 86470 30926 86522
rect 30926 86470 30938 86522
rect 30938 86470 30952 86522
rect 30976 86470 30990 86522
rect 30990 86470 31002 86522
rect 31002 86470 31032 86522
rect 31056 86470 31066 86522
rect 31066 86470 31112 86522
rect 30816 86468 30872 86470
rect 30896 86468 30952 86470
rect 30976 86468 31032 86470
rect 31056 86468 31112 86470
rect 32416 86522 32472 86524
rect 32496 86522 32552 86524
rect 32576 86522 32632 86524
rect 32656 86522 32712 86524
rect 32416 86470 32462 86522
rect 32462 86470 32472 86522
rect 32496 86470 32526 86522
rect 32526 86470 32538 86522
rect 32538 86470 32552 86522
rect 32576 86470 32590 86522
rect 32590 86470 32602 86522
rect 32602 86470 32632 86522
rect 32656 86470 32666 86522
rect 32666 86470 32712 86522
rect 32416 86468 32472 86470
rect 32496 86468 32552 86470
rect 32576 86468 32632 86470
rect 32656 86468 32712 86470
rect 34016 86522 34072 86524
rect 34096 86522 34152 86524
rect 34176 86522 34232 86524
rect 34256 86522 34312 86524
rect 34016 86470 34062 86522
rect 34062 86470 34072 86522
rect 34096 86470 34126 86522
rect 34126 86470 34138 86522
rect 34138 86470 34152 86522
rect 34176 86470 34190 86522
rect 34190 86470 34202 86522
rect 34202 86470 34232 86522
rect 34256 86470 34266 86522
rect 34266 86470 34312 86522
rect 34016 86468 34072 86470
rect 34096 86468 34152 86470
rect 34176 86468 34232 86470
rect 34256 86468 34312 86470
rect 30156 85978 30212 85980
rect 30236 85978 30292 85980
rect 30316 85978 30372 85980
rect 30396 85978 30452 85980
rect 30156 85926 30202 85978
rect 30202 85926 30212 85978
rect 30236 85926 30266 85978
rect 30266 85926 30278 85978
rect 30278 85926 30292 85978
rect 30316 85926 30330 85978
rect 30330 85926 30342 85978
rect 30342 85926 30372 85978
rect 30396 85926 30406 85978
rect 30406 85926 30452 85978
rect 30156 85924 30212 85926
rect 30236 85924 30292 85926
rect 30316 85924 30372 85926
rect 30396 85924 30452 85926
rect 31756 85978 31812 85980
rect 31836 85978 31892 85980
rect 31916 85978 31972 85980
rect 31996 85978 32052 85980
rect 31756 85926 31802 85978
rect 31802 85926 31812 85978
rect 31836 85926 31866 85978
rect 31866 85926 31878 85978
rect 31878 85926 31892 85978
rect 31916 85926 31930 85978
rect 31930 85926 31942 85978
rect 31942 85926 31972 85978
rect 31996 85926 32006 85978
rect 32006 85926 32052 85978
rect 31756 85924 31812 85926
rect 31836 85924 31892 85926
rect 31916 85924 31972 85926
rect 31996 85924 32052 85926
rect 33356 85978 33412 85980
rect 33436 85978 33492 85980
rect 33516 85978 33572 85980
rect 33596 85978 33652 85980
rect 33356 85926 33402 85978
rect 33402 85926 33412 85978
rect 33436 85926 33466 85978
rect 33466 85926 33478 85978
rect 33478 85926 33492 85978
rect 33516 85926 33530 85978
rect 33530 85926 33542 85978
rect 33542 85926 33572 85978
rect 33596 85926 33606 85978
rect 33606 85926 33652 85978
rect 33356 85924 33412 85926
rect 33436 85924 33492 85926
rect 33516 85924 33572 85926
rect 33596 85924 33652 85926
rect 35616 86522 35672 86524
rect 35696 86522 35752 86524
rect 35776 86522 35832 86524
rect 35856 86522 35912 86524
rect 35616 86470 35662 86522
rect 35662 86470 35672 86522
rect 35696 86470 35726 86522
rect 35726 86470 35738 86522
rect 35738 86470 35752 86522
rect 35776 86470 35790 86522
rect 35790 86470 35802 86522
rect 35802 86470 35832 86522
rect 35856 86470 35866 86522
rect 35866 86470 35912 86522
rect 35616 86468 35672 86470
rect 35696 86468 35752 86470
rect 35776 86468 35832 86470
rect 35856 86468 35912 86470
rect 37216 86522 37272 86524
rect 37296 86522 37352 86524
rect 37376 86522 37432 86524
rect 37456 86522 37512 86524
rect 37216 86470 37262 86522
rect 37262 86470 37272 86522
rect 37296 86470 37326 86522
rect 37326 86470 37338 86522
rect 37338 86470 37352 86522
rect 37376 86470 37390 86522
rect 37390 86470 37402 86522
rect 37402 86470 37432 86522
rect 37456 86470 37466 86522
rect 37466 86470 37512 86522
rect 37216 86468 37272 86470
rect 37296 86468 37352 86470
rect 37376 86468 37432 86470
rect 37456 86468 37512 86470
rect 34956 85978 35012 85980
rect 35036 85978 35092 85980
rect 35116 85978 35172 85980
rect 35196 85978 35252 85980
rect 34956 85926 35002 85978
rect 35002 85926 35012 85978
rect 35036 85926 35066 85978
rect 35066 85926 35078 85978
rect 35078 85926 35092 85978
rect 35116 85926 35130 85978
rect 35130 85926 35142 85978
rect 35142 85926 35172 85978
rect 35196 85926 35206 85978
rect 35206 85926 35252 85978
rect 34956 85924 35012 85926
rect 35036 85924 35092 85926
rect 35116 85924 35172 85926
rect 35196 85924 35252 85926
rect 36556 85978 36612 85980
rect 36636 85978 36692 85980
rect 36716 85978 36772 85980
rect 36796 85978 36852 85980
rect 36556 85926 36602 85978
rect 36602 85926 36612 85978
rect 36636 85926 36666 85978
rect 36666 85926 36678 85978
rect 36678 85926 36692 85978
rect 36716 85926 36730 85978
rect 36730 85926 36742 85978
rect 36742 85926 36772 85978
rect 36796 85926 36806 85978
rect 36806 85926 36852 85978
rect 36556 85924 36612 85926
rect 36636 85924 36692 85926
rect 36716 85924 36772 85926
rect 36796 85924 36852 85926
rect 38816 86522 38872 86524
rect 38896 86522 38952 86524
rect 38976 86522 39032 86524
rect 39056 86522 39112 86524
rect 38816 86470 38862 86522
rect 38862 86470 38872 86522
rect 38896 86470 38926 86522
rect 38926 86470 38938 86522
rect 38938 86470 38952 86522
rect 38976 86470 38990 86522
rect 38990 86470 39002 86522
rect 39002 86470 39032 86522
rect 39056 86470 39066 86522
rect 39066 86470 39112 86522
rect 38816 86468 38872 86470
rect 38896 86468 38952 86470
rect 38976 86468 39032 86470
rect 39056 86468 39112 86470
rect 40416 86522 40472 86524
rect 40496 86522 40552 86524
rect 40576 86522 40632 86524
rect 40656 86522 40712 86524
rect 40416 86470 40462 86522
rect 40462 86470 40472 86522
rect 40496 86470 40526 86522
rect 40526 86470 40538 86522
rect 40538 86470 40552 86522
rect 40576 86470 40590 86522
rect 40590 86470 40602 86522
rect 40602 86470 40632 86522
rect 40656 86470 40666 86522
rect 40666 86470 40712 86522
rect 40416 86468 40472 86470
rect 40496 86468 40552 86470
rect 40576 86468 40632 86470
rect 40656 86468 40712 86470
rect 38842 86148 38898 86184
rect 38842 86128 38844 86148
rect 38844 86128 38896 86148
rect 38896 86128 38898 86148
rect 38156 85978 38212 85980
rect 38236 85978 38292 85980
rect 38316 85978 38372 85980
rect 38396 85978 38452 85980
rect 38156 85926 38202 85978
rect 38202 85926 38212 85978
rect 38236 85926 38266 85978
rect 38266 85926 38278 85978
rect 38278 85926 38292 85978
rect 38316 85926 38330 85978
rect 38330 85926 38342 85978
rect 38342 85926 38372 85978
rect 38396 85926 38406 85978
rect 38406 85926 38452 85978
rect 38156 85924 38212 85926
rect 38236 85924 38292 85926
rect 38316 85924 38372 85926
rect 38396 85924 38452 85926
rect 39756 85978 39812 85980
rect 39836 85978 39892 85980
rect 39916 85978 39972 85980
rect 39996 85978 40052 85980
rect 39756 85926 39802 85978
rect 39802 85926 39812 85978
rect 39836 85926 39866 85978
rect 39866 85926 39878 85978
rect 39878 85926 39892 85978
rect 39916 85926 39930 85978
rect 39930 85926 39942 85978
rect 39942 85926 39972 85978
rect 39996 85926 40006 85978
rect 40006 85926 40052 85978
rect 39756 85924 39812 85926
rect 39836 85924 39892 85926
rect 39916 85924 39972 85926
rect 39996 85924 40052 85926
rect 41356 85978 41412 85980
rect 41436 85978 41492 85980
rect 41516 85978 41572 85980
rect 41596 85978 41652 85980
rect 41356 85926 41402 85978
rect 41402 85926 41412 85978
rect 41436 85926 41466 85978
rect 41466 85926 41478 85978
rect 41478 85926 41492 85978
rect 41516 85926 41530 85978
rect 41530 85926 41542 85978
rect 41542 85926 41572 85978
rect 41596 85926 41606 85978
rect 41606 85926 41652 85978
rect 41356 85924 41412 85926
rect 41436 85924 41492 85926
rect 41516 85924 41572 85926
rect 41596 85924 41652 85926
rect 40038 85584 40094 85640
rect 42016 86522 42072 86524
rect 42096 86522 42152 86524
rect 42176 86522 42232 86524
rect 42256 86522 42312 86524
rect 42016 86470 42062 86522
rect 42062 86470 42072 86522
rect 42096 86470 42126 86522
rect 42126 86470 42138 86522
rect 42138 86470 42152 86522
rect 42176 86470 42190 86522
rect 42190 86470 42202 86522
rect 42202 86470 42232 86522
rect 42256 86470 42266 86522
rect 42266 86470 42312 86522
rect 42016 86468 42072 86470
rect 42096 86468 42152 86470
rect 42176 86468 42232 86470
rect 42256 86468 42312 86470
rect 43616 86522 43672 86524
rect 43696 86522 43752 86524
rect 43776 86522 43832 86524
rect 43856 86522 43912 86524
rect 43616 86470 43662 86522
rect 43662 86470 43672 86522
rect 43696 86470 43726 86522
rect 43726 86470 43738 86522
rect 43738 86470 43752 86522
rect 43776 86470 43790 86522
rect 43790 86470 43802 86522
rect 43802 86470 43832 86522
rect 43856 86470 43866 86522
rect 43866 86470 43912 86522
rect 43616 86468 43672 86470
rect 43696 86468 43752 86470
rect 43776 86468 43832 86470
rect 43856 86468 43912 86470
rect 42956 85978 43012 85980
rect 43036 85978 43092 85980
rect 43116 85978 43172 85980
rect 43196 85978 43252 85980
rect 42956 85926 43002 85978
rect 43002 85926 43012 85978
rect 43036 85926 43066 85978
rect 43066 85926 43078 85978
rect 43078 85926 43092 85978
rect 43116 85926 43130 85978
rect 43130 85926 43142 85978
rect 43142 85926 43172 85978
rect 43196 85926 43206 85978
rect 43206 85926 43252 85978
rect 42956 85924 43012 85926
rect 43036 85924 43092 85926
rect 43116 85924 43172 85926
rect 43196 85924 43252 85926
rect 44556 85978 44612 85980
rect 44636 85978 44692 85980
rect 44716 85978 44772 85980
rect 44796 85978 44852 85980
rect 44556 85926 44602 85978
rect 44602 85926 44612 85978
rect 44636 85926 44666 85978
rect 44666 85926 44678 85978
rect 44678 85926 44692 85978
rect 44716 85926 44730 85978
rect 44730 85926 44742 85978
rect 44742 85926 44772 85978
rect 44796 85926 44806 85978
rect 44806 85926 44852 85978
rect 44556 85924 44612 85926
rect 44636 85924 44692 85926
rect 44716 85924 44772 85926
rect 44796 85924 44852 85926
rect 41786 85584 41842 85640
rect 42798 85604 42854 85640
rect 42798 85584 42800 85604
rect 42800 85584 42852 85604
rect 42852 85584 42854 85604
rect 42522 84360 42578 84416
rect 44730 84360 44786 84416
rect 45216 86522 45272 86524
rect 45296 86522 45352 86524
rect 45376 86522 45432 86524
rect 45456 86522 45512 86524
rect 45216 86470 45262 86522
rect 45262 86470 45272 86522
rect 45296 86470 45326 86522
rect 45326 86470 45338 86522
rect 45338 86470 45352 86522
rect 45376 86470 45390 86522
rect 45390 86470 45402 86522
rect 45402 86470 45432 86522
rect 45456 86470 45466 86522
rect 45466 86470 45512 86522
rect 45216 86468 45272 86470
rect 45296 86468 45352 86470
rect 45376 86468 45432 86470
rect 45456 86468 45512 86470
rect 46816 86522 46872 86524
rect 46896 86522 46952 86524
rect 46976 86522 47032 86524
rect 47056 86522 47112 86524
rect 46816 86470 46862 86522
rect 46862 86470 46872 86522
rect 46896 86470 46926 86522
rect 46926 86470 46938 86522
rect 46938 86470 46952 86522
rect 46976 86470 46990 86522
rect 46990 86470 47002 86522
rect 47002 86470 47032 86522
rect 47056 86470 47066 86522
rect 47066 86470 47112 86522
rect 46816 86468 46872 86470
rect 46896 86468 46952 86470
rect 46976 86468 47032 86470
rect 47056 86468 47112 86470
rect 46156 85978 46212 85980
rect 46236 85978 46292 85980
rect 46316 85978 46372 85980
rect 46396 85978 46452 85980
rect 46156 85926 46202 85978
rect 46202 85926 46212 85978
rect 46236 85926 46266 85978
rect 46266 85926 46278 85978
rect 46278 85926 46292 85978
rect 46316 85926 46330 85978
rect 46330 85926 46342 85978
rect 46342 85926 46372 85978
rect 46396 85926 46406 85978
rect 46406 85926 46452 85978
rect 46156 85924 46212 85926
rect 46236 85924 46292 85926
rect 46316 85924 46372 85926
rect 46396 85924 46452 85926
rect 48416 86522 48472 86524
rect 48496 86522 48552 86524
rect 48576 86522 48632 86524
rect 48656 86522 48712 86524
rect 48416 86470 48462 86522
rect 48462 86470 48472 86522
rect 48496 86470 48526 86522
rect 48526 86470 48538 86522
rect 48538 86470 48552 86522
rect 48576 86470 48590 86522
rect 48590 86470 48602 86522
rect 48602 86470 48632 86522
rect 48656 86470 48666 86522
rect 48666 86470 48712 86522
rect 48416 86468 48472 86470
rect 48496 86468 48552 86470
rect 48576 86468 48632 86470
rect 48656 86468 48712 86470
rect 50016 86522 50072 86524
rect 50096 86522 50152 86524
rect 50176 86522 50232 86524
rect 50256 86522 50312 86524
rect 50016 86470 50062 86522
rect 50062 86470 50072 86522
rect 50096 86470 50126 86522
rect 50126 86470 50138 86522
rect 50138 86470 50152 86522
rect 50176 86470 50190 86522
rect 50190 86470 50202 86522
rect 50202 86470 50232 86522
rect 50256 86470 50266 86522
rect 50266 86470 50312 86522
rect 50016 86468 50072 86470
rect 50096 86468 50152 86470
rect 50176 86468 50232 86470
rect 50256 86468 50312 86470
rect 51616 86522 51672 86524
rect 51696 86522 51752 86524
rect 51776 86522 51832 86524
rect 51856 86522 51912 86524
rect 51616 86470 51662 86522
rect 51662 86470 51672 86522
rect 51696 86470 51726 86522
rect 51726 86470 51738 86522
rect 51738 86470 51752 86522
rect 51776 86470 51790 86522
rect 51790 86470 51802 86522
rect 51802 86470 51832 86522
rect 51856 86470 51866 86522
rect 51866 86470 51912 86522
rect 51616 86468 51672 86470
rect 51696 86468 51752 86470
rect 51776 86468 51832 86470
rect 51856 86468 51912 86470
rect 53216 86522 53272 86524
rect 53296 86522 53352 86524
rect 53376 86522 53432 86524
rect 53456 86522 53512 86524
rect 53216 86470 53262 86522
rect 53262 86470 53272 86522
rect 53296 86470 53326 86522
rect 53326 86470 53338 86522
rect 53338 86470 53352 86522
rect 53376 86470 53390 86522
rect 53390 86470 53402 86522
rect 53402 86470 53432 86522
rect 53456 86470 53466 86522
rect 53466 86470 53512 86522
rect 53216 86468 53272 86470
rect 53296 86468 53352 86470
rect 53376 86468 53432 86470
rect 53456 86468 53512 86470
rect 48870 86148 48926 86184
rect 48870 86128 48872 86148
rect 48872 86128 48924 86148
rect 48924 86128 48926 86148
rect 47756 85978 47812 85980
rect 47836 85978 47892 85980
rect 47916 85978 47972 85980
rect 47996 85978 48052 85980
rect 47756 85926 47802 85978
rect 47802 85926 47812 85978
rect 47836 85926 47866 85978
rect 47866 85926 47878 85978
rect 47878 85926 47892 85978
rect 47916 85926 47930 85978
rect 47930 85926 47942 85978
rect 47942 85926 47972 85978
rect 47996 85926 48006 85978
rect 48006 85926 48052 85978
rect 47756 85924 47812 85926
rect 47836 85924 47892 85926
rect 47916 85924 47972 85926
rect 47996 85924 48052 85926
rect 49356 85978 49412 85980
rect 49436 85978 49492 85980
rect 49516 85978 49572 85980
rect 49596 85978 49652 85980
rect 49356 85926 49402 85978
rect 49402 85926 49412 85978
rect 49436 85926 49466 85978
rect 49466 85926 49478 85978
rect 49478 85926 49492 85978
rect 49516 85926 49530 85978
rect 49530 85926 49542 85978
rect 49542 85926 49572 85978
rect 49596 85926 49606 85978
rect 49606 85926 49652 85978
rect 49356 85924 49412 85926
rect 49436 85924 49492 85926
rect 49516 85924 49572 85926
rect 49596 85924 49652 85926
rect 54816 86522 54872 86524
rect 54896 86522 54952 86524
rect 54976 86522 55032 86524
rect 55056 86522 55112 86524
rect 54816 86470 54862 86522
rect 54862 86470 54872 86522
rect 54896 86470 54926 86522
rect 54926 86470 54938 86522
rect 54938 86470 54952 86522
rect 54976 86470 54990 86522
rect 54990 86470 55002 86522
rect 55002 86470 55032 86522
rect 55056 86470 55066 86522
rect 55066 86470 55112 86522
rect 54816 86468 54872 86470
rect 54896 86468 54952 86470
rect 54976 86468 55032 86470
rect 55056 86468 55112 86470
rect 56416 86522 56472 86524
rect 56496 86522 56552 86524
rect 56576 86522 56632 86524
rect 56656 86522 56712 86524
rect 56416 86470 56462 86522
rect 56462 86470 56472 86522
rect 56496 86470 56526 86522
rect 56526 86470 56538 86522
rect 56538 86470 56552 86522
rect 56576 86470 56590 86522
rect 56590 86470 56602 86522
rect 56602 86470 56632 86522
rect 56656 86470 56666 86522
rect 56666 86470 56712 86522
rect 56416 86468 56472 86470
rect 56496 86468 56552 86470
rect 56576 86468 56632 86470
rect 56656 86468 56712 86470
rect 58016 86522 58072 86524
rect 58096 86522 58152 86524
rect 58176 86522 58232 86524
rect 58256 86522 58312 86524
rect 58016 86470 58062 86522
rect 58062 86470 58072 86522
rect 58096 86470 58126 86522
rect 58126 86470 58138 86522
rect 58138 86470 58152 86522
rect 58176 86470 58190 86522
rect 58190 86470 58202 86522
rect 58202 86470 58232 86522
rect 58256 86470 58266 86522
rect 58266 86470 58312 86522
rect 58016 86468 58072 86470
rect 58096 86468 58152 86470
rect 58176 86468 58232 86470
rect 58256 86468 58312 86470
rect 59616 86522 59672 86524
rect 59696 86522 59752 86524
rect 59776 86522 59832 86524
rect 59856 86522 59912 86524
rect 59616 86470 59662 86522
rect 59662 86470 59672 86522
rect 59696 86470 59726 86522
rect 59726 86470 59738 86522
rect 59738 86470 59752 86522
rect 59776 86470 59790 86522
rect 59790 86470 59802 86522
rect 59802 86470 59832 86522
rect 59856 86470 59866 86522
rect 59866 86470 59912 86522
rect 59616 86468 59672 86470
rect 59696 86468 59752 86470
rect 59776 86468 59832 86470
rect 59856 86468 59912 86470
rect 55310 86164 55312 86184
rect 55312 86164 55364 86184
rect 55364 86164 55366 86184
rect 55310 86128 55366 86164
rect 50956 85978 51012 85980
rect 51036 85978 51092 85980
rect 51116 85978 51172 85980
rect 51196 85978 51252 85980
rect 50956 85926 51002 85978
rect 51002 85926 51012 85978
rect 51036 85926 51066 85978
rect 51066 85926 51078 85978
rect 51078 85926 51092 85978
rect 51116 85926 51130 85978
rect 51130 85926 51142 85978
rect 51142 85926 51172 85978
rect 51196 85926 51206 85978
rect 51206 85926 51252 85978
rect 50956 85924 51012 85926
rect 51036 85924 51092 85926
rect 51116 85924 51172 85926
rect 51196 85924 51252 85926
rect 52556 85978 52612 85980
rect 52636 85978 52692 85980
rect 52716 85978 52772 85980
rect 52796 85978 52852 85980
rect 52556 85926 52602 85978
rect 52602 85926 52612 85978
rect 52636 85926 52666 85978
rect 52666 85926 52678 85978
rect 52678 85926 52692 85978
rect 52716 85926 52730 85978
rect 52730 85926 52742 85978
rect 52742 85926 52772 85978
rect 52796 85926 52806 85978
rect 52806 85926 52852 85978
rect 52556 85924 52612 85926
rect 52636 85924 52692 85926
rect 52716 85924 52772 85926
rect 52796 85924 52852 85926
rect 46570 85584 46626 85640
rect 47306 85584 47362 85640
rect 49238 85584 49294 85640
rect 50802 85584 50858 85640
rect 54156 85978 54212 85980
rect 54236 85978 54292 85980
rect 54316 85978 54372 85980
rect 54396 85978 54452 85980
rect 54156 85926 54202 85978
rect 54202 85926 54212 85978
rect 54236 85926 54266 85978
rect 54266 85926 54278 85978
rect 54278 85926 54292 85978
rect 54316 85926 54330 85978
rect 54330 85926 54342 85978
rect 54342 85926 54372 85978
rect 54396 85926 54406 85978
rect 54406 85926 54452 85978
rect 54156 85924 54212 85926
rect 54236 85924 54292 85926
rect 54316 85924 54372 85926
rect 54396 85924 54452 85926
rect 55756 85978 55812 85980
rect 55836 85978 55892 85980
rect 55916 85978 55972 85980
rect 55996 85978 56052 85980
rect 55756 85926 55802 85978
rect 55802 85926 55812 85978
rect 55836 85926 55866 85978
rect 55866 85926 55878 85978
rect 55878 85926 55892 85978
rect 55916 85926 55930 85978
rect 55930 85926 55942 85978
rect 55942 85926 55972 85978
rect 55996 85926 56006 85978
rect 56006 85926 56052 85978
rect 55756 85924 55812 85926
rect 55836 85924 55892 85926
rect 55916 85924 55972 85926
rect 55996 85924 56052 85926
rect 57356 85978 57412 85980
rect 57436 85978 57492 85980
rect 57516 85978 57572 85980
rect 57596 85978 57652 85980
rect 57356 85926 57402 85978
rect 57402 85926 57412 85978
rect 57436 85926 57466 85978
rect 57466 85926 57478 85978
rect 57478 85926 57492 85978
rect 57516 85926 57530 85978
rect 57530 85926 57542 85978
rect 57542 85926 57572 85978
rect 57596 85926 57606 85978
rect 57606 85926 57652 85978
rect 57356 85924 57412 85926
rect 57436 85924 57492 85926
rect 57516 85924 57572 85926
rect 57596 85924 57652 85926
rect 58956 85978 59012 85980
rect 59036 85978 59092 85980
rect 59116 85978 59172 85980
rect 59196 85978 59252 85980
rect 58956 85926 59002 85978
rect 59002 85926 59012 85978
rect 59036 85926 59066 85978
rect 59066 85926 59078 85978
rect 59078 85926 59092 85978
rect 59116 85926 59130 85978
rect 59130 85926 59142 85978
rect 59142 85926 59172 85978
rect 59196 85926 59206 85978
rect 59206 85926 59252 85978
rect 58956 85924 59012 85926
rect 59036 85924 59092 85926
rect 59116 85924 59172 85926
rect 59196 85924 59252 85926
rect 60556 85978 60612 85980
rect 60636 85978 60692 85980
rect 60716 85978 60772 85980
rect 60796 85978 60852 85980
rect 60556 85926 60602 85978
rect 60602 85926 60612 85978
rect 60636 85926 60666 85978
rect 60666 85926 60678 85978
rect 60678 85926 60692 85978
rect 60716 85926 60730 85978
rect 60730 85926 60742 85978
rect 60742 85926 60772 85978
rect 60796 85926 60806 85978
rect 60806 85926 60852 85978
rect 60556 85924 60612 85926
rect 60636 85924 60692 85926
rect 60716 85924 60772 85926
rect 60796 85924 60852 85926
rect 61216 86522 61272 86524
rect 61296 86522 61352 86524
rect 61376 86522 61432 86524
rect 61456 86522 61512 86524
rect 61216 86470 61262 86522
rect 61262 86470 61272 86522
rect 61296 86470 61326 86522
rect 61326 86470 61338 86522
rect 61338 86470 61352 86522
rect 61376 86470 61390 86522
rect 61390 86470 61402 86522
rect 61402 86470 61432 86522
rect 61456 86470 61466 86522
rect 61466 86470 61512 86522
rect 61216 86468 61272 86470
rect 61296 86468 61352 86470
rect 61376 86468 61432 86470
rect 61456 86468 61512 86470
rect 62156 85978 62212 85980
rect 62236 85978 62292 85980
rect 62316 85978 62372 85980
rect 62396 85978 62452 85980
rect 62156 85926 62202 85978
rect 62202 85926 62212 85978
rect 62236 85926 62266 85978
rect 62266 85926 62278 85978
rect 62278 85926 62292 85978
rect 62316 85926 62330 85978
rect 62330 85926 62342 85978
rect 62342 85926 62372 85978
rect 62396 85926 62406 85978
rect 62406 85926 62452 85978
rect 62156 85924 62212 85926
rect 62236 85924 62292 85926
rect 62316 85924 62372 85926
rect 62396 85924 62452 85926
rect 61014 85856 61070 85912
rect 62816 86522 62872 86524
rect 62896 86522 62952 86524
rect 62976 86522 63032 86524
rect 63056 86522 63112 86524
rect 62816 86470 62862 86522
rect 62862 86470 62872 86522
rect 62896 86470 62926 86522
rect 62926 86470 62938 86522
rect 62938 86470 62952 86522
rect 62976 86470 62990 86522
rect 62990 86470 63002 86522
rect 63002 86470 63032 86522
rect 63056 86470 63066 86522
rect 63066 86470 63112 86522
rect 62816 86468 62872 86470
rect 62896 86468 62952 86470
rect 62976 86468 63032 86470
rect 63056 86468 63112 86470
rect 64416 86522 64472 86524
rect 64496 86522 64552 86524
rect 64576 86522 64632 86524
rect 64656 86522 64712 86524
rect 64416 86470 64462 86522
rect 64462 86470 64472 86522
rect 64496 86470 64526 86522
rect 64526 86470 64538 86522
rect 64538 86470 64552 86522
rect 64576 86470 64590 86522
rect 64590 86470 64602 86522
rect 64602 86470 64632 86522
rect 64656 86470 64666 86522
rect 64666 86470 64712 86522
rect 64416 86468 64472 86470
rect 64496 86468 64552 86470
rect 64576 86468 64632 86470
rect 64656 86468 64712 86470
rect 66016 86522 66072 86524
rect 66096 86522 66152 86524
rect 66176 86522 66232 86524
rect 66256 86522 66312 86524
rect 66016 86470 66062 86522
rect 66062 86470 66072 86522
rect 66096 86470 66126 86522
rect 66126 86470 66138 86522
rect 66138 86470 66152 86522
rect 66176 86470 66190 86522
rect 66190 86470 66202 86522
rect 66202 86470 66232 86522
rect 66256 86470 66266 86522
rect 66266 86470 66312 86522
rect 66016 86468 66072 86470
rect 66096 86468 66152 86470
rect 66176 86468 66232 86470
rect 66256 86468 66312 86470
rect 67616 86522 67672 86524
rect 67696 86522 67752 86524
rect 67776 86522 67832 86524
rect 67856 86522 67912 86524
rect 67616 86470 67662 86522
rect 67662 86470 67672 86522
rect 67696 86470 67726 86522
rect 67726 86470 67738 86522
rect 67738 86470 67752 86522
rect 67776 86470 67790 86522
rect 67790 86470 67802 86522
rect 67802 86470 67832 86522
rect 67856 86470 67866 86522
rect 67866 86470 67912 86522
rect 67616 86468 67672 86470
rect 67696 86468 67752 86470
rect 67776 86468 67832 86470
rect 67856 86468 67912 86470
rect 63756 85978 63812 85980
rect 63836 85978 63892 85980
rect 63916 85978 63972 85980
rect 63996 85978 64052 85980
rect 63756 85926 63802 85978
rect 63802 85926 63812 85978
rect 63836 85926 63866 85978
rect 63866 85926 63878 85978
rect 63878 85926 63892 85978
rect 63916 85926 63930 85978
rect 63930 85926 63942 85978
rect 63942 85926 63972 85978
rect 63996 85926 64006 85978
rect 64006 85926 64052 85978
rect 63756 85924 63812 85926
rect 63836 85924 63892 85926
rect 63916 85924 63972 85926
rect 63996 85924 64052 85926
rect 65356 85978 65412 85980
rect 65436 85978 65492 85980
rect 65516 85978 65572 85980
rect 65596 85978 65652 85980
rect 65356 85926 65402 85978
rect 65402 85926 65412 85978
rect 65436 85926 65466 85978
rect 65466 85926 65478 85978
rect 65478 85926 65492 85978
rect 65516 85926 65530 85978
rect 65530 85926 65542 85978
rect 65542 85926 65572 85978
rect 65596 85926 65606 85978
rect 65606 85926 65652 85978
rect 65356 85924 65412 85926
rect 65436 85924 65492 85926
rect 65516 85924 65572 85926
rect 65596 85924 65652 85926
rect 66956 85978 67012 85980
rect 67036 85978 67092 85980
rect 67116 85978 67172 85980
rect 67196 85978 67252 85980
rect 66956 85926 67002 85978
rect 67002 85926 67012 85978
rect 67036 85926 67066 85978
rect 67066 85926 67078 85978
rect 67078 85926 67092 85978
rect 67116 85926 67130 85978
rect 67130 85926 67142 85978
rect 67142 85926 67172 85978
rect 67196 85926 67206 85978
rect 67206 85926 67252 85978
rect 66956 85924 67012 85926
rect 67036 85924 67092 85926
rect 67116 85924 67172 85926
rect 67196 85924 67252 85926
rect 63498 85856 63554 85912
rect 69216 86522 69272 86524
rect 69296 86522 69352 86524
rect 69376 86522 69432 86524
rect 69456 86522 69512 86524
rect 69216 86470 69262 86522
rect 69262 86470 69272 86522
rect 69296 86470 69326 86522
rect 69326 86470 69338 86522
rect 69338 86470 69352 86522
rect 69376 86470 69390 86522
rect 69390 86470 69402 86522
rect 69402 86470 69432 86522
rect 69456 86470 69466 86522
rect 69466 86470 69512 86522
rect 69216 86468 69272 86470
rect 69296 86468 69352 86470
rect 69376 86468 69432 86470
rect 69456 86468 69512 86470
rect 70816 86522 70872 86524
rect 70896 86522 70952 86524
rect 70976 86522 71032 86524
rect 71056 86522 71112 86524
rect 70816 86470 70862 86522
rect 70862 86470 70872 86522
rect 70896 86470 70926 86522
rect 70926 86470 70938 86522
rect 70938 86470 70952 86522
rect 70976 86470 70990 86522
rect 70990 86470 71002 86522
rect 71002 86470 71032 86522
rect 71056 86470 71066 86522
rect 71066 86470 71112 86522
rect 70816 86468 70872 86470
rect 70896 86468 70952 86470
rect 70976 86468 71032 86470
rect 71056 86468 71112 86470
rect 68556 85978 68612 85980
rect 68636 85978 68692 85980
rect 68716 85978 68772 85980
rect 68796 85978 68852 85980
rect 68556 85926 68602 85978
rect 68602 85926 68612 85978
rect 68636 85926 68666 85978
rect 68666 85926 68678 85978
rect 68678 85926 68692 85978
rect 68716 85926 68730 85978
rect 68730 85926 68742 85978
rect 68742 85926 68772 85978
rect 68796 85926 68806 85978
rect 68806 85926 68852 85978
rect 68556 85924 68612 85926
rect 68636 85924 68692 85926
rect 68716 85924 68772 85926
rect 68796 85924 68852 85926
rect 70156 85978 70212 85980
rect 70236 85978 70292 85980
rect 70316 85978 70372 85980
rect 70396 85978 70452 85980
rect 70156 85926 70202 85978
rect 70202 85926 70212 85978
rect 70236 85926 70266 85978
rect 70266 85926 70278 85978
rect 70278 85926 70292 85978
rect 70316 85926 70330 85978
rect 70330 85926 70342 85978
rect 70342 85926 70372 85978
rect 70396 85926 70406 85978
rect 70406 85926 70452 85978
rect 70156 85924 70212 85926
rect 70236 85924 70292 85926
rect 70316 85924 70372 85926
rect 70396 85924 70452 85926
rect 71756 85978 71812 85980
rect 71836 85978 71892 85980
rect 71916 85978 71972 85980
rect 71996 85978 72052 85980
rect 71756 85926 71802 85978
rect 71802 85926 71812 85978
rect 71836 85926 71866 85978
rect 71866 85926 71878 85978
rect 71878 85926 71892 85978
rect 71916 85926 71930 85978
rect 71930 85926 71942 85978
rect 71942 85926 71972 85978
rect 71996 85926 72006 85978
rect 72006 85926 72052 85978
rect 71756 85924 71812 85926
rect 71836 85924 71892 85926
rect 71916 85924 71972 85926
rect 71996 85924 72052 85926
rect 72416 86522 72472 86524
rect 72496 86522 72552 86524
rect 72576 86522 72632 86524
rect 72656 86522 72712 86524
rect 72416 86470 72462 86522
rect 72462 86470 72472 86522
rect 72496 86470 72526 86522
rect 72526 86470 72538 86522
rect 72538 86470 72552 86522
rect 72576 86470 72590 86522
rect 72590 86470 72602 86522
rect 72602 86470 72632 86522
rect 72656 86470 72666 86522
rect 72666 86470 72712 86522
rect 72416 86468 72472 86470
rect 72496 86468 72552 86470
rect 72576 86468 72632 86470
rect 72656 86468 72712 86470
rect 74016 86522 74072 86524
rect 74096 86522 74152 86524
rect 74176 86522 74232 86524
rect 74256 86522 74312 86524
rect 74016 86470 74062 86522
rect 74062 86470 74072 86522
rect 74096 86470 74126 86522
rect 74126 86470 74138 86522
rect 74138 86470 74152 86522
rect 74176 86470 74190 86522
rect 74190 86470 74202 86522
rect 74202 86470 74232 86522
rect 74256 86470 74266 86522
rect 74266 86470 74312 86522
rect 74016 86468 74072 86470
rect 74096 86468 74152 86470
rect 74176 86468 74232 86470
rect 74256 86468 74312 86470
rect 75616 86522 75672 86524
rect 75696 86522 75752 86524
rect 75776 86522 75832 86524
rect 75856 86522 75912 86524
rect 75616 86470 75662 86522
rect 75662 86470 75672 86522
rect 75696 86470 75726 86522
rect 75726 86470 75738 86522
rect 75738 86470 75752 86522
rect 75776 86470 75790 86522
rect 75790 86470 75802 86522
rect 75802 86470 75832 86522
rect 75856 86470 75866 86522
rect 75866 86470 75912 86522
rect 75616 86468 75672 86470
rect 75696 86468 75752 86470
rect 75776 86468 75832 86470
rect 75856 86468 75912 86470
rect 77216 86522 77272 86524
rect 77296 86522 77352 86524
rect 77376 86522 77432 86524
rect 77456 86522 77512 86524
rect 77216 86470 77262 86522
rect 77262 86470 77272 86522
rect 77296 86470 77326 86522
rect 77326 86470 77338 86522
rect 77338 86470 77352 86522
rect 77376 86470 77390 86522
rect 77390 86470 77402 86522
rect 77402 86470 77432 86522
rect 77456 86470 77466 86522
rect 77466 86470 77512 86522
rect 77216 86468 77272 86470
rect 77296 86468 77352 86470
rect 77376 86468 77432 86470
rect 77456 86468 77512 86470
rect 73356 85978 73412 85980
rect 73436 85978 73492 85980
rect 73516 85978 73572 85980
rect 73596 85978 73652 85980
rect 73356 85926 73402 85978
rect 73402 85926 73412 85978
rect 73436 85926 73466 85978
rect 73466 85926 73478 85978
rect 73478 85926 73492 85978
rect 73516 85926 73530 85978
rect 73530 85926 73542 85978
rect 73542 85926 73572 85978
rect 73596 85926 73606 85978
rect 73606 85926 73652 85978
rect 73356 85924 73412 85926
rect 73436 85924 73492 85926
rect 73516 85924 73572 85926
rect 73596 85924 73652 85926
rect 68098 85856 68154 85912
rect 72146 85856 72202 85912
rect 68006 85720 68062 85776
rect 74956 85978 75012 85980
rect 75036 85978 75092 85980
rect 75116 85978 75172 85980
rect 75196 85978 75252 85980
rect 74956 85926 75002 85978
rect 75002 85926 75012 85978
rect 75036 85926 75066 85978
rect 75066 85926 75078 85978
rect 75078 85926 75092 85978
rect 75116 85926 75130 85978
rect 75130 85926 75142 85978
rect 75142 85926 75172 85978
rect 75196 85926 75206 85978
rect 75206 85926 75252 85978
rect 74956 85924 75012 85926
rect 75036 85924 75092 85926
rect 75116 85924 75172 85926
rect 75196 85924 75252 85926
rect 76556 85978 76612 85980
rect 76636 85978 76692 85980
rect 76716 85978 76772 85980
rect 76796 85978 76852 85980
rect 76556 85926 76602 85978
rect 76602 85926 76612 85978
rect 76636 85926 76666 85978
rect 76666 85926 76678 85978
rect 76678 85926 76692 85978
rect 76716 85926 76730 85978
rect 76730 85926 76742 85978
rect 76742 85926 76772 85978
rect 76796 85926 76806 85978
rect 76806 85926 76852 85978
rect 76556 85924 76612 85926
rect 76636 85924 76692 85926
rect 76716 85924 76772 85926
rect 76796 85924 76852 85926
rect 78816 86522 78872 86524
rect 78896 86522 78952 86524
rect 78976 86522 79032 86524
rect 79056 86522 79112 86524
rect 78816 86470 78862 86522
rect 78862 86470 78872 86522
rect 78896 86470 78926 86522
rect 78926 86470 78938 86522
rect 78938 86470 78952 86522
rect 78976 86470 78990 86522
rect 78990 86470 79002 86522
rect 79002 86470 79032 86522
rect 79056 86470 79066 86522
rect 79066 86470 79112 86522
rect 78816 86468 78872 86470
rect 78896 86468 78952 86470
rect 78976 86468 79032 86470
rect 79056 86468 79112 86470
rect 80416 86522 80472 86524
rect 80496 86522 80552 86524
rect 80576 86522 80632 86524
rect 80656 86522 80712 86524
rect 80416 86470 80462 86522
rect 80462 86470 80472 86522
rect 80496 86470 80526 86522
rect 80526 86470 80538 86522
rect 80538 86470 80552 86522
rect 80576 86470 80590 86522
rect 80590 86470 80602 86522
rect 80602 86470 80632 86522
rect 80656 86470 80666 86522
rect 80666 86470 80712 86522
rect 80416 86468 80472 86470
rect 80496 86468 80552 86470
rect 80576 86468 80632 86470
rect 80656 86468 80712 86470
rect 82016 86522 82072 86524
rect 82096 86522 82152 86524
rect 82176 86522 82232 86524
rect 82256 86522 82312 86524
rect 82016 86470 82062 86522
rect 82062 86470 82072 86522
rect 82096 86470 82126 86522
rect 82126 86470 82138 86522
rect 82138 86470 82152 86522
rect 82176 86470 82190 86522
rect 82190 86470 82202 86522
rect 82202 86470 82232 86522
rect 82256 86470 82266 86522
rect 82266 86470 82312 86522
rect 82016 86468 82072 86470
rect 82096 86468 82152 86470
rect 82176 86468 82232 86470
rect 82256 86468 82312 86470
rect 83616 86522 83672 86524
rect 83696 86522 83752 86524
rect 83776 86522 83832 86524
rect 83856 86522 83912 86524
rect 83616 86470 83662 86522
rect 83662 86470 83672 86522
rect 83696 86470 83726 86522
rect 83726 86470 83738 86522
rect 83738 86470 83752 86522
rect 83776 86470 83790 86522
rect 83790 86470 83802 86522
rect 83802 86470 83832 86522
rect 83856 86470 83866 86522
rect 83866 86470 83912 86522
rect 83616 86468 83672 86470
rect 83696 86468 83752 86470
rect 83776 86468 83832 86470
rect 83856 86468 83912 86470
rect 85216 86522 85272 86524
rect 85296 86522 85352 86524
rect 85376 86522 85432 86524
rect 85456 86522 85512 86524
rect 85216 86470 85262 86522
rect 85262 86470 85272 86522
rect 85296 86470 85326 86522
rect 85326 86470 85338 86522
rect 85338 86470 85352 86522
rect 85376 86470 85390 86522
rect 85390 86470 85402 86522
rect 85402 86470 85432 86522
rect 85456 86470 85466 86522
rect 85466 86470 85512 86522
rect 85216 86468 85272 86470
rect 85296 86468 85352 86470
rect 85376 86468 85432 86470
rect 85456 86468 85512 86470
rect 86816 86522 86872 86524
rect 86896 86522 86952 86524
rect 86976 86522 87032 86524
rect 87056 86522 87112 86524
rect 86816 86470 86862 86522
rect 86862 86470 86872 86522
rect 86896 86470 86926 86522
rect 86926 86470 86938 86522
rect 86938 86470 86952 86522
rect 86976 86470 86990 86522
rect 86990 86470 87002 86522
rect 87002 86470 87032 86522
rect 87056 86470 87066 86522
rect 87066 86470 87112 86522
rect 86816 86468 86872 86470
rect 86896 86468 86952 86470
rect 86976 86468 87032 86470
rect 87056 86468 87112 86470
rect 88416 86522 88472 86524
rect 88496 86522 88552 86524
rect 88576 86522 88632 86524
rect 88656 86522 88712 86524
rect 88416 86470 88462 86522
rect 88462 86470 88472 86522
rect 88496 86470 88526 86522
rect 88526 86470 88538 86522
rect 88538 86470 88552 86522
rect 88576 86470 88590 86522
rect 88590 86470 88602 86522
rect 88602 86470 88632 86522
rect 88656 86470 88666 86522
rect 88666 86470 88712 86522
rect 88416 86468 88472 86470
rect 88496 86468 88552 86470
rect 88576 86468 88632 86470
rect 88656 86468 88712 86470
rect 90016 86522 90072 86524
rect 90096 86522 90152 86524
rect 90176 86522 90232 86524
rect 90256 86522 90312 86524
rect 90016 86470 90062 86522
rect 90062 86470 90072 86522
rect 90096 86470 90126 86522
rect 90126 86470 90138 86522
rect 90138 86470 90152 86522
rect 90176 86470 90190 86522
rect 90190 86470 90202 86522
rect 90202 86470 90232 86522
rect 90256 86470 90266 86522
rect 90266 86470 90312 86522
rect 90016 86468 90072 86470
rect 90096 86468 90152 86470
rect 90176 86468 90232 86470
rect 90256 86468 90312 86470
rect 78156 85978 78212 85980
rect 78236 85978 78292 85980
rect 78316 85978 78372 85980
rect 78396 85978 78452 85980
rect 78156 85926 78202 85978
rect 78202 85926 78212 85978
rect 78236 85926 78266 85978
rect 78266 85926 78278 85978
rect 78278 85926 78292 85978
rect 78316 85926 78330 85978
rect 78330 85926 78342 85978
rect 78342 85926 78372 85978
rect 78396 85926 78406 85978
rect 78406 85926 78452 85978
rect 78156 85924 78212 85926
rect 78236 85924 78292 85926
rect 78316 85924 78372 85926
rect 78396 85924 78452 85926
rect 79756 85978 79812 85980
rect 79836 85978 79892 85980
rect 79916 85978 79972 85980
rect 79996 85978 80052 85980
rect 79756 85926 79802 85978
rect 79802 85926 79812 85978
rect 79836 85926 79866 85978
rect 79866 85926 79878 85978
rect 79878 85926 79892 85978
rect 79916 85926 79930 85978
rect 79930 85926 79942 85978
rect 79942 85926 79972 85978
rect 79996 85926 80006 85978
rect 80006 85926 80052 85978
rect 79756 85924 79812 85926
rect 79836 85924 79892 85926
rect 79916 85924 79972 85926
rect 79996 85924 80052 85926
rect 81356 85978 81412 85980
rect 81436 85978 81492 85980
rect 81516 85978 81572 85980
rect 81596 85978 81652 85980
rect 81356 85926 81402 85978
rect 81402 85926 81412 85978
rect 81436 85926 81466 85978
rect 81466 85926 81478 85978
rect 81478 85926 81492 85978
rect 81516 85926 81530 85978
rect 81530 85926 81542 85978
rect 81542 85926 81572 85978
rect 81596 85926 81606 85978
rect 81606 85926 81652 85978
rect 81356 85924 81412 85926
rect 81436 85924 81492 85926
rect 81516 85924 81572 85926
rect 81596 85924 81652 85926
rect 82956 85978 83012 85980
rect 83036 85978 83092 85980
rect 83116 85978 83172 85980
rect 83196 85978 83252 85980
rect 82956 85926 83002 85978
rect 83002 85926 83012 85978
rect 83036 85926 83066 85978
rect 83066 85926 83078 85978
rect 83078 85926 83092 85978
rect 83116 85926 83130 85978
rect 83130 85926 83142 85978
rect 83142 85926 83172 85978
rect 83196 85926 83206 85978
rect 83206 85926 83252 85978
rect 82956 85924 83012 85926
rect 83036 85924 83092 85926
rect 83116 85924 83172 85926
rect 83196 85924 83252 85926
rect 84556 85978 84612 85980
rect 84636 85978 84692 85980
rect 84716 85978 84772 85980
rect 84796 85978 84852 85980
rect 84556 85926 84602 85978
rect 84602 85926 84612 85978
rect 84636 85926 84666 85978
rect 84666 85926 84678 85978
rect 84678 85926 84692 85978
rect 84716 85926 84730 85978
rect 84730 85926 84742 85978
rect 84742 85926 84772 85978
rect 84796 85926 84806 85978
rect 84806 85926 84852 85978
rect 84556 85924 84612 85926
rect 84636 85924 84692 85926
rect 84716 85924 84772 85926
rect 84796 85924 84852 85926
rect 86156 85978 86212 85980
rect 86236 85978 86292 85980
rect 86316 85978 86372 85980
rect 86396 85978 86452 85980
rect 86156 85926 86202 85978
rect 86202 85926 86212 85978
rect 86236 85926 86266 85978
rect 86266 85926 86278 85978
rect 86278 85926 86292 85978
rect 86316 85926 86330 85978
rect 86330 85926 86342 85978
rect 86342 85926 86372 85978
rect 86396 85926 86406 85978
rect 86406 85926 86452 85978
rect 86156 85924 86212 85926
rect 86236 85924 86292 85926
rect 86316 85924 86372 85926
rect 86396 85924 86452 85926
rect 87756 85978 87812 85980
rect 87836 85978 87892 85980
rect 87916 85978 87972 85980
rect 87996 85978 88052 85980
rect 87756 85926 87802 85978
rect 87802 85926 87812 85978
rect 87836 85926 87866 85978
rect 87866 85926 87878 85978
rect 87878 85926 87892 85978
rect 87916 85926 87930 85978
rect 87930 85926 87942 85978
rect 87942 85926 87972 85978
rect 87996 85926 88006 85978
rect 88006 85926 88052 85978
rect 87756 85924 87812 85926
rect 87836 85924 87892 85926
rect 87916 85924 87972 85926
rect 87996 85924 88052 85926
rect 89356 85978 89412 85980
rect 89436 85978 89492 85980
rect 89516 85978 89572 85980
rect 89596 85978 89652 85980
rect 89356 85926 89402 85978
rect 89402 85926 89412 85978
rect 89436 85926 89466 85978
rect 89466 85926 89478 85978
rect 89478 85926 89492 85978
rect 89516 85926 89530 85978
rect 89530 85926 89542 85978
rect 89542 85926 89572 85978
rect 89596 85926 89606 85978
rect 89606 85926 89652 85978
rect 89356 85924 89412 85926
rect 89436 85924 89492 85926
rect 89516 85924 89572 85926
rect 89596 85924 89652 85926
rect 90956 85978 91012 85980
rect 91036 85978 91092 85980
rect 91116 85978 91172 85980
rect 91196 85978 91252 85980
rect 90956 85926 91002 85978
rect 91002 85926 91012 85978
rect 91036 85926 91066 85978
rect 91066 85926 91078 85978
rect 91078 85926 91092 85978
rect 91116 85926 91130 85978
rect 91130 85926 91142 85978
rect 91142 85926 91172 85978
rect 91196 85926 91206 85978
rect 91206 85926 91252 85978
rect 90956 85924 91012 85926
rect 91036 85924 91092 85926
rect 91116 85924 91172 85926
rect 91196 85924 91252 85926
rect 91616 86522 91672 86524
rect 91696 86522 91752 86524
rect 91776 86522 91832 86524
rect 91856 86522 91912 86524
rect 91616 86470 91662 86522
rect 91662 86470 91672 86522
rect 91696 86470 91726 86522
rect 91726 86470 91738 86522
rect 91738 86470 91752 86522
rect 91776 86470 91790 86522
rect 91790 86470 91802 86522
rect 91802 86470 91832 86522
rect 91856 86470 91866 86522
rect 91866 86470 91912 86522
rect 91616 86468 91672 86470
rect 91696 86468 91752 86470
rect 91776 86468 91832 86470
rect 91856 86468 91912 86470
rect 93216 86522 93272 86524
rect 93296 86522 93352 86524
rect 93376 86522 93432 86524
rect 93456 86522 93512 86524
rect 93216 86470 93262 86522
rect 93262 86470 93272 86522
rect 93296 86470 93326 86522
rect 93326 86470 93338 86522
rect 93338 86470 93352 86522
rect 93376 86470 93390 86522
rect 93390 86470 93402 86522
rect 93402 86470 93432 86522
rect 93456 86470 93466 86522
rect 93466 86470 93512 86522
rect 93216 86468 93272 86470
rect 93296 86468 93352 86470
rect 93376 86468 93432 86470
rect 93456 86468 93512 86470
rect 94816 86522 94872 86524
rect 94896 86522 94952 86524
rect 94976 86522 95032 86524
rect 95056 86522 95112 86524
rect 94816 86470 94862 86522
rect 94862 86470 94872 86522
rect 94896 86470 94926 86522
rect 94926 86470 94938 86522
rect 94938 86470 94952 86522
rect 94976 86470 94990 86522
rect 94990 86470 95002 86522
rect 95002 86470 95032 86522
rect 95056 86470 95066 86522
rect 95066 86470 95112 86522
rect 94816 86468 94872 86470
rect 94896 86468 94952 86470
rect 94976 86468 95032 86470
rect 95056 86468 95112 86470
rect 96416 86522 96472 86524
rect 96496 86522 96552 86524
rect 96576 86522 96632 86524
rect 96656 86522 96712 86524
rect 96416 86470 96462 86522
rect 96462 86470 96472 86522
rect 96496 86470 96526 86522
rect 96526 86470 96538 86522
rect 96538 86470 96552 86522
rect 96576 86470 96590 86522
rect 96590 86470 96602 86522
rect 96602 86470 96632 86522
rect 96656 86470 96666 86522
rect 96666 86470 96712 86522
rect 96416 86468 96472 86470
rect 96496 86468 96552 86470
rect 96576 86468 96632 86470
rect 96656 86468 96712 86470
rect 98016 86522 98072 86524
rect 98096 86522 98152 86524
rect 98176 86522 98232 86524
rect 98256 86522 98312 86524
rect 98016 86470 98062 86522
rect 98062 86470 98072 86522
rect 98096 86470 98126 86522
rect 98126 86470 98138 86522
rect 98138 86470 98152 86522
rect 98176 86470 98190 86522
rect 98190 86470 98202 86522
rect 98202 86470 98232 86522
rect 98256 86470 98266 86522
rect 98266 86470 98312 86522
rect 98016 86468 98072 86470
rect 98096 86468 98152 86470
rect 98176 86468 98232 86470
rect 98256 86468 98312 86470
rect 99616 86522 99672 86524
rect 99696 86522 99752 86524
rect 99776 86522 99832 86524
rect 99856 86522 99912 86524
rect 99616 86470 99662 86522
rect 99662 86470 99672 86522
rect 99696 86470 99726 86522
rect 99726 86470 99738 86522
rect 99738 86470 99752 86522
rect 99776 86470 99790 86522
rect 99790 86470 99802 86522
rect 99802 86470 99832 86522
rect 99856 86470 99866 86522
rect 99866 86470 99912 86522
rect 99616 86468 99672 86470
rect 99696 86468 99752 86470
rect 99776 86468 99832 86470
rect 99856 86468 99912 86470
rect 101216 86522 101272 86524
rect 101296 86522 101352 86524
rect 101376 86522 101432 86524
rect 101456 86522 101512 86524
rect 101216 86470 101262 86522
rect 101262 86470 101272 86522
rect 101296 86470 101326 86522
rect 101326 86470 101338 86522
rect 101338 86470 101352 86522
rect 101376 86470 101390 86522
rect 101390 86470 101402 86522
rect 101402 86470 101432 86522
rect 101456 86470 101466 86522
rect 101466 86470 101512 86522
rect 101216 86468 101272 86470
rect 101296 86468 101352 86470
rect 101376 86468 101432 86470
rect 101456 86468 101512 86470
rect 102816 86522 102872 86524
rect 102896 86522 102952 86524
rect 102976 86522 103032 86524
rect 103056 86522 103112 86524
rect 102816 86470 102862 86522
rect 102862 86470 102872 86522
rect 102896 86470 102926 86522
rect 102926 86470 102938 86522
rect 102938 86470 102952 86522
rect 102976 86470 102990 86522
rect 102990 86470 103002 86522
rect 103002 86470 103032 86522
rect 103056 86470 103066 86522
rect 103066 86470 103112 86522
rect 102816 86468 102872 86470
rect 102896 86468 102952 86470
rect 102976 86468 103032 86470
rect 103056 86468 103112 86470
rect 104416 86522 104472 86524
rect 104496 86522 104552 86524
rect 104576 86522 104632 86524
rect 104656 86522 104712 86524
rect 104416 86470 104462 86522
rect 104462 86470 104472 86522
rect 104496 86470 104526 86522
rect 104526 86470 104538 86522
rect 104538 86470 104552 86522
rect 104576 86470 104590 86522
rect 104590 86470 104602 86522
rect 104602 86470 104632 86522
rect 104656 86470 104666 86522
rect 104666 86470 104712 86522
rect 104416 86468 104472 86470
rect 104496 86468 104552 86470
rect 104576 86468 104632 86470
rect 104656 86468 104712 86470
rect 106016 86522 106072 86524
rect 106096 86522 106152 86524
rect 106176 86522 106232 86524
rect 106256 86522 106312 86524
rect 106016 86470 106062 86522
rect 106062 86470 106072 86522
rect 106096 86470 106126 86522
rect 106126 86470 106138 86522
rect 106138 86470 106152 86522
rect 106176 86470 106190 86522
rect 106190 86470 106202 86522
rect 106202 86470 106232 86522
rect 106256 86470 106266 86522
rect 106266 86470 106312 86522
rect 106016 86468 106072 86470
rect 106096 86468 106152 86470
rect 106176 86468 106232 86470
rect 106256 86468 106312 86470
rect 107616 86522 107672 86524
rect 107696 86522 107752 86524
rect 107776 86522 107832 86524
rect 107856 86522 107912 86524
rect 107616 86470 107662 86522
rect 107662 86470 107672 86522
rect 107696 86470 107726 86522
rect 107726 86470 107738 86522
rect 107738 86470 107752 86522
rect 107776 86470 107790 86522
rect 107790 86470 107802 86522
rect 107802 86470 107832 86522
rect 107856 86470 107866 86522
rect 107866 86470 107912 86522
rect 107616 86468 107672 86470
rect 107696 86468 107752 86470
rect 107776 86468 107832 86470
rect 107856 86468 107912 86470
rect 92556 85978 92612 85980
rect 92636 85978 92692 85980
rect 92716 85978 92772 85980
rect 92796 85978 92852 85980
rect 92556 85926 92602 85978
rect 92602 85926 92612 85978
rect 92636 85926 92666 85978
rect 92666 85926 92678 85978
rect 92678 85926 92692 85978
rect 92716 85926 92730 85978
rect 92730 85926 92742 85978
rect 92742 85926 92772 85978
rect 92796 85926 92806 85978
rect 92806 85926 92852 85978
rect 92556 85924 92612 85926
rect 92636 85924 92692 85926
rect 92716 85924 92772 85926
rect 92796 85924 92852 85926
rect 94156 85978 94212 85980
rect 94236 85978 94292 85980
rect 94316 85978 94372 85980
rect 94396 85978 94452 85980
rect 94156 85926 94202 85978
rect 94202 85926 94212 85978
rect 94236 85926 94266 85978
rect 94266 85926 94278 85978
rect 94278 85926 94292 85978
rect 94316 85926 94330 85978
rect 94330 85926 94342 85978
rect 94342 85926 94372 85978
rect 94396 85926 94406 85978
rect 94406 85926 94452 85978
rect 94156 85924 94212 85926
rect 94236 85924 94292 85926
rect 94316 85924 94372 85926
rect 94396 85924 94452 85926
rect 95756 85978 95812 85980
rect 95836 85978 95892 85980
rect 95916 85978 95972 85980
rect 95996 85978 96052 85980
rect 95756 85926 95802 85978
rect 95802 85926 95812 85978
rect 95836 85926 95866 85978
rect 95866 85926 95878 85978
rect 95878 85926 95892 85978
rect 95916 85926 95930 85978
rect 95930 85926 95942 85978
rect 95942 85926 95972 85978
rect 95996 85926 96006 85978
rect 96006 85926 96052 85978
rect 95756 85924 95812 85926
rect 95836 85924 95892 85926
rect 95916 85924 95972 85926
rect 95996 85924 96052 85926
rect 97356 85978 97412 85980
rect 97436 85978 97492 85980
rect 97516 85978 97572 85980
rect 97596 85978 97652 85980
rect 97356 85926 97402 85978
rect 97402 85926 97412 85978
rect 97436 85926 97466 85978
rect 97466 85926 97478 85978
rect 97478 85926 97492 85978
rect 97516 85926 97530 85978
rect 97530 85926 97542 85978
rect 97542 85926 97572 85978
rect 97596 85926 97606 85978
rect 97606 85926 97652 85978
rect 97356 85924 97412 85926
rect 97436 85924 97492 85926
rect 97516 85924 97572 85926
rect 97596 85924 97652 85926
rect 98956 85978 99012 85980
rect 99036 85978 99092 85980
rect 99116 85978 99172 85980
rect 99196 85978 99252 85980
rect 98956 85926 99002 85978
rect 99002 85926 99012 85978
rect 99036 85926 99066 85978
rect 99066 85926 99078 85978
rect 99078 85926 99092 85978
rect 99116 85926 99130 85978
rect 99130 85926 99142 85978
rect 99142 85926 99172 85978
rect 99196 85926 99206 85978
rect 99206 85926 99252 85978
rect 98956 85924 99012 85926
rect 99036 85924 99092 85926
rect 99116 85924 99172 85926
rect 99196 85924 99252 85926
rect 100556 85978 100612 85980
rect 100636 85978 100692 85980
rect 100716 85978 100772 85980
rect 100796 85978 100852 85980
rect 100556 85926 100602 85978
rect 100602 85926 100612 85978
rect 100636 85926 100666 85978
rect 100666 85926 100678 85978
rect 100678 85926 100692 85978
rect 100716 85926 100730 85978
rect 100730 85926 100742 85978
rect 100742 85926 100772 85978
rect 100796 85926 100806 85978
rect 100806 85926 100852 85978
rect 100556 85924 100612 85926
rect 100636 85924 100692 85926
rect 100716 85924 100772 85926
rect 100796 85924 100852 85926
rect 102156 85978 102212 85980
rect 102236 85978 102292 85980
rect 102316 85978 102372 85980
rect 102396 85978 102452 85980
rect 102156 85926 102202 85978
rect 102202 85926 102212 85978
rect 102236 85926 102266 85978
rect 102266 85926 102278 85978
rect 102278 85926 102292 85978
rect 102316 85926 102330 85978
rect 102330 85926 102342 85978
rect 102342 85926 102372 85978
rect 102396 85926 102406 85978
rect 102406 85926 102452 85978
rect 102156 85924 102212 85926
rect 102236 85924 102292 85926
rect 102316 85924 102372 85926
rect 102396 85924 102452 85926
rect 103756 85978 103812 85980
rect 103836 85978 103892 85980
rect 103916 85978 103972 85980
rect 103996 85978 104052 85980
rect 103756 85926 103802 85978
rect 103802 85926 103812 85978
rect 103836 85926 103866 85978
rect 103866 85926 103878 85978
rect 103878 85926 103892 85978
rect 103916 85926 103930 85978
rect 103930 85926 103942 85978
rect 103942 85926 103972 85978
rect 103996 85926 104006 85978
rect 104006 85926 104052 85978
rect 103756 85924 103812 85926
rect 103836 85924 103892 85926
rect 103916 85924 103972 85926
rect 103996 85924 104052 85926
rect 105356 85978 105412 85980
rect 105436 85978 105492 85980
rect 105516 85978 105572 85980
rect 105596 85978 105652 85980
rect 105356 85926 105402 85978
rect 105402 85926 105412 85978
rect 105436 85926 105466 85978
rect 105466 85926 105478 85978
rect 105478 85926 105492 85978
rect 105516 85926 105530 85978
rect 105530 85926 105542 85978
rect 105542 85926 105572 85978
rect 105596 85926 105606 85978
rect 105606 85926 105652 85978
rect 105356 85924 105412 85926
rect 105436 85924 105492 85926
rect 105516 85924 105572 85926
rect 105596 85924 105652 85926
rect 106956 85978 107012 85980
rect 107036 85978 107092 85980
rect 107116 85978 107172 85980
rect 107196 85978 107252 85980
rect 106956 85926 107002 85978
rect 107002 85926 107012 85978
rect 107036 85926 107066 85978
rect 107066 85926 107078 85978
rect 107078 85926 107092 85978
rect 107116 85926 107130 85978
rect 107130 85926 107142 85978
rect 107142 85926 107172 85978
rect 107196 85926 107206 85978
rect 107206 85926 107252 85978
rect 106956 85924 107012 85926
rect 107036 85924 107092 85926
rect 107116 85924 107172 85926
rect 107196 85924 107252 85926
rect 55218 85620 55220 85640
rect 55220 85620 55272 85640
rect 55272 85620 55274 85640
rect 55218 85584 55274 85620
rect 55678 85604 55734 85640
rect 55678 85584 55680 85604
rect 55680 85584 55732 85604
rect 55732 85584 55734 85604
rect 58346 85584 58402 85640
rect 62486 85584 62542 85640
rect 73158 85584 73214 85640
rect 74630 85584 74686 85640
rect 75918 85584 75974 85640
rect 77666 85584 77722 85640
rect 91282 85584 91338 85640
rect 100942 85584 100998 85640
rect 53010 85040 53066 85096
rect 52458 84768 52514 84824
rect 51170 84632 51226 84688
rect 53838 84632 53894 84688
rect 66258 84632 66314 84688
rect 71226 84632 71282 84688
rect 57610 84496 57666 84552
rect 78678 84496 78734 84552
rect 59910 83680 59966 83736
rect 70214 83680 70270 83736
rect 108556 85978 108612 85980
rect 108636 85978 108692 85980
rect 108716 85978 108772 85980
rect 108796 85978 108852 85980
rect 108556 85926 108602 85978
rect 108602 85926 108612 85978
rect 108636 85926 108666 85978
rect 108666 85926 108678 85978
rect 108678 85926 108692 85978
rect 108716 85926 108730 85978
rect 108730 85926 108742 85978
rect 108742 85926 108772 85978
rect 108796 85926 108806 85978
rect 108806 85926 108852 85978
rect 108556 85924 108612 85926
rect 108636 85924 108692 85926
rect 108716 85924 108772 85926
rect 108796 85924 108852 85926
rect 108026 80442 108082 80498
rect 11794 32434 11850 32490
rect 11616 1658 11672 1660
rect 11696 1658 11752 1660
rect 11776 1658 11832 1660
rect 11856 1658 11912 1660
rect 11616 1606 11662 1658
rect 11662 1606 11672 1658
rect 11696 1606 11726 1658
rect 11726 1606 11738 1658
rect 11738 1606 11752 1658
rect 11776 1606 11790 1658
rect 11790 1606 11802 1658
rect 11802 1606 11832 1658
rect 11856 1606 11866 1658
rect 11866 1606 11912 1658
rect 11616 1604 11672 1606
rect 11696 1604 11752 1606
rect 11776 1604 11832 1606
rect 11856 1604 11912 1606
rect 10956 1114 11012 1116
rect 11036 1114 11092 1116
rect 11116 1114 11172 1116
rect 11196 1114 11252 1116
rect 10956 1062 11002 1114
rect 11002 1062 11012 1114
rect 11036 1062 11066 1114
rect 11066 1062 11078 1114
rect 11078 1062 11092 1114
rect 11116 1062 11130 1114
rect 11130 1062 11142 1114
rect 11142 1062 11172 1114
rect 11196 1062 11206 1114
rect 11206 1062 11252 1114
rect 10956 1060 11012 1062
rect 11036 1060 11092 1062
rect 11116 1060 11172 1062
rect 11196 1060 11252 1062
rect 108026 20602 108082 20658
rect 107934 18400 107990 18456
rect 17866 3848 17922 3904
rect 39210 3848 39266 3904
rect 40314 3848 40370 3904
rect 45006 3848 45062 3904
rect 46110 3868 46166 3904
rect 46110 3848 46112 3868
rect 46112 3848 46164 3868
rect 46164 3848 46166 3868
rect 28722 3712 28778 3768
rect 29826 3712 29882 3768
rect 50894 3848 50950 3904
rect 54390 3884 54392 3904
rect 54392 3884 54444 3904
rect 54444 3884 54446 3904
rect 54390 3848 54446 3884
rect 47490 3712 47546 3768
rect 29642 3304 29698 3360
rect 13216 1658 13272 1660
rect 13296 1658 13352 1660
rect 13376 1658 13432 1660
rect 13456 1658 13512 1660
rect 13216 1606 13262 1658
rect 13262 1606 13272 1658
rect 13296 1606 13326 1658
rect 13326 1606 13338 1658
rect 13338 1606 13352 1658
rect 13376 1606 13390 1658
rect 13390 1606 13402 1658
rect 13402 1606 13432 1658
rect 13456 1606 13466 1658
rect 13466 1606 13512 1658
rect 13216 1604 13272 1606
rect 13296 1604 13352 1606
rect 13376 1604 13432 1606
rect 13456 1604 13512 1606
rect 14816 1658 14872 1660
rect 14896 1658 14952 1660
rect 14976 1658 15032 1660
rect 15056 1658 15112 1660
rect 14816 1606 14862 1658
rect 14862 1606 14872 1658
rect 14896 1606 14926 1658
rect 14926 1606 14938 1658
rect 14938 1606 14952 1658
rect 14976 1606 14990 1658
rect 14990 1606 15002 1658
rect 15002 1606 15032 1658
rect 15056 1606 15066 1658
rect 15066 1606 15112 1658
rect 14816 1604 14872 1606
rect 14896 1604 14952 1606
rect 14976 1604 15032 1606
rect 15056 1604 15112 1606
rect 16416 1658 16472 1660
rect 16496 1658 16552 1660
rect 16576 1658 16632 1660
rect 16656 1658 16712 1660
rect 16416 1606 16462 1658
rect 16462 1606 16472 1658
rect 16496 1606 16526 1658
rect 16526 1606 16538 1658
rect 16538 1606 16552 1658
rect 16576 1606 16590 1658
rect 16590 1606 16602 1658
rect 16602 1606 16632 1658
rect 16656 1606 16666 1658
rect 16666 1606 16712 1658
rect 16416 1604 16472 1606
rect 16496 1604 16552 1606
rect 16576 1604 16632 1606
rect 16656 1604 16712 1606
rect 18016 1658 18072 1660
rect 18096 1658 18152 1660
rect 18176 1658 18232 1660
rect 18256 1658 18312 1660
rect 18016 1606 18062 1658
rect 18062 1606 18072 1658
rect 18096 1606 18126 1658
rect 18126 1606 18138 1658
rect 18138 1606 18152 1658
rect 18176 1606 18190 1658
rect 18190 1606 18202 1658
rect 18202 1606 18232 1658
rect 18256 1606 18266 1658
rect 18266 1606 18312 1658
rect 18016 1604 18072 1606
rect 18096 1604 18152 1606
rect 18176 1604 18232 1606
rect 18256 1604 18312 1606
rect 19616 1658 19672 1660
rect 19696 1658 19752 1660
rect 19776 1658 19832 1660
rect 19856 1658 19912 1660
rect 19616 1606 19662 1658
rect 19662 1606 19672 1658
rect 19696 1606 19726 1658
rect 19726 1606 19738 1658
rect 19738 1606 19752 1658
rect 19776 1606 19790 1658
rect 19790 1606 19802 1658
rect 19802 1606 19832 1658
rect 19856 1606 19866 1658
rect 19866 1606 19912 1658
rect 19616 1604 19672 1606
rect 19696 1604 19752 1606
rect 19776 1604 19832 1606
rect 19856 1604 19912 1606
rect 21216 1658 21272 1660
rect 21296 1658 21352 1660
rect 21376 1658 21432 1660
rect 21456 1658 21512 1660
rect 21216 1606 21262 1658
rect 21262 1606 21272 1658
rect 21296 1606 21326 1658
rect 21326 1606 21338 1658
rect 21338 1606 21352 1658
rect 21376 1606 21390 1658
rect 21390 1606 21402 1658
rect 21402 1606 21432 1658
rect 21456 1606 21466 1658
rect 21466 1606 21512 1658
rect 21216 1604 21272 1606
rect 21296 1604 21352 1606
rect 21376 1604 21432 1606
rect 21456 1604 21512 1606
rect 22816 1658 22872 1660
rect 22896 1658 22952 1660
rect 22976 1658 23032 1660
rect 23056 1658 23112 1660
rect 22816 1606 22862 1658
rect 22862 1606 22872 1658
rect 22896 1606 22926 1658
rect 22926 1606 22938 1658
rect 22938 1606 22952 1658
rect 22976 1606 22990 1658
rect 22990 1606 23002 1658
rect 23002 1606 23032 1658
rect 23056 1606 23066 1658
rect 23066 1606 23112 1658
rect 22816 1604 22872 1606
rect 22896 1604 22952 1606
rect 22976 1604 23032 1606
rect 23056 1604 23112 1606
rect 24416 1658 24472 1660
rect 24496 1658 24552 1660
rect 24576 1658 24632 1660
rect 24656 1658 24712 1660
rect 24416 1606 24462 1658
rect 24462 1606 24472 1658
rect 24496 1606 24526 1658
rect 24526 1606 24538 1658
rect 24538 1606 24552 1658
rect 24576 1606 24590 1658
rect 24590 1606 24602 1658
rect 24602 1606 24632 1658
rect 24656 1606 24666 1658
rect 24666 1606 24712 1658
rect 24416 1604 24472 1606
rect 24496 1604 24552 1606
rect 24576 1604 24632 1606
rect 24656 1604 24712 1606
rect 26016 1658 26072 1660
rect 26096 1658 26152 1660
rect 26176 1658 26232 1660
rect 26256 1658 26312 1660
rect 26016 1606 26062 1658
rect 26062 1606 26072 1658
rect 26096 1606 26126 1658
rect 26126 1606 26138 1658
rect 26138 1606 26152 1658
rect 26176 1606 26190 1658
rect 26190 1606 26202 1658
rect 26202 1606 26232 1658
rect 26256 1606 26266 1658
rect 26266 1606 26312 1658
rect 26016 1604 26072 1606
rect 26096 1604 26152 1606
rect 26176 1604 26232 1606
rect 26256 1604 26312 1606
rect 12556 1114 12612 1116
rect 12636 1114 12692 1116
rect 12716 1114 12772 1116
rect 12796 1114 12852 1116
rect 12556 1062 12602 1114
rect 12602 1062 12612 1114
rect 12636 1062 12666 1114
rect 12666 1062 12678 1114
rect 12678 1062 12692 1114
rect 12716 1062 12730 1114
rect 12730 1062 12742 1114
rect 12742 1062 12772 1114
rect 12796 1062 12806 1114
rect 12806 1062 12852 1114
rect 12556 1060 12612 1062
rect 12636 1060 12692 1062
rect 12716 1060 12772 1062
rect 12796 1060 12852 1062
rect 14156 1114 14212 1116
rect 14236 1114 14292 1116
rect 14316 1114 14372 1116
rect 14396 1114 14452 1116
rect 14156 1062 14202 1114
rect 14202 1062 14212 1114
rect 14236 1062 14266 1114
rect 14266 1062 14278 1114
rect 14278 1062 14292 1114
rect 14316 1062 14330 1114
rect 14330 1062 14342 1114
rect 14342 1062 14372 1114
rect 14396 1062 14406 1114
rect 14406 1062 14452 1114
rect 14156 1060 14212 1062
rect 14236 1060 14292 1062
rect 14316 1060 14372 1062
rect 14396 1060 14452 1062
rect 15756 1114 15812 1116
rect 15836 1114 15892 1116
rect 15916 1114 15972 1116
rect 15996 1114 16052 1116
rect 15756 1062 15802 1114
rect 15802 1062 15812 1114
rect 15836 1062 15866 1114
rect 15866 1062 15878 1114
rect 15878 1062 15892 1114
rect 15916 1062 15930 1114
rect 15930 1062 15942 1114
rect 15942 1062 15972 1114
rect 15996 1062 16006 1114
rect 16006 1062 16052 1114
rect 15756 1060 15812 1062
rect 15836 1060 15892 1062
rect 15916 1060 15972 1062
rect 15996 1060 16052 1062
rect 17356 1114 17412 1116
rect 17436 1114 17492 1116
rect 17516 1114 17572 1116
rect 17596 1114 17652 1116
rect 17356 1062 17402 1114
rect 17402 1062 17412 1114
rect 17436 1062 17466 1114
rect 17466 1062 17478 1114
rect 17478 1062 17492 1114
rect 17516 1062 17530 1114
rect 17530 1062 17542 1114
rect 17542 1062 17572 1114
rect 17596 1062 17606 1114
rect 17606 1062 17652 1114
rect 17356 1060 17412 1062
rect 17436 1060 17492 1062
rect 17516 1060 17572 1062
rect 17596 1060 17652 1062
rect 18956 1114 19012 1116
rect 19036 1114 19092 1116
rect 19116 1114 19172 1116
rect 19196 1114 19252 1116
rect 18956 1062 19002 1114
rect 19002 1062 19012 1114
rect 19036 1062 19066 1114
rect 19066 1062 19078 1114
rect 19078 1062 19092 1114
rect 19116 1062 19130 1114
rect 19130 1062 19142 1114
rect 19142 1062 19172 1114
rect 19196 1062 19206 1114
rect 19206 1062 19252 1114
rect 18956 1060 19012 1062
rect 19036 1060 19092 1062
rect 19116 1060 19172 1062
rect 19196 1060 19252 1062
rect 20556 1114 20612 1116
rect 20636 1114 20692 1116
rect 20716 1114 20772 1116
rect 20796 1114 20852 1116
rect 20556 1062 20602 1114
rect 20602 1062 20612 1114
rect 20636 1062 20666 1114
rect 20666 1062 20678 1114
rect 20678 1062 20692 1114
rect 20716 1062 20730 1114
rect 20730 1062 20742 1114
rect 20742 1062 20772 1114
rect 20796 1062 20806 1114
rect 20806 1062 20852 1114
rect 20556 1060 20612 1062
rect 20636 1060 20692 1062
rect 20716 1060 20772 1062
rect 20796 1060 20852 1062
rect 22156 1114 22212 1116
rect 22236 1114 22292 1116
rect 22316 1114 22372 1116
rect 22396 1114 22452 1116
rect 22156 1062 22202 1114
rect 22202 1062 22212 1114
rect 22236 1062 22266 1114
rect 22266 1062 22278 1114
rect 22278 1062 22292 1114
rect 22316 1062 22330 1114
rect 22330 1062 22342 1114
rect 22342 1062 22372 1114
rect 22396 1062 22406 1114
rect 22406 1062 22452 1114
rect 22156 1060 22212 1062
rect 22236 1060 22292 1062
rect 22316 1060 22372 1062
rect 22396 1060 22452 1062
rect 10598 448 10654 504
rect 27616 1658 27672 1660
rect 27696 1658 27752 1660
rect 27776 1658 27832 1660
rect 27856 1658 27912 1660
rect 27616 1606 27662 1658
rect 27662 1606 27672 1658
rect 27696 1606 27726 1658
rect 27726 1606 27738 1658
rect 27738 1606 27752 1658
rect 27776 1606 27790 1658
rect 27790 1606 27802 1658
rect 27802 1606 27832 1658
rect 27856 1606 27866 1658
rect 27866 1606 27912 1658
rect 27616 1604 27672 1606
rect 27696 1604 27752 1606
rect 27776 1604 27832 1606
rect 27856 1604 27912 1606
rect 29216 1658 29272 1660
rect 29296 1658 29352 1660
rect 29376 1658 29432 1660
rect 29456 1658 29512 1660
rect 29216 1606 29262 1658
rect 29262 1606 29272 1658
rect 29296 1606 29326 1658
rect 29326 1606 29338 1658
rect 29338 1606 29352 1658
rect 29376 1606 29390 1658
rect 29390 1606 29402 1658
rect 29402 1606 29432 1658
rect 29456 1606 29466 1658
rect 29466 1606 29512 1658
rect 29216 1604 29272 1606
rect 29296 1604 29352 1606
rect 29376 1604 29432 1606
rect 29456 1604 29512 1606
rect 32034 2352 32090 2408
rect 30816 1658 30872 1660
rect 30896 1658 30952 1660
rect 30976 1658 31032 1660
rect 31056 1658 31112 1660
rect 30816 1606 30862 1658
rect 30862 1606 30872 1658
rect 30896 1606 30926 1658
rect 30926 1606 30938 1658
rect 30938 1606 30952 1658
rect 30976 1606 30990 1658
rect 30990 1606 31002 1658
rect 31002 1606 31032 1658
rect 31056 1606 31066 1658
rect 31066 1606 31112 1658
rect 30816 1604 30872 1606
rect 30896 1604 30952 1606
rect 30976 1604 31032 1606
rect 31056 1604 31112 1606
rect 32416 1658 32472 1660
rect 32496 1658 32552 1660
rect 32576 1658 32632 1660
rect 32656 1658 32712 1660
rect 32416 1606 32462 1658
rect 32462 1606 32472 1658
rect 32496 1606 32526 1658
rect 32526 1606 32538 1658
rect 32538 1606 32552 1658
rect 32576 1606 32590 1658
rect 32590 1606 32602 1658
rect 32602 1606 32632 1658
rect 32656 1606 32666 1658
rect 32666 1606 32712 1658
rect 32416 1604 32472 1606
rect 32496 1604 32552 1606
rect 32576 1604 32632 1606
rect 32656 1604 32712 1606
rect 34016 1658 34072 1660
rect 34096 1658 34152 1660
rect 34176 1658 34232 1660
rect 34256 1658 34312 1660
rect 34016 1606 34062 1658
rect 34062 1606 34072 1658
rect 34096 1606 34126 1658
rect 34126 1606 34138 1658
rect 34138 1606 34152 1658
rect 34176 1606 34190 1658
rect 34190 1606 34202 1658
rect 34202 1606 34232 1658
rect 34256 1606 34266 1658
rect 34266 1606 34312 1658
rect 34016 1604 34072 1606
rect 34096 1604 34152 1606
rect 34176 1604 34232 1606
rect 34256 1604 34312 1606
rect 37002 2624 37058 2680
rect 49698 2624 49754 2680
rect 42798 2352 42854 2408
rect 43810 2352 43866 2408
rect 48594 2352 48650 2408
rect 37462 2080 37518 2136
rect 35616 1658 35672 1660
rect 35696 1658 35752 1660
rect 35776 1658 35832 1660
rect 35856 1658 35912 1660
rect 35616 1606 35662 1658
rect 35662 1606 35672 1658
rect 35696 1606 35726 1658
rect 35726 1606 35738 1658
rect 35738 1606 35752 1658
rect 35776 1606 35790 1658
rect 35790 1606 35802 1658
rect 35802 1606 35832 1658
rect 35856 1606 35866 1658
rect 35866 1606 35912 1658
rect 35616 1604 35672 1606
rect 35696 1604 35752 1606
rect 35776 1604 35832 1606
rect 35856 1604 35912 1606
rect 37216 1658 37272 1660
rect 37296 1658 37352 1660
rect 37376 1658 37432 1660
rect 37456 1658 37512 1660
rect 37216 1606 37262 1658
rect 37262 1606 37272 1658
rect 37296 1606 37326 1658
rect 37326 1606 37338 1658
rect 37338 1606 37352 1658
rect 37376 1606 37390 1658
rect 37390 1606 37402 1658
rect 37402 1606 37432 1658
rect 37456 1606 37466 1658
rect 37466 1606 37512 1658
rect 37216 1604 37272 1606
rect 37296 1604 37352 1606
rect 37376 1604 37432 1606
rect 37456 1604 37512 1606
rect 38816 1658 38872 1660
rect 38896 1658 38952 1660
rect 38976 1658 39032 1660
rect 39056 1658 39112 1660
rect 38816 1606 38862 1658
rect 38862 1606 38872 1658
rect 38896 1606 38926 1658
rect 38926 1606 38938 1658
rect 38938 1606 38952 1658
rect 38976 1606 38990 1658
rect 38990 1606 39002 1658
rect 39002 1606 39032 1658
rect 39056 1606 39066 1658
rect 39066 1606 39112 1658
rect 38816 1604 38872 1606
rect 38896 1604 38952 1606
rect 38976 1604 39032 1606
rect 39056 1604 39112 1606
rect 40416 1658 40472 1660
rect 40496 1658 40552 1660
rect 40576 1658 40632 1660
rect 40656 1658 40712 1660
rect 40416 1606 40462 1658
rect 40462 1606 40472 1658
rect 40496 1606 40526 1658
rect 40526 1606 40538 1658
rect 40538 1606 40552 1658
rect 40576 1606 40590 1658
rect 40590 1606 40602 1658
rect 40602 1606 40632 1658
rect 40656 1606 40666 1658
rect 40666 1606 40712 1658
rect 40416 1604 40472 1606
rect 40496 1604 40552 1606
rect 40576 1604 40632 1606
rect 40656 1604 40712 1606
rect 42016 1658 42072 1660
rect 42096 1658 42152 1660
rect 42176 1658 42232 1660
rect 42256 1658 42312 1660
rect 42016 1606 42062 1658
rect 42062 1606 42072 1658
rect 42096 1606 42126 1658
rect 42126 1606 42138 1658
rect 42138 1606 42152 1658
rect 42176 1606 42190 1658
rect 42190 1606 42202 1658
rect 42202 1606 42232 1658
rect 42256 1606 42266 1658
rect 42266 1606 42312 1658
rect 42016 1604 42072 1606
rect 42096 1604 42152 1606
rect 42176 1604 42232 1606
rect 42256 1604 42312 1606
rect 43616 1658 43672 1660
rect 43696 1658 43752 1660
rect 43776 1658 43832 1660
rect 43856 1658 43912 1660
rect 43616 1606 43662 1658
rect 43662 1606 43672 1658
rect 43696 1606 43726 1658
rect 43726 1606 43738 1658
rect 43738 1606 43752 1658
rect 43776 1606 43790 1658
rect 43790 1606 43802 1658
rect 43802 1606 43832 1658
rect 43856 1606 43866 1658
rect 43866 1606 43912 1658
rect 43616 1604 43672 1606
rect 43696 1604 43752 1606
rect 43776 1604 43832 1606
rect 43856 1604 43912 1606
rect 45216 1658 45272 1660
rect 45296 1658 45352 1660
rect 45376 1658 45432 1660
rect 45456 1658 45512 1660
rect 45216 1606 45262 1658
rect 45262 1606 45272 1658
rect 45296 1606 45326 1658
rect 45326 1606 45338 1658
rect 45338 1606 45352 1658
rect 45376 1606 45390 1658
rect 45390 1606 45402 1658
rect 45402 1606 45432 1658
rect 45456 1606 45466 1658
rect 45466 1606 45512 1658
rect 45216 1604 45272 1606
rect 45296 1604 45352 1606
rect 45376 1604 45432 1606
rect 45456 1604 45512 1606
rect 46816 1658 46872 1660
rect 46896 1658 46952 1660
rect 46976 1658 47032 1660
rect 47056 1658 47112 1660
rect 46816 1606 46862 1658
rect 46862 1606 46872 1658
rect 46896 1606 46926 1658
rect 46926 1606 46938 1658
rect 46938 1606 46952 1658
rect 46976 1606 46990 1658
rect 46990 1606 47002 1658
rect 47002 1606 47032 1658
rect 47056 1606 47066 1658
rect 47066 1606 47112 1658
rect 46816 1604 46872 1606
rect 46896 1604 46952 1606
rect 46976 1604 47032 1606
rect 47056 1604 47112 1606
rect 48416 1658 48472 1660
rect 48496 1658 48552 1660
rect 48576 1658 48632 1660
rect 48656 1658 48712 1660
rect 48416 1606 48462 1658
rect 48462 1606 48472 1658
rect 48496 1606 48526 1658
rect 48526 1606 48538 1658
rect 48538 1606 48552 1658
rect 48576 1606 48590 1658
rect 48590 1606 48602 1658
rect 48602 1606 48632 1658
rect 48656 1606 48666 1658
rect 48666 1606 48712 1658
rect 48416 1604 48472 1606
rect 48496 1604 48552 1606
rect 48576 1604 48632 1606
rect 48656 1604 48712 1606
rect 50016 1658 50072 1660
rect 50096 1658 50152 1660
rect 50176 1658 50232 1660
rect 50256 1658 50312 1660
rect 50016 1606 50062 1658
rect 50062 1606 50072 1658
rect 50096 1606 50126 1658
rect 50126 1606 50138 1658
rect 50138 1606 50152 1658
rect 50176 1606 50190 1658
rect 50190 1606 50202 1658
rect 50202 1606 50232 1658
rect 50256 1606 50266 1658
rect 50266 1606 50312 1658
rect 50016 1604 50072 1606
rect 50096 1604 50152 1606
rect 50176 1604 50232 1606
rect 50256 1604 50312 1606
rect 51616 1658 51672 1660
rect 51696 1658 51752 1660
rect 51776 1658 51832 1660
rect 51856 1658 51912 1660
rect 51616 1606 51662 1658
rect 51662 1606 51672 1658
rect 51696 1606 51726 1658
rect 51726 1606 51738 1658
rect 51738 1606 51752 1658
rect 51776 1606 51790 1658
rect 51790 1606 51802 1658
rect 51802 1606 51832 1658
rect 51856 1606 51866 1658
rect 51866 1606 51912 1658
rect 51616 1604 51672 1606
rect 51696 1604 51752 1606
rect 51776 1604 51832 1606
rect 51856 1604 51912 1606
rect 53216 1658 53272 1660
rect 53296 1658 53352 1660
rect 53376 1658 53432 1660
rect 53456 1658 53512 1660
rect 53216 1606 53262 1658
rect 53262 1606 53272 1658
rect 53296 1606 53326 1658
rect 53326 1606 53338 1658
rect 53338 1606 53352 1658
rect 53376 1606 53390 1658
rect 53390 1606 53402 1658
rect 53402 1606 53432 1658
rect 53456 1606 53466 1658
rect 53466 1606 53512 1658
rect 53216 1604 53272 1606
rect 53296 1604 53352 1606
rect 53376 1604 53432 1606
rect 53456 1604 53512 1606
rect 23756 1114 23812 1116
rect 23836 1114 23892 1116
rect 23916 1114 23972 1116
rect 23996 1114 24052 1116
rect 23756 1062 23802 1114
rect 23802 1062 23812 1114
rect 23836 1062 23866 1114
rect 23866 1062 23878 1114
rect 23878 1062 23892 1114
rect 23916 1062 23930 1114
rect 23930 1062 23942 1114
rect 23942 1062 23972 1114
rect 23996 1062 24006 1114
rect 24006 1062 24052 1114
rect 23756 1060 23812 1062
rect 23836 1060 23892 1062
rect 23916 1060 23972 1062
rect 23996 1060 24052 1062
rect 25356 1114 25412 1116
rect 25436 1114 25492 1116
rect 25516 1114 25572 1116
rect 25596 1114 25652 1116
rect 25356 1062 25402 1114
rect 25402 1062 25412 1114
rect 25436 1062 25466 1114
rect 25466 1062 25478 1114
rect 25478 1062 25492 1114
rect 25516 1062 25530 1114
rect 25530 1062 25542 1114
rect 25542 1062 25572 1114
rect 25596 1062 25606 1114
rect 25606 1062 25652 1114
rect 25356 1060 25412 1062
rect 25436 1060 25492 1062
rect 25516 1060 25572 1062
rect 25596 1060 25652 1062
rect 26956 1114 27012 1116
rect 27036 1114 27092 1116
rect 27116 1114 27172 1116
rect 27196 1114 27252 1116
rect 26956 1062 27002 1114
rect 27002 1062 27012 1114
rect 27036 1062 27066 1114
rect 27066 1062 27078 1114
rect 27078 1062 27092 1114
rect 27116 1062 27130 1114
rect 27130 1062 27142 1114
rect 27142 1062 27172 1114
rect 27196 1062 27206 1114
rect 27206 1062 27252 1114
rect 26956 1060 27012 1062
rect 27036 1060 27092 1062
rect 27116 1060 27172 1062
rect 27196 1060 27252 1062
rect 26330 856 26386 912
rect 30562 1264 30618 1320
rect 28556 1114 28612 1116
rect 28636 1114 28692 1116
rect 28716 1114 28772 1116
rect 28796 1114 28852 1116
rect 28556 1062 28602 1114
rect 28602 1062 28612 1114
rect 28636 1062 28666 1114
rect 28666 1062 28678 1114
rect 28678 1062 28692 1114
rect 28716 1062 28730 1114
rect 28730 1062 28742 1114
rect 28742 1062 28772 1114
rect 28796 1062 28806 1114
rect 28806 1062 28852 1114
rect 28556 1060 28612 1062
rect 28636 1060 28692 1062
rect 28716 1060 28772 1062
rect 28796 1060 28852 1062
rect 30156 1114 30212 1116
rect 30236 1114 30292 1116
rect 30316 1114 30372 1116
rect 30396 1114 30452 1116
rect 30156 1062 30202 1114
rect 30202 1062 30212 1114
rect 30236 1062 30266 1114
rect 30266 1062 30278 1114
rect 30278 1062 30292 1114
rect 30316 1062 30330 1114
rect 30330 1062 30342 1114
rect 30342 1062 30372 1114
rect 30396 1062 30406 1114
rect 30406 1062 30452 1114
rect 30156 1060 30212 1062
rect 30236 1060 30292 1062
rect 30316 1060 30372 1062
rect 30396 1060 30452 1062
rect 31756 1114 31812 1116
rect 31836 1114 31892 1116
rect 31916 1114 31972 1116
rect 31996 1114 32052 1116
rect 31756 1062 31802 1114
rect 31802 1062 31812 1114
rect 31836 1062 31866 1114
rect 31866 1062 31878 1114
rect 31878 1062 31892 1114
rect 31916 1062 31930 1114
rect 31930 1062 31942 1114
rect 31942 1062 31972 1114
rect 31996 1062 32006 1114
rect 32006 1062 32052 1114
rect 31756 1060 31812 1062
rect 31836 1060 31892 1062
rect 31916 1060 31972 1062
rect 31996 1060 32052 1062
rect 32218 584 32274 640
rect 33230 1264 33286 1320
rect 33138 312 33194 368
rect 33356 1114 33412 1116
rect 33436 1114 33492 1116
rect 33516 1114 33572 1116
rect 33596 1114 33652 1116
rect 33356 1062 33402 1114
rect 33402 1062 33412 1114
rect 33436 1062 33466 1114
rect 33466 1062 33478 1114
rect 33478 1062 33492 1114
rect 33516 1062 33530 1114
rect 33530 1062 33542 1114
rect 33542 1062 33572 1114
rect 33596 1062 33606 1114
rect 33606 1062 33652 1114
rect 33356 1060 33412 1062
rect 33436 1060 33492 1062
rect 33516 1060 33572 1062
rect 33596 1060 33652 1062
rect 34518 1264 34574 1320
rect 37278 1264 37334 1320
rect 34956 1114 35012 1116
rect 35036 1114 35092 1116
rect 35116 1114 35172 1116
rect 35196 1114 35252 1116
rect 34956 1062 35002 1114
rect 35002 1062 35012 1114
rect 35036 1062 35066 1114
rect 35066 1062 35078 1114
rect 35078 1062 35092 1114
rect 35116 1062 35130 1114
rect 35130 1062 35142 1114
rect 35142 1062 35172 1114
rect 35196 1062 35206 1114
rect 35206 1062 35252 1114
rect 34956 1060 35012 1062
rect 35036 1060 35092 1062
rect 35116 1060 35172 1062
rect 35196 1060 35252 1062
rect 36556 1114 36612 1116
rect 36636 1114 36692 1116
rect 36716 1114 36772 1116
rect 36796 1114 36852 1116
rect 36556 1062 36602 1114
rect 36602 1062 36612 1114
rect 36636 1062 36666 1114
rect 36666 1062 36678 1114
rect 36678 1062 36692 1114
rect 36716 1062 36730 1114
rect 36730 1062 36742 1114
rect 36742 1062 36772 1114
rect 36796 1062 36806 1114
rect 36806 1062 36852 1114
rect 36556 1060 36612 1062
rect 36636 1060 36692 1062
rect 36716 1060 36772 1062
rect 36796 1060 36852 1062
rect 38156 1114 38212 1116
rect 38236 1114 38292 1116
rect 38316 1114 38372 1116
rect 38396 1114 38452 1116
rect 38156 1062 38202 1114
rect 38202 1062 38212 1114
rect 38236 1062 38266 1114
rect 38266 1062 38278 1114
rect 38278 1062 38292 1114
rect 38316 1062 38330 1114
rect 38330 1062 38342 1114
rect 38342 1062 38372 1114
rect 38396 1062 38406 1114
rect 38406 1062 38452 1114
rect 38156 1060 38212 1062
rect 38236 1060 38292 1062
rect 38316 1060 38372 1062
rect 38396 1060 38452 1062
rect 39756 1114 39812 1116
rect 39836 1114 39892 1116
rect 39916 1114 39972 1116
rect 39996 1114 40052 1116
rect 39756 1062 39802 1114
rect 39802 1062 39812 1114
rect 39836 1062 39866 1114
rect 39866 1062 39878 1114
rect 39878 1062 39892 1114
rect 39916 1062 39930 1114
rect 39930 1062 39942 1114
rect 39942 1062 39972 1114
rect 39996 1062 40006 1114
rect 40006 1062 40052 1114
rect 39756 1060 39812 1062
rect 39836 1060 39892 1062
rect 39916 1060 39972 1062
rect 39996 1060 40052 1062
rect 41356 1114 41412 1116
rect 41436 1114 41492 1116
rect 41516 1114 41572 1116
rect 41596 1114 41652 1116
rect 41356 1062 41402 1114
rect 41402 1062 41412 1114
rect 41436 1062 41466 1114
rect 41466 1062 41478 1114
rect 41478 1062 41492 1114
rect 41516 1062 41530 1114
rect 41530 1062 41542 1114
rect 41542 1062 41572 1114
rect 41596 1062 41606 1114
rect 41606 1062 41652 1114
rect 41356 1060 41412 1062
rect 41436 1060 41492 1062
rect 41516 1060 41572 1062
rect 41596 1060 41652 1062
rect 42956 1114 43012 1116
rect 43036 1114 43092 1116
rect 43116 1114 43172 1116
rect 43196 1114 43252 1116
rect 42956 1062 43002 1114
rect 43002 1062 43012 1114
rect 43036 1062 43066 1114
rect 43066 1062 43078 1114
rect 43078 1062 43092 1114
rect 43116 1062 43130 1114
rect 43130 1062 43142 1114
rect 43142 1062 43172 1114
rect 43196 1062 43206 1114
rect 43206 1062 43252 1114
rect 42956 1060 43012 1062
rect 43036 1060 43092 1062
rect 43116 1060 43172 1062
rect 43196 1060 43252 1062
rect 44556 1114 44612 1116
rect 44636 1114 44692 1116
rect 44716 1114 44772 1116
rect 44796 1114 44852 1116
rect 44556 1062 44602 1114
rect 44602 1062 44612 1114
rect 44636 1062 44666 1114
rect 44666 1062 44678 1114
rect 44678 1062 44692 1114
rect 44716 1062 44730 1114
rect 44730 1062 44742 1114
rect 44742 1062 44772 1114
rect 44796 1062 44806 1114
rect 44806 1062 44852 1114
rect 44556 1060 44612 1062
rect 44636 1060 44692 1062
rect 44716 1060 44772 1062
rect 44796 1060 44852 1062
rect 46156 1114 46212 1116
rect 46236 1114 46292 1116
rect 46316 1114 46372 1116
rect 46396 1114 46452 1116
rect 46156 1062 46202 1114
rect 46202 1062 46212 1114
rect 46236 1062 46266 1114
rect 46266 1062 46278 1114
rect 46278 1062 46292 1114
rect 46316 1062 46330 1114
rect 46330 1062 46342 1114
rect 46342 1062 46372 1114
rect 46396 1062 46406 1114
rect 46406 1062 46452 1114
rect 46156 1060 46212 1062
rect 46236 1060 46292 1062
rect 46316 1060 46372 1062
rect 46396 1060 46452 1062
rect 47756 1114 47812 1116
rect 47836 1114 47892 1116
rect 47916 1114 47972 1116
rect 47996 1114 48052 1116
rect 47756 1062 47802 1114
rect 47802 1062 47812 1114
rect 47836 1062 47866 1114
rect 47866 1062 47878 1114
rect 47878 1062 47892 1114
rect 47916 1062 47930 1114
rect 47930 1062 47942 1114
rect 47942 1062 47972 1114
rect 47996 1062 48006 1114
rect 48006 1062 48052 1114
rect 47756 1060 47812 1062
rect 47836 1060 47892 1062
rect 47916 1060 47972 1062
rect 47996 1060 48052 1062
rect 49356 1114 49412 1116
rect 49436 1114 49492 1116
rect 49516 1114 49572 1116
rect 49596 1114 49652 1116
rect 49356 1062 49402 1114
rect 49402 1062 49412 1114
rect 49436 1062 49466 1114
rect 49466 1062 49478 1114
rect 49478 1062 49492 1114
rect 49516 1062 49530 1114
rect 49530 1062 49542 1114
rect 49542 1062 49572 1114
rect 49596 1062 49606 1114
rect 49606 1062 49652 1114
rect 49356 1060 49412 1062
rect 49436 1060 49492 1062
rect 49516 1060 49572 1062
rect 49596 1060 49652 1062
rect 50956 1114 51012 1116
rect 51036 1114 51092 1116
rect 51116 1114 51172 1116
rect 51196 1114 51252 1116
rect 50956 1062 51002 1114
rect 51002 1062 51012 1114
rect 51036 1062 51066 1114
rect 51066 1062 51078 1114
rect 51078 1062 51092 1114
rect 51116 1062 51130 1114
rect 51130 1062 51142 1114
rect 51142 1062 51172 1114
rect 51196 1062 51206 1114
rect 51206 1062 51252 1114
rect 50956 1060 51012 1062
rect 51036 1060 51092 1062
rect 51116 1060 51172 1062
rect 51196 1060 51252 1062
rect 52556 1114 52612 1116
rect 52636 1114 52692 1116
rect 52716 1114 52772 1116
rect 52796 1114 52852 1116
rect 52556 1062 52602 1114
rect 52602 1062 52612 1114
rect 52636 1062 52666 1114
rect 52666 1062 52678 1114
rect 52678 1062 52692 1114
rect 52716 1062 52730 1114
rect 52730 1062 52742 1114
rect 52742 1062 52772 1114
rect 52796 1062 52806 1114
rect 52806 1062 52852 1114
rect 52556 1060 52612 1062
rect 52636 1060 52692 1062
rect 52716 1060 52772 1062
rect 52796 1060 52852 1062
rect 54156 1114 54212 1116
rect 54236 1114 54292 1116
rect 54316 1114 54372 1116
rect 54396 1114 54452 1116
rect 54156 1062 54202 1114
rect 54202 1062 54212 1114
rect 54236 1062 54266 1114
rect 54266 1062 54278 1114
rect 54278 1062 54292 1114
rect 54316 1062 54330 1114
rect 54330 1062 54342 1114
rect 54342 1062 54372 1114
rect 54396 1062 54406 1114
rect 54406 1062 54452 1114
rect 54156 1060 54212 1062
rect 54236 1060 54292 1062
rect 54316 1060 54372 1062
rect 54396 1060 54452 1062
rect 55402 2624 55458 2680
rect 57978 2624 58034 2680
rect 108118 17610 108174 17666
rect 108118 3576 108174 3632
rect 108026 3440 108082 3496
rect 94962 2488 95018 2544
rect 54816 1658 54872 1660
rect 54896 1658 54952 1660
rect 54976 1658 55032 1660
rect 55056 1658 55112 1660
rect 54816 1606 54862 1658
rect 54862 1606 54872 1658
rect 54896 1606 54926 1658
rect 54926 1606 54938 1658
rect 54938 1606 54952 1658
rect 54976 1606 54990 1658
rect 54990 1606 55002 1658
rect 55002 1606 55032 1658
rect 55056 1606 55066 1658
rect 55066 1606 55112 1658
rect 54816 1604 54872 1606
rect 54896 1604 54952 1606
rect 54976 1604 55032 1606
rect 55056 1604 55112 1606
rect 56416 1658 56472 1660
rect 56496 1658 56552 1660
rect 56576 1658 56632 1660
rect 56656 1658 56712 1660
rect 56416 1606 56462 1658
rect 56462 1606 56472 1658
rect 56496 1606 56526 1658
rect 56526 1606 56538 1658
rect 56538 1606 56552 1658
rect 56576 1606 56590 1658
rect 56590 1606 56602 1658
rect 56602 1606 56632 1658
rect 56656 1606 56666 1658
rect 56666 1606 56712 1658
rect 56416 1604 56472 1606
rect 56496 1604 56552 1606
rect 56576 1604 56632 1606
rect 56656 1604 56712 1606
rect 58016 1658 58072 1660
rect 58096 1658 58152 1660
rect 58176 1658 58232 1660
rect 58256 1658 58312 1660
rect 58016 1606 58062 1658
rect 58062 1606 58072 1658
rect 58096 1606 58126 1658
rect 58126 1606 58138 1658
rect 58138 1606 58152 1658
rect 58176 1606 58190 1658
rect 58190 1606 58202 1658
rect 58202 1606 58232 1658
rect 58256 1606 58266 1658
rect 58266 1606 58312 1658
rect 58016 1604 58072 1606
rect 58096 1604 58152 1606
rect 58176 1604 58232 1606
rect 58256 1604 58312 1606
rect 59616 1658 59672 1660
rect 59696 1658 59752 1660
rect 59776 1658 59832 1660
rect 59856 1658 59912 1660
rect 59616 1606 59662 1658
rect 59662 1606 59672 1658
rect 59696 1606 59726 1658
rect 59726 1606 59738 1658
rect 59738 1606 59752 1658
rect 59776 1606 59790 1658
rect 59790 1606 59802 1658
rect 59802 1606 59832 1658
rect 59856 1606 59866 1658
rect 59866 1606 59912 1658
rect 59616 1604 59672 1606
rect 59696 1604 59752 1606
rect 59776 1604 59832 1606
rect 59856 1604 59912 1606
rect 61216 1658 61272 1660
rect 61296 1658 61352 1660
rect 61376 1658 61432 1660
rect 61456 1658 61512 1660
rect 61216 1606 61262 1658
rect 61262 1606 61272 1658
rect 61296 1606 61326 1658
rect 61326 1606 61338 1658
rect 61338 1606 61352 1658
rect 61376 1606 61390 1658
rect 61390 1606 61402 1658
rect 61402 1606 61432 1658
rect 61456 1606 61466 1658
rect 61466 1606 61512 1658
rect 61216 1604 61272 1606
rect 61296 1604 61352 1606
rect 61376 1604 61432 1606
rect 61456 1604 61512 1606
rect 62816 1658 62872 1660
rect 62896 1658 62952 1660
rect 62976 1658 63032 1660
rect 63056 1658 63112 1660
rect 62816 1606 62862 1658
rect 62862 1606 62872 1658
rect 62896 1606 62926 1658
rect 62926 1606 62938 1658
rect 62938 1606 62952 1658
rect 62976 1606 62990 1658
rect 62990 1606 63002 1658
rect 63002 1606 63032 1658
rect 63056 1606 63066 1658
rect 63066 1606 63112 1658
rect 62816 1604 62872 1606
rect 62896 1604 62952 1606
rect 62976 1604 63032 1606
rect 63056 1604 63112 1606
rect 64416 1658 64472 1660
rect 64496 1658 64552 1660
rect 64576 1658 64632 1660
rect 64656 1658 64712 1660
rect 64416 1606 64462 1658
rect 64462 1606 64472 1658
rect 64496 1606 64526 1658
rect 64526 1606 64538 1658
rect 64538 1606 64552 1658
rect 64576 1606 64590 1658
rect 64590 1606 64602 1658
rect 64602 1606 64632 1658
rect 64656 1606 64666 1658
rect 64666 1606 64712 1658
rect 64416 1604 64472 1606
rect 64496 1604 64552 1606
rect 64576 1604 64632 1606
rect 64656 1604 64712 1606
rect 66016 1658 66072 1660
rect 66096 1658 66152 1660
rect 66176 1658 66232 1660
rect 66256 1658 66312 1660
rect 66016 1606 66062 1658
rect 66062 1606 66072 1658
rect 66096 1606 66126 1658
rect 66126 1606 66138 1658
rect 66138 1606 66152 1658
rect 66176 1606 66190 1658
rect 66190 1606 66202 1658
rect 66202 1606 66232 1658
rect 66256 1606 66266 1658
rect 66266 1606 66312 1658
rect 66016 1604 66072 1606
rect 66096 1604 66152 1606
rect 66176 1604 66232 1606
rect 66256 1604 66312 1606
rect 67616 1658 67672 1660
rect 67696 1658 67752 1660
rect 67776 1658 67832 1660
rect 67856 1658 67912 1660
rect 67616 1606 67662 1658
rect 67662 1606 67672 1658
rect 67696 1606 67726 1658
rect 67726 1606 67738 1658
rect 67738 1606 67752 1658
rect 67776 1606 67790 1658
rect 67790 1606 67802 1658
rect 67802 1606 67832 1658
rect 67856 1606 67866 1658
rect 67866 1606 67912 1658
rect 67616 1604 67672 1606
rect 67696 1604 67752 1606
rect 67776 1604 67832 1606
rect 67856 1604 67912 1606
rect 69216 1658 69272 1660
rect 69296 1658 69352 1660
rect 69376 1658 69432 1660
rect 69456 1658 69512 1660
rect 69216 1606 69262 1658
rect 69262 1606 69272 1658
rect 69296 1606 69326 1658
rect 69326 1606 69338 1658
rect 69338 1606 69352 1658
rect 69376 1606 69390 1658
rect 69390 1606 69402 1658
rect 69402 1606 69432 1658
rect 69456 1606 69466 1658
rect 69466 1606 69512 1658
rect 69216 1604 69272 1606
rect 69296 1604 69352 1606
rect 69376 1604 69432 1606
rect 69456 1604 69512 1606
rect 70816 1658 70872 1660
rect 70896 1658 70952 1660
rect 70976 1658 71032 1660
rect 71056 1658 71112 1660
rect 70816 1606 70862 1658
rect 70862 1606 70872 1658
rect 70896 1606 70926 1658
rect 70926 1606 70938 1658
rect 70938 1606 70952 1658
rect 70976 1606 70990 1658
rect 70990 1606 71002 1658
rect 71002 1606 71032 1658
rect 71056 1606 71066 1658
rect 71066 1606 71112 1658
rect 70816 1604 70872 1606
rect 70896 1604 70952 1606
rect 70976 1604 71032 1606
rect 71056 1604 71112 1606
rect 72416 1658 72472 1660
rect 72496 1658 72552 1660
rect 72576 1658 72632 1660
rect 72656 1658 72712 1660
rect 72416 1606 72462 1658
rect 72462 1606 72472 1658
rect 72496 1606 72526 1658
rect 72526 1606 72538 1658
rect 72538 1606 72552 1658
rect 72576 1606 72590 1658
rect 72590 1606 72602 1658
rect 72602 1606 72632 1658
rect 72656 1606 72666 1658
rect 72666 1606 72712 1658
rect 72416 1604 72472 1606
rect 72496 1604 72552 1606
rect 72576 1604 72632 1606
rect 72656 1604 72712 1606
rect 74016 1658 74072 1660
rect 74096 1658 74152 1660
rect 74176 1658 74232 1660
rect 74256 1658 74312 1660
rect 74016 1606 74062 1658
rect 74062 1606 74072 1658
rect 74096 1606 74126 1658
rect 74126 1606 74138 1658
rect 74138 1606 74152 1658
rect 74176 1606 74190 1658
rect 74190 1606 74202 1658
rect 74202 1606 74232 1658
rect 74256 1606 74266 1658
rect 74266 1606 74312 1658
rect 74016 1604 74072 1606
rect 74096 1604 74152 1606
rect 74176 1604 74232 1606
rect 74256 1604 74312 1606
rect 75616 1658 75672 1660
rect 75696 1658 75752 1660
rect 75776 1658 75832 1660
rect 75856 1658 75912 1660
rect 75616 1606 75662 1658
rect 75662 1606 75672 1658
rect 75696 1606 75726 1658
rect 75726 1606 75738 1658
rect 75738 1606 75752 1658
rect 75776 1606 75790 1658
rect 75790 1606 75802 1658
rect 75802 1606 75832 1658
rect 75856 1606 75866 1658
rect 75866 1606 75912 1658
rect 75616 1604 75672 1606
rect 75696 1604 75752 1606
rect 75776 1604 75832 1606
rect 75856 1604 75912 1606
rect 77216 1658 77272 1660
rect 77296 1658 77352 1660
rect 77376 1658 77432 1660
rect 77456 1658 77512 1660
rect 77216 1606 77262 1658
rect 77262 1606 77272 1658
rect 77296 1606 77326 1658
rect 77326 1606 77338 1658
rect 77338 1606 77352 1658
rect 77376 1606 77390 1658
rect 77390 1606 77402 1658
rect 77402 1606 77432 1658
rect 77456 1606 77466 1658
rect 77466 1606 77512 1658
rect 77216 1604 77272 1606
rect 77296 1604 77352 1606
rect 77376 1604 77432 1606
rect 77456 1604 77512 1606
rect 78816 1658 78872 1660
rect 78896 1658 78952 1660
rect 78976 1658 79032 1660
rect 79056 1658 79112 1660
rect 78816 1606 78862 1658
rect 78862 1606 78872 1658
rect 78896 1606 78926 1658
rect 78926 1606 78938 1658
rect 78938 1606 78952 1658
rect 78976 1606 78990 1658
rect 78990 1606 79002 1658
rect 79002 1606 79032 1658
rect 79056 1606 79066 1658
rect 79066 1606 79112 1658
rect 78816 1604 78872 1606
rect 78896 1604 78952 1606
rect 78976 1604 79032 1606
rect 79056 1604 79112 1606
rect 80416 1658 80472 1660
rect 80496 1658 80552 1660
rect 80576 1658 80632 1660
rect 80656 1658 80712 1660
rect 80416 1606 80462 1658
rect 80462 1606 80472 1658
rect 80496 1606 80526 1658
rect 80526 1606 80538 1658
rect 80538 1606 80552 1658
rect 80576 1606 80590 1658
rect 80590 1606 80602 1658
rect 80602 1606 80632 1658
rect 80656 1606 80666 1658
rect 80666 1606 80712 1658
rect 80416 1604 80472 1606
rect 80496 1604 80552 1606
rect 80576 1604 80632 1606
rect 80656 1604 80712 1606
rect 82016 1658 82072 1660
rect 82096 1658 82152 1660
rect 82176 1658 82232 1660
rect 82256 1658 82312 1660
rect 82016 1606 82062 1658
rect 82062 1606 82072 1658
rect 82096 1606 82126 1658
rect 82126 1606 82138 1658
rect 82138 1606 82152 1658
rect 82176 1606 82190 1658
rect 82190 1606 82202 1658
rect 82202 1606 82232 1658
rect 82256 1606 82266 1658
rect 82266 1606 82312 1658
rect 82016 1604 82072 1606
rect 82096 1604 82152 1606
rect 82176 1604 82232 1606
rect 82256 1604 82312 1606
rect 83616 1658 83672 1660
rect 83696 1658 83752 1660
rect 83776 1658 83832 1660
rect 83856 1658 83912 1660
rect 83616 1606 83662 1658
rect 83662 1606 83672 1658
rect 83696 1606 83726 1658
rect 83726 1606 83738 1658
rect 83738 1606 83752 1658
rect 83776 1606 83790 1658
rect 83790 1606 83802 1658
rect 83802 1606 83832 1658
rect 83856 1606 83866 1658
rect 83866 1606 83912 1658
rect 83616 1604 83672 1606
rect 83696 1604 83752 1606
rect 83776 1604 83832 1606
rect 83856 1604 83912 1606
rect 85216 1658 85272 1660
rect 85296 1658 85352 1660
rect 85376 1658 85432 1660
rect 85456 1658 85512 1660
rect 85216 1606 85262 1658
rect 85262 1606 85272 1658
rect 85296 1606 85326 1658
rect 85326 1606 85338 1658
rect 85338 1606 85352 1658
rect 85376 1606 85390 1658
rect 85390 1606 85402 1658
rect 85402 1606 85432 1658
rect 85456 1606 85466 1658
rect 85466 1606 85512 1658
rect 85216 1604 85272 1606
rect 85296 1604 85352 1606
rect 85376 1604 85432 1606
rect 85456 1604 85512 1606
rect 86816 1658 86872 1660
rect 86896 1658 86952 1660
rect 86976 1658 87032 1660
rect 87056 1658 87112 1660
rect 86816 1606 86862 1658
rect 86862 1606 86872 1658
rect 86896 1606 86926 1658
rect 86926 1606 86938 1658
rect 86938 1606 86952 1658
rect 86976 1606 86990 1658
rect 86990 1606 87002 1658
rect 87002 1606 87032 1658
rect 87056 1606 87066 1658
rect 87066 1606 87112 1658
rect 86816 1604 86872 1606
rect 86896 1604 86952 1606
rect 86976 1604 87032 1606
rect 87056 1604 87112 1606
rect 88416 1658 88472 1660
rect 88496 1658 88552 1660
rect 88576 1658 88632 1660
rect 88656 1658 88712 1660
rect 88416 1606 88462 1658
rect 88462 1606 88472 1658
rect 88496 1606 88526 1658
rect 88526 1606 88538 1658
rect 88538 1606 88552 1658
rect 88576 1606 88590 1658
rect 88590 1606 88602 1658
rect 88602 1606 88632 1658
rect 88656 1606 88666 1658
rect 88666 1606 88712 1658
rect 88416 1604 88472 1606
rect 88496 1604 88552 1606
rect 88576 1604 88632 1606
rect 88656 1604 88712 1606
rect 90016 1658 90072 1660
rect 90096 1658 90152 1660
rect 90176 1658 90232 1660
rect 90256 1658 90312 1660
rect 90016 1606 90062 1658
rect 90062 1606 90072 1658
rect 90096 1606 90126 1658
rect 90126 1606 90138 1658
rect 90138 1606 90152 1658
rect 90176 1606 90190 1658
rect 90190 1606 90202 1658
rect 90202 1606 90232 1658
rect 90256 1606 90266 1658
rect 90266 1606 90312 1658
rect 90016 1604 90072 1606
rect 90096 1604 90152 1606
rect 90176 1604 90232 1606
rect 90256 1604 90312 1606
rect 91616 1658 91672 1660
rect 91696 1658 91752 1660
rect 91776 1658 91832 1660
rect 91856 1658 91912 1660
rect 91616 1606 91662 1658
rect 91662 1606 91672 1658
rect 91696 1606 91726 1658
rect 91726 1606 91738 1658
rect 91738 1606 91752 1658
rect 91776 1606 91790 1658
rect 91790 1606 91802 1658
rect 91802 1606 91832 1658
rect 91856 1606 91866 1658
rect 91866 1606 91912 1658
rect 91616 1604 91672 1606
rect 91696 1604 91752 1606
rect 91776 1604 91832 1606
rect 91856 1604 91912 1606
rect 93216 1658 93272 1660
rect 93296 1658 93352 1660
rect 93376 1658 93432 1660
rect 93456 1658 93512 1660
rect 93216 1606 93262 1658
rect 93262 1606 93272 1658
rect 93296 1606 93326 1658
rect 93326 1606 93338 1658
rect 93338 1606 93352 1658
rect 93376 1606 93390 1658
rect 93390 1606 93402 1658
rect 93402 1606 93432 1658
rect 93456 1606 93466 1658
rect 93466 1606 93512 1658
rect 93216 1604 93272 1606
rect 93296 1604 93352 1606
rect 93376 1604 93432 1606
rect 93456 1604 93512 1606
rect 94816 1658 94872 1660
rect 94896 1658 94952 1660
rect 94976 1658 95032 1660
rect 95056 1658 95112 1660
rect 94816 1606 94862 1658
rect 94862 1606 94872 1658
rect 94896 1606 94926 1658
rect 94926 1606 94938 1658
rect 94938 1606 94952 1658
rect 94976 1606 94990 1658
rect 94990 1606 95002 1658
rect 95002 1606 95032 1658
rect 95056 1606 95066 1658
rect 95066 1606 95112 1658
rect 94816 1604 94872 1606
rect 94896 1604 94952 1606
rect 94976 1604 95032 1606
rect 95056 1604 95112 1606
rect 96416 1658 96472 1660
rect 96496 1658 96552 1660
rect 96576 1658 96632 1660
rect 96656 1658 96712 1660
rect 96416 1606 96462 1658
rect 96462 1606 96472 1658
rect 96496 1606 96526 1658
rect 96526 1606 96538 1658
rect 96538 1606 96552 1658
rect 96576 1606 96590 1658
rect 96590 1606 96602 1658
rect 96602 1606 96632 1658
rect 96656 1606 96666 1658
rect 96666 1606 96712 1658
rect 96416 1604 96472 1606
rect 96496 1604 96552 1606
rect 96576 1604 96632 1606
rect 96656 1604 96712 1606
rect 98016 1658 98072 1660
rect 98096 1658 98152 1660
rect 98176 1658 98232 1660
rect 98256 1658 98312 1660
rect 98016 1606 98062 1658
rect 98062 1606 98072 1658
rect 98096 1606 98126 1658
rect 98126 1606 98138 1658
rect 98138 1606 98152 1658
rect 98176 1606 98190 1658
rect 98190 1606 98202 1658
rect 98202 1606 98232 1658
rect 98256 1606 98266 1658
rect 98266 1606 98312 1658
rect 98016 1604 98072 1606
rect 98096 1604 98152 1606
rect 98176 1604 98232 1606
rect 98256 1604 98312 1606
rect 99616 1658 99672 1660
rect 99696 1658 99752 1660
rect 99776 1658 99832 1660
rect 99856 1658 99912 1660
rect 99616 1606 99662 1658
rect 99662 1606 99672 1658
rect 99696 1606 99726 1658
rect 99726 1606 99738 1658
rect 99738 1606 99752 1658
rect 99776 1606 99790 1658
rect 99790 1606 99802 1658
rect 99802 1606 99832 1658
rect 99856 1606 99866 1658
rect 99866 1606 99912 1658
rect 99616 1604 99672 1606
rect 99696 1604 99752 1606
rect 99776 1604 99832 1606
rect 99856 1604 99912 1606
rect 101216 1658 101272 1660
rect 101296 1658 101352 1660
rect 101376 1658 101432 1660
rect 101456 1658 101512 1660
rect 101216 1606 101262 1658
rect 101262 1606 101272 1658
rect 101296 1606 101326 1658
rect 101326 1606 101338 1658
rect 101338 1606 101352 1658
rect 101376 1606 101390 1658
rect 101390 1606 101402 1658
rect 101402 1606 101432 1658
rect 101456 1606 101466 1658
rect 101466 1606 101512 1658
rect 101216 1604 101272 1606
rect 101296 1604 101352 1606
rect 101376 1604 101432 1606
rect 101456 1604 101512 1606
rect 102816 1658 102872 1660
rect 102896 1658 102952 1660
rect 102976 1658 103032 1660
rect 103056 1658 103112 1660
rect 102816 1606 102862 1658
rect 102862 1606 102872 1658
rect 102896 1606 102926 1658
rect 102926 1606 102938 1658
rect 102938 1606 102952 1658
rect 102976 1606 102990 1658
rect 102990 1606 103002 1658
rect 103002 1606 103032 1658
rect 103056 1606 103066 1658
rect 103066 1606 103112 1658
rect 102816 1604 102872 1606
rect 102896 1604 102952 1606
rect 102976 1604 103032 1606
rect 103056 1604 103112 1606
rect 104416 1658 104472 1660
rect 104496 1658 104552 1660
rect 104576 1658 104632 1660
rect 104656 1658 104712 1660
rect 104416 1606 104462 1658
rect 104462 1606 104472 1658
rect 104496 1606 104526 1658
rect 104526 1606 104538 1658
rect 104538 1606 104552 1658
rect 104576 1606 104590 1658
rect 104590 1606 104602 1658
rect 104602 1606 104632 1658
rect 104656 1606 104666 1658
rect 104666 1606 104712 1658
rect 104416 1604 104472 1606
rect 104496 1604 104552 1606
rect 104576 1604 104632 1606
rect 104656 1604 104712 1606
rect 106016 1658 106072 1660
rect 106096 1658 106152 1660
rect 106176 1658 106232 1660
rect 106256 1658 106312 1660
rect 106016 1606 106062 1658
rect 106062 1606 106072 1658
rect 106096 1606 106126 1658
rect 106126 1606 106138 1658
rect 106138 1606 106152 1658
rect 106176 1606 106190 1658
rect 106190 1606 106202 1658
rect 106202 1606 106232 1658
rect 106256 1606 106266 1658
rect 106266 1606 106312 1658
rect 106016 1604 106072 1606
rect 106096 1604 106152 1606
rect 106176 1604 106232 1606
rect 106256 1604 106312 1606
rect 107616 1658 107672 1660
rect 107696 1658 107752 1660
rect 107776 1658 107832 1660
rect 107856 1658 107912 1660
rect 107616 1606 107662 1658
rect 107662 1606 107672 1658
rect 107696 1606 107726 1658
rect 107726 1606 107738 1658
rect 107738 1606 107752 1658
rect 107776 1606 107790 1658
rect 107790 1606 107802 1658
rect 107802 1606 107832 1658
rect 107856 1606 107866 1658
rect 107866 1606 107912 1658
rect 107616 1604 107672 1606
rect 107696 1604 107752 1606
rect 107776 1604 107832 1606
rect 107856 1604 107912 1606
rect 56598 1264 56654 1320
rect 57978 1264 58034 1320
rect 59358 1284 59414 1320
rect 59358 1264 59360 1284
rect 59360 1264 59412 1284
rect 59412 1264 59414 1284
rect 55756 1114 55812 1116
rect 55836 1114 55892 1116
rect 55916 1114 55972 1116
rect 55996 1114 56052 1116
rect 55756 1062 55802 1114
rect 55802 1062 55812 1114
rect 55836 1062 55866 1114
rect 55866 1062 55878 1114
rect 55878 1062 55892 1114
rect 55916 1062 55930 1114
rect 55930 1062 55942 1114
rect 55942 1062 55972 1114
rect 55996 1062 56006 1114
rect 56006 1062 56052 1114
rect 55756 1060 55812 1062
rect 55836 1060 55892 1062
rect 55916 1060 55972 1062
rect 55996 1060 56052 1062
rect 57356 1114 57412 1116
rect 57436 1114 57492 1116
rect 57516 1114 57572 1116
rect 57596 1114 57652 1116
rect 57356 1062 57402 1114
rect 57402 1062 57412 1114
rect 57436 1062 57466 1114
rect 57466 1062 57478 1114
rect 57478 1062 57492 1114
rect 57516 1062 57530 1114
rect 57530 1062 57542 1114
rect 57542 1062 57572 1114
rect 57596 1062 57606 1114
rect 57606 1062 57652 1114
rect 57356 1060 57412 1062
rect 57436 1060 57492 1062
rect 57516 1060 57572 1062
rect 57596 1060 57652 1062
rect 60922 1264 60978 1320
rect 62486 1264 62542 1320
rect 63498 1264 63554 1320
rect 64878 1264 64934 1320
rect 65154 1264 65210 1320
rect 66258 1264 66314 1320
rect 67638 1264 67694 1320
rect 69018 1264 69074 1320
rect 58956 1114 59012 1116
rect 59036 1114 59092 1116
rect 59116 1114 59172 1116
rect 59196 1114 59252 1116
rect 58956 1062 59002 1114
rect 59002 1062 59012 1114
rect 59036 1062 59066 1114
rect 59066 1062 59078 1114
rect 59078 1062 59092 1114
rect 59116 1062 59130 1114
rect 59130 1062 59142 1114
rect 59142 1062 59172 1114
rect 59196 1062 59206 1114
rect 59206 1062 59252 1114
rect 58956 1060 59012 1062
rect 59036 1060 59092 1062
rect 59116 1060 59172 1062
rect 59196 1060 59252 1062
rect 60556 1114 60612 1116
rect 60636 1114 60692 1116
rect 60716 1114 60772 1116
rect 60796 1114 60852 1116
rect 60556 1062 60602 1114
rect 60602 1062 60612 1114
rect 60636 1062 60666 1114
rect 60666 1062 60678 1114
rect 60678 1062 60692 1114
rect 60716 1062 60730 1114
rect 60730 1062 60742 1114
rect 60742 1062 60772 1114
rect 60796 1062 60806 1114
rect 60806 1062 60852 1114
rect 60556 1060 60612 1062
rect 60636 1060 60692 1062
rect 60716 1060 60772 1062
rect 60796 1060 60852 1062
rect 62156 1114 62212 1116
rect 62236 1114 62292 1116
rect 62316 1114 62372 1116
rect 62396 1114 62452 1116
rect 62156 1062 62202 1114
rect 62202 1062 62212 1114
rect 62236 1062 62266 1114
rect 62266 1062 62278 1114
rect 62278 1062 62292 1114
rect 62316 1062 62330 1114
rect 62330 1062 62342 1114
rect 62342 1062 62372 1114
rect 62396 1062 62406 1114
rect 62406 1062 62452 1114
rect 62156 1060 62212 1062
rect 62236 1060 62292 1062
rect 62316 1060 62372 1062
rect 62396 1060 62452 1062
rect 63756 1114 63812 1116
rect 63836 1114 63892 1116
rect 63916 1114 63972 1116
rect 63996 1114 64052 1116
rect 63756 1062 63802 1114
rect 63802 1062 63812 1114
rect 63836 1062 63866 1114
rect 63866 1062 63878 1114
rect 63878 1062 63892 1114
rect 63916 1062 63930 1114
rect 63930 1062 63942 1114
rect 63942 1062 63972 1114
rect 63996 1062 64006 1114
rect 64006 1062 64052 1114
rect 63756 1060 63812 1062
rect 63836 1060 63892 1062
rect 63916 1060 63972 1062
rect 63996 1060 64052 1062
rect 65356 1114 65412 1116
rect 65436 1114 65492 1116
rect 65516 1114 65572 1116
rect 65596 1114 65652 1116
rect 65356 1062 65402 1114
rect 65402 1062 65412 1114
rect 65436 1062 65466 1114
rect 65466 1062 65478 1114
rect 65478 1062 65492 1114
rect 65516 1062 65530 1114
rect 65530 1062 65542 1114
rect 65542 1062 65572 1114
rect 65596 1062 65606 1114
rect 65606 1062 65652 1114
rect 65356 1060 65412 1062
rect 65436 1060 65492 1062
rect 65516 1060 65572 1062
rect 65596 1060 65652 1062
rect 66956 1114 67012 1116
rect 67036 1114 67092 1116
rect 67116 1114 67172 1116
rect 67196 1114 67252 1116
rect 66956 1062 67002 1114
rect 67002 1062 67012 1114
rect 67036 1062 67066 1114
rect 67066 1062 67078 1114
rect 67078 1062 67092 1114
rect 67116 1062 67130 1114
rect 67130 1062 67142 1114
rect 67142 1062 67172 1114
rect 67196 1062 67206 1114
rect 67206 1062 67252 1114
rect 66956 1060 67012 1062
rect 67036 1060 67092 1062
rect 67116 1060 67172 1062
rect 67196 1060 67252 1062
rect 68556 1114 68612 1116
rect 68636 1114 68692 1116
rect 68716 1114 68772 1116
rect 68796 1114 68852 1116
rect 68556 1062 68602 1114
rect 68602 1062 68612 1114
rect 68636 1062 68666 1114
rect 68666 1062 68678 1114
rect 68678 1062 68692 1114
rect 68716 1062 68730 1114
rect 68730 1062 68742 1114
rect 68742 1062 68772 1114
rect 68796 1062 68806 1114
rect 68806 1062 68852 1114
rect 68556 1060 68612 1062
rect 68636 1060 68692 1062
rect 68716 1060 68772 1062
rect 68796 1060 68852 1062
rect 70156 1114 70212 1116
rect 70236 1114 70292 1116
rect 70316 1114 70372 1116
rect 70396 1114 70452 1116
rect 70156 1062 70202 1114
rect 70202 1062 70212 1114
rect 70236 1062 70266 1114
rect 70266 1062 70278 1114
rect 70278 1062 70292 1114
rect 70316 1062 70330 1114
rect 70330 1062 70342 1114
rect 70342 1062 70372 1114
rect 70396 1062 70406 1114
rect 70406 1062 70452 1114
rect 70156 1060 70212 1062
rect 70236 1060 70292 1062
rect 70316 1060 70372 1062
rect 70396 1060 70452 1062
rect 71756 1114 71812 1116
rect 71836 1114 71892 1116
rect 71916 1114 71972 1116
rect 71996 1114 72052 1116
rect 71756 1062 71802 1114
rect 71802 1062 71812 1114
rect 71836 1062 71866 1114
rect 71866 1062 71878 1114
rect 71878 1062 71892 1114
rect 71916 1062 71930 1114
rect 71930 1062 71942 1114
rect 71942 1062 71972 1114
rect 71996 1062 72006 1114
rect 72006 1062 72052 1114
rect 71756 1060 71812 1062
rect 71836 1060 71892 1062
rect 71916 1060 71972 1062
rect 71996 1060 72052 1062
rect 73356 1114 73412 1116
rect 73436 1114 73492 1116
rect 73516 1114 73572 1116
rect 73596 1114 73652 1116
rect 73356 1062 73402 1114
rect 73402 1062 73412 1114
rect 73436 1062 73466 1114
rect 73466 1062 73478 1114
rect 73478 1062 73492 1114
rect 73516 1062 73530 1114
rect 73530 1062 73542 1114
rect 73542 1062 73572 1114
rect 73596 1062 73606 1114
rect 73606 1062 73652 1114
rect 73356 1060 73412 1062
rect 73436 1060 73492 1062
rect 73516 1060 73572 1062
rect 73596 1060 73652 1062
rect 74956 1114 75012 1116
rect 75036 1114 75092 1116
rect 75116 1114 75172 1116
rect 75196 1114 75252 1116
rect 74956 1062 75002 1114
rect 75002 1062 75012 1114
rect 75036 1062 75066 1114
rect 75066 1062 75078 1114
rect 75078 1062 75092 1114
rect 75116 1062 75130 1114
rect 75130 1062 75142 1114
rect 75142 1062 75172 1114
rect 75196 1062 75206 1114
rect 75206 1062 75252 1114
rect 74956 1060 75012 1062
rect 75036 1060 75092 1062
rect 75116 1060 75172 1062
rect 75196 1060 75252 1062
rect 76556 1114 76612 1116
rect 76636 1114 76692 1116
rect 76716 1114 76772 1116
rect 76796 1114 76852 1116
rect 76556 1062 76602 1114
rect 76602 1062 76612 1114
rect 76636 1062 76666 1114
rect 76666 1062 76678 1114
rect 76678 1062 76692 1114
rect 76716 1062 76730 1114
rect 76730 1062 76742 1114
rect 76742 1062 76772 1114
rect 76796 1062 76806 1114
rect 76806 1062 76852 1114
rect 76556 1060 76612 1062
rect 76636 1060 76692 1062
rect 76716 1060 76772 1062
rect 76796 1060 76852 1062
rect 78156 1114 78212 1116
rect 78236 1114 78292 1116
rect 78316 1114 78372 1116
rect 78396 1114 78452 1116
rect 78156 1062 78202 1114
rect 78202 1062 78212 1114
rect 78236 1062 78266 1114
rect 78266 1062 78278 1114
rect 78278 1062 78292 1114
rect 78316 1062 78330 1114
rect 78330 1062 78342 1114
rect 78342 1062 78372 1114
rect 78396 1062 78406 1114
rect 78406 1062 78452 1114
rect 78156 1060 78212 1062
rect 78236 1060 78292 1062
rect 78316 1060 78372 1062
rect 78396 1060 78452 1062
rect 79756 1114 79812 1116
rect 79836 1114 79892 1116
rect 79916 1114 79972 1116
rect 79996 1114 80052 1116
rect 79756 1062 79802 1114
rect 79802 1062 79812 1114
rect 79836 1062 79866 1114
rect 79866 1062 79878 1114
rect 79878 1062 79892 1114
rect 79916 1062 79930 1114
rect 79930 1062 79942 1114
rect 79942 1062 79972 1114
rect 79996 1062 80006 1114
rect 80006 1062 80052 1114
rect 79756 1060 79812 1062
rect 79836 1060 79892 1062
rect 79916 1060 79972 1062
rect 79996 1060 80052 1062
rect 81356 1114 81412 1116
rect 81436 1114 81492 1116
rect 81516 1114 81572 1116
rect 81596 1114 81652 1116
rect 81356 1062 81402 1114
rect 81402 1062 81412 1114
rect 81436 1062 81466 1114
rect 81466 1062 81478 1114
rect 81478 1062 81492 1114
rect 81516 1062 81530 1114
rect 81530 1062 81542 1114
rect 81542 1062 81572 1114
rect 81596 1062 81606 1114
rect 81606 1062 81652 1114
rect 81356 1060 81412 1062
rect 81436 1060 81492 1062
rect 81516 1060 81572 1062
rect 81596 1060 81652 1062
rect 82956 1114 83012 1116
rect 83036 1114 83092 1116
rect 83116 1114 83172 1116
rect 83196 1114 83252 1116
rect 82956 1062 83002 1114
rect 83002 1062 83012 1114
rect 83036 1062 83066 1114
rect 83066 1062 83078 1114
rect 83078 1062 83092 1114
rect 83116 1062 83130 1114
rect 83130 1062 83142 1114
rect 83142 1062 83172 1114
rect 83196 1062 83206 1114
rect 83206 1062 83252 1114
rect 82956 1060 83012 1062
rect 83036 1060 83092 1062
rect 83116 1060 83172 1062
rect 83196 1060 83252 1062
rect 84556 1114 84612 1116
rect 84636 1114 84692 1116
rect 84716 1114 84772 1116
rect 84796 1114 84852 1116
rect 84556 1062 84602 1114
rect 84602 1062 84612 1114
rect 84636 1062 84666 1114
rect 84666 1062 84678 1114
rect 84678 1062 84692 1114
rect 84716 1062 84730 1114
rect 84730 1062 84742 1114
rect 84742 1062 84772 1114
rect 84796 1062 84806 1114
rect 84806 1062 84852 1114
rect 84556 1060 84612 1062
rect 84636 1060 84692 1062
rect 84716 1060 84772 1062
rect 84796 1060 84852 1062
rect 86156 1114 86212 1116
rect 86236 1114 86292 1116
rect 86316 1114 86372 1116
rect 86396 1114 86452 1116
rect 86156 1062 86202 1114
rect 86202 1062 86212 1114
rect 86236 1062 86266 1114
rect 86266 1062 86278 1114
rect 86278 1062 86292 1114
rect 86316 1062 86330 1114
rect 86330 1062 86342 1114
rect 86342 1062 86372 1114
rect 86396 1062 86406 1114
rect 86406 1062 86452 1114
rect 86156 1060 86212 1062
rect 86236 1060 86292 1062
rect 86316 1060 86372 1062
rect 86396 1060 86452 1062
rect 87756 1114 87812 1116
rect 87836 1114 87892 1116
rect 87916 1114 87972 1116
rect 87996 1114 88052 1116
rect 87756 1062 87802 1114
rect 87802 1062 87812 1114
rect 87836 1062 87866 1114
rect 87866 1062 87878 1114
rect 87878 1062 87892 1114
rect 87916 1062 87930 1114
rect 87930 1062 87942 1114
rect 87942 1062 87972 1114
rect 87996 1062 88006 1114
rect 88006 1062 88052 1114
rect 87756 1060 87812 1062
rect 87836 1060 87892 1062
rect 87916 1060 87972 1062
rect 87996 1060 88052 1062
rect 89356 1114 89412 1116
rect 89436 1114 89492 1116
rect 89516 1114 89572 1116
rect 89596 1114 89652 1116
rect 89356 1062 89402 1114
rect 89402 1062 89412 1114
rect 89436 1062 89466 1114
rect 89466 1062 89478 1114
rect 89478 1062 89492 1114
rect 89516 1062 89530 1114
rect 89530 1062 89542 1114
rect 89542 1062 89572 1114
rect 89596 1062 89606 1114
rect 89606 1062 89652 1114
rect 89356 1060 89412 1062
rect 89436 1060 89492 1062
rect 89516 1060 89572 1062
rect 89596 1060 89652 1062
rect 90956 1114 91012 1116
rect 91036 1114 91092 1116
rect 91116 1114 91172 1116
rect 91196 1114 91252 1116
rect 90956 1062 91002 1114
rect 91002 1062 91012 1114
rect 91036 1062 91066 1114
rect 91066 1062 91078 1114
rect 91078 1062 91092 1114
rect 91116 1062 91130 1114
rect 91130 1062 91142 1114
rect 91142 1062 91172 1114
rect 91196 1062 91206 1114
rect 91206 1062 91252 1114
rect 90956 1060 91012 1062
rect 91036 1060 91092 1062
rect 91116 1060 91172 1062
rect 91196 1060 91252 1062
rect 92556 1114 92612 1116
rect 92636 1114 92692 1116
rect 92716 1114 92772 1116
rect 92796 1114 92852 1116
rect 92556 1062 92602 1114
rect 92602 1062 92612 1114
rect 92636 1062 92666 1114
rect 92666 1062 92678 1114
rect 92678 1062 92692 1114
rect 92716 1062 92730 1114
rect 92730 1062 92742 1114
rect 92742 1062 92772 1114
rect 92796 1062 92806 1114
rect 92806 1062 92852 1114
rect 92556 1060 92612 1062
rect 92636 1060 92692 1062
rect 92716 1060 92772 1062
rect 92796 1060 92852 1062
rect 94156 1114 94212 1116
rect 94236 1114 94292 1116
rect 94316 1114 94372 1116
rect 94396 1114 94452 1116
rect 94156 1062 94202 1114
rect 94202 1062 94212 1114
rect 94236 1062 94266 1114
rect 94266 1062 94278 1114
rect 94278 1062 94292 1114
rect 94316 1062 94330 1114
rect 94330 1062 94342 1114
rect 94342 1062 94372 1114
rect 94396 1062 94406 1114
rect 94406 1062 94452 1114
rect 94156 1060 94212 1062
rect 94236 1060 94292 1062
rect 94316 1060 94372 1062
rect 94396 1060 94452 1062
rect 95756 1114 95812 1116
rect 95836 1114 95892 1116
rect 95916 1114 95972 1116
rect 95996 1114 96052 1116
rect 95756 1062 95802 1114
rect 95802 1062 95812 1114
rect 95836 1062 95866 1114
rect 95866 1062 95878 1114
rect 95878 1062 95892 1114
rect 95916 1062 95930 1114
rect 95930 1062 95942 1114
rect 95942 1062 95972 1114
rect 95996 1062 96006 1114
rect 96006 1062 96052 1114
rect 95756 1060 95812 1062
rect 95836 1060 95892 1062
rect 95916 1060 95972 1062
rect 95996 1060 96052 1062
rect 97356 1114 97412 1116
rect 97436 1114 97492 1116
rect 97516 1114 97572 1116
rect 97596 1114 97652 1116
rect 97356 1062 97402 1114
rect 97402 1062 97412 1114
rect 97436 1062 97466 1114
rect 97466 1062 97478 1114
rect 97478 1062 97492 1114
rect 97516 1062 97530 1114
rect 97530 1062 97542 1114
rect 97542 1062 97572 1114
rect 97596 1062 97606 1114
rect 97606 1062 97652 1114
rect 97356 1060 97412 1062
rect 97436 1060 97492 1062
rect 97516 1060 97572 1062
rect 97596 1060 97652 1062
rect 98956 1114 99012 1116
rect 99036 1114 99092 1116
rect 99116 1114 99172 1116
rect 99196 1114 99252 1116
rect 98956 1062 99002 1114
rect 99002 1062 99012 1114
rect 99036 1062 99066 1114
rect 99066 1062 99078 1114
rect 99078 1062 99092 1114
rect 99116 1062 99130 1114
rect 99130 1062 99142 1114
rect 99142 1062 99172 1114
rect 99196 1062 99206 1114
rect 99206 1062 99252 1114
rect 98956 1060 99012 1062
rect 99036 1060 99092 1062
rect 99116 1060 99172 1062
rect 99196 1060 99252 1062
rect 100556 1114 100612 1116
rect 100636 1114 100692 1116
rect 100716 1114 100772 1116
rect 100796 1114 100852 1116
rect 100556 1062 100602 1114
rect 100602 1062 100612 1114
rect 100636 1062 100666 1114
rect 100666 1062 100678 1114
rect 100678 1062 100692 1114
rect 100716 1062 100730 1114
rect 100730 1062 100742 1114
rect 100742 1062 100772 1114
rect 100796 1062 100806 1114
rect 100806 1062 100852 1114
rect 100556 1060 100612 1062
rect 100636 1060 100692 1062
rect 100716 1060 100772 1062
rect 100796 1060 100852 1062
rect 102156 1114 102212 1116
rect 102236 1114 102292 1116
rect 102316 1114 102372 1116
rect 102396 1114 102452 1116
rect 102156 1062 102202 1114
rect 102202 1062 102212 1114
rect 102236 1062 102266 1114
rect 102266 1062 102278 1114
rect 102278 1062 102292 1114
rect 102316 1062 102330 1114
rect 102330 1062 102342 1114
rect 102342 1062 102372 1114
rect 102396 1062 102406 1114
rect 102406 1062 102452 1114
rect 102156 1060 102212 1062
rect 102236 1060 102292 1062
rect 102316 1060 102372 1062
rect 102396 1060 102452 1062
rect 103756 1114 103812 1116
rect 103836 1114 103892 1116
rect 103916 1114 103972 1116
rect 103996 1114 104052 1116
rect 103756 1062 103802 1114
rect 103802 1062 103812 1114
rect 103836 1062 103866 1114
rect 103866 1062 103878 1114
rect 103878 1062 103892 1114
rect 103916 1062 103930 1114
rect 103930 1062 103942 1114
rect 103942 1062 103972 1114
rect 103996 1062 104006 1114
rect 104006 1062 104052 1114
rect 103756 1060 103812 1062
rect 103836 1060 103892 1062
rect 103916 1060 103972 1062
rect 103996 1060 104052 1062
rect 105356 1114 105412 1116
rect 105436 1114 105492 1116
rect 105516 1114 105572 1116
rect 105596 1114 105652 1116
rect 105356 1062 105402 1114
rect 105402 1062 105412 1114
rect 105436 1062 105466 1114
rect 105466 1062 105478 1114
rect 105478 1062 105492 1114
rect 105516 1062 105530 1114
rect 105530 1062 105542 1114
rect 105542 1062 105572 1114
rect 105596 1062 105606 1114
rect 105606 1062 105652 1114
rect 105356 1060 105412 1062
rect 105436 1060 105492 1062
rect 105516 1060 105572 1062
rect 105596 1060 105652 1062
rect 106956 1114 107012 1116
rect 107036 1114 107092 1116
rect 107116 1114 107172 1116
rect 107196 1114 107252 1116
rect 106956 1062 107002 1114
rect 107002 1062 107012 1114
rect 107036 1062 107066 1114
rect 107066 1062 107078 1114
rect 107078 1062 107092 1114
rect 107116 1062 107130 1114
rect 107130 1062 107142 1114
rect 107142 1062 107172 1114
rect 107196 1062 107206 1114
rect 107206 1062 107252 1114
rect 106956 1060 107012 1062
rect 107036 1060 107092 1062
rect 107116 1060 107172 1062
rect 107196 1060 107252 1062
rect 108556 1114 108612 1116
rect 108636 1114 108692 1116
rect 108716 1114 108772 1116
rect 108796 1114 108852 1116
rect 108556 1062 108602 1114
rect 108602 1062 108612 1114
rect 108636 1062 108666 1114
rect 108666 1062 108678 1114
rect 108678 1062 108692 1114
rect 108716 1062 108730 1114
rect 108730 1062 108742 1114
rect 108742 1062 108772 1114
rect 108796 1062 108806 1114
rect 108806 1062 108852 1114
rect 108556 1060 108612 1062
rect 108636 1060 108692 1062
rect 108716 1060 108772 1062
rect 108796 1060 108852 1062
<< metal3 >>
rect 3606 86528 3922 86529
rect 3606 86464 3612 86528
rect 3676 86464 3692 86528
rect 3756 86464 3772 86528
rect 3836 86464 3852 86528
rect 3916 86464 3922 86528
rect 3606 86463 3922 86464
rect 5206 86528 5522 86529
rect 5206 86464 5212 86528
rect 5276 86464 5292 86528
rect 5356 86464 5372 86528
rect 5436 86464 5452 86528
rect 5516 86464 5522 86528
rect 5206 86463 5522 86464
rect 6806 86528 7122 86529
rect 6806 86464 6812 86528
rect 6876 86464 6892 86528
rect 6956 86464 6972 86528
rect 7036 86464 7052 86528
rect 7116 86464 7122 86528
rect 6806 86463 7122 86464
rect 8406 86528 8722 86529
rect 8406 86464 8412 86528
rect 8476 86464 8492 86528
rect 8556 86464 8572 86528
rect 8636 86464 8652 86528
rect 8716 86464 8722 86528
rect 8406 86463 8722 86464
rect 10006 86528 10322 86529
rect 10006 86464 10012 86528
rect 10076 86464 10092 86528
rect 10156 86464 10172 86528
rect 10236 86464 10252 86528
rect 10316 86464 10322 86528
rect 10006 86463 10322 86464
rect 11606 86528 11922 86529
rect 11606 86464 11612 86528
rect 11676 86464 11692 86528
rect 11756 86464 11772 86528
rect 11836 86464 11852 86528
rect 11916 86464 11922 86528
rect 11606 86463 11922 86464
rect 13206 86528 13522 86529
rect 13206 86464 13212 86528
rect 13276 86464 13292 86528
rect 13356 86464 13372 86528
rect 13436 86464 13452 86528
rect 13516 86464 13522 86528
rect 13206 86463 13522 86464
rect 14806 86528 15122 86529
rect 14806 86464 14812 86528
rect 14876 86464 14892 86528
rect 14956 86464 14972 86528
rect 15036 86464 15052 86528
rect 15116 86464 15122 86528
rect 14806 86463 15122 86464
rect 16406 86528 16722 86529
rect 16406 86464 16412 86528
rect 16476 86464 16492 86528
rect 16556 86464 16572 86528
rect 16636 86464 16652 86528
rect 16716 86464 16722 86528
rect 16406 86463 16722 86464
rect 18006 86528 18322 86529
rect 18006 86464 18012 86528
rect 18076 86464 18092 86528
rect 18156 86464 18172 86528
rect 18236 86464 18252 86528
rect 18316 86464 18322 86528
rect 18006 86463 18322 86464
rect 19606 86528 19922 86529
rect 19606 86464 19612 86528
rect 19676 86464 19692 86528
rect 19756 86464 19772 86528
rect 19836 86464 19852 86528
rect 19916 86464 19922 86528
rect 19606 86463 19922 86464
rect 21206 86528 21522 86529
rect 21206 86464 21212 86528
rect 21276 86464 21292 86528
rect 21356 86464 21372 86528
rect 21436 86464 21452 86528
rect 21516 86464 21522 86528
rect 21206 86463 21522 86464
rect 22806 86528 23122 86529
rect 22806 86464 22812 86528
rect 22876 86464 22892 86528
rect 22956 86464 22972 86528
rect 23036 86464 23052 86528
rect 23116 86464 23122 86528
rect 22806 86463 23122 86464
rect 24406 86528 24722 86529
rect 24406 86464 24412 86528
rect 24476 86464 24492 86528
rect 24556 86464 24572 86528
rect 24636 86464 24652 86528
rect 24716 86464 24722 86528
rect 24406 86463 24722 86464
rect 26006 86528 26322 86529
rect 26006 86464 26012 86528
rect 26076 86464 26092 86528
rect 26156 86464 26172 86528
rect 26236 86464 26252 86528
rect 26316 86464 26322 86528
rect 26006 86463 26322 86464
rect 27606 86528 27922 86529
rect 27606 86464 27612 86528
rect 27676 86464 27692 86528
rect 27756 86464 27772 86528
rect 27836 86464 27852 86528
rect 27916 86464 27922 86528
rect 27606 86463 27922 86464
rect 29206 86528 29522 86529
rect 29206 86464 29212 86528
rect 29276 86464 29292 86528
rect 29356 86464 29372 86528
rect 29436 86464 29452 86528
rect 29516 86464 29522 86528
rect 29206 86463 29522 86464
rect 30806 86528 31122 86529
rect 30806 86464 30812 86528
rect 30876 86464 30892 86528
rect 30956 86464 30972 86528
rect 31036 86464 31052 86528
rect 31116 86464 31122 86528
rect 30806 86463 31122 86464
rect 32406 86528 32722 86529
rect 32406 86464 32412 86528
rect 32476 86464 32492 86528
rect 32556 86464 32572 86528
rect 32636 86464 32652 86528
rect 32716 86464 32722 86528
rect 32406 86463 32722 86464
rect 34006 86528 34322 86529
rect 34006 86464 34012 86528
rect 34076 86464 34092 86528
rect 34156 86464 34172 86528
rect 34236 86464 34252 86528
rect 34316 86464 34322 86528
rect 34006 86463 34322 86464
rect 35606 86528 35922 86529
rect 35606 86464 35612 86528
rect 35676 86464 35692 86528
rect 35756 86464 35772 86528
rect 35836 86464 35852 86528
rect 35916 86464 35922 86528
rect 35606 86463 35922 86464
rect 37206 86528 37522 86529
rect 37206 86464 37212 86528
rect 37276 86464 37292 86528
rect 37356 86464 37372 86528
rect 37436 86464 37452 86528
rect 37516 86464 37522 86528
rect 37206 86463 37522 86464
rect 38806 86528 39122 86529
rect 38806 86464 38812 86528
rect 38876 86464 38892 86528
rect 38956 86464 38972 86528
rect 39036 86464 39052 86528
rect 39116 86464 39122 86528
rect 38806 86463 39122 86464
rect 40406 86528 40722 86529
rect 40406 86464 40412 86528
rect 40476 86464 40492 86528
rect 40556 86464 40572 86528
rect 40636 86464 40652 86528
rect 40716 86464 40722 86528
rect 40406 86463 40722 86464
rect 42006 86528 42322 86529
rect 42006 86464 42012 86528
rect 42076 86464 42092 86528
rect 42156 86464 42172 86528
rect 42236 86464 42252 86528
rect 42316 86464 42322 86528
rect 42006 86463 42322 86464
rect 43606 86528 43922 86529
rect 43606 86464 43612 86528
rect 43676 86464 43692 86528
rect 43756 86464 43772 86528
rect 43836 86464 43852 86528
rect 43916 86464 43922 86528
rect 43606 86463 43922 86464
rect 45206 86528 45522 86529
rect 45206 86464 45212 86528
rect 45276 86464 45292 86528
rect 45356 86464 45372 86528
rect 45436 86464 45452 86528
rect 45516 86464 45522 86528
rect 45206 86463 45522 86464
rect 46806 86528 47122 86529
rect 46806 86464 46812 86528
rect 46876 86464 46892 86528
rect 46956 86464 46972 86528
rect 47036 86464 47052 86528
rect 47116 86464 47122 86528
rect 46806 86463 47122 86464
rect 48406 86528 48722 86529
rect 48406 86464 48412 86528
rect 48476 86464 48492 86528
rect 48556 86464 48572 86528
rect 48636 86464 48652 86528
rect 48716 86464 48722 86528
rect 48406 86463 48722 86464
rect 50006 86528 50322 86529
rect 50006 86464 50012 86528
rect 50076 86464 50092 86528
rect 50156 86464 50172 86528
rect 50236 86464 50252 86528
rect 50316 86464 50322 86528
rect 50006 86463 50322 86464
rect 51606 86528 51922 86529
rect 51606 86464 51612 86528
rect 51676 86464 51692 86528
rect 51756 86464 51772 86528
rect 51836 86464 51852 86528
rect 51916 86464 51922 86528
rect 51606 86463 51922 86464
rect 53206 86528 53522 86529
rect 53206 86464 53212 86528
rect 53276 86464 53292 86528
rect 53356 86464 53372 86528
rect 53436 86464 53452 86528
rect 53516 86464 53522 86528
rect 53206 86463 53522 86464
rect 54806 86528 55122 86529
rect 54806 86464 54812 86528
rect 54876 86464 54892 86528
rect 54956 86464 54972 86528
rect 55036 86464 55052 86528
rect 55116 86464 55122 86528
rect 54806 86463 55122 86464
rect 56406 86528 56722 86529
rect 56406 86464 56412 86528
rect 56476 86464 56492 86528
rect 56556 86464 56572 86528
rect 56636 86464 56652 86528
rect 56716 86464 56722 86528
rect 56406 86463 56722 86464
rect 58006 86528 58322 86529
rect 58006 86464 58012 86528
rect 58076 86464 58092 86528
rect 58156 86464 58172 86528
rect 58236 86464 58252 86528
rect 58316 86464 58322 86528
rect 58006 86463 58322 86464
rect 59606 86528 59922 86529
rect 59606 86464 59612 86528
rect 59676 86464 59692 86528
rect 59756 86464 59772 86528
rect 59836 86464 59852 86528
rect 59916 86464 59922 86528
rect 59606 86463 59922 86464
rect 61206 86528 61522 86529
rect 61206 86464 61212 86528
rect 61276 86464 61292 86528
rect 61356 86464 61372 86528
rect 61436 86464 61452 86528
rect 61516 86464 61522 86528
rect 61206 86463 61522 86464
rect 62806 86528 63122 86529
rect 62806 86464 62812 86528
rect 62876 86464 62892 86528
rect 62956 86464 62972 86528
rect 63036 86464 63052 86528
rect 63116 86464 63122 86528
rect 62806 86463 63122 86464
rect 64406 86528 64722 86529
rect 64406 86464 64412 86528
rect 64476 86464 64492 86528
rect 64556 86464 64572 86528
rect 64636 86464 64652 86528
rect 64716 86464 64722 86528
rect 64406 86463 64722 86464
rect 66006 86528 66322 86529
rect 66006 86464 66012 86528
rect 66076 86464 66092 86528
rect 66156 86464 66172 86528
rect 66236 86464 66252 86528
rect 66316 86464 66322 86528
rect 66006 86463 66322 86464
rect 67606 86528 67922 86529
rect 67606 86464 67612 86528
rect 67676 86464 67692 86528
rect 67756 86464 67772 86528
rect 67836 86464 67852 86528
rect 67916 86464 67922 86528
rect 67606 86463 67922 86464
rect 69206 86528 69522 86529
rect 69206 86464 69212 86528
rect 69276 86464 69292 86528
rect 69356 86464 69372 86528
rect 69436 86464 69452 86528
rect 69516 86464 69522 86528
rect 69206 86463 69522 86464
rect 70806 86528 71122 86529
rect 70806 86464 70812 86528
rect 70876 86464 70892 86528
rect 70956 86464 70972 86528
rect 71036 86464 71052 86528
rect 71116 86464 71122 86528
rect 70806 86463 71122 86464
rect 72406 86528 72722 86529
rect 72406 86464 72412 86528
rect 72476 86464 72492 86528
rect 72556 86464 72572 86528
rect 72636 86464 72652 86528
rect 72716 86464 72722 86528
rect 72406 86463 72722 86464
rect 74006 86528 74322 86529
rect 74006 86464 74012 86528
rect 74076 86464 74092 86528
rect 74156 86464 74172 86528
rect 74236 86464 74252 86528
rect 74316 86464 74322 86528
rect 74006 86463 74322 86464
rect 75606 86528 75922 86529
rect 75606 86464 75612 86528
rect 75676 86464 75692 86528
rect 75756 86464 75772 86528
rect 75836 86464 75852 86528
rect 75916 86464 75922 86528
rect 75606 86463 75922 86464
rect 77206 86528 77522 86529
rect 77206 86464 77212 86528
rect 77276 86464 77292 86528
rect 77356 86464 77372 86528
rect 77436 86464 77452 86528
rect 77516 86464 77522 86528
rect 77206 86463 77522 86464
rect 78806 86528 79122 86529
rect 78806 86464 78812 86528
rect 78876 86464 78892 86528
rect 78956 86464 78972 86528
rect 79036 86464 79052 86528
rect 79116 86464 79122 86528
rect 78806 86463 79122 86464
rect 80406 86528 80722 86529
rect 80406 86464 80412 86528
rect 80476 86464 80492 86528
rect 80556 86464 80572 86528
rect 80636 86464 80652 86528
rect 80716 86464 80722 86528
rect 80406 86463 80722 86464
rect 82006 86528 82322 86529
rect 82006 86464 82012 86528
rect 82076 86464 82092 86528
rect 82156 86464 82172 86528
rect 82236 86464 82252 86528
rect 82316 86464 82322 86528
rect 82006 86463 82322 86464
rect 83606 86528 83922 86529
rect 83606 86464 83612 86528
rect 83676 86464 83692 86528
rect 83756 86464 83772 86528
rect 83836 86464 83852 86528
rect 83916 86464 83922 86528
rect 83606 86463 83922 86464
rect 85206 86528 85522 86529
rect 85206 86464 85212 86528
rect 85276 86464 85292 86528
rect 85356 86464 85372 86528
rect 85436 86464 85452 86528
rect 85516 86464 85522 86528
rect 85206 86463 85522 86464
rect 86806 86528 87122 86529
rect 86806 86464 86812 86528
rect 86876 86464 86892 86528
rect 86956 86464 86972 86528
rect 87036 86464 87052 86528
rect 87116 86464 87122 86528
rect 86806 86463 87122 86464
rect 88406 86528 88722 86529
rect 88406 86464 88412 86528
rect 88476 86464 88492 86528
rect 88556 86464 88572 86528
rect 88636 86464 88652 86528
rect 88716 86464 88722 86528
rect 88406 86463 88722 86464
rect 90006 86528 90322 86529
rect 90006 86464 90012 86528
rect 90076 86464 90092 86528
rect 90156 86464 90172 86528
rect 90236 86464 90252 86528
rect 90316 86464 90322 86528
rect 90006 86463 90322 86464
rect 91606 86528 91922 86529
rect 91606 86464 91612 86528
rect 91676 86464 91692 86528
rect 91756 86464 91772 86528
rect 91836 86464 91852 86528
rect 91916 86464 91922 86528
rect 91606 86463 91922 86464
rect 93206 86528 93522 86529
rect 93206 86464 93212 86528
rect 93276 86464 93292 86528
rect 93356 86464 93372 86528
rect 93436 86464 93452 86528
rect 93516 86464 93522 86528
rect 93206 86463 93522 86464
rect 94806 86528 95122 86529
rect 94806 86464 94812 86528
rect 94876 86464 94892 86528
rect 94956 86464 94972 86528
rect 95036 86464 95052 86528
rect 95116 86464 95122 86528
rect 94806 86463 95122 86464
rect 96406 86528 96722 86529
rect 96406 86464 96412 86528
rect 96476 86464 96492 86528
rect 96556 86464 96572 86528
rect 96636 86464 96652 86528
rect 96716 86464 96722 86528
rect 96406 86463 96722 86464
rect 98006 86528 98322 86529
rect 98006 86464 98012 86528
rect 98076 86464 98092 86528
rect 98156 86464 98172 86528
rect 98236 86464 98252 86528
rect 98316 86464 98322 86528
rect 98006 86463 98322 86464
rect 99606 86528 99922 86529
rect 99606 86464 99612 86528
rect 99676 86464 99692 86528
rect 99756 86464 99772 86528
rect 99836 86464 99852 86528
rect 99916 86464 99922 86528
rect 99606 86463 99922 86464
rect 101206 86528 101522 86529
rect 101206 86464 101212 86528
rect 101276 86464 101292 86528
rect 101356 86464 101372 86528
rect 101436 86464 101452 86528
rect 101516 86464 101522 86528
rect 101206 86463 101522 86464
rect 102806 86528 103122 86529
rect 102806 86464 102812 86528
rect 102876 86464 102892 86528
rect 102956 86464 102972 86528
rect 103036 86464 103052 86528
rect 103116 86464 103122 86528
rect 102806 86463 103122 86464
rect 104406 86528 104722 86529
rect 104406 86464 104412 86528
rect 104476 86464 104492 86528
rect 104556 86464 104572 86528
rect 104636 86464 104652 86528
rect 104716 86464 104722 86528
rect 104406 86463 104722 86464
rect 106006 86528 106322 86529
rect 106006 86464 106012 86528
rect 106076 86464 106092 86528
rect 106156 86464 106172 86528
rect 106236 86464 106252 86528
rect 106316 86464 106322 86528
rect 106006 86463 106322 86464
rect 107606 86528 107922 86529
rect 107606 86464 107612 86528
rect 107676 86464 107692 86528
rect 107756 86464 107772 86528
rect 107836 86464 107852 86528
rect 107916 86464 107922 86528
rect 107606 86463 107922 86464
rect 11462 86124 11468 86188
rect 11532 86186 11538 86188
rect 38837 86186 38903 86189
rect 11532 86184 38903 86186
rect 11532 86128 38842 86184
rect 38898 86128 38903 86184
rect 11532 86126 38903 86128
rect 11532 86124 11538 86126
rect 38837 86123 38903 86126
rect 48865 86186 48931 86189
rect 55305 86186 55371 86189
rect 48865 86184 55371 86186
rect 48865 86128 48870 86184
rect 48926 86128 55310 86184
rect 55366 86128 55371 86184
rect 48865 86126 55371 86128
rect 48865 86123 48931 86126
rect 55305 86123 55371 86126
rect 2946 85984 3262 85985
rect 2946 85920 2952 85984
rect 3016 85920 3032 85984
rect 3096 85920 3112 85984
rect 3176 85920 3192 85984
rect 3256 85920 3262 85984
rect 2946 85919 3262 85920
rect 4546 85984 4862 85985
rect 4546 85920 4552 85984
rect 4616 85920 4632 85984
rect 4696 85920 4712 85984
rect 4776 85920 4792 85984
rect 4856 85920 4862 85984
rect 4546 85919 4862 85920
rect 6146 85984 6462 85985
rect 6146 85920 6152 85984
rect 6216 85920 6232 85984
rect 6296 85920 6312 85984
rect 6376 85920 6392 85984
rect 6456 85920 6462 85984
rect 6146 85919 6462 85920
rect 7746 85984 8062 85985
rect 7746 85920 7752 85984
rect 7816 85920 7832 85984
rect 7896 85920 7912 85984
rect 7976 85920 7992 85984
rect 8056 85920 8062 85984
rect 7746 85919 8062 85920
rect 9346 85984 9662 85985
rect 9346 85920 9352 85984
rect 9416 85920 9432 85984
rect 9496 85920 9512 85984
rect 9576 85920 9592 85984
rect 9656 85920 9662 85984
rect 9346 85919 9662 85920
rect 10946 85984 11262 85985
rect 10946 85920 10952 85984
rect 11016 85920 11032 85984
rect 11096 85920 11112 85984
rect 11176 85920 11192 85984
rect 11256 85920 11262 85984
rect 10946 85919 11262 85920
rect 12546 85984 12862 85985
rect 12546 85920 12552 85984
rect 12616 85920 12632 85984
rect 12696 85920 12712 85984
rect 12776 85920 12792 85984
rect 12856 85920 12862 85984
rect 12546 85919 12862 85920
rect 14146 85984 14462 85985
rect 14146 85920 14152 85984
rect 14216 85920 14232 85984
rect 14296 85920 14312 85984
rect 14376 85920 14392 85984
rect 14456 85920 14462 85984
rect 14146 85919 14462 85920
rect 15746 85984 16062 85985
rect 15746 85920 15752 85984
rect 15816 85920 15832 85984
rect 15896 85920 15912 85984
rect 15976 85920 15992 85984
rect 16056 85920 16062 85984
rect 15746 85919 16062 85920
rect 17346 85984 17662 85985
rect 17346 85920 17352 85984
rect 17416 85920 17432 85984
rect 17496 85920 17512 85984
rect 17576 85920 17592 85984
rect 17656 85920 17662 85984
rect 17346 85919 17662 85920
rect 18946 85984 19262 85985
rect 18946 85920 18952 85984
rect 19016 85920 19032 85984
rect 19096 85920 19112 85984
rect 19176 85920 19192 85984
rect 19256 85920 19262 85984
rect 18946 85919 19262 85920
rect 20546 85984 20862 85985
rect 20546 85920 20552 85984
rect 20616 85920 20632 85984
rect 20696 85920 20712 85984
rect 20776 85920 20792 85984
rect 20856 85920 20862 85984
rect 20546 85919 20862 85920
rect 22146 85984 22462 85985
rect 22146 85920 22152 85984
rect 22216 85920 22232 85984
rect 22296 85920 22312 85984
rect 22376 85920 22392 85984
rect 22456 85920 22462 85984
rect 22146 85919 22462 85920
rect 23746 85984 24062 85985
rect 23746 85920 23752 85984
rect 23816 85920 23832 85984
rect 23896 85920 23912 85984
rect 23976 85920 23992 85984
rect 24056 85920 24062 85984
rect 23746 85919 24062 85920
rect 25346 85984 25662 85985
rect 25346 85920 25352 85984
rect 25416 85920 25432 85984
rect 25496 85920 25512 85984
rect 25576 85920 25592 85984
rect 25656 85920 25662 85984
rect 25346 85919 25662 85920
rect 26946 85984 27262 85985
rect 26946 85920 26952 85984
rect 27016 85920 27032 85984
rect 27096 85920 27112 85984
rect 27176 85920 27192 85984
rect 27256 85920 27262 85984
rect 26946 85919 27262 85920
rect 28546 85984 28862 85985
rect 28546 85920 28552 85984
rect 28616 85920 28632 85984
rect 28696 85920 28712 85984
rect 28776 85920 28792 85984
rect 28856 85920 28862 85984
rect 28546 85919 28862 85920
rect 30146 85984 30462 85985
rect 30146 85920 30152 85984
rect 30216 85920 30232 85984
rect 30296 85920 30312 85984
rect 30376 85920 30392 85984
rect 30456 85920 30462 85984
rect 30146 85919 30462 85920
rect 31746 85984 32062 85985
rect 31746 85920 31752 85984
rect 31816 85920 31832 85984
rect 31896 85920 31912 85984
rect 31976 85920 31992 85984
rect 32056 85920 32062 85984
rect 31746 85919 32062 85920
rect 33346 85984 33662 85985
rect 33346 85920 33352 85984
rect 33416 85920 33432 85984
rect 33496 85920 33512 85984
rect 33576 85920 33592 85984
rect 33656 85920 33662 85984
rect 33346 85919 33662 85920
rect 34946 85984 35262 85985
rect 34946 85920 34952 85984
rect 35016 85920 35032 85984
rect 35096 85920 35112 85984
rect 35176 85920 35192 85984
rect 35256 85920 35262 85984
rect 34946 85919 35262 85920
rect 36546 85984 36862 85985
rect 36546 85920 36552 85984
rect 36616 85920 36632 85984
rect 36696 85920 36712 85984
rect 36776 85920 36792 85984
rect 36856 85920 36862 85984
rect 36546 85919 36862 85920
rect 38146 85984 38462 85985
rect 38146 85920 38152 85984
rect 38216 85920 38232 85984
rect 38296 85920 38312 85984
rect 38376 85920 38392 85984
rect 38456 85920 38462 85984
rect 38146 85919 38462 85920
rect 39746 85984 40062 85985
rect 39746 85920 39752 85984
rect 39816 85920 39832 85984
rect 39896 85920 39912 85984
rect 39976 85920 39992 85984
rect 40056 85920 40062 85984
rect 39746 85919 40062 85920
rect 41346 85984 41662 85985
rect 41346 85920 41352 85984
rect 41416 85920 41432 85984
rect 41496 85920 41512 85984
rect 41576 85920 41592 85984
rect 41656 85920 41662 85984
rect 41346 85919 41662 85920
rect 42946 85984 43262 85985
rect 42946 85920 42952 85984
rect 43016 85920 43032 85984
rect 43096 85920 43112 85984
rect 43176 85920 43192 85984
rect 43256 85920 43262 85984
rect 42946 85919 43262 85920
rect 44546 85984 44862 85985
rect 44546 85920 44552 85984
rect 44616 85920 44632 85984
rect 44696 85920 44712 85984
rect 44776 85920 44792 85984
rect 44856 85920 44862 85984
rect 44546 85919 44862 85920
rect 46146 85984 46462 85985
rect 46146 85920 46152 85984
rect 46216 85920 46232 85984
rect 46296 85920 46312 85984
rect 46376 85920 46392 85984
rect 46456 85920 46462 85984
rect 46146 85919 46462 85920
rect 47746 85984 48062 85985
rect 47746 85920 47752 85984
rect 47816 85920 47832 85984
rect 47896 85920 47912 85984
rect 47976 85920 47992 85984
rect 48056 85920 48062 85984
rect 47746 85919 48062 85920
rect 49346 85984 49662 85985
rect 49346 85920 49352 85984
rect 49416 85920 49432 85984
rect 49496 85920 49512 85984
rect 49576 85920 49592 85984
rect 49656 85920 49662 85984
rect 49346 85919 49662 85920
rect 50946 85984 51262 85985
rect 50946 85920 50952 85984
rect 51016 85920 51032 85984
rect 51096 85920 51112 85984
rect 51176 85920 51192 85984
rect 51256 85920 51262 85984
rect 50946 85919 51262 85920
rect 52546 85984 52862 85985
rect 52546 85920 52552 85984
rect 52616 85920 52632 85984
rect 52696 85920 52712 85984
rect 52776 85920 52792 85984
rect 52856 85920 52862 85984
rect 52546 85919 52862 85920
rect 54146 85984 54462 85985
rect 54146 85920 54152 85984
rect 54216 85920 54232 85984
rect 54296 85920 54312 85984
rect 54376 85920 54392 85984
rect 54456 85920 54462 85984
rect 54146 85919 54462 85920
rect 55746 85984 56062 85985
rect 55746 85920 55752 85984
rect 55816 85920 55832 85984
rect 55896 85920 55912 85984
rect 55976 85920 55992 85984
rect 56056 85920 56062 85984
rect 55746 85919 56062 85920
rect 57346 85984 57662 85985
rect 57346 85920 57352 85984
rect 57416 85920 57432 85984
rect 57496 85920 57512 85984
rect 57576 85920 57592 85984
rect 57656 85920 57662 85984
rect 57346 85919 57662 85920
rect 58946 85984 59262 85985
rect 58946 85920 58952 85984
rect 59016 85920 59032 85984
rect 59096 85920 59112 85984
rect 59176 85920 59192 85984
rect 59256 85920 59262 85984
rect 58946 85919 59262 85920
rect 60546 85984 60862 85985
rect 60546 85920 60552 85984
rect 60616 85920 60632 85984
rect 60696 85920 60712 85984
rect 60776 85920 60792 85984
rect 60856 85920 60862 85984
rect 60546 85919 60862 85920
rect 62146 85984 62462 85985
rect 62146 85920 62152 85984
rect 62216 85920 62232 85984
rect 62296 85920 62312 85984
rect 62376 85920 62392 85984
rect 62456 85920 62462 85984
rect 62146 85919 62462 85920
rect 63746 85984 64062 85985
rect 63746 85920 63752 85984
rect 63816 85920 63832 85984
rect 63896 85920 63912 85984
rect 63976 85920 63992 85984
rect 64056 85920 64062 85984
rect 63746 85919 64062 85920
rect 65346 85984 65662 85985
rect 65346 85920 65352 85984
rect 65416 85920 65432 85984
rect 65496 85920 65512 85984
rect 65576 85920 65592 85984
rect 65656 85920 65662 85984
rect 65346 85919 65662 85920
rect 66946 85984 67262 85985
rect 66946 85920 66952 85984
rect 67016 85920 67032 85984
rect 67096 85920 67112 85984
rect 67176 85920 67192 85984
rect 67256 85920 67262 85984
rect 66946 85919 67262 85920
rect 68546 85984 68862 85985
rect 68546 85920 68552 85984
rect 68616 85920 68632 85984
rect 68696 85920 68712 85984
rect 68776 85920 68792 85984
rect 68856 85920 68862 85984
rect 68546 85919 68862 85920
rect 70146 85984 70462 85985
rect 70146 85920 70152 85984
rect 70216 85920 70232 85984
rect 70296 85920 70312 85984
rect 70376 85920 70392 85984
rect 70456 85920 70462 85984
rect 70146 85919 70462 85920
rect 71746 85984 72062 85985
rect 71746 85920 71752 85984
rect 71816 85920 71832 85984
rect 71896 85920 71912 85984
rect 71976 85920 71992 85984
rect 72056 85920 72062 85984
rect 71746 85919 72062 85920
rect 73346 85984 73662 85985
rect 73346 85920 73352 85984
rect 73416 85920 73432 85984
rect 73496 85920 73512 85984
rect 73576 85920 73592 85984
rect 73656 85920 73662 85984
rect 73346 85919 73662 85920
rect 74946 85984 75262 85985
rect 74946 85920 74952 85984
rect 75016 85920 75032 85984
rect 75096 85920 75112 85984
rect 75176 85920 75192 85984
rect 75256 85920 75262 85984
rect 74946 85919 75262 85920
rect 76546 85984 76862 85985
rect 76546 85920 76552 85984
rect 76616 85920 76632 85984
rect 76696 85920 76712 85984
rect 76776 85920 76792 85984
rect 76856 85920 76862 85984
rect 76546 85919 76862 85920
rect 78146 85984 78462 85985
rect 78146 85920 78152 85984
rect 78216 85920 78232 85984
rect 78296 85920 78312 85984
rect 78376 85920 78392 85984
rect 78456 85920 78462 85984
rect 78146 85919 78462 85920
rect 79746 85984 80062 85985
rect 79746 85920 79752 85984
rect 79816 85920 79832 85984
rect 79896 85920 79912 85984
rect 79976 85920 79992 85984
rect 80056 85920 80062 85984
rect 79746 85919 80062 85920
rect 81346 85984 81662 85985
rect 81346 85920 81352 85984
rect 81416 85920 81432 85984
rect 81496 85920 81512 85984
rect 81576 85920 81592 85984
rect 81656 85920 81662 85984
rect 81346 85919 81662 85920
rect 82946 85984 83262 85985
rect 82946 85920 82952 85984
rect 83016 85920 83032 85984
rect 83096 85920 83112 85984
rect 83176 85920 83192 85984
rect 83256 85920 83262 85984
rect 82946 85919 83262 85920
rect 84546 85984 84862 85985
rect 84546 85920 84552 85984
rect 84616 85920 84632 85984
rect 84696 85920 84712 85984
rect 84776 85920 84792 85984
rect 84856 85920 84862 85984
rect 84546 85919 84862 85920
rect 86146 85984 86462 85985
rect 86146 85920 86152 85984
rect 86216 85920 86232 85984
rect 86296 85920 86312 85984
rect 86376 85920 86392 85984
rect 86456 85920 86462 85984
rect 86146 85919 86462 85920
rect 87746 85984 88062 85985
rect 87746 85920 87752 85984
rect 87816 85920 87832 85984
rect 87896 85920 87912 85984
rect 87976 85920 87992 85984
rect 88056 85920 88062 85984
rect 87746 85919 88062 85920
rect 89346 85984 89662 85985
rect 89346 85920 89352 85984
rect 89416 85920 89432 85984
rect 89496 85920 89512 85984
rect 89576 85920 89592 85984
rect 89656 85920 89662 85984
rect 89346 85919 89662 85920
rect 90946 85984 91262 85985
rect 90946 85920 90952 85984
rect 91016 85920 91032 85984
rect 91096 85920 91112 85984
rect 91176 85920 91192 85984
rect 91256 85920 91262 85984
rect 90946 85919 91262 85920
rect 92546 85984 92862 85985
rect 92546 85920 92552 85984
rect 92616 85920 92632 85984
rect 92696 85920 92712 85984
rect 92776 85920 92792 85984
rect 92856 85920 92862 85984
rect 92546 85919 92862 85920
rect 94146 85984 94462 85985
rect 94146 85920 94152 85984
rect 94216 85920 94232 85984
rect 94296 85920 94312 85984
rect 94376 85920 94392 85984
rect 94456 85920 94462 85984
rect 94146 85919 94462 85920
rect 95746 85984 96062 85985
rect 95746 85920 95752 85984
rect 95816 85920 95832 85984
rect 95896 85920 95912 85984
rect 95976 85920 95992 85984
rect 96056 85920 96062 85984
rect 95746 85919 96062 85920
rect 97346 85984 97662 85985
rect 97346 85920 97352 85984
rect 97416 85920 97432 85984
rect 97496 85920 97512 85984
rect 97576 85920 97592 85984
rect 97656 85920 97662 85984
rect 97346 85919 97662 85920
rect 98946 85984 99262 85985
rect 98946 85920 98952 85984
rect 99016 85920 99032 85984
rect 99096 85920 99112 85984
rect 99176 85920 99192 85984
rect 99256 85920 99262 85984
rect 98946 85919 99262 85920
rect 100546 85984 100862 85985
rect 100546 85920 100552 85984
rect 100616 85920 100632 85984
rect 100696 85920 100712 85984
rect 100776 85920 100792 85984
rect 100856 85920 100862 85984
rect 100546 85919 100862 85920
rect 102146 85984 102462 85985
rect 102146 85920 102152 85984
rect 102216 85920 102232 85984
rect 102296 85920 102312 85984
rect 102376 85920 102392 85984
rect 102456 85920 102462 85984
rect 102146 85919 102462 85920
rect 103746 85984 104062 85985
rect 103746 85920 103752 85984
rect 103816 85920 103832 85984
rect 103896 85920 103912 85984
rect 103976 85920 103992 85984
rect 104056 85920 104062 85984
rect 103746 85919 104062 85920
rect 105346 85984 105662 85985
rect 105346 85920 105352 85984
rect 105416 85920 105432 85984
rect 105496 85920 105512 85984
rect 105576 85920 105592 85984
rect 105656 85920 105662 85984
rect 105346 85919 105662 85920
rect 106946 85984 107262 85985
rect 106946 85920 106952 85984
rect 107016 85920 107032 85984
rect 107096 85920 107112 85984
rect 107176 85920 107192 85984
rect 107256 85920 107262 85984
rect 106946 85919 107262 85920
rect 108546 85984 108862 85985
rect 108546 85920 108552 85984
rect 108616 85920 108632 85984
rect 108696 85920 108712 85984
rect 108776 85920 108792 85984
rect 108856 85920 108862 85984
rect 108546 85919 108862 85920
rect 61009 85916 61075 85917
rect 60958 85852 60964 85916
rect 61028 85914 61075 85916
rect 63493 85916 63559 85917
rect 68093 85916 68159 85917
rect 72141 85916 72207 85917
rect 63493 85914 63540 85916
rect 61028 85912 61120 85914
rect 61070 85856 61120 85912
rect 61028 85854 61120 85856
rect 63448 85912 63540 85914
rect 63448 85856 63498 85912
rect 63448 85854 63540 85856
rect 61028 85852 61075 85854
rect 61009 85851 61075 85852
rect 63493 85852 63540 85854
rect 63604 85852 63610 85916
rect 68093 85914 68140 85916
rect 68048 85912 68140 85914
rect 68048 85856 68098 85912
rect 68048 85854 68140 85856
rect 68093 85852 68140 85854
rect 68204 85852 68210 85916
rect 72141 85912 72188 85916
rect 72252 85914 72258 85916
rect 72141 85856 72146 85912
rect 72141 85852 72188 85856
rect 72252 85854 72298 85914
rect 72252 85852 72258 85854
rect 63493 85851 63559 85852
rect 68093 85851 68159 85852
rect 72141 85851 72207 85852
rect 68001 85778 68067 85781
rect 68318 85778 68324 85780
rect 68001 85776 68324 85778
rect 68001 85720 68006 85776
rect 68062 85720 68324 85776
rect 68001 85718 68324 85720
rect 68001 85715 68067 85718
rect 68318 85716 68324 85718
rect 68388 85716 68394 85780
rect 40033 85642 40099 85645
rect 41781 85644 41847 85645
rect 40166 85642 40172 85644
rect 40033 85640 40172 85642
rect 40033 85584 40038 85640
rect 40094 85584 40172 85640
rect 40033 85582 40172 85584
rect 40033 85579 40099 85582
rect 40166 85580 40172 85582
rect 40236 85580 40242 85644
rect 41781 85640 41828 85644
rect 41892 85642 41898 85644
rect 42793 85642 42859 85645
rect 46565 85644 46631 85645
rect 47301 85644 47367 85645
rect 44030 85642 44036 85644
rect 41781 85584 41786 85640
rect 41781 85580 41828 85584
rect 41892 85582 41938 85642
rect 42793 85640 44036 85642
rect 42793 85584 42798 85640
rect 42854 85584 44036 85640
rect 42793 85582 44036 85584
rect 41892 85580 41898 85582
rect 41781 85579 41847 85580
rect 42793 85579 42859 85582
rect 44030 85580 44036 85582
rect 44100 85580 44106 85644
rect 46565 85640 46612 85644
rect 46676 85642 46682 85644
rect 46565 85584 46570 85640
rect 46565 85580 46612 85584
rect 46676 85582 46722 85642
rect 47301 85640 47348 85644
rect 47412 85642 47418 85644
rect 47301 85584 47306 85640
rect 46676 85580 46682 85582
rect 47301 85580 47348 85584
rect 47412 85582 47458 85642
rect 47412 85580 47418 85582
rect 48998 85580 49004 85644
rect 49068 85642 49074 85644
rect 49233 85642 49299 85645
rect 49068 85640 49299 85642
rect 49068 85584 49238 85640
rect 49294 85584 49299 85640
rect 49068 85582 49299 85584
rect 49068 85580 49074 85582
rect 46565 85579 46631 85580
rect 47301 85579 47367 85580
rect 49233 85579 49299 85582
rect 50470 85580 50476 85644
rect 50540 85642 50546 85644
rect 50797 85642 50863 85645
rect 50540 85640 50863 85642
rect 50540 85584 50802 85640
rect 50858 85584 50863 85640
rect 50540 85582 50863 85584
rect 50540 85580 50546 85582
rect 50797 85579 50863 85582
rect 55213 85644 55279 85645
rect 55213 85640 55260 85644
rect 55324 85642 55330 85644
rect 55673 85642 55739 85645
rect 56174 85642 56180 85644
rect 55213 85584 55218 85640
rect 55213 85580 55260 85584
rect 55324 85582 55370 85642
rect 55673 85640 56180 85642
rect 55673 85584 55678 85640
rect 55734 85584 56180 85640
rect 55673 85582 56180 85584
rect 55324 85580 55330 85582
rect 55213 85579 55279 85580
rect 55673 85579 55739 85582
rect 56174 85580 56180 85582
rect 56244 85580 56250 85644
rect 58341 85642 58407 85645
rect 58750 85642 58756 85644
rect 58341 85640 58756 85642
rect 58341 85584 58346 85640
rect 58402 85584 58756 85640
rect 58341 85582 58756 85584
rect 58341 85579 58407 85582
rect 58750 85580 58756 85582
rect 58820 85580 58826 85644
rect 62481 85642 62547 85645
rect 62614 85642 62620 85644
rect 62481 85640 62620 85642
rect 62481 85584 62486 85640
rect 62542 85584 62620 85640
rect 62481 85582 62620 85584
rect 62481 85579 62547 85582
rect 62614 85580 62620 85582
rect 62684 85580 62690 85644
rect 73153 85642 73219 85645
rect 73838 85642 73844 85644
rect 73153 85640 73844 85642
rect 73153 85584 73158 85640
rect 73214 85584 73844 85640
rect 73153 85582 73844 85584
rect 73153 85579 73219 85582
rect 73838 85580 73844 85582
rect 73908 85580 73914 85644
rect 74625 85642 74691 85645
rect 75913 85642 75979 85645
rect 77661 85644 77727 85645
rect 76230 85642 76236 85644
rect 74625 85640 75378 85642
rect 74625 85584 74630 85640
rect 74686 85584 75378 85640
rect 74625 85582 75378 85584
rect 74625 85579 74691 85582
rect 75318 85508 75378 85582
rect 75913 85640 76236 85642
rect 75913 85584 75918 85640
rect 75974 85584 76236 85640
rect 75913 85582 76236 85584
rect 75913 85579 75979 85582
rect 76230 85580 76236 85582
rect 76300 85580 76306 85644
rect 77661 85642 77708 85644
rect 77616 85640 77708 85642
rect 77616 85584 77666 85640
rect 77616 85582 77708 85584
rect 77661 85580 77708 85582
rect 77772 85580 77778 85644
rect 91277 85642 91343 85645
rect 100937 85642 101003 85645
rect 101990 85642 101996 85644
rect 91277 85640 91570 85642
rect 91277 85584 91282 85640
rect 91338 85584 91570 85640
rect 91277 85582 91570 85584
rect 77661 85579 77727 85580
rect 91277 85579 91343 85582
rect 91510 85508 91570 85582
rect 100937 85640 101996 85642
rect 100937 85584 100942 85640
rect 100998 85584 101996 85640
rect 100937 85582 101996 85584
rect 100937 85579 101003 85582
rect 101990 85580 101996 85582
rect 102060 85580 102066 85644
rect 75310 85444 75316 85508
rect 75380 85444 75386 85508
rect 91502 85444 91508 85508
rect 91572 85444 91578 85508
rect 3606 85440 3922 85441
rect 3606 85376 3612 85440
rect 3676 85376 3692 85440
rect 3756 85376 3772 85440
rect 3836 85376 3852 85440
rect 3916 85376 3922 85440
rect 3606 85375 3922 85376
rect 5206 85440 5522 85441
rect 5206 85376 5212 85440
rect 5276 85376 5292 85440
rect 5356 85376 5372 85440
rect 5436 85376 5452 85440
rect 5516 85376 5522 85440
rect 5206 85375 5522 85376
rect 6806 85440 7122 85441
rect 6806 85376 6812 85440
rect 6876 85376 6892 85440
rect 6956 85376 6972 85440
rect 7036 85376 7052 85440
rect 7116 85376 7122 85440
rect 6806 85375 7122 85376
rect 8406 85440 8722 85441
rect 8406 85376 8412 85440
rect 8476 85376 8492 85440
rect 8556 85376 8572 85440
rect 8636 85376 8652 85440
rect 8716 85376 8722 85440
rect 8406 85375 8722 85376
rect 5073 85098 5139 85101
rect 53005 85098 53071 85101
rect 5073 85096 53071 85098
rect 5073 85040 5078 85096
rect 5134 85040 53010 85096
rect 53066 85040 53071 85096
rect 5073 85038 53071 85040
rect 5073 85035 5139 85038
rect 53005 85035 53071 85038
rect 2946 84896 3262 84897
rect 2946 84832 2952 84896
rect 3016 84832 3032 84896
rect 3096 84832 3112 84896
rect 3176 84832 3192 84896
rect 3256 84832 3262 84896
rect 2946 84831 3262 84832
rect 4546 84896 4862 84897
rect 4546 84832 4552 84896
rect 4616 84832 4632 84896
rect 4696 84832 4712 84896
rect 4776 84832 4792 84896
rect 4856 84832 4862 84896
rect 4546 84831 4862 84832
rect 6146 84896 6462 84897
rect 6146 84832 6152 84896
rect 6216 84832 6232 84896
rect 6296 84832 6312 84896
rect 6376 84832 6392 84896
rect 6456 84832 6462 84896
rect 6146 84831 6462 84832
rect 7746 84896 8062 84897
rect 7746 84832 7752 84896
rect 7816 84832 7832 84896
rect 7896 84832 7912 84896
rect 7976 84832 7992 84896
rect 8056 84832 8062 84896
rect 7746 84831 8062 84832
rect 9346 84896 9662 84897
rect 9346 84832 9352 84896
rect 9416 84832 9432 84896
rect 9496 84832 9512 84896
rect 9576 84832 9592 84896
rect 9656 84832 9662 84896
rect 9346 84831 9662 84832
rect 52453 84828 52519 84829
rect 52453 84826 52500 84828
rect 52408 84824 52500 84826
rect 52408 84768 52458 84824
rect 52408 84766 52500 84768
rect 52453 84764 52500 84766
rect 52564 84764 52570 84828
rect 52453 84763 52519 84764
rect 51165 84692 51231 84693
rect 53833 84692 53899 84693
rect 51165 84690 51212 84692
rect 51120 84688 51212 84690
rect 51120 84632 51170 84688
rect 51120 84630 51212 84632
rect 51165 84628 51212 84630
rect 51276 84628 51282 84692
rect 53782 84628 53788 84692
rect 53852 84690 53899 84692
rect 66253 84692 66319 84693
rect 71221 84692 71287 84693
rect 66253 84690 66300 84692
rect 53852 84688 53944 84690
rect 53894 84632 53944 84688
rect 53852 84630 53944 84632
rect 66208 84688 66300 84690
rect 66208 84632 66258 84688
rect 66208 84630 66300 84632
rect 53852 84628 53899 84630
rect 51165 84627 51231 84628
rect 53833 84627 53899 84628
rect 66253 84628 66300 84630
rect 66364 84628 66370 84692
rect 71221 84690 71268 84692
rect 71176 84688 71268 84690
rect 71176 84632 71226 84688
rect 71176 84630 71268 84632
rect 71221 84628 71268 84630
rect 71332 84628 71338 84692
rect 66253 84627 66319 84628
rect 71221 84627 71287 84628
rect 57605 84556 57671 84557
rect 78673 84556 78739 84557
rect 57605 84554 57652 84556
rect 57560 84552 57652 84554
rect 57560 84496 57610 84552
rect 57560 84494 57652 84496
rect 57605 84492 57652 84494
rect 57716 84492 57722 84556
rect 78622 84492 78628 84556
rect 78692 84554 78739 84556
rect 78692 84552 78784 84554
rect 78734 84496 78784 84552
rect 78692 84494 78784 84496
rect 78692 84492 78739 84494
rect 57605 84491 57671 84492
rect 78673 84491 78739 84492
rect 933 84418 999 84421
rect 0 84416 999 84418
rect 0 84360 938 84416
rect 994 84360 999 84416
rect 0 84358 999 84360
rect 933 84355 999 84358
rect 42517 84420 42583 84421
rect 44725 84420 44791 84421
rect 42517 84416 42564 84420
rect 42628 84418 42634 84420
rect 42517 84360 42522 84416
rect 42517 84356 42564 84360
rect 42628 84358 42674 84418
rect 44725 84416 44772 84420
rect 44836 84418 44842 84420
rect 44725 84360 44730 84416
rect 42628 84356 42634 84358
rect 44725 84356 44772 84360
rect 44836 84358 44882 84418
rect 44836 84356 44842 84358
rect 42517 84355 42583 84356
rect 44725 84355 44791 84356
rect 3606 84352 3922 84353
rect 3606 84288 3612 84352
rect 3676 84288 3692 84352
rect 3756 84288 3772 84352
rect 3836 84288 3852 84352
rect 3916 84288 3922 84352
rect 3606 84287 3922 84288
rect 5206 84352 5522 84353
rect 5206 84288 5212 84352
rect 5276 84288 5292 84352
rect 5356 84288 5372 84352
rect 5436 84288 5452 84352
rect 5516 84288 5522 84352
rect 5206 84287 5522 84288
rect 6806 84352 7122 84353
rect 6806 84288 6812 84352
rect 6876 84288 6892 84352
rect 6956 84288 6972 84352
rect 7036 84288 7052 84352
rect 7116 84288 7122 84352
rect 6806 84287 7122 84288
rect 8406 84352 8722 84353
rect 8406 84288 8412 84352
rect 8476 84288 8492 84352
rect 8556 84288 8572 84352
rect 8636 84288 8652 84352
rect 8716 84288 8722 84352
rect 8406 84287 8722 84288
rect 10910 84220 10916 84284
rect 10980 84282 10986 84284
rect 65006 84282 65012 84284
rect 10980 84222 65012 84282
rect 10980 84220 10986 84222
rect 65006 84220 65012 84222
rect 65076 84220 65082 84284
rect 2946 83808 3262 83809
rect 2946 83744 2952 83808
rect 3016 83744 3032 83808
rect 3096 83744 3112 83808
rect 3176 83744 3192 83808
rect 3256 83744 3262 83808
rect 2946 83743 3262 83744
rect 4546 83808 4862 83809
rect 4546 83744 4552 83808
rect 4616 83744 4632 83808
rect 4696 83744 4712 83808
rect 4776 83744 4792 83808
rect 4856 83744 4862 83808
rect 4546 83743 4862 83744
rect 6146 83808 6462 83809
rect 6146 83744 6152 83808
rect 6216 83744 6232 83808
rect 6296 83744 6312 83808
rect 6376 83744 6392 83808
rect 6456 83744 6462 83808
rect 6146 83743 6462 83744
rect 7746 83808 8062 83809
rect 7746 83744 7752 83808
rect 7816 83744 7832 83808
rect 7896 83744 7912 83808
rect 7976 83744 7992 83808
rect 8056 83744 8062 83808
rect 7746 83743 8062 83744
rect 9346 83808 9662 83809
rect 9346 83744 9352 83808
rect 9416 83744 9432 83808
rect 9496 83744 9512 83808
rect 9576 83744 9592 83808
rect 9656 83744 9662 83808
rect 9346 83743 9662 83744
rect 59905 83738 59971 83741
rect 70209 83740 70275 83741
rect 60144 83738 60150 83740
rect 59905 83736 60150 83738
rect 59905 83680 59910 83736
rect 59966 83680 60150 83736
rect 59905 83678 60150 83680
rect 59905 83675 59971 83678
rect 60144 83676 60150 83678
rect 60214 83676 60220 83740
rect 70208 83676 70214 83740
rect 70278 83738 70284 83740
rect 70278 83678 70366 83738
rect 70278 83676 70284 83678
rect 70209 83675 70275 83676
rect 933 83466 999 83469
rect 0 83464 999 83466
rect 0 83408 938 83464
rect 994 83408 999 83464
rect 0 83406 999 83408
rect 933 83403 999 83406
rect 3606 83264 3922 83265
rect 3606 83200 3612 83264
rect 3676 83200 3692 83264
rect 3756 83200 3772 83264
rect 3836 83200 3852 83264
rect 3916 83200 3922 83264
rect 3606 83199 3922 83200
rect 5206 83264 5522 83265
rect 5206 83200 5212 83264
rect 5276 83200 5292 83264
rect 5356 83200 5372 83264
rect 5436 83200 5452 83264
rect 5516 83200 5522 83264
rect 5206 83199 5522 83200
rect 6806 83264 7122 83265
rect 6806 83200 6812 83264
rect 6876 83200 6892 83264
rect 6956 83200 6972 83264
rect 7036 83200 7052 83264
rect 7116 83200 7122 83264
rect 6806 83199 7122 83200
rect 8406 83264 8722 83265
rect 8406 83200 8412 83264
rect 8476 83200 8492 83264
rect 8556 83200 8572 83264
rect 8636 83200 8652 83264
rect 8716 83200 8722 83264
rect 8406 83199 8722 83200
rect 1485 82786 1551 82789
rect 798 82784 1551 82786
rect 798 82728 1490 82784
rect 1546 82728 1551 82784
rect 798 82726 1551 82728
rect 798 82514 858 82726
rect 1485 82723 1551 82726
rect 2946 82720 3262 82721
rect 2946 82656 2952 82720
rect 3016 82656 3032 82720
rect 3096 82656 3112 82720
rect 3176 82656 3192 82720
rect 3256 82656 3262 82720
rect 2946 82655 3262 82656
rect 4546 82720 4862 82721
rect 4546 82656 4552 82720
rect 4616 82656 4632 82720
rect 4696 82656 4712 82720
rect 4776 82656 4792 82720
rect 4856 82656 4862 82720
rect 4546 82655 4862 82656
rect 6146 82720 6462 82721
rect 6146 82656 6152 82720
rect 6216 82656 6232 82720
rect 6296 82656 6312 82720
rect 6376 82656 6392 82720
rect 6456 82656 6462 82720
rect 6146 82655 6462 82656
rect 7746 82720 8062 82721
rect 7746 82656 7752 82720
rect 7816 82656 7832 82720
rect 7896 82656 7912 82720
rect 7976 82656 7992 82720
rect 8056 82656 8062 82720
rect 7746 82655 8062 82656
rect 9346 82720 9662 82721
rect 9346 82656 9352 82720
rect 9416 82656 9432 82720
rect 9496 82656 9512 82720
rect 9576 82656 9592 82720
rect 9656 82656 9662 82720
rect 9346 82655 9662 82656
rect 0 82454 858 82514
rect 3606 82176 3922 82177
rect 3606 82112 3612 82176
rect 3676 82112 3692 82176
rect 3756 82112 3772 82176
rect 3836 82112 3852 82176
rect 3916 82112 3922 82176
rect 3606 82111 3922 82112
rect 5206 82176 5522 82177
rect 5206 82112 5212 82176
rect 5276 82112 5292 82176
rect 5356 82112 5372 82176
rect 5436 82112 5452 82176
rect 5516 82112 5522 82176
rect 5206 82111 5522 82112
rect 6806 82176 7122 82177
rect 6806 82112 6812 82176
rect 6876 82112 6892 82176
rect 6956 82112 6972 82176
rect 7036 82112 7052 82176
rect 7116 82112 7122 82176
rect 6806 82111 7122 82112
rect 8406 82176 8722 82177
rect 8406 82112 8412 82176
rect 8476 82112 8492 82176
rect 8556 82112 8572 82176
rect 8636 82112 8652 82176
rect 8716 82112 8722 82176
rect 8406 82111 8722 82112
rect 2946 81632 3262 81633
rect 2946 81568 2952 81632
rect 3016 81568 3032 81632
rect 3096 81568 3112 81632
rect 3176 81568 3192 81632
rect 3256 81568 3262 81632
rect 2946 81567 3262 81568
rect 4546 81632 4862 81633
rect 4546 81568 4552 81632
rect 4616 81568 4632 81632
rect 4696 81568 4712 81632
rect 4776 81568 4792 81632
rect 4856 81568 4862 81632
rect 4546 81567 4862 81568
rect 6146 81632 6462 81633
rect 6146 81568 6152 81632
rect 6216 81568 6232 81632
rect 6296 81568 6312 81632
rect 6376 81568 6392 81632
rect 6456 81568 6462 81632
rect 6146 81567 6462 81568
rect 7746 81632 8062 81633
rect 7746 81568 7752 81632
rect 7816 81568 7832 81632
rect 7896 81568 7912 81632
rect 7976 81568 7992 81632
rect 8056 81568 8062 81632
rect 7746 81567 8062 81568
rect 9346 81632 9662 81633
rect 9346 81568 9352 81632
rect 9416 81568 9432 81632
rect 9496 81568 9512 81632
rect 9576 81568 9592 81632
rect 9656 81568 9662 81632
rect 9346 81567 9662 81568
rect 933 81562 999 81565
rect 0 81560 999 81562
rect 0 81504 938 81560
rect 994 81504 999 81560
rect 0 81502 999 81504
rect 933 81499 999 81502
rect 3606 81088 3922 81089
rect 3606 81024 3612 81088
rect 3676 81024 3692 81088
rect 3756 81024 3772 81088
rect 3836 81024 3852 81088
rect 3916 81024 3922 81088
rect 3606 81023 3922 81024
rect 5206 81088 5522 81089
rect 5206 81024 5212 81088
rect 5276 81024 5292 81088
rect 5356 81024 5372 81088
rect 5436 81024 5452 81088
rect 5516 81024 5522 81088
rect 5206 81023 5522 81024
rect 6806 81088 7122 81089
rect 6806 81024 6812 81088
rect 6876 81024 6892 81088
rect 6956 81024 6972 81088
rect 7036 81024 7052 81088
rect 7116 81024 7122 81088
rect 6806 81023 7122 81024
rect 8406 81088 8722 81089
rect 8406 81024 8412 81088
rect 8476 81024 8492 81088
rect 8556 81024 8572 81088
rect 8636 81024 8652 81088
rect 8716 81024 8722 81088
rect 8406 81023 8722 81024
rect 933 80610 999 80613
rect 0 80608 999 80610
rect 0 80552 938 80608
rect 994 80552 999 80608
rect 0 80550 999 80552
rect 933 80547 999 80550
rect 2946 80544 3262 80545
rect 2946 80480 2952 80544
rect 3016 80480 3032 80544
rect 3096 80480 3112 80544
rect 3176 80480 3192 80544
rect 3256 80480 3262 80544
rect 2946 80479 3262 80480
rect 4546 80544 4862 80545
rect 4546 80480 4552 80544
rect 4616 80480 4632 80544
rect 4696 80480 4712 80544
rect 4776 80480 4792 80544
rect 4856 80480 4862 80544
rect 4546 80479 4862 80480
rect 6146 80544 6462 80545
rect 6146 80480 6152 80544
rect 6216 80480 6232 80544
rect 6296 80480 6312 80544
rect 6376 80480 6392 80544
rect 6456 80480 6462 80544
rect 6146 80479 6462 80480
rect 7746 80544 8062 80545
rect 7746 80480 7752 80544
rect 7816 80480 7832 80544
rect 7896 80480 7912 80544
rect 7976 80480 7992 80544
rect 8056 80480 8062 80544
rect 7746 80479 8062 80480
rect 9346 80544 9662 80545
rect 9346 80480 9352 80544
rect 9416 80480 9432 80544
rect 9496 80480 9512 80544
rect 9576 80480 9592 80544
rect 9656 80480 9662 80544
rect 108021 80500 108087 80503
rect 9346 80479 9662 80480
rect 107924 80498 108087 80500
rect 107924 80442 108026 80498
rect 108082 80442 108087 80498
rect 107924 80440 108087 80442
rect 108021 80437 108087 80440
rect 3606 80000 3922 80001
rect 3606 79936 3612 80000
rect 3676 79936 3692 80000
rect 3756 79936 3772 80000
rect 3836 79936 3852 80000
rect 3916 79936 3922 80000
rect 3606 79935 3922 79936
rect 5206 80000 5522 80001
rect 5206 79936 5212 80000
rect 5276 79936 5292 80000
rect 5356 79936 5372 80000
rect 5436 79936 5452 80000
rect 5516 79936 5522 80000
rect 5206 79935 5522 79936
rect 6806 80000 7122 80001
rect 6806 79936 6812 80000
rect 6876 79936 6892 80000
rect 6956 79936 6972 80000
rect 7036 79936 7052 80000
rect 7116 79936 7122 80000
rect 6806 79935 7122 79936
rect 8406 80000 8722 80001
rect 8406 79936 8412 80000
rect 8476 79936 8492 80000
rect 8556 79936 8572 80000
rect 8636 79936 8652 80000
rect 8716 79936 8722 80000
rect 8406 79935 8722 79936
rect 933 79658 999 79661
rect 0 79656 999 79658
rect 0 79600 938 79656
rect 994 79600 999 79656
rect 0 79598 999 79600
rect 933 79595 999 79598
rect 2946 79456 3262 79457
rect 2946 79392 2952 79456
rect 3016 79392 3032 79456
rect 3096 79392 3112 79456
rect 3176 79392 3192 79456
rect 3256 79392 3262 79456
rect 2946 79391 3262 79392
rect 4546 79456 4862 79457
rect 4546 79392 4552 79456
rect 4616 79392 4632 79456
rect 4696 79392 4712 79456
rect 4776 79392 4792 79456
rect 4856 79392 4862 79456
rect 4546 79391 4862 79392
rect 6146 79456 6462 79457
rect 6146 79392 6152 79456
rect 6216 79392 6232 79456
rect 6296 79392 6312 79456
rect 6376 79392 6392 79456
rect 6456 79392 6462 79456
rect 6146 79391 6462 79392
rect 7746 79456 8062 79457
rect 7746 79392 7752 79456
rect 7816 79392 7832 79456
rect 7896 79392 7912 79456
rect 7976 79392 7992 79456
rect 8056 79392 8062 79456
rect 7746 79391 8062 79392
rect 9346 79456 9662 79457
rect 9346 79392 9352 79456
rect 9416 79392 9432 79456
rect 9496 79392 9512 79456
rect 9576 79392 9592 79456
rect 9656 79392 9662 79456
rect 9346 79391 9662 79392
rect 3606 78912 3922 78913
rect 3606 78848 3612 78912
rect 3676 78848 3692 78912
rect 3756 78848 3772 78912
rect 3836 78848 3852 78912
rect 3916 78848 3922 78912
rect 3606 78847 3922 78848
rect 5206 78912 5522 78913
rect 5206 78848 5212 78912
rect 5276 78848 5292 78912
rect 5356 78848 5372 78912
rect 5436 78848 5452 78912
rect 5516 78848 5522 78912
rect 5206 78847 5522 78848
rect 6806 78912 7122 78913
rect 6806 78848 6812 78912
rect 6876 78848 6892 78912
rect 6956 78848 6972 78912
rect 7036 78848 7052 78912
rect 7116 78848 7122 78912
rect 6806 78847 7122 78848
rect 8406 78912 8722 78913
rect 8406 78848 8412 78912
rect 8476 78848 8492 78912
rect 8556 78848 8572 78912
rect 8636 78848 8652 78912
rect 8716 78848 8722 78912
rect 8406 78847 8722 78848
rect 933 78706 999 78709
rect 0 78704 999 78706
rect 0 78648 938 78704
rect 994 78648 999 78704
rect 0 78646 999 78648
rect 933 78643 999 78646
rect 2946 78368 3262 78369
rect 2946 78304 2952 78368
rect 3016 78304 3032 78368
rect 3096 78304 3112 78368
rect 3176 78304 3192 78368
rect 3256 78304 3262 78368
rect 2946 78303 3262 78304
rect 4546 78368 4862 78369
rect 4546 78304 4552 78368
rect 4616 78304 4632 78368
rect 4696 78304 4712 78368
rect 4776 78304 4792 78368
rect 4856 78304 4862 78368
rect 4546 78303 4862 78304
rect 6146 78368 6462 78369
rect 6146 78304 6152 78368
rect 6216 78304 6232 78368
rect 6296 78304 6312 78368
rect 6376 78304 6392 78368
rect 6456 78304 6462 78368
rect 6146 78303 6462 78304
rect 7746 78368 8062 78369
rect 7746 78304 7752 78368
rect 7816 78304 7832 78368
rect 7896 78304 7912 78368
rect 7976 78304 7992 78368
rect 8056 78304 8062 78368
rect 7746 78303 8062 78304
rect 9346 78368 9662 78369
rect 9346 78304 9352 78368
rect 9416 78304 9432 78368
rect 9496 78304 9512 78368
rect 9576 78304 9592 78368
rect 9656 78304 9662 78368
rect 9346 78303 9662 78304
rect 3606 77824 3922 77825
rect 3606 77760 3612 77824
rect 3676 77760 3692 77824
rect 3756 77760 3772 77824
rect 3836 77760 3852 77824
rect 3916 77760 3922 77824
rect 3606 77759 3922 77760
rect 5206 77824 5522 77825
rect 5206 77760 5212 77824
rect 5276 77760 5292 77824
rect 5356 77760 5372 77824
rect 5436 77760 5452 77824
rect 5516 77760 5522 77824
rect 5206 77759 5522 77760
rect 6806 77824 7122 77825
rect 6806 77760 6812 77824
rect 6876 77760 6892 77824
rect 6956 77760 6972 77824
rect 7036 77760 7052 77824
rect 7116 77760 7122 77824
rect 6806 77759 7122 77760
rect 8406 77824 8722 77825
rect 8406 77760 8412 77824
rect 8476 77760 8492 77824
rect 8556 77760 8572 77824
rect 8636 77760 8652 77824
rect 8716 77760 8722 77824
rect 8406 77759 8722 77760
rect 933 77754 999 77757
rect 0 77752 999 77754
rect 0 77696 938 77752
rect 994 77696 999 77752
rect 0 77694 999 77696
rect 933 77691 999 77694
rect 2946 77280 3262 77281
rect 2946 77216 2952 77280
rect 3016 77216 3032 77280
rect 3096 77216 3112 77280
rect 3176 77216 3192 77280
rect 3256 77216 3262 77280
rect 2946 77215 3262 77216
rect 4546 77280 4862 77281
rect 4546 77216 4552 77280
rect 4616 77216 4632 77280
rect 4696 77216 4712 77280
rect 4776 77216 4792 77280
rect 4856 77216 4862 77280
rect 4546 77215 4862 77216
rect 6146 77280 6462 77281
rect 6146 77216 6152 77280
rect 6216 77216 6232 77280
rect 6296 77216 6312 77280
rect 6376 77216 6392 77280
rect 6456 77216 6462 77280
rect 6146 77215 6462 77216
rect 7746 77280 8062 77281
rect 7746 77216 7752 77280
rect 7816 77216 7832 77280
rect 7896 77216 7912 77280
rect 7976 77216 7992 77280
rect 8056 77216 8062 77280
rect 7746 77215 8062 77216
rect 9346 77280 9662 77281
rect 9346 77216 9352 77280
rect 9416 77216 9432 77280
rect 9496 77216 9512 77280
rect 9576 77216 9592 77280
rect 9656 77216 9662 77280
rect 9346 77215 9662 77216
rect 933 76802 999 76805
rect 0 76800 999 76802
rect 0 76744 938 76800
rect 994 76744 999 76800
rect 0 76742 999 76744
rect 933 76739 999 76742
rect 3606 76736 3922 76737
rect 3606 76672 3612 76736
rect 3676 76672 3692 76736
rect 3756 76672 3772 76736
rect 3836 76672 3852 76736
rect 3916 76672 3922 76736
rect 3606 76671 3922 76672
rect 5206 76736 5522 76737
rect 5206 76672 5212 76736
rect 5276 76672 5292 76736
rect 5356 76672 5372 76736
rect 5436 76672 5452 76736
rect 5516 76672 5522 76736
rect 5206 76671 5522 76672
rect 6806 76736 7122 76737
rect 6806 76672 6812 76736
rect 6876 76672 6892 76736
rect 6956 76672 6972 76736
rect 7036 76672 7052 76736
rect 7116 76672 7122 76736
rect 6806 76671 7122 76672
rect 8406 76736 8722 76737
rect 8406 76672 8412 76736
rect 8476 76672 8492 76736
rect 8556 76672 8572 76736
rect 8636 76672 8652 76736
rect 8716 76672 8722 76736
rect 8406 76671 8722 76672
rect 2946 76192 3262 76193
rect 2946 76128 2952 76192
rect 3016 76128 3032 76192
rect 3096 76128 3112 76192
rect 3176 76128 3192 76192
rect 3256 76128 3262 76192
rect 2946 76127 3262 76128
rect 4546 76192 4862 76193
rect 4546 76128 4552 76192
rect 4616 76128 4632 76192
rect 4696 76128 4712 76192
rect 4776 76128 4792 76192
rect 4856 76128 4862 76192
rect 4546 76127 4862 76128
rect 6146 76192 6462 76193
rect 6146 76128 6152 76192
rect 6216 76128 6232 76192
rect 6296 76128 6312 76192
rect 6376 76128 6392 76192
rect 6456 76128 6462 76192
rect 6146 76127 6462 76128
rect 7746 76192 8062 76193
rect 7746 76128 7752 76192
rect 7816 76128 7832 76192
rect 7896 76128 7912 76192
rect 7976 76128 7992 76192
rect 8056 76128 8062 76192
rect 7746 76127 8062 76128
rect 9346 76192 9662 76193
rect 9346 76128 9352 76192
rect 9416 76128 9432 76192
rect 9496 76128 9512 76192
rect 9576 76128 9592 76192
rect 9656 76128 9662 76192
rect 9346 76127 9662 76128
rect 1485 75850 1551 75853
rect 0 75848 1551 75850
rect 0 75792 1490 75848
rect 1546 75792 1551 75848
rect 0 75790 1551 75792
rect 1485 75787 1551 75790
rect 3606 75648 3922 75649
rect 3606 75584 3612 75648
rect 3676 75584 3692 75648
rect 3756 75584 3772 75648
rect 3836 75584 3852 75648
rect 3916 75584 3922 75648
rect 3606 75583 3922 75584
rect 5206 75648 5522 75649
rect 5206 75584 5212 75648
rect 5276 75584 5292 75648
rect 5356 75584 5372 75648
rect 5436 75584 5452 75648
rect 5516 75584 5522 75648
rect 5206 75583 5522 75584
rect 6806 75648 7122 75649
rect 6806 75584 6812 75648
rect 6876 75584 6892 75648
rect 6956 75584 6972 75648
rect 7036 75584 7052 75648
rect 7116 75584 7122 75648
rect 6806 75583 7122 75584
rect 8406 75648 8722 75649
rect 8406 75584 8412 75648
rect 8476 75584 8492 75648
rect 8556 75584 8572 75648
rect 8636 75584 8652 75648
rect 8716 75584 8722 75648
rect 8406 75583 8722 75584
rect 2946 75104 3262 75105
rect 2946 75040 2952 75104
rect 3016 75040 3032 75104
rect 3096 75040 3112 75104
rect 3176 75040 3192 75104
rect 3256 75040 3262 75104
rect 2946 75039 3262 75040
rect 4546 75104 4862 75105
rect 4546 75040 4552 75104
rect 4616 75040 4632 75104
rect 4696 75040 4712 75104
rect 4776 75040 4792 75104
rect 4856 75040 4862 75104
rect 4546 75039 4862 75040
rect 6146 75104 6462 75105
rect 6146 75040 6152 75104
rect 6216 75040 6232 75104
rect 6296 75040 6312 75104
rect 6376 75040 6392 75104
rect 6456 75040 6462 75104
rect 6146 75039 6462 75040
rect 7746 75104 8062 75105
rect 7746 75040 7752 75104
rect 7816 75040 7832 75104
rect 7896 75040 7912 75104
rect 7976 75040 7992 75104
rect 8056 75040 8062 75104
rect 7746 75039 8062 75040
rect 9346 75104 9662 75105
rect 9346 75040 9352 75104
rect 9416 75040 9432 75104
rect 9496 75040 9512 75104
rect 9576 75040 9592 75104
rect 9656 75040 9662 75104
rect 9346 75039 9662 75040
rect 933 74898 999 74901
rect 0 74896 999 74898
rect 0 74840 938 74896
rect 994 74840 999 74896
rect 0 74838 999 74840
rect 933 74835 999 74838
rect 7281 74624 7347 74629
rect 7281 74568 7286 74624
rect 7342 74568 7347 74624
rect 7281 74563 7347 74568
rect 3606 74560 3922 74561
rect 3606 74496 3612 74560
rect 3676 74496 3692 74560
rect 3756 74496 3772 74560
rect 3836 74496 3852 74560
rect 3916 74496 3922 74560
rect 3606 74495 3922 74496
rect 5206 74560 5522 74561
rect 5206 74496 5212 74560
rect 5276 74496 5292 74560
rect 5356 74496 5372 74560
rect 5436 74496 5452 74560
rect 5516 74496 5522 74560
rect 5206 74495 5522 74496
rect 6806 74560 7122 74561
rect 6806 74496 6812 74560
rect 6876 74496 6892 74560
rect 6956 74496 6972 74560
rect 7036 74496 7052 74560
rect 7116 74496 7122 74560
rect 6806 74495 7122 74496
rect 2946 74016 3262 74017
rect 2946 73952 2952 74016
rect 3016 73952 3032 74016
rect 3096 73952 3112 74016
rect 3176 73952 3192 74016
rect 3256 73952 3262 74016
rect 2946 73951 3262 73952
rect 4546 74016 4862 74017
rect 4546 73952 4552 74016
rect 4616 73952 4632 74016
rect 4696 73952 4712 74016
rect 4776 73952 4792 74016
rect 4856 73952 4862 74016
rect 4546 73951 4862 73952
rect 6146 74016 6462 74017
rect 6146 73952 6152 74016
rect 6216 73952 6232 74016
rect 6296 73952 6312 74016
rect 6376 73952 6392 74016
rect 6456 73952 6462 74016
rect 6146 73951 6462 73952
rect 933 73946 999 73949
rect 0 73944 999 73946
rect 0 73888 938 73944
rect 994 73888 999 73944
rect 0 73886 999 73888
rect 933 73883 999 73886
rect 7284 73538 7344 74563
rect 8406 74560 8722 74561
rect 8406 74496 8412 74560
rect 8476 74496 8492 74560
rect 8556 74496 8572 74560
rect 8636 74496 8652 74560
rect 8716 74496 8722 74560
rect 8406 74495 8722 74496
rect 9949 74354 10015 74357
rect 10910 74354 10916 74356
rect 9949 74352 10916 74354
rect 9949 74296 9954 74352
rect 10010 74296 10916 74352
rect 9949 74294 10916 74296
rect 9949 74291 10015 74294
rect 10910 74292 10916 74294
rect 10980 74292 10986 74356
rect 7746 74016 8062 74017
rect 7746 73952 7752 74016
rect 7816 73952 7832 74016
rect 7896 73952 7912 74016
rect 7976 73952 7992 74016
rect 8056 73952 8062 74016
rect 7746 73951 8062 73952
rect 9346 74016 9662 74017
rect 9346 73952 9352 74016
rect 9416 73952 9432 74016
rect 9496 73952 9512 74016
rect 9576 73952 9592 74016
rect 9656 73952 9662 74016
rect 9346 73951 9662 73952
rect 9121 73674 9187 73677
rect 7606 73672 9187 73674
rect 7606 73616 9126 73672
rect 9182 73616 9187 73672
rect 7606 73614 9187 73616
rect 7465 73538 7531 73541
rect 7284 73536 7531 73538
rect 7284 73480 7470 73536
rect 7526 73480 7531 73536
rect 7284 73478 7531 73480
rect 7465 73475 7531 73478
rect 3606 73472 3922 73473
rect 3606 73408 3612 73472
rect 3676 73408 3692 73472
rect 3756 73408 3772 73472
rect 3836 73408 3852 73472
rect 3916 73408 3922 73472
rect 3606 73407 3922 73408
rect 5206 73472 5522 73473
rect 5206 73408 5212 73472
rect 5276 73408 5292 73472
rect 5356 73408 5372 73472
rect 5436 73408 5452 73472
rect 5516 73408 5522 73472
rect 5206 73407 5522 73408
rect 6806 73472 7122 73473
rect 6806 73408 6812 73472
rect 6876 73408 6892 73472
rect 6956 73408 6972 73472
rect 7036 73408 7052 73472
rect 7116 73408 7122 73472
rect 6806 73407 7122 73408
rect 7005 73266 7071 73269
rect 7606 73266 7666 73614
rect 9121 73611 9187 73614
rect 7741 73538 7807 73541
rect 8201 73538 8267 73541
rect 7741 73536 8267 73538
rect 7741 73480 7746 73536
rect 7802 73480 8206 73536
rect 8262 73480 8267 73536
rect 7741 73478 8267 73480
rect 7741 73475 7807 73478
rect 8201 73475 8267 73478
rect 8406 73472 8722 73473
rect 8406 73408 8412 73472
rect 8476 73408 8492 73472
rect 8556 73408 8572 73472
rect 8636 73408 8652 73472
rect 8716 73408 8722 73472
rect 8406 73407 8722 73408
rect 7005 73264 7666 73266
rect 7005 73208 7010 73264
rect 7066 73208 7666 73264
rect 7005 73206 7666 73208
rect 8109 73266 8175 73269
rect 8661 73266 8727 73269
rect 8109 73264 8727 73266
rect 8109 73208 8114 73264
rect 8170 73208 8666 73264
rect 8722 73208 8727 73264
rect 8109 73206 8727 73208
rect 7005 73203 7071 73206
rect 8109 73203 8175 73206
rect 8661 73203 8727 73206
rect 6729 73130 6795 73133
rect 8477 73130 8543 73133
rect 6729 73128 8543 73130
rect 6729 73072 6734 73128
rect 6790 73072 8482 73128
rect 8538 73072 8543 73128
rect 6729 73070 8543 73072
rect 6729 73067 6795 73070
rect 8477 73067 8543 73070
rect 933 72994 999 72997
rect 0 72992 999 72994
rect 0 72936 938 72992
rect 994 72936 999 72992
rect 0 72934 999 72936
rect 933 72931 999 72934
rect 2946 72928 3262 72929
rect 2946 72864 2952 72928
rect 3016 72864 3032 72928
rect 3096 72864 3112 72928
rect 3176 72864 3192 72928
rect 3256 72864 3262 72928
rect 2946 72863 3262 72864
rect 4546 72928 4862 72929
rect 4546 72864 4552 72928
rect 4616 72864 4632 72928
rect 4696 72864 4712 72928
rect 4776 72864 4792 72928
rect 4856 72864 4862 72928
rect 4546 72863 4862 72864
rect 6146 72928 6462 72929
rect 6146 72864 6152 72928
rect 6216 72864 6232 72928
rect 6296 72864 6312 72928
rect 6376 72864 6392 72928
rect 6456 72864 6462 72928
rect 6146 72863 6462 72864
rect 7746 72928 8062 72929
rect 7746 72864 7752 72928
rect 7816 72864 7832 72928
rect 7896 72864 7912 72928
rect 7976 72864 7992 72928
rect 8056 72864 8062 72928
rect 7746 72863 8062 72864
rect 9346 72928 9662 72929
rect 9346 72864 9352 72928
rect 9416 72864 9432 72928
rect 9496 72864 9512 72928
rect 9576 72864 9592 72928
rect 9656 72864 9662 72928
rect 9346 72863 9662 72864
rect 7189 72858 7255 72861
rect 7557 72858 7623 72861
rect 7189 72856 7623 72858
rect 7189 72800 7194 72856
rect 7250 72800 7562 72856
rect 7618 72800 7623 72856
rect 7189 72798 7623 72800
rect 7189 72795 7255 72798
rect 7557 72795 7623 72798
rect 6269 72722 6335 72725
rect 8385 72722 8451 72725
rect 6269 72720 8451 72722
rect 6269 72664 6274 72720
rect 6330 72664 8390 72720
rect 8446 72664 8451 72720
rect 6269 72662 8451 72664
rect 6269 72659 6335 72662
rect 8385 72659 8451 72662
rect 6821 72586 6887 72589
rect 9397 72586 9463 72589
rect 6821 72584 9463 72586
rect 6821 72528 6826 72584
rect 6882 72528 9402 72584
rect 9458 72528 9463 72584
rect 6821 72526 9463 72528
rect 6821 72523 6887 72526
rect 9397 72523 9463 72526
rect 3606 72384 3922 72385
rect 3606 72320 3612 72384
rect 3676 72320 3692 72384
rect 3756 72320 3772 72384
rect 3836 72320 3852 72384
rect 3916 72320 3922 72384
rect 3606 72319 3922 72320
rect 5206 72384 5522 72385
rect 5206 72320 5212 72384
rect 5276 72320 5292 72384
rect 5356 72320 5372 72384
rect 5436 72320 5452 72384
rect 5516 72320 5522 72384
rect 5206 72319 5522 72320
rect 6806 72384 7122 72385
rect 6806 72320 6812 72384
rect 6876 72320 6892 72384
rect 6956 72320 6972 72384
rect 7036 72320 7052 72384
rect 7116 72320 7122 72384
rect 6806 72319 7122 72320
rect 8406 72384 8722 72385
rect 8406 72320 8412 72384
rect 8476 72320 8492 72384
rect 8556 72320 8572 72384
rect 8636 72320 8652 72384
rect 8716 72320 8722 72384
rect 8406 72319 8722 72320
rect 5717 72176 5783 72181
rect 5717 72120 5722 72176
rect 5778 72120 5783 72176
rect 5717 72115 5783 72120
rect 7189 72178 7255 72181
rect 7925 72178 7991 72181
rect 7189 72176 7991 72178
rect 7189 72120 7194 72176
rect 7250 72120 7930 72176
rect 7986 72120 7991 72176
rect 7189 72118 7991 72120
rect 7189 72115 7255 72118
rect 7925 72115 7991 72118
rect 933 72042 999 72045
rect 0 72040 999 72042
rect 0 71984 938 72040
rect 994 71984 999 72040
rect 0 71982 999 71984
rect 933 71979 999 71982
rect 790 71844 796 71908
rect 860 71906 866 71908
rect 1577 71906 1643 71909
rect 860 71904 1643 71906
rect 860 71848 1582 71904
rect 1638 71848 1643 71904
rect 860 71846 1643 71848
rect 860 71844 866 71846
rect 1577 71843 1643 71846
rect 2946 71840 3262 71841
rect 2946 71776 2952 71840
rect 3016 71776 3032 71840
rect 3096 71776 3112 71840
rect 3176 71776 3192 71840
rect 3256 71776 3262 71840
rect 2946 71775 3262 71776
rect 4546 71840 4862 71841
rect 4546 71776 4552 71840
rect 4616 71776 4632 71840
rect 4696 71776 4712 71840
rect 4776 71776 4792 71840
rect 4856 71776 4862 71840
rect 4546 71775 4862 71776
rect 5720 71634 5780 72115
rect 6821 72042 6887 72045
rect 9397 72042 9463 72045
rect 6821 72040 9463 72042
rect 6821 71984 6826 72040
rect 6882 71984 9402 72040
rect 9458 71984 9463 72040
rect 6821 71982 9463 71984
rect 6821 71979 6887 71982
rect 9397 71979 9463 71982
rect 6146 71840 6462 71841
rect 6146 71776 6152 71840
rect 6216 71776 6232 71840
rect 6296 71776 6312 71840
rect 6376 71776 6392 71840
rect 6456 71776 6462 71840
rect 6146 71775 6462 71776
rect 7746 71840 8062 71841
rect 7746 71776 7752 71840
rect 7816 71776 7832 71840
rect 7896 71776 7912 71840
rect 7976 71776 7992 71840
rect 8056 71776 8062 71840
rect 7746 71775 8062 71776
rect 9346 71840 9662 71841
rect 9346 71776 9352 71840
rect 9416 71776 9432 71840
rect 9496 71776 9512 71840
rect 9576 71776 9592 71840
rect 9656 71776 9662 71840
rect 9346 71775 9662 71776
rect 7833 71634 7899 71637
rect 5720 71632 7899 71634
rect 5720 71576 7838 71632
rect 7894 71576 7899 71632
rect 5720 71574 7899 71576
rect 7833 71571 7899 71574
rect 2865 71498 2931 71501
rect 8385 71498 8451 71501
rect 2865 71496 8451 71498
rect 2865 71440 2870 71496
rect 2926 71440 8390 71496
rect 8446 71440 8451 71496
rect 2865 71438 8451 71440
rect 2865 71435 2931 71438
rect 8385 71435 8451 71438
rect 3606 71296 3922 71297
rect 3606 71232 3612 71296
rect 3676 71232 3692 71296
rect 3756 71232 3772 71296
rect 3836 71232 3852 71296
rect 3916 71232 3922 71296
rect 3606 71231 3922 71232
rect 5206 71296 5522 71297
rect 5206 71232 5212 71296
rect 5276 71232 5292 71296
rect 5356 71232 5372 71296
rect 5436 71232 5452 71296
rect 5516 71232 5522 71296
rect 5206 71231 5522 71232
rect 6806 71296 7122 71297
rect 6806 71232 6812 71296
rect 6876 71232 6892 71296
rect 6956 71232 6972 71296
rect 7036 71232 7052 71296
rect 7116 71232 7122 71296
rect 6806 71231 7122 71232
rect 8406 71296 8722 71297
rect 8406 71232 8412 71296
rect 8476 71232 8492 71296
rect 8556 71232 8572 71296
rect 8636 71232 8652 71296
rect 8716 71232 8722 71296
rect 8406 71231 8722 71232
rect 933 71090 999 71093
rect 0 71088 999 71090
rect 0 71032 938 71088
rect 994 71032 999 71088
rect 0 71030 999 71032
rect 933 71027 999 71030
rect 8477 71090 8543 71093
rect 10225 71090 10291 71093
rect 8477 71088 10291 71090
rect 8477 71032 8482 71088
rect 8538 71032 10230 71088
rect 10286 71032 10291 71088
rect 8477 71030 10291 71032
rect 8477 71027 8543 71030
rect 10225 71027 10291 71030
rect 6545 70954 6611 70957
rect 8201 70954 8267 70957
rect 9213 70954 9279 70957
rect 6545 70952 8267 70954
rect 6545 70896 6550 70952
rect 6606 70896 8206 70952
rect 8262 70896 8267 70952
rect 6545 70894 8267 70896
rect 6545 70891 6611 70894
rect 8201 70891 8267 70894
rect 9078 70952 9279 70954
rect 9078 70896 9218 70952
rect 9274 70896 9279 70952
rect 9078 70894 9279 70896
rect 2946 70752 3262 70753
rect 2946 70688 2952 70752
rect 3016 70688 3032 70752
rect 3096 70688 3112 70752
rect 3176 70688 3192 70752
rect 3256 70688 3262 70752
rect 2946 70687 3262 70688
rect 4546 70752 4862 70753
rect 4546 70688 4552 70752
rect 4616 70688 4632 70752
rect 4696 70688 4712 70752
rect 4776 70688 4792 70752
rect 4856 70688 4862 70752
rect 4546 70687 4862 70688
rect 6146 70752 6462 70753
rect 6146 70688 6152 70752
rect 6216 70688 6232 70752
rect 6296 70688 6312 70752
rect 6376 70688 6392 70752
rect 6456 70688 6462 70752
rect 6146 70687 6462 70688
rect 7746 70752 8062 70753
rect 7746 70688 7752 70752
rect 7816 70688 7832 70752
rect 7896 70688 7912 70752
rect 7976 70688 7992 70752
rect 8056 70688 8062 70752
rect 7746 70687 8062 70688
rect 5809 70546 5875 70549
rect 5766 70544 5875 70546
rect 5766 70488 5814 70544
rect 5870 70488 5875 70544
rect 5766 70483 5875 70488
rect 6913 70546 6979 70549
rect 7741 70546 7807 70549
rect 6913 70544 7807 70546
rect 6913 70488 6918 70544
rect 6974 70488 7746 70544
rect 7802 70488 7807 70544
rect 6913 70486 7807 70488
rect 6913 70483 6979 70486
rect 7741 70483 7807 70486
rect 8017 70546 8083 70549
rect 8477 70546 8543 70549
rect 8017 70544 8954 70546
rect 8017 70488 8022 70544
rect 8078 70488 8482 70544
rect 8538 70488 8954 70544
rect 8017 70486 8954 70488
rect 8017 70483 8083 70486
rect 8477 70483 8543 70486
rect 1393 70410 1459 70413
rect 1350 70408 1459 70410
rect 1350 70352 1398 70408
rect 1454 70352 1459 70408
rect 1350 70347 1459 70352
rect 4705 70410 4771 70413
rect 5766 70410 5826 70483
rect 8569 70410 8635 70413
rect 4705 70408 5642 70410
rect 4705 70352 4710 70408
rect 4766 70352 5642 70408
rect 4705 70350 5642 70352
rect 5766 70408 8635 70410
rect 5766 70352 8574 70408
rect 8630 70352 8635 70408
rect 5766 70350 8635 70352
rect 4705 70347 4771 70350
rect 1350 70138 1410 70347
rect 3606 70208 3922 70209
rect 3606 70144 3612 70208
rect 3676 70144 3692 70208
rect 3756 70144 3772 70208
rect 3836 70144 3852 70208
rect 3916 70144 3922 70208
rect 3606 70143 3922 70144
rect 5206 70208 5522 70209
rect 5206 70144 5212 70208
rect 5276 70144 5292 70208
rect 5356 70144 5372 70208
rect 5436 70144 5452 70208
rect 5516 70144 5522 70208
rect 5206 70143 5522 70144
rect 0 70078 1410 70138
rect 2681 70002 2747 70005
rect 5349 70002 5415 70005
rect 2681 70000 5415 70002
rect 2681 69944 2686 70000
rect 2742 69944 5354 70000
rect 5410 69944 5415 70000
rect 2681 69942 5415 69944
rect 5582 70002 5642 70350
rect 8569 70347 8635 70350
rect 6806 70208 7122 70209
rect 6806 70144 6812 70208
rect 6876 70144 6892 70208
rect 6956 70144 6972 70208
rect 7036 70144 7052 70208
rect 7116 70144 7122 70208
rect 6806 70143 7122 70144
rect 8406 70208 8722 70209
rect 8406 70144 8412 70208
rect 8476 70144 8492 70208
rect 8556 70144 8572 70208
rect 8636 70144 8652 70208
rect 8716 70144 8722 70208
rect 8406 70143 8722 70144
rect 8894 70138 8954 70486
rect 9078 70277 9138 70894
rect 9213 70891 9279 70894
rect 9346 70752 9662 70753
rect 9346 70688 9352 70752
rect 9416 70688 9432 70752
rect 9496 70688 9512 70752
rect 9576 70688 9592 70752
rect 9656 70688 9662 70752
rect 9346 70687 9662 70688
rect 9078 70272 9187 70277
rect 9078 70216 9126 70272
rect 9182 70216 9187 70272
rect 9078 70214 9187 70216
rect 9121 70211 9187 70214
rect 9305 70138 9371 70141
rect 8894 70136 9371 70138
rect 8894 70080 9310 70136
rect 9366 70080 9371 70136
rect 8894 70078 9371 70080
rect 9305 70075 9371 70078
rect 9581 70002 9647 70005
rect 5582 70000 9647 70002
rect 5582 69944 9586 70000
rect 9642 69944 9647 70000
rect 5582 69942 9647 69944
rect 2681 69939 2747 69942
rect 5349 69939 5415 69942
rect 9581 69939 9647 69942
rect 2589 69866 2655 69869
rect 10542 69866 10548 69868
rect 2589 69864 10548 69866
rect 2589 69808 2594 69864
rect 2650 69808 10548 69864
rect 2589 69806 10548 69808
rect 2589 69803 2655 69806
rect 10542 69804 10548 69806
rect 10612 69804 10618 69868
rect 2946 69664 3262 69665
rect 2946 69600 2952 69664
rect 3016 69600 3032 69664
rect 3096 69600 3112 69664
rect 3176 69600 3192 69664
rect 3256 69600 3262 69664
rect 2946 69599 3262 69600
rect 4546 69664 4862 69665
rect 4546 69600 4552 69664
rect 4616 69600 4632 69664
rect 4696 69600 4712 69664
rect 4776 69600 4792 69664
rect 4856 69600 4862 69664
rect 4546 69599 4862 69600
rect 6146 69664 6462 69665
rect 6146 69600 6152 69664
rect 6216 69600 6232 69664
rect 6296 69600 6312 69664
rect 6376 69600 6392 69664
rect 6456 69600 6462 69664
rect 6146 69599 6462 69600
rect 7746 69664 8062 69665
rect 7746 69600 7752 69664
rect 7816 69600 7832 69664
rect 7896 69600 7912 69664
rect 7976 69600 7992 69664
rect 8056 69600 8062 69664
rect 7746 69599 8062 69600
rect 9346 69664 9662 69665
rect 9346 69600 9352 69664
rect 9416 69600 9432 69664
rect 9496 69600 9512 69664
rect 9576 69600 9592 69664
rect 9656 69600 9662 69664
rect 9346 69599 9662 69600
rect 5349 69458 5415 69461
rect 11094 69458 11100 69460
rect 5349 69456 11100 69458
rect 5349 69400 5354 69456
rect 5410 69400 11100 69456
rect 5349 69398 11100 69400
rect 5349 69395 5415 69398
rect 11094 69396 11100 69398
rect 11164 69396 11170 69460
rect 2129 69322 2195 69325
rect 10501 69322 10567 69325
rect 2129 69320 10567 69322
rect 2129 69264 2134 69320
rect 2190 69264 10506 69320
rect 10562 69264 10567 69320
rect 2129 69262 10567 69264
rect 2129 69259 2195 69262
rect 10501 69259 10567 69262
rect 933 69186 999 69189
rect 0 69184 999 69186
rect 0 69128 938 69184
rect 994 69128 999 69184
rect 0 69126 999 69128
rect 933 69123 999 69126
rect 3606 69120 3922 69121
rect 3606 69056 3612 69120
rect 3676 69056 3692 69120
rect 3756 69056 3772 69120
rect 3836 69056 3852 69120
rect 3916 69056 3922 69120
rect 3606 69055 3922 69056
rect 5206 69120 5522 69121
rect 5206 69056 5212 69120
rect 5276 69056 5292 69120
rect 5356 69056 5372 69120
rect 5436 69056 5452 69120
rect 5516 69056 5522 69120
rect 5206 69055 5522 69056
rect 6806 69120 7122 69121
rect 6806 69056 6812 69120
rect 6876 69056 6892 69120
rect 6956 69056 6972 69120
rect 7036 69056 7052 69120
rect 7116 69056 7122 69120
rect 6806 69055 7122 69056
rect 8406 69120 8722 69121
rect 8406 69056 8412 69120
rect 8476 69056 8492 69120
rect 8556 69056 8572 69120
rect 8636 69056 8652 69120
rect 8716 69056 8722 69120
rect 8406 69055 8722 69056
rect 4153 68914 4219 68917
rect 8385 68914 8451 68917
rect 4153 68912 8451 68914
rect 4153 68856 4158 68912
rect 4214 68856 8390 68912
rect 8446 68856 8451 68912
rect 4153 68854 8451 68856
rect 4153 68851 4219 68854
rect 8385 68851 8451 68854
rect 8569 68914 8635 68917
rect 11462 68914 11468 68916
rect 8569 68912 11468 68914
rect 8569 68856 8574 68912
rect 8630 68856 11468 68912
rect 8569 68854 11468 68856
rect 8569 68851 8635 68854
rect 11462 68852 11468 68854
rect 11532 68852 11538 68916
rect 5717 68778 5783 68781
rect 5901 68778 5967 68781
rect 7373 68778 7439 68781
rect 5717 68776 5826 68778
rect 5717 68720 5722 68776
rect 5778 68720 5826 68776
rect 5717 68715 5826 68720
rect 5901 68776 7439 68778
rect 5901 68720 5906 68776
rect 5962 68720 7378 68776
rect 7434 68720 7439 68776
rect 5901 68718 7439 68720
rect 5901 68715 5967 68718
rect 7373 68715 7439 68718
rect 2946 68576 3262 68577
rect 2946 68512 2952 68576
rect 3016 68512 3032 68576
rect 3096 68512 3112 68576
rect 3176 68512 3192 68576
rect 3256 68512 3262 68576
rect 2946 68511 3262 68512
rect 4546 68576 4862 68577
rect 4546 68512 4552 68576
rect 4616 68512 4632 68576
rect 4696 68512 4712 68576
rect 4776 68512 4792 68576
rect 4856 68512 4862 68576
rect 4546 68511 4862 68512
rect 5766 68370 5826 68715
rect 6146 68576 6462 68577
rect 6146 68512 6152 68576
rect 6216 68512 6232 68576
rect 6296 68512 6312 68576
rect 6376 68512 6392 68576
rect 6456 68512 6462 68576
rect 6146 68511 6462 68512
rect 7746 68576 8062 68577
rect 7746 68512 7752 68576
rect 7816 68512 7832 68576
rect 7896 68512 7912 68576
rect 7976 68512 7992 68576
rect 8056 68512 8062 68576
rect 7746 68511 8062 68512
rect 9346 68576 9662 68577
rect 9346 68512 9352 68576
rect 9416 68512 9432 68576
rect 9496 68512 9512 68576
rect 9576 68512 9592 68576
rect 9656 68512 9662 68576
rect 9346 68511 9662 68512
rect 6085 68370 6151 68373
rect 9121 68370 9187 68373
rect 5766 68368 6151 68370
rect 5766 68312 6090 68368
rect 6146 68312 6151 68368
rect 5766 68310 6151 68312
rect 6085 68307 6151 68310
rect 6318 68368 9187 68370
rect 6318 68312 9126 68368
rect 9182 68312 9187 68368
rect 6318 68310 9187 68312
rect 933 68234 999 68237
rect 0 68232 999 68234
rect 0 68176 938 68232
rect 994 68176 999 68232
rect 0 68174 999 68176
rect 933 68171 999 68174
rect 2773 68234 2839 68237
rect 6318 68234 6378 68310
rect 9121 68307 9187 68310
rect 6913 68234 6979 68237
rect 2773 68232 6378 68234
rect 2773 68176 2778 68232
rect 2834 68176 6378 68232
rect 2773 68174 6378 68176
rect 6502 68232 6979 68234
rect 6502 68176 6918 68232
rect 6974 68176 6979 68232
rect 6502 68174 6979 68176
rect 2773 68171 2839 68174
rect 3606 68032 3922 68033
rect 3606 67968 3612 68032
rect 3676 67968 3692 68032
rect 3756 67968 3772 68032
rect 3836 67968 3852 68032
rect 3916 67968 3922 68032
rect 3606 67967 3922 67968
rect 5206 68032 5522 68033
rect 5206 67968 5212 68032
rect 5276 67968 5292 68032
rect 5356 67968 5372 68032
rect 5436 67968 5452 68032
rect 5516 67968 5522 68032
rect 5206 67967 5522 67968
rect 6502 67962 6562 68174
rect 6913 68171 6979 68174
rect 7925 68234 7991 68237
rect 8477 68234 8543 68237
rect 7925 68232 8543 68234
rect 7925 68176 7930 68232
rect 7986 68176 8482 68232
rect 8538 68176 8543 68232
rect 7925 68174 8543 68176
rect 7925 68171 7991 68174
rect 8477 68171 8543 68174
rect 6806 68032 7122 68033
rect 6806 67968 6812 68032
rect 6876 67968 6892 68032
rect 6956 67968 6972 68032
rect 7036 67968 7052 68032
rect 7116 67968 7122 68032
rect 6806 67967 7122 67968
rect 8406 68032 8722 68033
rect 8406 67968 8412 68032
rect 8476 67968 8492 68032
rect 8556 67968 8572 68032
rect 8636 67968 8652 68032
rect 8716 67968 8722 68032
rect 8406 67967 8722 67968
rect 5582 67902 6562 67962
rect 3877 67826 3943 67829
rect 4337 67826 4403 67829
rect 3877 67824 4403 67826
rect 3877 67768 3882 67824
rect 3938 67768 4342 67824
rect 4398 67768 4403 67824
rect 3877 67766 4403 67768
rect 3877 67763 3943 67766
rect 4337 67763 4403 67766
rect 4613 67826 4679 67829
rect 5582 67826 5642 67902
rect 4613 67824 5642 67826
rect 4613 67768 4618 67824
rect 4674 67768 5642 67824
rect 4613 67766 5642 67768
rect 4613 67763 4679 67766
rect 4521 67690 4587 67693
rect 4340 67688 4587 67690
rect 4340 67632 4526 67688
rect 4582 67632 4587 67688
rect 4340 67630 4587 67632
rect 1485 67554 1551 67557
rect 798 67552 1551 67554
rect 798 67496 1490 67552
rect 1546 67496 1551 67552
rect 798 67494 1551 67496
rect 798 67282 858 67494
rect 1485 67491 1551 67494
rect 2946 67488 3262 67489
rect 2946 67424 2952 67488
rect 3016 67424 3032 67488
rect 3096 67424 3112 67488
rect 3176 67424 3192 67488
rect 3256 67424 3262 67488
rect 2946 67423 3262 67424
rect 4340 67285 4400 67630
rect 4521 67627 4587 67630
rect 6177 67690 6243 67693
rect 9305 67690 9371 67693
rect 6177 67688 9371 67690
rect 6177 67632 6182 67688
rect 6238 67632 9310 67688
rect 9366 67632 9371 67688
rect 6177 67630 9371 67632
rect 6177 67627 6243 67630
rect 9305 67627 9371 67630
rect 4546 67488 4862 67489
rect 4546 67424 4552 67488
rect 4616 67424 4632 67488
rect 4696 67424 4712 67488
rect 4776 67424 4792 67488
rect 4856 67424 4862 67488
rect 4546 67423 4862 67424
rect 6146 67488 6462 67489
rect 6146 67424 6152 67488
rect 6216 67424 6232 67488
rect 6296 67424 6312 67488
rect 6376 67424 6392 67488
rect 6456 67424 6462 67488
rect 6146 67423 6462 67424
rect 7746 67488 8062 67489
rect 7746 67424 7752 67488
rect 7816 67424 7832 67488
rect 7896 67424 7912 67488
rect 7976 67424 7992 67488
rect 8056 67424 8062 67488
rect 7746 67423 8062 67424
rect 9346 67488 9662 67489
rect 9346 67424 9352 67488
rect 9416 67424 9432 67488
rect 9496 67424 9512 67488
rect 9576 67424 9592 67488
rect 9656 67424 9662 67488
rect 9346 67423 9662 67424
rect 8477 67418 8543 67421
rect 8158 67416 8543 67418
rect 8158 67360 8482 67416
rect 8538 67360 8543 67416
rect 8158 67358 8543 67360
rect 0 67222 858 67282
rect 4337 67280 4403 67285
rect 4337 67224 4342 67280
rect 4398 67224 4403 67280
rect 4337 67219 4403 67224
rect 6913 67282 6979 67285
rect 8158 67282 8218 67358
rect 8477 67355 8543 67358
rect 6913 67280 8218 67282
rect 6913 67224 6918 67280
rect 6974 67224 8218 67280
rect 6913 67222 8218 67224
rect 8569 67282 8635 67285
rect 9305 67282 9371 67285
rect 8569 67280 9371 67282
rect 8569 67224 8574 67280
rect 8630 67224 9310 67280
rect 9366 67224 9371 67280
rect 8569 67222 9371 67224
rect 6913 67219 6979 67222
rect 8569 67219 8635 67222
rect 9305 67219 9371 67222
rect 5349 67146 5415 67149
rect 9121 67146 9187 67149
rect 9397 67146 9463 67149
rect 5349 67144 9463 67146
rect 5349 67088 5354 67144
rect 5410 67088 9126 67144
rect 9182 67088 9402 67144
rect 9458 67088 9463 67144
rect 5349 67086 9463 67088
rect 5349 67083 5415 67086
rect 9121 67083 9187 67086
rect 9397 67083 9463 67086
rect 3606 66944 3922 66945
rect 3606 66880 3612 66944
rect 3676 66880 3692 66944
rect 3756 66880 3772 66944
rect 3836 66880 3852 66944
rect 3916 66880 3922 66944
rect 3606 66879 3922 66880
rect 5206 66944 5522 66945
rect 5206 66880 5212 66944
rect 5276 66880 5292 66944
rect 5356 66880 5372 66944
rect 5436 66880 5452 66944
rect 5516 66880 5522 66944
rect 5206 66879 5522 66880
rect 6806 66944 7122 66945
rect 6806 66880 6812 66944
rect 6876 66880 6892 66944
rect 6956 66880 6972 66944
rect 7036 66880 7052 66944
rect 7116 66880 7122 66944
rect 6806 66879 7122 66880
rect 8406 66944 8722 66945
rect 8406 66880 8412 66944
rect 8476 66880 8492 66944
rect 8556 66880 8572 66944
rect 8636 66880 8652 66944
rect 8716 66880 8722 66944
rect 8406 66879 8722 66880
rect 4521 66738 4587 66741
rect 4521 66736 8080 66738
rect 4521 66680 4526 66736
rect 4582 66680 8080 66736
rect 4521 66678 8080 66680
rect 4521 66675 4587 66678
rect 4705 66602 4771 66605
rect 4705 66600 5044 66602
rect 4705 66544 4710 66600
rect 4766 66544 5044 66600
rect 4705 66542 5044 66544
rect 4705 66539 4771 66542
rect 4337 66466 4403 66469
rect 4294 66464 4403 66466
rect 4294 66408 4342 66464
rect 4398 66408 4403 66464
rect 4294 66403 4403 66408
rect 2946 66400 3262 66401
rect 2946 66336 2952 66400
rect 3016 66336 3032 66400
rect 3096 66336 3112 66400
rect 3176 66336 3192 66400
rect 3256 66336 3262 66400
rect 2946 66335 3262 66336
rect 933 66330 999 66333
rect 0 66328 999 66330
rect 0 66272 938 66328
rect 994 66272 999 66328
rect 0 66270 999 66272
rect 933 66267 999 66270
rect 4294 66194 4354 66403
rect 4546 66400 4862 66401
rect 4546 66336 4552 66400
rect 4616 66336 4632 66400
rect 4696 66336 4712 66400
rect 4776 66336 4792 66400
rect 4856 66336 4862 66400
rect 4546 66335 4862 66336
rect 4613 66194 4679 66197
rect 4294 66192 4679 66194
rect 4294 66136 4618 66192
rect 4674 66136 4679 66192
rect 4294 66134 4679 66136
rect 4613 66131 4679 66134
rect 3606 65856 3922 65857
rect 3606 65792 3612 65856
rect 3676 65792 3692 65856
rect 3756 65792 3772 65856
rect 3836 65792 3852 65856
rect 3916 65792 3922 65856
rect 3606 65791 3922 65792
rect 2773 65784 2839 65789
rect 2773 65728 2778 65784
rect 2834 65728 2839 65784
rect 2773 65723 2839 65728
rect 2776 65381 2836 65723
rect 4984 65650 5044 66542
rect 8020 66568 8080 66678
rect 8342 66678 11898 66738
rect 8342 66568 8402 66678
rect 11838 66604 11898 66678
rect 8020 66508 8402 66568
rect 11830 66540 11836 66604
rect 11900 66540 11906 66604
rect 6146 66400 6462 66401
rect 6146 66336 6152 66400
rect 6216 66336 6232 66400
rect 6296 66336 6312 66400
rect 6376 66336 6392 66400
rect 6456 66336 6462 66400
rect 6146 66335 6462 66336
rect 7746 66400 8062 66401
rect 7746 66336 7752 66400
rect 7816 66336 7832 66400
rect 7896 66336 7912 66400
rect 7976 66336 7992 66400
rect 8056 66336 8062 66400
rect 7746 66335 8062 66336
rect 9346 66400 9662 66401
rect 9346 66336 9352 66400
rect 9416 66336 9432 66400
rect 9496 66336 9512 66400
rect 9576 66336 9592 66400
rect 9656 66336 9662 66400
rect 9346 66335 9662 66336
rect 7373 66058 7439 66061
rect 8477 66058 8543 66061
rect 7373 66056 8543 66058
rect 7373 66000 7378 66056
rect 7434 66000 8482 66056
rect 8538 66000 8543 66056
rect 7373 65998 8543 66000
rect 7373 65995 7439 65998
rect 8477 65995 8543 65998
rect 5206 65856 5522 65857
rect 5206 65792 5212 65856
rect 5276 65792 5292 65856
rect 5356 65792 5372 65856
rect 5436 65792 5452 65856
rect 5516 65792 5522 65856
rect 5206 65791 5522 65792
rect 6806 65856 7122 65857
rect 6806 65792 6812 65856
rect 6876 65792 6892 65856
rect 6956 65792 6972 65856
rect 7036 65792 7052 65856
rect 7116 65792 7122 65856
rect 6806 65791 7122 65792
rect 8406 65856 8722 65857
rect 8406 65792 8412 65856
rect 8476 65792 8492 65856
rect 8556 65792 8572 65856
rect 8636 65792 8652 65856
rect 8716 65792 8722 65856
rect 8406 65791 8722 65792
rect 5349 65650 5415 65653
rect 4984 65648 5415 65650
rect 4984 65592 5354 65648
rect 5410 65592 5415 65648
rect 4984 65590 5415 65592
rect 5349 65587 5415 65590
rect 933 65378 999 65381
rect 0 65376 999 65378
rect 0 65320 938 65376
rect 994 65320 999 65376
rect 0 65318 999 65320
rect 933 65315 999 65318
rect 2773 65376 2839 65381
rect 2773 65320 2778 65376
rect 2834 65320 2839 65376
rect 2773 65315 2839 65320
rect 2946 65312 3262 65313
rect 2946 65248 2952 65312
rect 3016 65248 3032 65312
rect 3096 65248 3112 65312
rect 3176 65248 3192 65312
rect 3256 65248 3262 65312
rect 2946 65247 3262 65248
rect 4546 65312 4862 65313
rect 4546 65248 4552 65312
rect 4616 65248 4632 65312
rect 4696 65248 4712 65312
rect 4776 65248 4792 65312
rect 4856 65248 4862 65312
rect 4546 65247 4862 65248
rect 6146 65312 6462 65313
rect 6146 65248 6152 65312
rect 6216 65248 6232 65312
rect 6296 65248 6312 65312
rect 6376 65248 6392 65312
rect 6456 65248 6462 65312
rect 6146 65247 6462 65248
rect 7746 65312 8062 65313
rect 7746 65248 7752 65312
rect 7816 65248 7832 65312
rect 7896 65248 7912 65312
rect 7976 65248 7992 65312
rect 8056 65248 8062 65312
rect 7746 65247 8062 65248
rect 9346 65312 9662 65313
rect 9346 65248 9352 65312
rect 9416 65248 9432 65312
rect 9496 65248 9512 65312
rect 9576 65248 9592 65312
rect 9656 65248 9662 65312
rect 9346 65247 9662 65248
rect 1117 65106 1183 65109
rect 1577 65106 1643 65109
rect 1117 65104 1643 65106
rect 1117 65048 1122 65104
rect 1178 65048 1582 65104
rect 1638 65048 1643 65104
rect 1117 65046 1643 65048
rect 1117 65043 1183 65046
rect 1577 65043 1643 65046
rect 2129 65106 2195 65109
rect 11881 65106 11947 65109
rect 2129 65104 11947 65106
rect 2129 65048 2134 65104
rect 2190 65048 11886 65104
rect 11942 65048 11947 65104
rect 2129 65046 11947 65048
rect 2129 65043 2195 65046
rect 11881 65043 11947 65046
rect 7005 64970 7071 64973
rect 6686 64968 7071 64970
rect 6686 64912 7010 64968
rect 7066 64912 7071 64968
rect 6686 64910 7071 64912
rect 3606 64768 3922 64769
rect 3606 64704 3612 64768
rect 3676 64704 3692 64768
rect 3756 64704 3772 64768
rect 3836 64704 3852 64768
rect 3916 64704 3922 64768
rect 3606 64703 3922 64704
rect 5206 64768 5522 64769
rect 5206 64704 5212 64768
rect 5276 64704 5292 64768
rect 5356 64704 5372 64768
rect 5436 64704 5452 64768
rect 5516 64704 5522 64768
rect 5206 64703 5522 64704
rect 6686 64562 6746 64910
rect 7005 64907 7071 64910
rect 6806 64768 7122 64769
rect 6806 64704 6812 64768
rect 6876 64704 6892 64768
rect 6956 64704 6972 64768
rect 7036 64704 7052 64768
rect 7116 64704 7122 64768
rect 6806 64703 7122 64704
rect 8406 64768 8722 64769
rect 8406 64704 8412 64768
rect 8476 64704 8492 64768
rect 8556 64704 8572 64768
rect 8636 64704 8652 64768
rect 8716 64704 8722 64768
rect 8406 64703 8722 64704
rect 6821 64562 6887 64565
rect 6686 64560 6887 64562
rect 6686 64504 6826 64560
rect 6882 64504 6887 64560
rect 6686 64502 6887 64504
rect 6821 64499 6887 64502
rect 933 64426 999 64429
rect 0 64424 999 64426
rect 0 64368 938 64424
rect 994 64368 999 64424
rect 0 64366 999 64368
rect 933 64363 999 64366
rect 2946 64224 3262 64225
rect 2946 64160 2952 64224
rect 3016 64160 3032 64224
rect 3096 64160 3112 64224
rect 3176 64160 3192 64224
rect 3256 64160 3262 64224
rect 2946 64159 3262 64160
rect 4546 64224 4862 64225
rect 4546 64160 4552 64224
rect 4616 64160 4632 64224
rect 4696 64160 4712 64224
rect 4776 64160 4792 64224
rect 4856 64160 4862 64224
rect 4546 64159 4862 64160
rect 6146 64224 6462 64225
rect 6146 64160 6152 64224
rect 6216 64160 6232 64224
rect 6296 64160 6312 64224
rect 6376 64160 6392 64224
rect 6456 64160 6462 64224
rect 6146 64159 6462 64160
rect 7746 64224 8062 64225
rect 7746 64160 7752 64224
rect 7816 64160 7832 64224
rect 7896 64160 7912 64224
rect 7976 64160 7992 64224
rect 8056 64160 8062 64224
rect 7746 64159 8062 64160
rect 9346 64224 9662 64225
rect 9346 64160 9352 64224
rect 9416 64160 9432 64224
rect 9496 64160 9512 64224
rect 9576 64160 9592 64224
rect 9656 64160 9662 64224
rect 9346 64159 9662 64160
rect 3606 63680 3922 63681
rect 3606 63616 3612 63680
rect 3676 63616 3692 63680
rect 3756 63616 3772 63680
rect 3836 63616 3852 63680
rect 3916 63616 3922 63680
rect 3606 63615 3922 63616
rect 5206 63680 5522 63681
rect 5206 63616 5212 63680
rect 5276 63616 5292 63680
rect 5356 63616 5372 63680
rect 5436 63616 5452 63680
rect 5516 63616 5522 63680
rect 5206 63615 5522 63616
rect 6806 63680 7122 63681
rect 6806 63616 6812 63680
rect 6876 63616 6892 63680
rect 6956 63616 6972 63680
rect 7036 63616 7052 63680
rect 7116 63616 7122 63680
rect 6806 63615 7122 63616
rect 8406 63680 8722 63681
rect 8406 63616 8412 63680
rect 8476 63616 8492 63680
rect 8556 63616 8572 63680
rect 8636 63616 8652 63680
rect 8716 63616 8722 63680
rect 8406 63615 8722 63616
rect 1485 63474 1551 63477
rect 0 63472 1551 63474
rect 0 63416 1490 63472
rect 1546 63416 1551 63472
rect 0 63414 1551 63416
rect 1485 63411 1551 63414
rect 8201 63474 8267 63477
rect 8201 63472 8954 63474
rect 8201 63416 8206 63472
rect 8262 63416 8954 63472
rect 8201 63414 8954 63416
rect 8201 63411 8267 63414
rect 8894 63341 8954 63414
rect 6545 63338 6611 63341
rect 8385 63338 8451 63341
rect 6545 63336 8451 63338
rect 6545 63280 6550 63336
rect 6606 63280 8390 63336
rect 8446 63280 8451 63336
rect 6545 63278 8451 63280
rect 8894 63336 9003 63341
rect 8894 63280 8942 63336
rect 8998 63280 9003 63336
rect 8894 63278 9003 63280
rect 6545 63275 6611 63278
rect 8385 63275 8451 63278
rect 8937 63275 9003 63278
rect 2946 63136 3262 63137
rect 2946 63072 2952 63136
rect 3016 63072 3032 63136
rect 3096 63072 3112 63136
rect 3176 63072 3192 63136
rect 3256 63072 3262 63136
rect 2946 63071 3262 63072
rect 4546 63136 4862 63137
rect 4546 63072 4552 63136
rect 4616 63072 4632 63136
rect 4696 63072 4712 63136
rect 4776 63072 4792 63136
rect 4856 63072 4862 63136
rect 4546 63071 4862 63072
rect 6146 63136 6462 63137
rect 6146 63072 6152 63136
rect 6216 63072 6232 63136
rect 6296 63072 6312 63136
rect 6376 63072 6392 63136
rect 6456 63072 6462 63136
rect 6146 63071 6462 63072
rect 7746 63136 8062 63137
rect 7746 63072 7752 63136
rect 7816 63072 7832 63136
rect 7896 63072 7912 63136
rect 7976 63072 7992 63136
rect 8056 63072 8062 63136
rect 7746 63071 8062 63072
rect 9346 63136 9662 63137
rect 9346 63072 9352 63136
rect 9416 63072 9432 63136
rect 9496 63072 9512 63136
rect 9576 63072 9592 63136
rect 9656 63072 9662 63136
rect 9346 63071 9662 63072
rect 3601 62930 3667 62933
rect 8661 62930 8727 62933
rect 3601 62928 8727 62930
rect 3601 62872 3606 62928
rect 3662 62872 8666 62928
rect 8722 62872 8727 62928
rect 3601 62870 8727 62872
rect 3601 62867 3667 62870
rect 8661 62867 8727 62870
rect 6821 62794 6887 62797
rect 6821 62792 7298 62794
rect 6821 62736 6826 62792
rect 6882 62736 7298 62792
rect 6821 62734 7298 62736
rect 6821 62731 6887 62734
rect 3606 62592 3922 62593
rect 3606 62528 3612 62592
rect 3676 62528 3692 62592
rect 3756 62528 3772 62592
rect 3836 62528 3852 62592
rect 3916 62528 3922 62592
rect 3606 62527 3922 62528
rect 5206 62592 5522 62593
rect 5206 62528 5212 62592
rect 5276 62528 5292 62592
rect 5356 62528 5372 62592
rect 5436 62528 5452 62592
rect 5516 62528 5522 62592
rect 5206 62527 5522 62528
rect 6806 62592 7122 62593
rect 6806 62528 6812 62592
rect 6876 62528 6892 62592
rect 6956 62528 6972 62592
rect 7036 62528 7052 62592
rect 7116 62528 7122 62592
rect 6806 62527 7122 62528
rect 933 62522 999 62525
rect 0 62520 999 62522
rect 0 62464 938 62520
rect 994 62464 999 62520
rect 0 62462 999 62464
rect 933 62459 999 62462
rect 7238 62253 7298 62734
rect 8406 62592 8722 62593
rect 8406 62528 8412 62592
rect 8476 62528 8492 62592
rect 8556 62528 8572 62592
rect 8636 62528 8652 62592
rect 8716 62528 8722 62592
rect 8406 62527 8722 62528
rect 7238 62248 7347 62253
rect 7238 62192 7286 62248
rect 7342 62192 7347 62248
rect 7238 62190 7347 62192
rect 7281 62187 7347 62190
rect 2946 62048 3262 62049
rect 2946 61984 2952 62048
rect 3016 61984 3032 62048
rect 3096 61984 3112 62048
rect 3176 61984 3192 62048
rect 3256 61984 3262 62048
rect 2946 61983 3262 61984
rect 4546 62048 4862 62049
rect 4546 61984 4552 62048
rect 4616 61984 4632 62048
rect 4696 61984 4712 62048
rect 4776 61984 4792 62048
rect 4856 61984 4862 62048
rect 4546 61983 4862 61984
rect 6146 62048 6462 62049
rect 6146 61984 6152 62048
rect 6216 61984 6232 62048
rect 6296 61984 6312 62048
rect 6376 61984 6392 62048
rect 6456 61984 6462 62048
rect 6146 61983 6462 61984
rect 7746 62048 8062 62049
rect 7746 61984 7752 62048
rect 7816 61984 7832 62048
rect 7896 61984 7912 62048
rect 7976 61984 7992 62048
rect 8056 61984 8062 62048
rect 7746 61983 8062 61984
rect 9346 62048 9662 62049
rect 9346 61984 9352 62048
rect 9416 61984 9432 62048
rect 9496 61984 9512 62048
rect 9576 61984 9592 62048
rect 9656 61984 9662 62048
rect 9346 61983 9662 61984
rect 933 61570 999 61573
rect 0 61568 999 61570
rect 0 61512 938 61568
rect 994 61512 999 61568
rect 0 61510 999 61512
rect 933 61507 999 61510
rect 3606 61504 3922 61505
rect 3606 61440 3612 61504
rect 3676 61440 3692 61504
rect 3756 61440 3772 61504
rect 3836 61440 3852 61504
rect 3916 61440 3922 61504
rect 3606 61439 3922 61440
rect 5206 61504 5522 61505
rect 5206 61440 5212 61504
rect 5276 61440 5292 61504
rect 5356 61440 5372 61504
rect 5436 61440 5452 61504
rect 5516 61440 5522 61504
rect 5206 61439 5522 61440
rect 6806 61504 7122 61505
rect 6806 61440 6812 61504
rect 6876 61440 6892 61504
rect 6956 61440 6972 61504
rect 7036 61440 7052 61504
rect 7116 61440 7122 61504
rect 6806 61439 7122 61440
rect 8406 61504 8722 61505
rect 8406 61440 8412 61504
rect 8476 61440 8492 61504
rect 8556 61440 8572 61504
rect 8636 61440 8652 61504
rect 8716 61440 8722 61504
rect 8406 61439 8722 61440
rect 2946 60960 3262 60961
rect 2946 60896 2952 60960
rect 3016 60896 3032 60960
rect 3096 60896 3112 60960
rect 3176 60896 3192 60960
rect 3256 60896 3262 60960
rect 2946 60895 3262 60896
rect 4546 60960 4862 60961
rect 4546 60896 4552 60960
rect 4616 60896 4632 60960
rect 4696 60896 4712 60960
rect 4776 60896 4792 60960
rect 4856 60896 4862 60960
rect 4546 60895 4862 60896
rect 6146 60960 6462 60961
rect 6146 60896 6152 60960
rect 6216 60896 6232 60960
rect 6296 60896 6312 60960
rect 6376 60896 6392 60960
rect 6456 60896 6462 60960
rect 6146 60895 6462 60896
rect 7746 60960 8062 60961
rect 7746 60896 7752 60960
rect 7816 60896 7832 60960
rect 7896 60896 7912 60960
rect 7976 60896 7992 60960
rect 8056 60896 8062 60960
rect 7746 60895 8062 60896
rect 9346 60960 9662 60961
rect 9346 60896 9352 60960
rect 9416 60896 9432 60960
rect 9496 60896 9512 60960
rect 9576 60896 9592 60960
rect 9656 60896 9662 60960
rect 9346 60895 9662 60896
rect 933 60618 999 60621
rect 0 60616 999 60618
rect 0 60560 938 60616
rect 994 60560 999 60616
rect 0 60558 999 60560
rect 933 60555 999 60558
rect 9029 60482 9095 60485
rect 8894 60480 9095 60482
rect 8894 60424 9034 60480
rect 9090 60424 9095 60480
rect 8894 60422 9095 60424
rect 3606 60416 3922 60417
rect 3606 60352 3612 60416
rect 3676 60352 3692 60416
rect 3756 60352 3772 60416
rect 3836 60352 3852 60416
rect 3916 60352 3922 60416
rect 3606 60351 3922 60352
rect 5206 60416 5522 60417
rect 5206 60352 5212 60416
rect 5276 60352 5292 60416
rect 5356 60352 5372 60416
rect 5436 60352 5452 60416
rect 5516 60352 5522 60416
rect 5206 60351 5522 60352
rect 6806 60416 7122 60417
rect 6806 60352 6812 60416
rect 6876 60352 6892 60416
rect 6956 60352 6972 60416
rect 7036 60352 7052 60416
rect 7116 60352 7122 60416
rect 6806 60351 7122 60352
rect 8406 60416 8722 60417
rect 8406 60352 8412 60416
rect 8476 60352 8492 60416
rect 8556 60352 8572 60416
rect 8636 60352 8652 60416
rect 8716 60352 8722 60416
rect 8406 60351 8722 60352
rect 8894 60213 8954 60422
rect 9029 60419 9095 60422
rect 8894 60208 9003 60213
rect 8894 60152 8942 60208
rect 8998 60152 9003 60208
rect 8894 60150 9003 60152
rect 8937 60147 9003 60150
rect 2946 59872 3262 59873
rect 2946 59808 2952 59872
rect 3016 59808 3032 59872
rect 3096 59808 3112 59872
rect 3176 59808 3192 59872
rect 3256 59808 3262 59872
rect 2946 59807 3262 59808
rect 4546 59872 4862 59873
rect 4546 59808 4552 59872
rect 4616 59808 4632 59872
rect 4696 59808 4712 59872
rect 4776 59808 4792 59872
rect 4856 59808 4862 59872
rect 4546 59807 4862 59808
rect 6146 59872 6462 59873
rect 6146 59808 6152 59872
rect 6216 59808 6232 59872
rect 6296 59808 6312 59872
rect 6376 59808 6392 59872
rect 6456 59808 6462 59872
rect 6146 59807 6462 59808
rect 7746 59872 8062 59873
rect 7746 59808 7752 59872
rect 7816 59808 7832 59872
rect 7896 59808 7912 59872
rect 7976 59808 7992 59872
rect 8056 59808 8062 59872
rect 7746 59807 8062 59808
rect 9346 59872 9662 59873
rect 9346 59808 9352 59872
rect 9416 59808 9432 59872
rect 9496 59808 9512 59872
rect 9576 59808 9592 59872
rect 9656 59808 9662 59872
rect 9346 59807 9662 59808
rect 933 59666 999 59669
rect 0 59664 999 59666
rect 0 59608 938 59664
rect 994 59608 999 59664
rect 0 59606 999 59608
rect 933 59603 999 59606
rect 3606 59328 3922 59329
rect 3606 59264 3612 59328
rect 3676 59264 3692 59328
rect 3756 59264 3772 59328
rect 3836 59264 3852 59328
rect 3916 59264 3922 59328
rect 3606 59263 3922 59264
rect 5206 59328 5522 59329
rect 5206 59264 5212 59328
rect 5276 59264 5292 59328
rect 5356 59264 5372 59328
rect 5436 59264 5452 59328
rect 5516 59264 5522 59328
rect 5206 59263 5522 59264
rect 6806 59328 7122 59329
rect 6806 59264 6812 59328
rect 6876 59264 6892 59328
rect 6956 59264 6972 59328
rect 7036 59264 7052 59328
rect 7116 59264 7122 59328
rect 6806 59263 7122 59264
rect 8406 59328 8722 59329
rect 8406 59264 8412 59328
rect 8476 59264 8492 59328
rect 8556 59264 8572 59328
rect 8636 59264 8652 59328
rect 8716 59264 8722 59328
rect 8406 59263 8722 59264
rect 2946 58784 3262 58785
rect 2946 58720 2952 58784
rect 3016 58720 3032 58784
rect 3096 58720 3112 58784
rect 3176 58720 3192 58784
rect 3256 58720 3262 58784
rect 2946 58719 3262 58720
rect 4546 58784 4862 58785
rect 4546 58720 4552 58784
rect 4616 58720 4632 58784
rect 4696 58720 4712 58784
rect 4776 58720 4792 58784
rect 4856 58720 4862 58784
rect 4546 58719 4862 58720
rect 6146 58784 6462 58785
rect 6146 58720 6152 58784
rect 6216 58720 6232 58784
rect 6296 58720 6312 58784
rect 6376 58720 6392 58784
rect 6456 58720 6462 58784
rect 6146 58719 6462 58720
rect 7746 58784 8062 58785
rect 7746 58720 7752 58784
rect 7816 58720 7832 58784
rect 7896 58720 7912 58784
rect 7976 58720 7992 58784
rect 8056 58720 8062 58784
rect 7746 58719 8062 58720
rect 9346 58784 9662 58785
rect 9346 58720 9352 58784
rect 9416 58720 9432 58784
rect 9496 58720 9512 58784
rect 9576 58720 9592 58784
rect 9656 58720 9662 58784
rect 9346 58719 9662 58720
rect 933 58714 999 58717
rect 0 58712 999 58714
rect 0 58656 938 58712
rect 994 58656 999 58712
rect 0 58654 999 58656
rect 933 58651 999 58654
rect 3606 58240 3922 58241
rect 3606 58176 3612 58240
rect 3676 58176 3692 58240
rect 3756 58176 3772 58240
rect 3836 58176 3852 58240
rect 3916 58176 3922 58240
rect 3606 58175 3922 58176
rect 5206 58240 5522 58241
rect 5206 58176 5212 58240
rect 5276 58176 5292 58240
rect 5356 58176 5372 58240
rect 5436 58176 5452 58240
rect 5516 58176 5522 58240
rect 5206 58175 5522 58176
rect 6806 58240 7122 58241
rect 6806 58176 6812 58240
rect 6876 58176 6892 58240
rect 6956 58176 6972 58240
rect 7036 58176 7052 58240
rect 7116 58176 7122 58240
rect 6806 58175 7122 58176
rect 8406 58240 8722 58241
rect 8406 58176 8412 58240
rect 8476 58176 8492 58240
rect 8556 58176 8572 58240
rect 8636 58176 8652 58240
rect 8716 58176 8722 58240
rect 8406 58175 8722 58176
rect 6453 57898 6519 57901
rect 8293 57898 8359 57901
rect 8845 57898 8911 57901
rect 9305 57898 9371 57901
rect 6453 57896 6746 57898
rect 6453 57840 6458 57896
rect 6514 57840 6746 57896
rect 6453 57838 6746 57840
rect 6453 57835 6519 57838
rect 1577 57762 1643 57765
rect 0 57760 1643 57762
rect 0 57704 1582 57760
rect 1638 57704 1643 57760
rect 0 57702 1643 57704
rect 1577 57699 1643 57702
rect 2946 57696 3262 57697
rect 2946 57632 2952 57696
rect 3016 57632 3032 57696
rect 3096 57632 3112 57696
rect 3176 57632 3192 57696
rect 3256 57632 3262 57696
rect 2946 57631 3262 57632
rect 4546 57696 4862 57697
rect 4546 57632 4552 57696
rect 4616 57632 4632 57696
rect 4696 57632 4712 57696
rect 4776 57632 4792 57696
rect 4856 57632 4862 57696
rect 4546 57631 4862 57632
rect 6146 57696 6462 57697
rect 6146 57632 6152 57696
rect 6216 57632 6232 57696
rect 6296 57632 6312 57696
rect 6376 57632 6392 57696
rect 6456 57632 6462 57696
rect 6146 57631 6462 57632
rect 6545 57490 6611 57493
rect 6686 57490 6746 57838
rect 8293 57896 8911 57898
rect 8293 57840 8298 57896
rect 8354 57840 8850 57896
rect 8906 57840 8911 57896
rect 8293 57838 8911 57840
rect 8293 57835 8359 57838
rect 8845 57835 8911 57838
rect 9078 57896 9371 57898
rect 9078 57840 9310 57896
rect 9366 57840 9371 57896
rect 9078 57838 9371 57840
rect 8201 57762 8267 57765
rect 9078 57762 9138 57838
rect 9305 57835 9371 57838
rect 8201 57760 9138 57762
rect 8201 57704 8206 57760
rect 8262 57704 9138 57760
rect 8201 57702 9138 57704
rect 8201 57699 8267 57702
rect 7746 57696 8062 57697
rect 7746 57632 7752 57696
rect 7816 57632 7832 57696
rect 7896 57632 7912 57696
rect 7976 57632 7992 57696
rect 8056 57632 8062 57696
rect 7746 57631 8062 57632
rect 9346 57696 9662 57697
rect 9346 57632 9352 57696
rect 9416 57632 9432 57696
rect 9496 57632 9512 57696
rect 9576 57632 9592 57696
rect 9656 57632 9662 57696
rect 9346 57631 9662 57632
rect 6545 57488 6746 57490
rect 6545 57432 6550 57488
rect 6606 57432 6746 57488
rect 6545 57430 6746 57432
rect 6545 57427 6611 57430
rect 3606 57152 3922 57153
rect 3606 57088 3612 57152
rect 3676 57088 3692 57152
rect 3756 57088 3772 57152
rect 3836 57088 3852 57152
rect 3916 57088 3922 57152
rect 3606 57087 3922 57088
rect 5206 57152 5522 57153
rect 5206 57088 5212 57152
rect 5276 57088 5292 57152
rect 5356 57088 5372 57152
rect 5436 57088 5452 57152
rect 5516 57088 5522 57152
rect 5206 57087 5522 57088
rect 6806 57152 7122 57153
rect 6806 57088 6812 57152
rect 6876 57088 6892 57152
rect 6956 57088 6972 57152
rect 7036 57088 7052 57152
rect 7116 57088 7122 57152
rect 6806 57087 7122 57088
rect 8406 57152 8722 57153
rect 8406 57088 8412 57152
rect 8476 57088 8492 57152
rect 8556 57088 8572 57152
rect 8636 57088 8652 57152
rect 8716 57088 8722 57152
rect 8406 57087 8722 57088
rect 933 56810 999 56813
rect 0 56808 999 56810
rect 0 56752 938 56808
rect 994 56752 999 56808
rect 0 56750 999 56752
rect 933 56747 999 56750
rect 2946 56608 3262 56609
rect 2946 56544 2952 56608
rect 3016 56544 3032 56608
rect 3096 56544 3112 56608
rect 3176 56544 3192 56608
rect 3256 56544 3262 56608
rect 2946 56543 3262 56544
rect 4546 56608 4862 56609
rect 4546 56544 4552 56608
rect 4616 56544 4632 56608
rect 4696 56544 4712 56608
rect 4776 56544 4792 56608
rect 4856 56544 4862 56608
rect 4546 56543 4862 56544
rect 6146 56608 6462 56609
rect 6146 56544 6152 56608
rect 6216 56544 6232 56608
rect 6296 56544 6312 56608
rect 6376 56544 6392 56608
rect 6456 56544 6462 56608
rect 6146 56543 6462 56544
rect 7746 56608 8062 56609
rect 7746 56544 7752 56608
rect 7816 56544 7832 56608
rect 7896 56544 7912 56608
rect 7976 56544 7992 56608
rect 8056 56544 8062 56608
rect 7746 56543 8062 56544
rect 9346 56608 9662 56609
rect 9346 56544 9352 56608
rect 9416 56544 9432 56608
rect 9496 56544 9512 56608
rect 9576 56544 9592 56608
rect 9656 56544 9662 56608
rect 9346 56543 9662 56544
rect 3606 56064 3922 56065
rect 3606 56000 3612 56064
rect 3676 56000 3692 56064
rect 3756 56000 3772 56064
rect 3836 56000 3852 56064
rect 3916 56000 3922 56064
rect 3606 55999 3922 56000
rect 5206 56064 5522 56065
rect 5206 56000 5212 56064
rect 5276 56000 5292 56064
rect 5356 56000 5372 56064
rect 5436 56000 5452 56064
rect 5516 56000 5522 56064
rect 5206 55999 5522 56000
rect 6806 56064 7122 56065
rect 6806 56000 6812 56064
rect 6876 56000 6892 56064
rect 6956 56000 6972 56064
rect 7036 56000 7052 56064
rect 7116 56000 7122 56064
rect 6806 55999 7122 56000
rect 8406 56064 8722 56065
rect 8406 56000 8412 56064
rect 8476 56000 8492 56064
rect 8556 56000 8572 56064
rect 8636 56000 8652 56064
rect 8716 56000 8722 56064
rect 8406 55999 8722 56000
rect 933 55858 999 55861
rect 0 55856 999 55858
rect 0 55800 938 55856
rect 994 55800 999 55856
rect 0 55798 999 55800
rect 933 55795 999 55798
rect 2946 55520 3262 55521
rect 2946 55456 2952 55520
rect 3016 55456 3032 55520
rect 3096 55456 3112 55520
rect 3176 55456 3192 55520
rect 3256 55456 3262 55520
rect 2946 55455 3262 55456
rect 4546 55520 4862 55521
rect 4546 55456 4552 55520
rect 4616 55456 4632 55520
rect 4696 55456 4712 55520
rect 4776 55456 4792 55520
rect 4856 55456 4862 55520
rect 4546 55455 4862 55456
rect 6146 55520 6462 55521
rect 6146 55456 6152 55520
rect 6216 55456 6232 55520
rect 6296 55456 6312 55520
rect 6376 55456 6392 55520
rect 6456 55456 6462 55520
rect 6146 55455 6462 55456
rect 7746 55520 8062 55521
rect 7746 55456 7752 55520
rect 7816 55456 7832 55520
rect 7896 55456 7912 55520
rect 7976 55456 7992 55520
rect 8056 55456 8062 55520
rect 7746 55455 8062 55456
rect 9346 55520 9662 55521
rect 9346 55456 9352 55520
rect 9416 55456 9432 55520
rect 9496 55456 9512 55520
rect 9576 55456 9592 55520
rect 9656 55456 9662 55520
rect 9346 55455 9662 55456
rect 3606 54976 3922 54977
rect 3606 54912 3612 54976
rect 3676 54912 3692 54976
rect 3756 54912 3772 54976
rect 3836 54912 3852 54976
rect 3916 54912 3922 54976
rect 3606 54911 3922 54912
rect 5206 54976 5522 54977
rect 5206 54912 5212 54976
rect 5276 54912 5292 54976
rect 5356 54912 5372 54976
rect 5436 54912 5452 54976
rect 5516 54912 5522 54976
rect 5206 54911 5522 54912
rect 6806 54976 7122 54977
rect 6806 54912 6812 54976
rect 6876 54912 6892 54976
rect 6956 54912 6972 54976
rect 7036 54912 7052 54976
rect 7116 54912 7122 54976
rect 6806 54911 7122 54912
rect 8406 54976 8722 54977
rect 8406 54912 8412 54976
rect 8476 54912 8492 54976
rect 8556 54912 8572 54976
rect 8636 54912 8652 54976
rect 8716 54912 8722 54976
rect 8406 54911 8722 54912
rect 933 54906 999 54909
rect 0 54904 999 54906
rect 0 54848 938 54904
rect 994 54848 999 54904
rect 0 54846 999 54848
rect 933 54843 999 54846
rect 2946 54432 3262 54433
rect 2946 54368 2952 54432
rect 3016 54368 3032 54432
rect 3096 54368 3112 54432
rect 3176 54368 3192 54432
rect 3256 54368 3262 54432
rect 2946 54367 3262 54368
rect 4546 54432 4862 54433
rect 4546 54368 4552 54432
rect 4616 54368 4632 54432
rect 4696 54368 4712 54432
rect 4776 54368 4792 54432
rect 4856 54368 4862 54432
rect 4546 54367 4862 54368
rect 6146 54432 6462 54433
rect 6146 54368 6152 54432
rect 6216 54368 6232 54432
rect 6296 54368 6312 54432
rect 6376 54368 6392 54432
rect 6456 54368 6462 54432
rect 6146 54367 6462 54368
rect 7746 54432 8062 54433
rect 7746 54368 7752 54432
rect 7816 54368 7832 54432
rect 7896 54368 7912 54432
rect 7976 54368 7992 54432
rect 8056 54368 8062 54432
rect 7746 54367 8062 54368
rect 9346 54432 9662 54433
rect 9346 54368 9352 54432
rect 9416 54368 9432 54432
rect 9496 54368 9512 54432
rect 9576 54368 9592 54432
rect 9656 54368 9662 54432
rect 9346 54367 9662 54368
rect 4153 54226 4219 54229
rect 7833 54226 7899 54229
rect 4153 54224 7899 54226
rect 4153 54168 4158 54224
rect 4214 54168 7838 54224
rect 7894 54168 7899 54224
rect 4153 54166 7899 54168
rect 4153 54163 4219 54166
rect 7833 54163 7899 54166
rect 933 53954 999 53957
rect 0 53952 999 53954
rect 0 53896 938 53952
rect 994 53896 999 53952
rect 0 53894 999 53896
rect 933 53891 999 53894
rect 3606 53888 3922 53889
rect 3606 53824 3612 53888
rect 3676 53824 3692 53888
rect 3756 53824 3772 53888
rect 3836 53824 3852 53888
rect 3916 53824 3922 53888
rect 3606 53823 3922 53824
rect 5206 53888 5522 53889
rect 5206 53824 5212 53888
rect 5276 53824 5292 53888
rect 5356 53824 5372 53888
rect 5436 53824 5452 53888
rect 5516 53824 5522 53888
rect 5206 53823 5522 53824
rect 6806 53888 7122 53889
rect 6806 53824 6812 53888
rect 6876 53824 6892 53888
rect 6956 53824 6972 53888
rect 7036 53824 7052 53888
rect 7116 53824 7122 53888
rect 6806 53823 7122 53824
rect 8406 53888 8722 53889
rect 8406 53824 8412 53888
rect 8476 53824 8492 53888
rect 8556 53824 8572 53888
rect 8636 53824 8652 53888
rect 8716 53824 8722 53888
rect 8406 53823 8722 53824
rect 5993 53546 6059 53549
rect 7097 53546 7163 53549
rect 5993 53544 7163 53546
rect 5993 53488 5998 53544
rect 6054 53488 7102 53544
rect 7158 53488 7163 53544
rect 5993 53486 7163 53488
rect 5993 53483 6059 53486
rect 7097 53483 7163 53486
rect 2946 53344 3262 53345
rect 2946 53280 2952 53344
rect 3016 53280 3032 53344
rect 3096 53280 3112 53344
rect 3176 53280 3192 53344
rect 3256 53280 3262 53344
rect 2946 53279 3262 53280
rect 4546 53344 4862 53345
rect 4546 53280 4552 53344
rect 4616 53280 4632 53344
rect 4696 53280 4712 53344
rect 4776 53280 4792 53344
rect 4856 53280 4862 53344
rect 4546 53279 4862 53280
rect 6146 53344 6462 53345
rect 6146 53280 6152 53344
rect 6216 53280 6232 53344
rect 6296 53280 6312 53344
rect 6376 53280 6392 53344
rect 6456 53280 6462 53344
rect 6146 53279 6462 53280
rect 7746 53344 8062 53345
rect 7746 53280 7752 53344
rect 7816 53280 7832 53344
rect 7896 53280 7912 53344
rect 7976 53280 7992 53344
rect 8056 53280 8062 53344
rect 7746 53279 8062 53280
rect 9346 53344 9662 53345
rect 9346 53280 9352 53344
rect 9416 53280 9432 53344
rect 9496 53280 9512 53344
rect 9576 53280 9592 53344
rect 9656 53280 9662 53344
rect 9346 53279 9662 53280
rect 933 53002 999 53005
rect 0 53000 999 53002
rect 0 52944 938 53000
rect 994 52944 999 53000
rect 0 52942 999 52944
rect 933 52939 999 52942
rect 7189 53002 7255 53005
rect 7465 53002 7531 53005
rect 7189 53000 7531 53002
rect 7189 52944 7194 53000
rect 7250 52944 7470 53000
rect 7526 52944 7531 53000
rect 7189 52942 7531 52944
rect 7189 52939 7255 52942
rect 7465 52939 7531 52942
rect 3606 52800 3922 52801
rect 3606 52736 3612 52800
rect 3676 52736 3692 52800
rect 3756 52736 3772 52800
rect 3836 52736 3852 52800
rect 3916 52736 3922 52800
rect 3606 52735 3922 52736
rect 5206 52800 5522 52801
rect 5206 52736 5212 52800
rect 5276 52736 5292 52800
rect 5356 52736 5372 52800
rect 5436 52736 5452 52800
rect 5516 52736 5522 52800
rect 5206 52735 5522 52736
rect 6806 52800 7122 52801
rect 6806 52736 6812 52800
rect 6876 52736 6892 52800
rect 6956 52736 6972 52800
rect 7036 52736 7052 52800
rect 7116 52736 7122 52800
rect 6806 52735 7122 52736
rect 8406 52800 8722 52801
rect 8406 52736 8412 52800
rect 8476 52736 8492 52800
rect 8556 52736 8572 52800
rect 8636 52736 8652 52800
rect 8716 52736 8722 52800
rect 8406 52735 8722 52736
rect 1577 52322 1643 52325
rect 798 52320 1643 52322
rect 798 52264 1582 52320
rect 1638 52264 1643 52320
rect 798 52262 1643 52264
rect 798 52050 858 52262
rect 1577 52259 1643 52262
rect 2946 52256 3262 52257
rect 2946 52192 2952 52256
rect 3016 52192 3032 52256
rect 3096 52192 3112 52256
rect 3176 52192 3192 52256
rect 3256 52192 3262 52256
rect 2946 52191 3262 52192
rect 4546 52256 4862 52257
rect 4546 52192 4552 52256
rect 4616 52192 4632 52256
rect 4696 52192 4712 52256
rect 4776 52192 4792 52256
rect 4856 52192 4862 52256
rect 4546 52191 4862 52192
rect 6146 52256 6462 52257
rect 6146 52192 6152 52256
rect 6216 52192 6232 52256
rect 6296 52192 6312 52256
rect 6376 52192 6392 52256
rect 6456 52192 6462 52256
rect 6146 52191 6462 52192
rect 7746 52256 8062 52257
rect 7746 52192 7752 52256
rect 7816 52192 7832 52256
rect 7896 52192 7912 52256
rect 7976 52192 7992 52256
rect 8056 52192 8062 52256
rect 7746 52191 8062 52192
rect 9346 52256 9662 52257
rect 9346 52192 9352 52256
rect 9416 52192 9432 52256
rect 9496 52192 9512 52256
rect 9576 52192 9592 52256
rect 9656 52192 9662 52256
rect 9346 52191 9662 52192
rect 7373 52186 7439 52189
rect 7373 52184 7482 52186
rect 7373 52128 7378 52184
rect 7434 52128 7482 52184
rect 7373 52123 7482 52128
rect 0 51990 858 52050
rect 7422 51914 7482 52123
rect 7557 51914 7623 51917
rect 7422 51912 7623 51914
rect 7422 51856 7562 51912
rect 7618 51856 7623 51912
rect 7422 51854 7623 51856
rect 7557 51851 7623 51854
rect 3606 51712 3922 51713
rect 3606 51648 3612 51712
rect 3676 51648 3692 51712
rect 3756 51648 3772 51712
rect 3836 51648 3852 51712
rect 3916 51648 3922 51712
rect 3606 51647 3922 51648
rect 5206 51712 5522 51713
rect 5206 51648 5212 51712
rect 5276 51648 5292 51712
rect 5356 51648 5372 51712
rect 5436 51648 5452 51712
rect 5516 51648 5522 51712
rect 5206 51647 5522 51648
rect 6806 51712 7122 51713
rect 6806 51648 6812 51712
rect 6876 51648 6892 51712
rect 6956 51648 6972 51712
rect 7036 51648 7052 51712
rect 7116 51648 7122 51712
rect 6806 51647 7122 51648
rect 8406 51712 8722 51713
rect 8406 51648 8412 51712
rect 8476 51648 8492 51712
rect 8556 51648 8572 51712
rect 8636 51648 8652 51712
rect 8716 51648 8722 51712
rect 8406 51647 8722 51648
rect 6085 51370 6151 51373
rect 5950 51368 6151 51370
rect 5950 51312 6090 51368
rect 6146 51312 6151 51368
rect 5950 51310 6151 51312
rect 2946 51168 3262 51169
rect 2946 51104 2952 51168
rect 3016 51104 3032 51168
rect 3096 51104 3112 51168
rect 3176 51104 3192 51168
rect 3256 51104 3262 51168
rect 2946 51103 3262 51104
rect 4546 51168 4862 51169
rect 4546 51104 4552 51168
rect 4616 51104 4632 51168
rect 4696 51104 4712 51168
rect 4776 51104 4792 51168
rect 4856 51104 4862 51168
rect 4546 51103 4862 51104
rect 933 51098 999 51101
rect 0 51096 999 51098
rect 0 51040 938 51096
rect 994 51040 999 51096
rect 0 51038 999 51040
rect 933 51035 999 51038
rect 5950 50962 6010 51310
rect 6085 51307 6151 51310
rect 6146 51168 6462 51169
rect 6146 51104 6152 51168
rect 6216 51104 6232 51168
rect 6296 51104 6312 51168
rect 6376 51104 6392 51168
rect 6456 51104 6462 51168
rect 6146 51103 6462 51104
rect 7746 51168 8062 51169
rect 7746 51104 7752 51168
rect 7816 51104 7832 51168
rect 7896 51104 7912 51168
rect 7976 51104 7992 51168
rect 8056 51104 8062 51168
rect 7746 51103 8062 51104
rect 9346 51168 9662 51169
rect 9346 51104 9352 51168
rect 9416 51104 9432 51168
rect 9496 51104 9512 51168
rect 9576 51104 9592 51168
rect 9656 51104 9662 51168
rect 9346 51103 9662 51104
rect 6085 50962 6151 50965
rect 5950 50960 6151 50962
rect 5950 50904 6090 50960
rect 6146 50904 6151 50960
rect 5950 50902 6151 50904
rect 6085 50899 6151 50902
rect 3606 50624 3922 50625
rect 3606 50560 3612 50624
rect 3676 50560 3692 50624
rect 3756 50560 3772 50624
rect 3836 50560 3852 50624
rect 3916 50560 3922 50624
rect 3606 50559 3922 50560
rect 5206 50624 5522 50625
rect 5206 50560 5212 50624
rect 5276 50560 5292 50624
rect 5356 50560 5372 50624
rect 5436 50560 5452 50624
rect 5516 50560 5522 50624
rect 5206 50559 5522 50560
rect 6806 50624 7122 50625
rect 6806 50560 6812 50624
rect 6876 50560 6892 50624
rect 6956 50560 6972 50624
rect 7036 50560 7052 50624
rect 7116 50560 7122 50624
rect 6806 50559 7122 50560
rect 8406 50624 8722 50625
rect 8406 50560 8412 50624
rect 8476 50560 8492 50624
rect 8556 50560 8572 50624
rect 8636 50560 8652 50624
rect 8716 50560 8722 50624
rect 8406 50559 8722 50560
rect 9489 50282 9555 50285
rect 9078 50280 9555 50282
rect 9078 50224 9494 50280
rect 9550 50224 9555 50280
rect 9078 50222 9555 50224
rect 933 50146 999 50149
rect 0 50144 999 50146
rect 0 50088 938 50144
rect 994 50088 999 50144
rect 0 50086 999 50088
rect 933 50083 999 50086
rect 2946 50080 3262 50081
rect 2946 50016 2952 50080
rect 3016 50016 3032 50080
rect 3096 50016 3112 50080
rect 3176 50016 3192 50080
rect 3256 50016 3262 50080
rect 2946 50015 3262 50016
rect 4546 50080 4862 50081
rect 4546 50016 4552 50080
rect 4616 50016 4632 50080
rect 4696 50016 4712 50080
rect 4776 50016 4792 50080
rect 4856 50016 4862 50080
rect 4546 50015 4862 50016
rect 6146 50080 6462 50081
rect 6146 50016 6152 50080
rect 6216 50016 6232 50080
rect 6296 50016 6312 50080
rect 6376 50016 6392 50080
rect 6456 50016 6462 50080
rect 6146 50015 6462 50016
rect 7746 50080 8062 50081
rect 7746 50016 7752 50080
rect 7816 50016 7832 50080
rect 7896 50016 7912 50080
rect 7976 50016 7992 50080
rect 8056 50016 8062 50080
rect 7746 50015 8062 50016
rect 3606 49536 3922 49537
rect 3606 49472 3612 49536
rect 3676 49472 3692 49536
rect 3756 49472 3772 49536
rect 3836 49472 3852 49536
rect 3916 49472 3922 49536
rect 3606 49471 3922 49472
rect 5206 49536 5522 49537
rect 5206 49472 5212 49536
rect 5276 49472 5292 49536
rect 5356 49472 5372 49536
rect 5436 49472 5452 49536
rect 5516 49472 5522 49536
rect 5206 49471 5522 49472
rect 6806 49536 7122 49537
rect 6806 49472 6812 49536
rect 6876 49472 6892 49536
rect 6956 49472 6972 49536
rect 7036 49472 7052 49536
rect 7116 49472 7122 49536
rect 6806 49471 7122 49472
rect 8406 49536 8722 49537
rect 8406 49472 8412 49536
rect 8476 49472 8492 49536
rect 8556 49472 8572 49536
rect 8636 49472 8652 49536
rect 8716 49472 8722 49536
rect 8406 49471 8722 49472
rect 933 49194 999 49197
rect 0 49192 999 49194
rect 0 49136 938 49192
rect 994 49136 999 49192
rect 0 49134 999 49136
rect 933 49131 999 49134
rect 2946 48992 3262 48993
rect 2946 48928 2952 48992
rect 3016 48928 3032 48992
rect 3096 48928 3112 48992
rect 3176 48928 3192 48992
rect 3256 48928 3262 48992
rect 2946 48927 3262 48928
rect 4546 48992 4862 48993
rect 4546 48928 4552 48992
rect 4616 48928 4632 48992
rect 4696 48928 4712 48992
rect 4776 48928 4792 48992
rect 4856 48928 4862 48992
rect 4546 48927 4862 48928
rect 6146 48992 6462 48993
rect 6146 48928 6152 48992
rect 6216 48928 6232 48992
rect 6296 48928 6312 48992
rect 6376 48928 6392 48992
rect 6456 48928 6462 48992
rect 6146 48927 6462 48928
rect 7746 48992 8062 48993
rect 7746 48928 7752 48992
rect 7816 48928 7832 48992
rect 7896 48928 7912 48992
rect 7976 48928 7992 48992
rect 8056 48928 8062 48992
rect 7746 48927 8062 48928
rect 9078 48786 9138 50222
rect 9489 50219 9555 50222
rect 9346 50080 9662 50081
rect 9346 50016 9352 50080
rect 9416 50016 9432 50080
rect 9496 50016 9512 50080
rect 9576 50016 9592 50080
rect 9656 50016 9662 50080
rect 9346 50015 9662 50016
rect 9346 48992 9662 48993
rect 9346 48928 9352 48992
rect 9416 48928 9432 48992
rect 9496 48928 9512 48992
rect 9576 48928 9592 48992
rect 9656 48928 9662 48992
rect 9346 48927 9662 48928
rect 9305 48786 9371 48789
rect 9078 48784 9371 48786
rect 9078 48728 9310 48784
rect 9366 48728 9371 48784
rect 9078 48726 9371 48728
rect 9305 48723 9371 48726
rect 3606 48448 3922 48449
rect 3606 48384 3612 48448
rect 3676 48384 3692 48448
rect 3756 48384 3772 48448
rect 3836 48384 3852 48448
rect 3916 48384 3922 48448
rect 3606 48383 3922 48384
rect 5206 48448 5522 48449
rect 5206 48384 5212 48448
rect 5276 48384 5292 48448
rect 5356 48384 5372 48448
rect 5436 48384 5452 48448
rect 5516 48384 5522 48448
rect 5206 48383 5522 48384
rect 6806 48448 7122 48449
rect 6806 48384 6812 48448
rect 6876 48384 6892 48448
rect 6956 48384 6972 48448
rect 7036 48384 7052 48448
rect 7116 48384 7122 48448
rect 6806 48383 7122 48384
rect 8406 48448 8722 48449
rect 8406 48384 8412 48448
rect 8476 48384 8492 48448
rect 8556 48384 8572 48448
rect 8636 48384 8652 48448
rect 8716 48384 8722 48448
rect 8406 48383 8722 48384
rect 1577 48242 1643 48245
rect 0 48240 1643 48242
rect 0 48184 1582 48240
rect 1638 48184 1643 48240
rect 0 48182 1643 48184
rect 1577 48179 1643 48182
rect 9305 48106 9371 48109
rect 9078 48104 9371 48106
rect 9078 48048 9310 48104
rect 9366 48048 9371 48104
rect 9078 48046 9371 48048
rect 2946 47904 3262 47905
rect 2946 47840 2952 47904
rect 3016 47840 3032 47904
rect 3096 47840 3112 47904
rect 3176 47840 3192 47904
rect 3256 47840 3262 47904
rect 2946 47839 3262 47840
rect 4546 47904 4862 47905
rect 4546 47840 4552 47904
rect 4616 47840 4632 47904
rect 4696 47840 4712 47904
rect 4776 47840 4792 47904
rect 4856 47840 4862 47904
rect 4546 47839 4862 47840
rect 6146 47904 6462 47905
rect 6146 47840 6152 47904
rect 6216 47840 6232 47904
rect 6296 47840 6312 47904
rect 6376 47840 6392 47904
rect 6456 47840 6462 47904
rect 6146 47839 6462 47840
rect 7746 47904 8062 47905
rect 7746 47840 7752 47904
rect 7816 47840 7832 47904
rect 7896 47840 7912 47904
rect 7976 47840 7992 47904
rect 8056 47840 8062 47904
rect 7746 47839 8062 47840
rect 3606 47360 3922 47361
rect 3606 47296 3612 47360
rect 3676 47296 3692 47360
rect 3756 47296 3772 47360
rect 3836 47296 3852 47360
rect 3916 47296 3922 47360
rect 3606 47295 3922 47296
rect 5206 47360 5522 47361
rect 5206 47296 5212 47360
rect 5276 47296 5292 47360
rect 5356 47296 5372 47360
rect 5436 47296 5452 47360
rect 5516 47296 5522 47360
rect 5206 47295 5522 47296
rect 6806 47360 7122 47361
rect 6806 47296 6812 47360
rect 6876 47296 6892 47360
rect 6956 47296 6972 47360
rect 7036 47296 7052 47360
rect 7116 47296 7122 47360
rect 6806 47295 7122 47296
rect 8406 47360 8722 47361
rect 8406 47296 8412 47360
rect 8476 47296 8492 47360
rect 8556 47296 8572 47360
rect 8636 47296 8652 47360
rect 8716 47296 8722 47360
rect 8406 47295 8722 47296
rect 933 47290 999 47293
rect 0 47288 999 47290
rect 0 47232 938 47288
rect 994 47232 999 47288
rect 0 47230 999 47232
rect 933 47227 999 47230
rect 4429 47018 4495 47021
rect 4294 47016 4495 47018
rect 4294 46960 4434 47016
rect 4490 46960 4495 47016
rect 4294 46958 4495 46960
rect 2946 46816 3262 46817
rect 2946 46752 2952 46816
rect 3016 46752 3032 46816
rect 3096 46752 3112 46816
rect 3176 46752 3192 46816
rect 3256 46752 3262 46816
rect 2946 46751 3262 46752
rect 4294 46610 4354 46958
rect 4429 46955 4495 46958
rect 4546 46816 4862 46817
rect 4546 46752 4552 46816
rect 4616 46752 4632 46816
rect 4696 46752 4712 46816
rect 4776 46752 4792 46816
rect 4856 46752 4862 46816
rect 4546 46751 4862 46752
rect 6146 46816 6462 46817
rect 6146 46752 6152 46816
rect 6216 46752 6232 46816
rect 6296 46752 6312 46816
rect 6376 46752 6392 46816
rect 6456 46752 6462 46816
rect 6146 46751 6462 46752
rect 7746 46816 8062 46817
rect 7746 46752 7752 46816
rect 7816 46752 7832 46816
rect 7896 46752 7912 46816
rect 7976 46752 7992 46816
rect 8056 46752 8062 46816
rect 7746 46751 8062 46752
rect 4429 46610 4495 46613
rect 4294 46608 4495 46610
rect 4294 46552 4434 46608
rect 4490 46552 4495 46608
rect 4294 46550 4495 46552
rect 9078 46610 9138 48046
rect 9305 48043 9371 48046
rect 9346 47904 9662 47905
rect 9346 47840 9352 47904
rect 9416 47840 9432 47904
rect 9496 47840 9512 47904
rect 9576 47840 9592 47904
rect 9656 47840 9662 47904
rect 9346 47839 9662 47840
rect 9346 46816 9662 46817
rect 9346 46752 9352 46816
rect 9416 46752 9432 46816
rect 9496 46752 9512 46816
rect 9576 46752 9592 46816
rect 9656 46752 9662 46816
rect 9346 46751 9662 46752
rect 9305 46610 9371 46613
rect 9078 46608 9371 46610
rect 9078 46552 9310 46608
rect 9366 46552 9371 46608
rect 9078 46550 9371 46552
rect 4429 46547 4495 46550
rect 9305 46547 9371 46550
rect 7097 46474 7163 46477
rect 7097 46472 8264 46474
rect 7097 46416 7102 46472
rect 7158 46416 8264 46472
rect 7097 46414 8264 46416
rect 7097 46411 7163 46414
rect 933 46338 999 46341
rect 0 46336 999 46338
rect 0 46280 938 46336
rect 994 46280 999 46336
rect 0 46278 999 46280
rect 933 46275 999 46278
rect 3606 46272 3922 46273
rect 3606 46208 3612 46272
rect 3676 46208 3692 46272
rect 3756 46208 3772 46272
rect 3836 46208 3852 46272
rect 3916 46208 3922 46272
rect 3606 46207 3922 46208
rect 5206 46272 5522 46273
rect 5206 46208 5212 46272
rect 5276 46208 5292 46272
rect 5356 46208 5372 46272
rect 5436 46208 5452 46272
rect 5516 46208 5522 46272
rect 5206 46207 5522 46208
rect 6806 46272 7122 46273
rect 6806 46208 6812 46272
rect 6876 46208 6892 46272
rect 6956 46208 6972 46272
rect 7036 46208 7052 46272
rect 7116 46208 7122 46272
rect 6806 46207 7122 46208
rect 5993 45930 6059 45933
rect 5950 45928 6059 45930
rect 5950 45872 5998 45928
rect 6054 45872 6059 45928
rect 5950 45867 6059 45872
rect 2946 45728 3262 45729
rect 2946 45664 2952 45728
rect 3016 45664 3032 45728
rect 3096 45664 3112 45728
rect 3176 45664 3192 45728
rect 3256 45664 3262 45728
rect 2946 45663 3262 45664
rect 4546 45728 4862 45729
rect 4546 45664 4552 45728
rect 4616 45664 4632 45728
rect 4696 45664 4712 45728
rect 4776 45664 4792 45728
rect 4856 45664 4862 45728
rect 4546 45663 4862 45664
rect 4061 45522 4127 45525
rect 5950 45522 6010 45867
rect 6146 45728 6462 45729
rect 6146 45664 6152 45728
rect 6216 45664 6232 45728
rect 6296 45664 6312 45728
rect 6376 45664 6392 45728
rect 6456 45664 6462 45728
rect 6146 45663 6462 45664
rect 7746 45728 8062 45729
rect 7746 45664 7752 45728
rect 7816 45664 7832 45728
rect 7896 45664 7912 45728
rect 7976 45664 7992 45728
rect 8056 45664 8062 45728
rect 7746 45663 8062 45664
rect 8204 45661 8264 46414
rect 8406 46272 8722 46273
rect 8406 46208 8412 46272
rect 8476 46208 8492 46272
rect 8556 46208 8572 46272
rect 8636 46208 8652 46272
rect 8716 46208 8722 46272
rect 8406 46207 8722 46208
rect 9346 45728 9662 45729
rect 9346 45664 9352 45728
rect 9416 45664 9432 45728
rect 9496 45664 9512 45728
rect 9576 45664 9592 45728
rect 9656 45664 9662 45728
rect 9346 45663 9662 45664
rect 8201 45656 8267 45661
rect 8201 45600 8206 45656
rect 8262 45600 8267 45656
rect 8201 45595 8267 45600
rect 6085 45522 6151 45525
rect 4061 45520 5688 45522
rect 4061 45464 4066 45520
rect 4122 45464 5688 45520
rect 4061 45462 5688 45464
rect 5950 45520 6151 45522
rect 5950 45464 6090 45520
rect 6146 45464 6151 45520
rect 5950 45462 6151 45464
rect 4061 45459 4127 45462
rect 933 45386 999 45389
rect 5165 45386 5231 45389
rect 0 45384 999 45386
rect 0 45328 938 45384
rect 994 45328 999 45384
rect 0 45326 999 45328
rect 933 45323 999 45326
rect 5030 45384 5231 45386
rect 5030 45328 5170 45384
rect 5226 45328 5231 45384
rect 5030 45326 5231 45328
rect 3606 45184 3922 45185
rect 3606 45120 3612 45184
rect 3676 45120 3692 45184
rect 3756 45120 3772 45184
rect 3836 45120 3852 45184
rect 3916 45120 3922 45184
rect 3606 45119 3922 45120
rect 3969 44978 4035 44981
rect 5030 44978 5090 45326
rect 5165 45323 5231 45326
rect 5206 45184 5522 45185
rect 5206 45120 5212 45184
rect 5276 45120 5292 45184
rect 5356 45120 5372 45184
rect 5436 45120 5452 45184
rect 5516 45120 5522 45184
rect 5206 45119 5522 45120
rect 5165 44978 5231 44981
rect 3969 44976 4722 44978
rect 3969 44920 3974 44976
rect 4030 44920 4722 44976
rect 3969 44918 4722 44920
rect 5030 44976 5231 44978
rect 5030 44920 5170 44976
rect 5226 44920 5231 44976
rect 5030 44918 5231 44920
rect 3969 44915 4035 44918
rect 4662 44842 4722 44918
rect 5165 44915 5231 44918
rect 5628 44845 5688 45462
rect 6085 45459 6151 45462
rect 6806 45184 7122 45185
rect 6806 45120 6812 45184
rect 6876 45120 6892 45184
rect 6956 45120 6972 45184
rect 7036 45120 7052 45184
rect 7116 45120 7122 45184
rect 6806 45119 7122 45120
rect 8406 45184 8722 45185
rect 8406 45120 8412 45184
rect 8476 45120 8492 45184
rect 8556 45120 8572 45184
rect 8636 45120 8652 45184
rect 8716 45120 8722 45184
rect 8406 45119 8722 45120
rect 5441 44842 5507 44845
rect 4662 44840 5507 44842
rect 4662 44784 5446 44840
rect 5502 44784 5507 44840
rect 4662 44782 5507 44784
rect 5441 44779 5507 44782
rect 5625 44840 5691 44845
rect 5625 44784 5630 44840
rect 5686 44784 5691 44840
rect 5625 44779 5691 44784
rect 2946 44640 3262 44641
rect 2946 44576 2952 44640
rect 3016 44576 3032 44640
rect 3096 44576 3112 44640
rect 3176 44576 3192 44640
rect 3256 44576 3262 44640
rect 2946 44575 3262 44576
rect 4546 44640 4862 44641
rect 4546 44576 4552 44640
rect 4616 44576 4632 44640
rect 4696 44576 4712 44640
rect 4776 44576 4792 44640
rect 4856 44576 4862 44640
rect 4546 44575 4862 44576
rect 6146 44640 6462 44641
rect 6146 44576 6152 44640
rect 6216 44576 6232 44640
rect 6296 44576 6312 44640
rect 6376 44576 6392 44640
rect 6456 44576 6462 44640
rect 6146 44575 6462 44576
rect 7746 44640 8062 44641
rect 7746 44576 7752 44640
rect 7816 44576 7832 44640
rect 7896 44576 7912 44640
rect 7976 44576 7992 44640
rect 8056 44576 8062 44640
rect 7746 44575 8062 44576
rect 9346 44640 9662 44641
rect 9346 44576 9352 44640
rect 9416 44576 9432 44640
rect 9496 44576 9512 44640
rect 9576 44576 9592 44640
rect 9656 44576 9662 44640
rect 9346 44575 9662 44576
rect 933 44434 999 44437
rect 0 44432 999 44434
rect 0 44376 938 44432
rect 994 44376 999 44432
rect 0 44374 999 44376
rect 933 44371 999 44374
rect 3606 44096 3922 44097
rect 3606 44032 3612 44096
rect 3676 44032 3692 44096
rect 3756 44032 3772 44096
rect 3836 44032 3852 44096
rect 3916 44032 3922 44096
rect 3606 44031 3922 44032
rect 5206 44096 5522 44097
rect 5206 44032 5212 44096
rect 5276 44032 5292 44096
rect 5356 44032 5372 44096
rect 5436 44032 5452 44096
rect 5516 44032 5522 44096
rect 5206 44031 5522 44032
rect 6806 44096 7122 44097
rect 6806 44032 6812 44096
rect 6876 44032 6892 44096
rect 6956 44032 6972 44096
rect 7036 44032 7052 44096
rect 7116 44032 7122 44096
rect 6806 44031 7122 44032
rect 8406 44096 8722 44097
rect 8406 44032 8412 44096
rect 8476 44032 8492 44096
rect 8556 44032 8572 44096
rect 8636 44032 8652 44096
rect 8716 44032 8722 44096
rect 8406 44031 8722 44032
rect 6729 43890 6795 43893
rect 7189 43890 7255 43893
rect 6729 43888 7255 43890
rect 6729 43832 6734 43888
rect 6790 43832 7194 43888
rect 7250 43832 7255 43888
rect 6729 43830 7255 43832
rect 6729 43827 6795 43830
rect 7189 43827 7255 43830
rect 2946 43552 3262 43553
rect 2946 43488 2952 43552
rect 3016 43488 3032 43552
rect 3096 43488 3112 43552
rect 3176 43488 3192 43552
rect 3256 43488 3262 43552
rect 2946 43487 3262 43488
rect 4546 43552 4862 43553
rect 4546 43488 4552 43552
rect 4616 43488 4632 43552
rect 4696 43488 4712 43552
rect 4776 43488 4792 43552
rect 4856 43488 4862 43552
rect 4546 43487 4862 43488
rect 6146 43552 6462 43553
rect 6146 43488 6152 43552
rect 6216 43488 6232 43552
rect 6296 43488 6312 43552
rect 6376 43488 6392 43552
rect 6456 43488 6462 43552
rect 6146 43487 6462 43488
rect 7746 43552 8062 43553
rect 7746 43488 7752 43552
rect 7816 43488 7832 43552
rect 7896 43488 7912 43552
rect 7976 43488 7992 43552
rect 8056 43488 8062 43552
rect 7746 43487 8062 43488
rect 9346 43552 9662 43553
rect 9346 43488 9352 43552
rect 9416 43488 9432 43552
rect 9496 43488 9512 43552
rect 9576 43488 9592 43552
rect 9656 43488 9662 43552
rect 9346 43487 9662 43488
rect 933 43482 999 43485
rect 0 43480 999 43482
rect 0 43424 938 43480
rect 994 43424 999 43480
rect 0 43422 999 43424
rect 933 43419 999 43422
rect 3606 43008 3922 43009
rect 3606 42944 3612 43008
rect 3676 42944 3692 43008
rect 3756 42944 3772 43008
rect 3836 42944 3852 43008
rect 3916 42944 3922 43008
rect 3606 42943 3922 42944
rect 5206 43008 5522 43009
rect 5206 42944 5212 43008
rect 5276 42944 5292 43008
rect 5356 42944 5372 43008
rect 5436 42944 5452 43008
rect 5516 42944 5522 43008
rect 5206 42943 5522 42944
rect 6806 43008 7122 43009
rect 6806 42944 6812 43008
rect 6876 42944 6892 43008
rect 6956 42944 6972 43008
rect 7036 42944 7052 43008
rect 7116 42944 7122 43008
rect 6806 42943 7122 42944
rect 8406 43008 8722 43009
rect 8406 42944 8412 43008
rect 8476 42944 8492 43008
rect 8556 42944 8572 43008
rect 8636 42944 8652 43008
rect 8716 42944 8722 43008
rect 8406 42943 8722 42944
rect 5257 42666 5323 42669
rect 8937 42666 9003 42669
rect 5257 42664 9003 42666
rect 5257 42608 5262 42664
rect 5318 42608 8942 42664
rect 8998 42608 9003 42664
rect 5257 42606 9003 42608
rect 5257 42603 5323 42606
rect 8937 42603 9003 42606
rect 933 42530 999 42533
rect 0 42528 999 42530
rect 0 42472 938 42528
rect 994 42472 999 42528
rect 0 42470 999 42472
rect 933 42467 999 42470
rect 2946 42464 3262 42465
rect 2946 42400 2952 42464
rect 3016 42400 3032 42464
rect 3096 42400 3112 42464
rect 3176 42400 3192 42464
rect 3256 42400 3262 42464
rect 2946 42399 3262 42400
rect 4546 42464 4862 42465
rect 4546 42400 4552 42464
rect 4616 42400 4632 42464
rect 4696 42400 4712 42464
rect 4776 42400 4792 42464
rect 4856 42400 4862 42464
rect 4546 42399 4862 42400
rect 6146 42464 6462 42465
rect 6146 42400 6152 42464
rect 6216 42400 6232 42464
rect 6296 42400 6312 42464
rect 6376 42400 6392 42464
rect 6456 42400 6462 42464
rect 6146 42399 6462 42400
rect 7746 42464 8062 42465
rect 7746 42400 7752 42464
rect 7816 42400 7832 42464
rect 7896 42400 7912 42464
rect 7976 42400 7992 42464
rect 8056 42400 8062 42464
rect 7746 42399 8062 42400
rect 9346 42464 9662 42465
rect 9346 42400 9352 42464
rect 9416 42400 9432 42464
rect 9496 42400 9512 42464
rect 9576 42400 9592 42464
rect 9656 42400 9662 42464
rect 9346 42399 9662 42400
rect 4061 42258 4127 42261
rect 4613 42258 4679 42261
rect 4061 42256 4679 42258
rect 4061 42200 4066 42256
rect 4122 42200 4618 42256
rect 4674 42200 4679 42256
rect 4061 42198 4679 42200
rect 4061 42195 4127 42198
rect 4613 42195 4679 42198
rect 3606 41920 3922 41921
rect 3606 41856 3612 41920
rect 3676 41856 3692 41920
rect 3756 41856 3772 41920
rect 3836 41856 3852 41920
rect 3916 41856 3922 41920
rect 3606 41855 3922 41856
rect 5206 41920 5522 41921
rect 5206 41856 5212 41920
rect 5276 41856 5292 41920
rect 5356 41856 5372 41920
rect 5436 41856 5452 41920
rect 5516 41856 5522 41920
rect 5206 41855 5522 41856
rect 6806 41920 7122 41921
rect 6806 41856 6812 41920
rect 6876 41856 6892 41920
rect 6956 41856 6972 41920
rect 7036 41856 7052 41920
rect 7116 41856 7122 41920
rect 6806 41855 7122 41856
rect 8406 41920 8722 41921
rect 8406 41856 8412 41920
rect 8476 41856 8492 41920
rect 8556 41856 8572 41920
rect 8636 41856 8652 41920
rect 8716 41856 8722 41920
rect 8406 41855 8722 41856
rect 933 41578 999 41581
rect 0 41576 999 41578
rect 0 41520 938 41576
rect 994 41520 999 41576
rect 0 41518 999 41520
rect 933 41515 999 41518
rect 2946 41376 3262 41377
rect 2946 41312 2952 41376
rect 3016 41312 3032 41376
rect 3096 41312 3112 41376
rect 3176 41312 3192 41376
rect 3256 41312 3262 41376
rect 2946 41311 3262 41312
rect 4546 41376 4862 41377
rect 4546 41312 4552 41376
rect 4616 41312 4632 41376
rect 4696 41312 4712 41376
rect 4776 41312 4792 41376
rect 4856 41312 4862 41376
rect 4546 41311 4862 41312
rect 6146 41376 6462 41377
rect 6146 41312 6152 41376
rect 6216 41312 6232 41376
rect 6296 41312 6312 41376
rect 6376 41312 6392 41376
rect 6456 41312 6462 41376
rect 6146 41311 6462 41312
rect 7746 41376 8062 41377
rect 7746 41312 7752 41376
rect 7816 41312 7832 41376
rect 7896 41312 7912 41376
rect 7976 41312 7992 41376
rect 8056 41312 8062 41376
rect 7746 41311 8062 41312
rect 9346 41376 9662 41377
rect 9346 41312 9352 41376
rect 9416 41312 9432 41376
rect 9496 41312 9512 41376
rect 9576 41312 9592 41376
rect 9656 41312 9662 41376
rect 9346 41311 9662 41312
rect 3606 40832 3922 40833
rect 3606 40768 3612 40832
rect 3676 40768 3692 40832
rect 3756 40768 3772 40832
rect 3836 40768 3852 40832
rect 3916 40768 3922 40832
rect 3606 40767 3922 40768
rect 5206 40832 5522 40833
rect 5206 40768 5212 40832
rect 5276 40768 5292 40832
rect 5356 40768 5372 40832
rect 5436 40768 5452 40832
rect 5516 40768 5522 40832
rect 5206 40767 5522 40768
rect 6806 40832 7122 40833
rect 6806 40768 6812 40832
rect 6876 40768 6892 40832
rect 6956 40768 6972 40832
rect 7036 40768 7052 40832
rect 7116 40768 7122 40832
rect 6806 40767 7122 40768
rect 8406 40832 8722 40833
rect 8406 40768 8412 40832
rect 8476 40768 8492 40832
rect 8556 40768 8572 40832
rect 8636 40768 8652 40832
rect 8716 40768 8722 40832
rect 8406 40767 8722 40768
rect 1025 40626 1091 40629
rect 0 40624 1091 40626
rect 0 40568 1030 40624
rect 1086 40568 1091 40624
rect 0 40566 1091 40568
rect 1025 40563 1091 40566
rect 2946 40288 3262 40289
rect 2946 40224 2952 40288
rect 3016 40224 3032 40288
rect 3096 40224 3112 40288
rect 3176 40224 3192 40288
rect 3256 40224 3262 40288
rect 2946 40223 3262 40224
rect 4546 40288 4862 40289
rect 4546 40224 4552 40288
rect 4616 40224 4632 40288
rect 4696 40224 4712 40288
rect 4776 40224 4792 40288
rect 4856 40224 4862 40288
rect 4546 40223 4862 40224
rect 6146 40288 6462 40289
rect 6146 40224 6152 40288
rect 6216 40224 6232 40288
rect 6296 40224 6312 40288
rect 6376 40224 6392 40288
rect 6456 40224 6462 40288
rect 6146 40223 6462 40224
rect 7746 40288 8062 40289
rect 7746 40224 7752 40288
rect 7816 40224 7832 40288
rect 7896 40224 7912 40288
rect 7976 40224 7992 40288
rect 8056 40224 8062 40288
rect 7746 40223 8062 40224
rect 9346 40288 9662 40289
rect 9346 40224 9352 40288
rect 9416 40224 9432 40288
rect 9496 40224 9512 40288
rect 9576 40224 9592 40288
rect 9656 40224 9662 40288
rect 9346 40223 9662 40224
rect 1485 39946 1551 39949
rect 798 39944 1551 39946
rect 798 39888 1490 39944
rect 1546 39888 1551 39944
rect 798 39886 1551 39888
rect 798 39674 858 39886
rect 1485 39883 1551 39886
rect 7833 39946 7899 39949
rect 11094 39946 11100 39948
rect 7833 39944 11100 39946
rect 7833 39888 7838 39944
rect 7894 39888 11100 39944
rect 7833 39886 11100 39888
rect 7833 39883 7899 39886
rect 11094 39884 11100 39886
rect 11164 39884 11170 39948
rect 3606 39744 3922 39745
rect 3606 39680 3612 39744
rect 3676 39680 3692 39744
rect 3756 39680 3772 39744
rect 3836 39680 3852 39744
rect 3916 39680 3922 39744
rect 3606 39679 3922 39680
rect 5206 39744 5522 39745
rect 5206 39680 5212 39744
rect 5276 39680 5292 39744
rect 5356 39680 5372 39744
rect 5436 39680 5452 39744
rect 5516 39680 5522 39744
rect 5206 39679 5522 39680
rect 6806 39744 7122 39745
rect 6806 39680 6812 39744
rect 6876 39680 6892 39744
rect 6956 39680 6972 39744
rect 7036 39680 7052 39744
rect 7116 39680 7122 39744
rect 6806 39679 7122 39680
rect 8406 39744 8722 39745
rect 8406 39680 8412 39744
rect 8476 39680 8492 39744
rect 8556 39680 8572 39744
rect 8636 39680 8652 39744
rect 8716 39680 8722 39744
rect 8406 39679 8722 39680
rect 0 39614 858 39674
rect 2946 39200 3262 39201
rect 2946 39136 2952 39200
rect 3016 39136 3032 39200
rect 3096 39136 3112 39200
rect 3176 39136 3192 39200
rect 3256 39136 3262 39200
rect 2946 39135 3262 39136
rect 4546 39200 4862 39201
rect 4546 39136 4552 39200
rect 4616 39136 4632 39200
rect 4696 39136 4712 39200
rect 4776 39136 4792 39200
rect 4856 39136 4862 39200
rect 4546 39135 4862 39136
rect 6146 39200 6462 39201
rect 6146 39136 6152 39200
rect 6216 39136 6232 39200
rect 6296 39136 6312 39200
rect 6376 39136 6392 39200
rect 6456 39136 6462 39200
rect 6146 39135 6462 39136
rect 7746 39200 8062 39201
rect 7746 39136 7752 39200
rect 7816 39136 7832 39200
rect 7896 39136 7912 39200
rect 7976 39136 7992 39200
rect 8056 39136 8062 39200
rect 7746 39135 8062 39136
rect 9346 39200 9662 39201
rect 9346 39136 9352 39200
rect 9416 39136 9432 39200
rect 9496 39136 9512 39200
rect 9576 39136 9592 39200
rect 9656 39136 9662 39200
rect 9346 39135 9662 39136
rect 1025 38722 1091 38725
rect 0 38720 1091 38722
rect 0 38664 1030 38720
rect 1086 38664 1091 38720
rect 0 38662 1091 38664
rect 1025 38659 1091 38662
rect 3606 38656 3922 38657
rect 3606 38592 3612 38656
rect 3676 38592 3692 38656
rect 3756 38592 3772 38656
rect 3836 38592 3852 38656
rect 3916 38592 3922 38656
rect 3606 38591 3922 38592
rect 5206 38656 5522 38657
rect 5206 38592 5212 38656
rect 5276 38592 5292 38656
rect 5356 38592 5372 38656
rect 5436 38592 5452 38656
rect 5516 38592 5522 38656
rect 5206 38591 5522 38592
rect 6806 38656 7122 38657
rect 6806 38592 6812 38656
rect 6876 38592 6892 38656
rect 6956 38592 6972 38656
rect 7036 38592 7052 38656
rect 7116 38592 7122 38656
rect 6806 38591 7122 38592
rect 8406 38656 8722 38657
rect 8406 38592 8412 38656
rect 8476 38592 8492 38656
rect 8556 38592 8572 38656
rect 8636 38592 8652 38656
rect 8716 38592 8722 38656
rect 8406 38591 8722 38592
rect 8201 38450 8267 38453
rect 10542 38450 10548 38452
rect 8201 38448 10548 38450
rect 8201 38392 8206 38448
rect 8262 38392 10548 38448
rect 8201 38390 10548 38392
rect 8201 38387 8267 38390
rect 10542 38388 10548 38390
rect 10612 38388 10618 38452
rect 10501 38178 10567 38181
rect 11470 38178 12052 38204
rect 10501 38176 12052 38178
rect 10501 38120 10506 38176
rect 10562 38144 12052 38176
rect 10562 38120 11530 38144
rect 10501 38118 11530 38120
rect 10501 38115 10567 38118
rect 2946 38112 3262 38113
rect 2946 38048 2952 38112
rect 3016 38048 3032 38112
rect 3096 38048 3112 38112
rect 3176 38048 3192 38112
rect 3256 38048 3262 38112
rect 2946 38047 3262 38048
rect 4546 38112 4862 38113
rect 4546 38048 4552 38112
rect 4616 38048 4632 38112
rect 4696 38048 4712 38112
rect 4776 38048 4792 38112
rect 4856 38048 4862 38112
rect 4546 38047 4862 38048
rect 6146 38112 6462 38113
rect 6146 38048 6152 38112
rect 6216 38048 6232 38112
rect 6296 38048 6312 38112
rect 6376 38048 6392 38112
rect 6456 38048 6462 38112
rect 6146 38047 6462 38048
rect 7746 38112 8062 38113
rect 7746 38048 7752 38112
rect 7816 38048 7832 38112
rect 7896 38048 7912 38112
rect 7976 38048 7992 38112
rect 8056 38048 8062 38112
rect 7746 38047 8062 38048
rect 9346 38112 9662 38113
rect 9346 38048 9352 38112
rect 9416 38048 9432 38112
rect 9496 38048 9512 38112
rect 9576 38048 9592 38112
rect 9656 38048 9662 38112
rect 9346 38047 9662 38048
rect 1025 37770 1091 37773
rect 0 37768 1091 37770
rect 0 37712 1030 37768
rect 1086 37712 1091 37768
rect 0 37710 1091 37712
rect 1025 37707 1091 37710
rect 3606 37568 3922 37569
rect 3606 37504 3612 37568
rect 3676 37504 3692 37568
rect 3756 37504 3772 37568
rect 3836 37504 3852 37568
rect 3916 37504 3922 37568
rect 3606 37503 3922 37504
rect 5206 37568 5522 37569
rect 5206 37504 5212 37568
rect 5276 37504 5292 37568
rect 5356 37504 5372 37568
rect 5436 37504 5452 37568
rect 5516 37504 5522 37568
rect 5206 37503 5522 37504
rect 6806 37568 7122 37569
rect 6806 37504 6812 37568
rect 6876 37504 6892 37568
rect 6956 37504 6972 37568
rect 7036 37504 7052 37568
rect 7116 37504 7122 37568
rect 6806 37503 7122 37504
rect 8406 37568 8722 37569
rect 8406 37504 8412 37568
rect 8476 37504 8492 37568
rect 8556 37504 8572 37568
rect 8636 37504 8652 37568
rect 8716 37504 8722 37568
rect 8406 37503 8722 37504
rect 790 37300 796 37364
rect 860 37362 866 37364
rect 6913 37362 6979 37365
rect 860 37360 6979 37362
rect 860 37304 6918 37360
rect 6974 37304 6979 37360
rect 860 37302 6979 37304
rect 860 37300 866 37302
rect 6913 37299 6979 37302
rect 9765 37362 9831 37365
rect 10726 37362 10732 37364
rect 9765 37360 10732 37362
rect 9765 37304 9770 37360
rect 9826 37304 10732 37360
rect 9765 37302 10732 37304
rect 9765 37299 9831 37302
rect 10726 37300 10732 37302
rect 10796 37300 10802 37364
rect 2946 37024 3262 37025
rect 2946 36960 2952 37024
rect 3016 36960 3032 37024
rect 3096 36960 3112 37024
rect 3176 36960 3192 37024
rect 3256 36960 3262 37024
rect 2946 36959 3262 36960
rect 4546 37024 4862 37025
rect 4546 36960 4552 37024
rect 4616 36960 4632 37024
rect 4696 36960 4712 37024
rect 4776 36960 4792 37024
rect 4856 36960 4862 37024
rect 4546 36959 4862 36960
rect 6146 37024 6462 37025
rect 6146 36960 6152 37024
rect 6216 36960 6232 37024
rect 6296 36960 6312 37024
rect 6376 36960 6392 37024
rect 6456 36960 6462 37024
rect 6146 36959 6462 36960
rect 7746 37024 8062 37025
rect 7746 36960 7752 37024
rect 7816 36960 7832 37024
rect 7896 36960 7912 37024
rect 7976 36960 7992 37024
rect 8056 36960 8062 37024
rect 7746 36959 8062 36960
rect 9346 37024 9662 37025
rect 9346 36960 9352 37024
rect 9416 36960 9432 37024
rect 9496 36960 9512 37024
rect 9576 36960 9592 37024
rect 9656 36960 9662 37024
rect 9346 36959 9662 36960
rect 11470 36920 12052 36980
rect 1025 36818 1091 36821
rect 0 36816 1091 36818
rect 0 36760 1030 36816
rect 1086 36760 1091 36816
rect 0 36758 1091 36760
rect 1025 36755 1091 36758
rect 8293 36818 8359 36821
rect 11470 36818 11530 36920
rect 8293 36816 11530 36818
rect 8293 36760 8298 36816
rect 8354 36760 11530 36816
rect 8293 36758 11530 36760
rect 8293 36755 8359 36758
rect 4337 36682 4403 36685
rect 4294 36680 4403 36682
rect 4294 36624 4342 36680
rect 4398 36624 4403 36680
rect 4294 36619 4403 36624
rect 3606 36480 3922 36481
rect 3606 36416 3612 36480
rect 3676 36416 3692 36480
rect 3756 36416 3772 36480
rect 3836 36416 3852 36480
rect 3916 36416 3922 36480
rect 3606 36415 3922 36416
rect 4294 36413 4354 36619
rect 5206 36480 5522 36481
rect 5206 36416 5212 36480
rect 5276 36416 5292 36480
rect 5356 36416 5372 36480
rect 5436 36416 5452 36480
rect 5516 36416 5522 36480
rect 5206 36415 5522 36416
rect 6806 36480 7122 36481
rect 6806 36416 6812 36480
rect 6876 36416 6892 36480
rect 6956 36416 6972 36480
rect 7036 36416 7052 36480
rect 7116 36416 7122 36480
rect 6806 36415 7122 36416
rect 8406 36480 8722 36481
rect 8406 36416 8412 36480
rect 8476 36416 8492 36480
rect 8556 36416 8572 36480
rect 8636 36416 8652 36480
rect 8716 36416 8722 36480
rect 8406 36415 8722 36416
rect 4245 36408 4354 36413
rect 4245 36352 4250 36408
rect 4306 36352 4354 36408
rect 4245 36350 4354 36352
rect 8845 36410 8911 36413
rect 11646 36410 11652 36412
rect 8845 36408 11652 36410
rect 8845 36352 8850 36408
rect 8906 36352 11652 36408
rect 8845 36350 11652 36352
rect 4245 36347 4311 36350
rect 8845 36347 8911 36350
rect 11646 36348 11652 36350
rect 11716 36348 11722 36412
rect 2946 35936 3262 35937
rect 2946 35872 2952 35936
rect 3016 35872 3032 35936
rect 3096 35872 3112 35936
rect 3176 35872 3192 35936
rect 3256 35872 3262 35936
rect 2946 35871 3262 35872
rect 4546 35936 4862 35937
rect 4546 35872 4552 35936
rect 4616 35872 4632 35936
rect 4696 35872 4712 35936
rect 4776 35872 4792 35936
rect 4856 35872 4862 35936
rect 4546 35871 4862 35872
rect 6146 35936 6462 35937
rect 6146 35872 6152 35936
rect 6216 35872 6232 35936
rect 6296 35872 6312 35936
rect 6376 35872 6392 35936
rect 6456 35872 6462 35936
rect 6146 35871 6462 35872
rect 7746 35936 8062 35937
rect 7746 35872 7752 35936
rect 7816 35872 7832 35936
rect 7896 35872 7912 35936
rect 7976 35872 7992 35936
rect 8056 35872 8062 35936
rect 7746 35871 8062 35872
rect 9346 35936 9662 35937
rect 9346 35872 9352 35936
rect 9416 35872 9432 35936
rect 9496 35872 9512 35936
rect 9576 35872 9592 35936
rect 9656 35872 9662 35936
rect 9346 35871 9662 35872
rect 1393 35866 1459 35869
rect 0 35864 1459 35866
rect 0 35808 1398 35864
rect 1454 35808 1459 35864
rect 0 35806 1459 35808
rect 1393 35803 1459 35806
rect 3606 35392 3922 35393
rect 3606 35328 3612 35392
rect 3676 35328 3692 35392
rect 3756 35328 3772 35392
rect 3836 35328 3852 35392
rect 3916 35328 3922 35392
rect 3606 35327 3922 35328
rect 5206 35392 5522 35393
rect 5206 35328 5212 35392
rect 5276 35328 5292 35392
rect 5356 35328 5372 35392
rect 5436 35328 5452 35392
rect 5516 35328 5522 35392
rect 5206 35327 5522 35328
rect 6806 35392 7122 35393
rect 6806 35328 6812 35392
rect 6876 35328 6892 35392
rect 6956 35328 6972 35392
rect 7036 35328 7052 35392
rect 7116 35328 7122 35392
rect 6806 35327 7122 35328
rect 8406 35392 8722 35393
rect 8406 35328 8412 35392
rect 8476 35328 8492 35392
rect 8556 35328 8572 35392
rect 8636 35328 8652 35392
rect 8716 35328 8722 35392
rect 8406 35327 8722 35328
rect 8293 35186 8359 35189
rect 11470 35186 12052 35212
rect 8293 35184 12052 35186
rect 8293 35128 8298 35184
rect 8354 35152 12052 35184
rect 8354 35128 11530 35152
rect 8293 35126 11530 35128
rect 8293 35123 8359 35126
rect 933 34914 999 34917
rect 0 34912 999 34914
rect 0 34856 938 34912
rect 994 34856 999 34912
rect 0 34854 999 34856
rect 933 34851 999 34854
rect 2946 34848 3262 34849
rect 2946 34784 2952 34848
rect 3016 34784 3032 34848
rect 3096 34784 3112 34848
rect 3176 34784 3192 34848
rect 3256 34784 3262 34848
rect 2946 34783 3262 34784
rect 4546 34848 4862 34849
rect 4546 34784 4552 34848
rect 4616 34784 4632 34848
rect 4696 34784 4712 34848
rect 4776 34784 4792 34848
rect 4856 34784 4862 34848
rect 4546 34783 4862 34784
rect 6146 34848 6462 34849
rect 6146 34784 6152 34848
rect 6216 34784 6232 34848
rect 6296 34784 6312 34848
rect 6376 34784 6392 34848
rect 6456 34784 6462 34848
rect 6146 34783 6462 34784
rect 7746 34848 8062 34849
rect 7746 34784 7752 34848
rect 7816 34784 7832 34848
rect 7896 34784 7912 34848
rect 7976 34784 7992 34848
rect 8056 34784 8062 34848
rect 7746 34783 8062 34784
rect 9346 34848 9662 34849
rect 9346 34784 9352 34848
rect 9416 34784 9432 34848
rect 9496 34784 9512 34848
rect 9576 34784 9592 34848
rect 9656 34784 9662 34848
rect 9346 34783 9662 34784
rect 3606 34304 3922 34305
rect 3606 34240 3612 34304
rect 3676 34240 3692 34304
rect 3756 34240 3772 34304
rect 3836 34240 3852 34304
rect 3916 34240 3922 34304
rect 3606 34239 3922 34240
rect 5206 34304 5522 34305
rect 5206 34240 5212 34304
rect 5276 34240 5292 34304
rect 5356 34240 5372 34304
rect 5436 34240 5452 34304
rect 5516 34240 5522 34304
rect 5206 34239 5522 34240
rect 6806 34304 7122 34305
rect 6806 34240 6812 34304
rect 6876 34240 6892 34304
rect 6956 34240 6972 34304
rect 7036 34240 7052 34304
rect 7116 34240 7122 34304
rect 6806 34239 7122 34240
rect 8406 34304 8722 34305
rect 8406 34240 8412 34304
rect 8476 34240 8492 34304
rect 8556 34240 8572 34304
rect 8636 34240 8652 34304
rect 8716 34240 8722 34304
rect 8406 34239 8722 34240
rect 11830 34062 11836 34126
rect 11900 34124 11906 34126
rect 11900 34064 12052 34124
rect 11900 34062 11906 34064
rect 933 33962 999 33965
rect 0 33960 999 33962
rect 0 33904 938 33960
rect 994 33904 999 33960
rect 0 33902 999 33904
rect 933 33899 999 33902
rect 2946 33760 3262 33761
rect 2946 33696 2952 33760
rect 3016 33696 3032 33760
rect 3096 33696 3112 33760
rect 3176 33696 3192 33760
rect 3256 33696 3262 33760
rect 2946 33695 3262 33696
rect 4546 33760 4862 33761
rect 4546 33696 4552 33760
rect 4616 33696 4632 33760
rect 4696 33696 4712 33760
rect 4776 33696 4792 33760
rect 4856 33696 4862 33760
rect 4546 33695 4862 33696
rect 6146 33760 6462 33761
rect 6146 33696 6152 33760
rect 6216 33696 6232 33760
rect 6296 33696 6312 33760
rect 6376 33696 6392 33760
rect 6456 33696 6462 33760
rect 6146 33695 6462 33696
rect 7746 33760 8062 33761
rect 7746 33696 7752 33760
rect 7816 33696 7832 33760
rect 7896 33696 7912 33760
rect 7976 33696 7992 33760
rect 8056 33696 8062 33760
rect 7746 33695 8062 33696
rect 9346 33760 9662 33761
rect 9346 33696 9352 33760
rect 9416 33696 9432 33760
rect 9496 33696 9512 33760
rect 9576 33696 9592 33760
rect 9656 33696 9662 33760
rect 9346 33695 9662 33696
rect 3606 33216 3922 33217
rect 3606 33152 3612 33216
rect 3676 33152 3692 33216
rect 3756 33152 3772 33216
rect 3836 33152 3852 33216
rect 3916 33152 3922 33216
rect 3606 33151 3922 33152
rect 5206 33216 5522 33217
rect 5206 33152 5212 33216
rect 5276 33152 5292 33216
rect 5356 33152 5372 33216
rect 5436 33152 5452 33216
rect 5516 33152 5522 33216
rect 5206 33151 5522 33152
rect 6806 33216 7122 33217
rect 6806 33152 6812 33216
rect 6876 33152 6892 33216
rect 6956 33152 6972 33216
rect 7036 33152 7052 33216
rect 7116 33152 7122 33216
rect 6806 33151 7122 33152
rect 8406 33216 8722 33217
rect 8406 33152 8412 33216
rect 8476 33152 8492 33216
rect 8556 33152 8572 33216
rect 8636 33152 8652 33216
rect 8716 33152 8722 33216
rect 8406 33151 8722 33152
rect 1485 33146 1551 33149
rect 798 33144 1551 33146
rect 798 33088 1490 33144
rect 1546 33088 1551 33144
rect 798 33086 1551 33088
rect 798 33010 858 33086
rect 1485 33083 1551 33086
rect 0 32950 858 33010
rect 2946 32672 3262 32673
rect 2946 32608 2952 32672
rect 3016 32608 3032 32672
rect 3096 32608 3112 32672
rect 3176 32608 3192 32672
rect 3256 32608 3262 32672
rect 2946 32607 3262 32608
rect 4546 32672 4862 32673
rect 4546 32608 4552 32672
rect 4616 32608 4632 32672
rect 4696 32608 4712 32672
rect 4776 32608 4792 32672
rect 4856 32608 4862 32672
rect 4546 32607 4862 32608
rect 6146 32672 6462 32673
rect 6146 32608 6152 32672
rect 6216 32608 6232 32672
rect 6296 32608 6312 32672
rect 6376 32608 6392 32672
rect 6456 32608 6462 32672
rect 6146 32607 6462 32608
rect 7746 32672 8062 32673
rect 7746 32608 7752 32672
rect 7816 32608 7832 32672
rect 7896 32608 7912 32672
rect 7976 32608 7992 32672
rect 8056 32608 8062 32672
rect 7746 32607 8062 32608
rect 9346 32672 9662 32673
rect 9346 32608 9352 32672
rect 9416 32608 9432 32672
rect 9496 32608 9512 32672
rect 9576 32608 9592 32672
rect 9656 32608 9662 32672
rect 9346 32607 9662 32608
rect 11789 32492 11855 32495
rect 11789 32490 12052 32492
rect 11789 32434 11794 32490
rect 11850 32434 12052 32490
rect 11789 32432 12052 32434
rect 11789 32429 11855 32432
rect 7281 32330 7347 32333
rect 7238 32328 7347 32330
rect 7238 32272 7286 32328
rect 7342 32272 7347 32328
rect 7238 32267 7347 32272
rect 3606 32128 3922 32129
rect 3606 32064 3612 32128
rect 3676 32064 3692 32128
rect 3756 32064 3772 32128
rect 3836 32064 3852 32128
rect 3916 32064 3922 32128
rect 3606 32063 3922 32064
rect 5206 32128 5522 32129
rect 5206 32064 5212 32128
rect 5276 32064 5292 32128
rect 5356 32064 5372 32128
rect 5436 32064 5452 32128
rect 5516 32064 5522 32128
rect 5206 32063 5522 32064
rect 6806 32128 7122 32129
rect 6806 32064 6812 32128
rect 6876 32064 6892 32128
rect 6956 32064 6972 32128
rect 7036 32064 7052 32128
rect 7116 32064 7122 32128
rect 6806 32063 7122 32064
rect 933 32058 999 32061
rect 0 32056 999 32058
rect 0 32000 938 32056
rect 994 32000 999 32056
rect 0 31998 999 32000
rect 933 31995 999 31998
rect 5993 31922 6059 31925
rect 5950 31920 6059 31922
rect 5950 31864 5998 31920
rect 6054 31864 6059 31920
rect 5950 31859 6059 31864
rect 7005 31922 7071 31925
rect 7238 31922 7298 32267
rect 8406 32128 8722 32129
rect 8406 32064 8412 32128
rect 8476 32064 8492 32128
rect 8556 32064 8572 32128
rect 8636 32064 8652 32128
rect 8716 32064 8722 32128
rect 8406 32063 8722 32064
rect 7005 31920 7298 31922
rect 7005 31864 7010 31920
rect 7066 31864 7298 31920
rect 7005 31862 7298 31864
rect 7005 31859 7071 31862
rect 2946 31584 3262 31585
rect 2946 31520 2952 31584
rect 3016 31520 3032 31584
rect 3096 31520 3112 31584
rect 3176 31520 3192 31584
rect 3256 31520 3262 31584
rect 2946 31519 3262 31520
rect 4546 31584 4862 31585
rect 4546 31520 4552 31584
rect 4616 31520 4632 31584
rect 4696 31520 4712 31584
rect 4776 31520 4792 31584
rect 4856 31520 4862 31584
rect 4546 31519 4862 31520
rect 5950 31381 6010 31859
rect 8937 31786 9003 31789
rect 9489 31786 9555 31789
rect 8937 31784 9555 31786
rect 8937 31728 8942 31784
rect 8998 31728 9494 31784
rect 9550 31728 9555 31784
rect 8937 31726 9555 31728
rect 8937 31723 9003 31726
rect 9489 31723 9555 31726
rect 6146 31584 6462 31585
rect 6146 31520 6152 31584
rect 6216 31520 6232 31584
rect 6296 31520 6312 31584
rect 6376 31520 6392 31584
rect 6456 31520 6462 31584
rect 6146 31519 6462 31520
rect 7746 31584 8062 31585
rect 7746 31520 7752 31584
rect 7816 31520 7832 31584
rect 7896 31520 7912 31584
rect 7976 31520 7992 31584
rect 8056 31520 8062 31584
rect 7746 31519 8062 31520
rect 9346 31584 9662 31585
rect 9346 31520 9352 31584
rect 9416 31520 9432 31584
rect 9496 31520 9512 31584
rect 9576 31520 9592 31584
rect 9656 31520 9662 31584
rect 9346 31519 9662 31520
rect 10409 31514 10475 31517
rect 11470 31514 12052 31540
rect 10409 31512 12052 31514
rect 10409 31456 10414 31512
rect 10470 31480 12052 31512
rect 10470 31456 11530 31480
rect 10409 31454 11530 31456
rect 10409 31451 10475 31454
rect 5950 31376 6059 31381
rect 5950 31320 5998 31376
rect 6054 31320 6059 31376
rect 5950 31318 6059 31320
rect 5993 31315 6059 31318
rect 933 31106 999 31109
rect 0 31104 999 31106
rect 0 31048 938 31104
rect 994 31048 999 31104
rect 0 31046 999 31048
rect 933 31043 999 31046
rect 3606 31040 3922 31041
rect 3606 30976 3612 31040
rect 3676 30976 3692 31040
rect 3756 30976 3772 31040
rect 3836 30976 3852 31040
rect 3916 30976 3922 31040
rect 3606 30975 3922 30976
rect 5206 31040 5522 31041
rect 5206 30976 5212 31040
rect 5276 30976 5292 31040
rect 5356 30976 5372 31040
rect 5436 30976 5452 31040
rect 5516 30976 5522 31040
rect 5206 30975 5522 30976
rect 6806 31040 7122 31041
rect 6806 30976 6812 31040
rect 6876 30976 6892 31040
rect 6956 30976 6972 31040
rect 7036 30976 7052 31040
rect 7116 30976 7122 31040
rect 6806 30975 7122 30976
rect 8406 31040 8722 31041
rect 8406 30976 8412 31040
rect 8476 30976 8492 31040
rect 8556 30976 8572 31040
rect 8636 30976 8652 31040
rect 8716 30976 8722 31040
rect 8406 30975 8722 30976
rect 6085 30698 6151 30701
rect 5950 30696 6151 30698
rect 5950 30640 6090 30696
rect 6146 30640 6151 30696
rect 5950 30638 6151 30640
rect 2946 30496 3262 30497
rect 2946 30432 2952 30496
rect 3016 30432 3032 30496
rect 3096 30432 3112 30496
rect 3176 30432 3192 30496
rect 3256 30432 3262 30496
rect 2946 30431 3262 30432
rect 4546 30496 4862 30497
rect 4546 30432 4552 30496
rect 4616 30432 4632 30496
rect 4696 30432 4712 30496
rect 4776 30432 4792 30496
rect 4856 30432 4862 30496
rect 4546 30431 4862 30432
rect 933 30154 999 30157
rect 0 30152 999 30154
rect 0 30096 938 30152
rect 994 30096 999 30152
rect 0 30094 999 30096
rect 933 30091 999 30094
rect 3606 29952 3922 29953
rect 3606 29888 3612 29952
rect 3676 29888 3692 29952
rect 3756 29888 3772 29952
rect 3836 29888 3852 29952
rect 3916 29888 3922 29952
rect 3606 29887 3922 29888
rect 5206 29952 5522 29953
rect 5206 29888 5212 29952
rect 5276 29888 5292 29952
rect 5356 29888 5372 29952
rect 5436 29888 5452 29952
rect 5516 29888 5522 29952
rect 5206 29887 5522 29888
rect 2946 29408 3262 29409
rect 2946 29344 2952 29408
rect 3016 29344 3032 29408
rect 3096 29344 3112 29408
rect 3176 29344 3192 29408
rect 3256 29344 3262 29408
rect 2946 29343 3262 29344
rect 4546 29408 4862 29409
rect 4546 29344 4552 29408
rect 4616 29344 4632 29408
rect 4696 29344 4712 29408
rect 4776 29344 4792 29408
rect 4856 29344 4862 29408
rect 4546 29343 4862 29344
rect 933 29202 999 29205
rect 0 29200 999 29202
rect 0 29144 938 29200
rect 994 29144 999 29200
rect 0 29142 999 29144
rect 5950 29202 6010 30638
rect 6085 30635 6151 30638
rect 6146 30496 6462 30497
rect 6146 30432 6152 30496
rect 6216 30432 6232 30496
rect 6296 30432 6312 30496
rect 6376 30432 6392 30496
rect 6456 30432 6462 30496
rect 6146 30431 6462 30432
rect 7746 30496 8062 30497
rect 7746 30432 7752 30496
rect 7816 30432 7832 30496
rect 7896 30432 7912 30496
rect 7976 30432 7992 30496
rect 8056 30432 8062 30496
rect 7746 30431 8062 30432
rect 9346 30496 9662 30497
rect 9346 30432 9352 30496
rect 9416 30432 9432 30496
rect 9496 30432 9512 30496
rect 9576 30432 9592 30496
rect 9656 30432 9662 30496
rect 9346 30431 9662 30432
rect 6806 29952 7122 29953
rect 6806 29888 6812 29952
rect 6876 29888 6892 29952
rect 6956 29888 6972 29952
rect 7036 29888 7052 29952
rect 7116 29888 7122 29952
rect 6806 29887 7122 29888
rect 8406 29952 8722 29953
rect 8406 29888 8412 29952
rect 8476 29888 8492 29952
rect 8556 29888 8572 29952
rect 8636 29888 8652 29952
rect 8716 29888 8722 29952
rect 8406 29887 8722 29888
rect 10317 29746 10383 29749
rect 11470 29746 12052 29772
rect 10317 29744 12052 29746
rect 10317 29688 10322 29744
rect 10378 29712 12052 29744
rect 10378 29688 11530 29712
rect 10317 29686 11530 29688
rect 10317 29683 10383 29686
rect 6146 29408 6462 29409
rect 6146 29344 6152 29408
rect 6216 29344 6232 29408
rect 6296 29344 6312 29408
rect 6376 29344 6392 29408
rect 6456 29344 6462 29408
rect 6146 29343 6462 29344
rect 7746 29408 8062 29409
rect 7746 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8062 29408
rect 7746 29343 8062 29344
rect 9346 29408 9662 29409
rect 9346 29344 9352 29408
rect 9416 29344 9432 29408
rect 9496 29344 9512 29408
rect 9576 29344 9592 29408
rect 9656 29344 9662 29408
rect 9346 29343 9662 29344
rect 6085 29202 6151 29205
rect 5950 29200 6151 29202
rect 5950 29144 6090 29200
rect 6146 29144 6151 29200
rect 5950 29142 6151 29144
rect 933 29139 999 29142
rect 6085 29139 6151 29142
rect 3606 28864 3922 28865
rect 3606 28800 3612 28864
rect 3676 28800 3692 28864
rect 3756 28800 3772 28864
rect 3836 28800 3852 28864
rect 3916 28800 3922 28864
rect 3606 28799 3922 28800
rect 5206 28864 5522 28865
rect 5206 28800 5212 28864
rect 5276 28800 5292 28864
rect 5356 28800 5372 28864
rect 5436 28800 5452 28864
rect 5516 28800 5522 28864
rect 5206 28799 5522 28800
rect 6806 28864 7122 28865
rect 6806 28800 6812 28864
rect 6876 28800 6892 28864
rect 6956 28800 6972 28864
rect 7036 28800 7052 28864
rect 7116 28800 7122 28864
rect 6806 28799 7122 28800
rect 8406 28864 8722 28865
rect 8406 28800 8412 28864
rect 8476 28800 8492 28864
rect 8556 28800 8572 28864
rect 8636 28800 8652 28864
rect 8716 28800 8722 28864
rect 8406 28799 8722 28800
rect 5901 28522 5967 28525
rect 7925 28522 7991 28525
rect 5901 28520 6010 28522
rect 5901 28464 5906 28520
rect 5962 28464 6010 28520
rect 5901 28459 6010 28464
rect 2946 28320 3262 28321
rect 2946 28256 2952 28320
rect 3016 28256 3032 28320
rect 3096 28256 3112 28320
rect 3176 28256 3192 28320
rect 3256 28256 3262 28320
rect 2946 28255 3262 28256
rect 4546 28320 4862 28321
rect 4546 28256 4552 28320
rect 4616 28256 4632 28320
rect 4696 28256 4712 28320
rect 4776 28256 4792 28320
rect 4856 28256 4862 28320
rect 4546 28255 4862 28256
rect 5950 28253 6010 28459
rect 7468 28520 7991 28522
rect 7468 28464 7930 28520
rect 7986 28464 7991 28520
rect 7468 28462 7991 28464
rect 7468 28389 7528 28462
rect 7925 28459 7991 28462
rect 7465 28384 7531 28389
rect 7465 28328 7470 28384
rect 7526 28328 7531 28384
rect 7465 28323 7531 28328
rect 6146 28320 6462 28321
rect 6146 28256 6152 28320
rect 6216 28256 6232 28320
rect 6296 28256 6312 28320
rect 6376 28256 6392 28320
rect 6456 28256 6462 28320
rect 6146 28255 6462 28256
rect 7746 28320 8062 28321
rect 7746 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8062 28320
rect 7746 28255 8062 28256
rect 9346 28320 9662 28321
rect 9346 28256 9352 28320
rect 9416 28256 9432 28320
rect 9496 28256 9512 28320
rect 9576 28256 9592 28320
rect 9656 28256 9662 28320
rect 9346 28255 9662 28256
rect 933 28250 999 28253
rect 0 28248 999 28250
rect 0 28192 938 28248
rect 994 28192 999 28248
rect 0 28190 999 28192
rect 933 28187 999 28190
rect 5901 28248 6010 28253
rect 5901 28192 5906 28248
rect 5962 28192 6010 28248
rect 5901 28190 6010 28192
rect 5901 28187 5967 28190
rect 5441 27978 5507 27981
rect 7005 27978 7071 27981
rect 5441 27976 5642 27978
rect 5441 27920 5446 27976
rect 5502 27920 5642 27976
rect 5441 27918 5642 27920
rect 5441 27915 5507 27918
rect 3606 27776 3922 27777
rect 3606 27712 3612 27776
rect 3676 27712 3692 27776
rect 3756 27712 3772 27776
rect 3836 27712 3852 27776
rect 3916 27712 3922 27776
rect 3606 27711 3922 27712
rect 5206 27776 5522 27777
rect 5206 27712 5212 27776
rect 5276 27712 5292 27776
rect 5356 27712 5372 27776
rect 5436 27712 5452 27776
rect 5516 27712 5522 27776
rect 5206 27711 5522 27712
rect 5441 27570 5507 27573
rect 5582 27570 5642 27918
rect 7005 27976 7298 27978
rect 7005 27920 7010 27976
rect 7066 27920 7298 27976
rect 7005 27918 7298 27920
rect 7005 27915 7071 27918
rect 6806 27776 7122 27777
rect 6806 27712 6812 27776
rect 6876 27712 6892 27776
rect 6956 27712 6972 27776
rect 7036 27712 7052 27776
rect 7116 27712 7122 27776
rect 6806 27711 7122 27712
rect 7238 27573 7298 27918
rect 8406 27776 8722 27777
rect 8406 27712 8412 27776
rect 8476 27712 8492 27776
rect 8556 27712 8572 27776
rect 8636 27712 8652 27776
rect 8716 27712 8722 27776
rect 8406 27711 8722 27712
rect 5441 27568 5642 27570
rect 5441 27512 5446 27568
rect 5502 27512 5642 27568
rect 5441 27510 5642 27512
rect 7189 27568 7298 27573
rect 7189 27512 7194 27568
rect 7250 27512 7298 27568
rect 7189 27510 7298 27512
rect 5441 27507 5507 27510
rect 7189 27507 7255 27510
rect 933 27298 999 27301
rect 0 27296 999 27298
rect 0 27240 938 27296
rect 994 27240 999 27296
rect 0 27238 999 27240
rect 933 27235 999 27238
rect 2946 27232 3262 27233
rect 2946 27168 2952 27232
rect 3016 27168 3032 27232
rect 3096 27168 3112 27232
rect 3176 27168 3192 27232
rect 3256 27168 3262 27232
rect 2946 27167 3262 27168
rect 4546 27232 4862 27233
rect 4546 27168 4552 27232
rect 4616 27168 4632 27232
rect 4696 27168 4712 27232
rect 4776 27168 4792 27232
rect 4856 27168 4862 27232
rect 4546 27167 4862 27168
rect 6146 27232 6462 27233
rect 6146 27168 6152 27232
rect 6216 27168 6232 27232
rect 6296 27168 6312 27232
rect 6376 27168 6392 27232
rect 6456 27168 6462 27232
rect 6146 27167 6462 27168
rect 7746 27232 8062 27233
rect 7746 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8062 27232
rect 7746 27167 8062 27168
rect 9346 27232 9662 27233
rect 9346 27168 9352 27232
rect 9416 27168 9432 27232
rect 9496 27168 9512 27232
rect 9576 27168 9592 27232
rect 9656 27168 9662 27232
rect 9346 27167 9662 27168
rect 3606 26688 3922 26689
rect 3606 26624 3612 26688
rect 3676 26624 3692 26688
rect 3756 26624 3772 26688
rect 3836 26624 3852 26688
rect 3916 26624 3922 26688
rect 3606 26623 3922 26624
rect 5206 26688 5522 26689
rect 5206 26624 5212 26688
rect 5276 26624 5292 26688
rect 5356 26624 5372 26688
rect 5436 26624 5452 26688
rect 5516 26624 5522 26688
rect 5206 26623 5522 26624
rect 6806 26688 7122 26689
rect 6806 26624 6812 26688
rect 6876 26624 6892 26688
rect 6956 26624 6972 26688
rect 7036 26624 7052 26688
rect 7116 26624 7122 26688
rect 6806 26623 7122 26624
rect 8406 26688 8722 26689
rect 8406 26624 8412 26688
rect 8476 26624 8492 26688
rect 8556 26624 8572 26688
rect 8636 26624 8652 26688
rect 8716 26624 8722 26688
rect 8406 26623 8722 26624
rect 933 26346 999 26349
rect 6085 26346 6151 26349
rect 0 26344 999 26346
rect 0 26288 938 26344
rect 994 26288 999 26344
rect 0 26286 999 26288
rect 933 26283 999 26286
rect 5950 26344 6151 26346
rect 5950 26288 6090 26344
rect 6146 26288 6151 26344
rect 5950 26286 6151 26288
rect 2946 26144 3262 26145
rect 2946 26080 2952 26144
rect 3016 26080 3032 26144
rect 3096 26080 3112 26144
rect 3176 26080 3192 26144
rect 3256 26080 3262 26144
rect 2946 26079 3262 26080
rect 4546 26144 4862 26145
rect 4546 26080 4552 26144
rect 4616 26080 4632 26144
rect 4696 26080 4712 26144
rect 4776 26080 4792 26144
rect 4856 26080 4862 26144
rect 4546 26079 4862 26080
rect 5809 25938 5875 25941
rect 5950 25938 6010 26286
rect 6085 26283 6151 26286
rect 6146 26144 6462 26145
rect 6146 26080 6152 26144
rect 6216 26080 6232 26144
rect 6296 26080 6312 26144
rect 6376 26080 6392 26144
rect 6456 26080 6462 26144
rect 6146 26079 6462 26080
rect 7746 26144 8062 26145
rect 7746 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8062 26144
rect 7746 26079 8062 26080
rect 9346 26144 9662 26145
rect 9346 26080 9352 26144
rect 9416 26080 9432 26144
rect 9496 26080 9512 26144
rect 9576 26080 9592 26144
rect 9656 26080 9662 26144
rect 9346 26079 9662 26080
rect 5809 25936 6010 25938
rect 5809 25880 5814 25936
rect 5870 25880 6010 25936
rect 5809 25878 6010 25880
rect 5809 25875 5875 25878
rect 7649 25802 7715 25805
rect 11830 25802 11836 25804
rect 7649 25800 11836 25802
rect 7649 25744 7654 25800
rect 7710 25744 11836 25800
rect 7649 25742 11836 25744
rect 7649 25739 7715 25742
rect 11830 25740 11836 25742
rect 11900 25740 11906 25804
rect 3606 25600 3922 25601
rect 3606 25536 3612 25600
rect 3676 25536 3692 25600
rect 3756 25536 3772 25600
rect 3836 25536 3852 25600
rect 3916 25536 3922 25600
rect 3606 25535 3922 25536
rect 5206 25600 5522 25601
rect 5206 25536 5212 25600
rect 5276 25536 5292 25600
rect 5356 25536 5372 25600
rect 5436 25536 5452 25600
rect 5516 25536 5522 25600
rect 5206 25535 5522 25536
rect 6806 25600 7122 25601
rect 6806 25536 6812 25600
rect 6876 25536 6892 25600
rect 6956 25536 6972 25600
rect 7036 25536 7052 25600
rect 7116 25536 7122 25600
rect 6806 25535 7122 25536
rect 8406 25600 8722 25601
rect 8406 25536 8412 25600
rect 8476 25536 8492 25600
rect 8556 25536 8572 25600
rect 8636 25536 8652 25600
rect 8716 25536 8722 25600
rect 8406 25535 8722 25536
rect 933 25394 999 25397
rect 0 25392 999 25394
rect 0 25336 938 25392
rect 994 25336 999 25392
rect 0 25334 999 25336
rect 933 25331 999 25334
rect 2946 25056 3262 25057
rect 2946 24992 2952 25056
rect 3016 24992 3032 25056
rect 3096 24992 3112 25056
rect 3176 24992 3192 25056
rect 3256 24992 3262 25056
rect 2946 24991 3262 24992
rect 4546 25056 4862 25057
rect 4546 24992 4552 25056
rect 4616 24992 4632 25056
rect 4696 24992 4712 25056
rect 4776 24992 4792 25056
rect 4856 24992 4862 25056
rect 4546 24991 4862 24992
rect 6146 25056 6462 25057
rect 6146 24992 6152 25056
rect 6216 24992 6232 25056
rect 6296 24992 6312 25056
rect 6376 24992 6392 25056
rect 6456 24992 6462 25056
rect 6146 24991 6462 24992
rect 7746 25056 8062 25057
rect 7746 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8062 25056
rect 7746 24991 8062 24992
rect 9346 25056 9662 25057
rect 9346 24992 9352 25056
rect 9416 24992 9432 25056
rect 9496 24992 9512 25056
rect 9576 24992 9592 25056
rect 9656 24992 9662 25056
rect 9346 24991 9662 24992
rect 3606 24512 3922 24513
rect 3606 24448 3612 24512
rect 3676 24448 3692 24512
rect 3756 24448 3772 24512
rect 3836 24448 3852 24512
rect 3916 24448 3922 24512
rect 3606 24447 3922 24448
rect 5206 24512 5522 24513
rect 5206 24448 5212 24512
rect 5276 24448 5292 24512
rect 5356 24448 5372 24512
rect 5436 24448 5452 24512
rect 5516 24448 5522 24512
rect 5206 24447 5522 24448
rect 6806 24512 7122 24513
rect 6806 24448 6812 24512
rect 6876 24448 6892 24512
rect 6956 24448 6972 24512
rect 7036 24448 7052 24512
rect 7116 24448 7122 24512
rect 6806 24447 7122 24448
rect 8406 24512 8722 24513
rect 8406 24448 8412 24512
rect 8476 24448 8492 24512
rect 8556 24448 8572 24512
rect 8636 24448 8652 24512
rect 8716 24448 8722 24512
rect 8406 24447 8722 24448
rect 933 24442 999 24445
rect 0 24440 999 24442
rect 0 24384 938 24440
rect 994 24384 999 24440
rect 0 24382 999 24384
rect 933 24379 999 24382
rect 2946 23968 3262 23969
rect 2946 23904 2952 23968
rect 3016 23904 3032 23968
rect 3096 23904 3112 23968
rect 3176 23904 3192 23968
rect 3256 23904 3262 23968
rect 2946 23903 3262 23904
rect 4546 23968 4862 23969
rect 4546 23904 4552 23968
rect 4616 23904 4632 23968
rect 4696 23904 4712 23968
rect 4776 23904 4792 23968
rect 4856 23904 4862 23968
rect 4546 23903 4862 23904
rect 6146 23968 6462 23969
rect 6146 23904 6152 23968
rect 6216 23904 6232 23968
rect 6296 23904 6312 23968
rect 6376 23904 6392 23968
rect 6456 23904 6462 23968
rect 6146 23903 6462 23904
rect 7746 23968 8062 23969
rect 7746 23904 7752 23968
rect 7816 23904 7832 23968
rect 7896 23904 7912 23968
rect 7976 23904 7992 23968
rect 8056 23904 8062 23968
rect 7746 23903 8062 23904
rect 9346 23968 9662 23969
rect 9346 23904 9352 23968
rect 9416 23904 9432 23968
rect 9496 23904 9512 23968
rect 9576 23904 9592 23968
rect 9656 23904 9662 23968
rect 9346 23903 9662 23904
rect 933 23490 999 23493
rect 0 23488 999 23490
rect 0 23432 938 23488
rect 994 23432 999 23488
rect 0 23430 999 23432
rect 933 23427 999 23430
rect 3606 23424 3922 23425
rect 3606 23360 3612 23424
rect 3676 23360 3692 23424
rect 3756 23360 3772 23424
rect 3836 23360 3852 23424
rect 3916 23360 3922 23424
rect 3606 23359 3922 23360
rect 5206 23424 5522 23425
rect 5206 23360 5212 23424
rect 5276 23360 5292 23424
rect 5356 23360 5372 23424
rect 5436 23360 5452 23424
rect 5516 23360 5522 23424
rect 5206 23359 5522 23360
rect 6806 23424 7122 23425
rect 6806 23360 6812 23424
rect 6876 23360 6892 23424
rect 6956 23360 6972 23424
rect 7036 23360 7052 23424
rect 7116 23360 7122 23424
rect 6806 23359 7122 23360
rect 8406 23424 8722 23425
rect 8406 23360 8412 23424
rect 8476 23360 8492 23424
rect 8556 23360 8572 23424
rect 8636 23360 8652 23424
rect 8716 23360 8722 23424
rect 8406 23359 8722 23360
rect 4337 22946 4403 22949
rect 4294 22944 4403 22946
rect 4294 22888 4342 22944
rect 4398 22888 4403 22944
rect 4294 22883 4403 22888
rect 2946 22880 3262 22881
rect 2946 22816 2952 22880
rect 3016 22816 3032 22880
rect 3096 22816 3112 22880
rect 3176 22816 3192 22880
rect 3256 22816 3262 22880
rect 2946 22815 3262 22816
rect 4294 22677 4354 22883
rect 4546 22880 4862 22881
rect 4546 22816 4552 22880
rect 4616 22816 4632 22880
rect 4696 22816 4712 22880
rect 4776 22816 4792 22880
rect 4856 22816 4862 22880
rect 4546 22815 4862 22816
rect 6146 22880 6462 22881
rect 6146 22816 6152 22880
rect 6216 22816 6232 22880
rect 6296 22816 6312 22880
rect 6376 22816 6392 22880
rect 6456 22816 6462 22880
rect 6146 22815 6462 22816
rect 7746 22880 8062 22881
rect 7746 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8062 22880
rect 7746 22815 8062 22816
rect 9346 22880 9662 22881
rect 9346 22816 9352 22880
rect 9416 22816 9432 22880
rect 9496 22816 9512 22880
rect 9576 22816 9592 22880
rect 9656 22816 9662 22880
rect 9346 22815 9662 22816
rect 4245 22672 4354 22677
rect 4245 22616 4250 22672
rect 4306 22616 4354 22672
rect 4245 22614 4354 22616
rect 4245 22611 4311 22614
rect 933 22538 999 22541
rect 0 22536 999 22538
rect 0 22480 938 22536
rect 994 22480 999 22536
rect 0 22478 999 22480
rect 933 22475 999 22478
rect 3606 22336 3922 22337
rect 3606 22272 3612 22336
rect 3676 22272 3692 22336
rect 3756 22272 3772 22336
rect 3836 22272 3852 22336
rect 3916 22272 3922 22336
rect 3606 22271 3922 22272
rect 5206 22336 5522 22337
rect 5206 22272 5212 22336
rect 5276 22272 5292 22336
rect 5356 22272 5372 22336
rect 5436 22272 5452 22336
rect 5516 22272 5522 22336
rect 5206 22271 5522 22272
rect 6806 22336 7122 22337
rect 6806 22272 6812 22336
rect 6876 22272 6892 22336
rect 6956 22272 6972 22336
rect 7036 22272 7052 22336
rect 7116 22272 7122 22336
rect 6806 22271 7122 22272
rect 8406 22336 8722 22337
rect 8406 22272 8412 22336
rect 8476 22272 8492 22336
rect 8556 22272 8572 22336
rect 8636 22272 8652 22336
rect 8716 22272 8722 22336
rect 8406 22271 8722 22272
rect 2946 21792 3262 21793
rect 2946 21728 2952 21792
rect 3016 21728 3032 21792
rect 3096 21728 3112 21792
rect 3176 21728 3192 21792
rect 3256 21728 3262 21792
rect 2946 21727 3262 21728
rect 4546 21792 4862 21793
rect 4546 21728 4552 21792
rect 4616 21728 4632 21792
rect 4696 21728 4712 21792
rect 4776 21728 4792 21792
rect 4856 21728 4862 21792
rect 4546 21727 4862 21728
rect 6146 21792 6462 21793
rect 6146 21728 6152 21792
rect 6216 21728 6232 21792
rect 6296 21728 6312 21792
rect 6376 21728 6392 21792
rect 6456 21728 6462 21792
rect 6146 21727 6462 21728
rect 7746 21792 8062 21793
rect 7746 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8062 21792
rect 7746 21727 8062 21728
rect 9346 21792 9662 21793
rect 9346 21728 9352 21792
rect 9416 21728 9432 21792
rect 9496 21728 9512 21792
rect 9576 21728 9592 21792
rect 9656 21728 9662 21792
rect 9346 21727 9662 21728
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 933 21523 999 21526
rect 3606 21248 3922 21249
rect 3606 21184 3612 21248
rect 3676 21184 3692 21248
rect 3756 21184 3772 21248
rect 3836 21184 3852 21248
rect 3916 21184 3922 21248
rect 3606 21183 3922 21184
rect 5206 21248 5522 21249
rect 5206 21184 5212 21248
rect 5276 21184 5292 21248
rect 5356 21184 5372 21248
rect 5436 21184 5452 21248
rect 5516 21184 5522 21248
rect 5206 21183 5522 21184
rect 6806 21248 7122 21249
rect 6806 21184 6812 21248
rect 6876 21184 6892 21248
rect 6956 21184 6972 21248
rect 7036 21184 7052 21248
rect 7116 21184 7122 21248
rect 6806 21183 7122 21184
rect 8406 21248 8722 21249
rect 8406 21184 8412 21248
rect 8476 21184 8492 21248
rect 8556 21184 8572 21248
rect 8636 21184 8652 21248
rect 8716 21184 8722 21248
rect 8406 21183 8722 21184
rect 2946 20704 3262 20705
rect 2946 20640 2952 20704
rect 3016 20640 3032 20704
rect 3096 20640 3112 20704
rect 3176 20640 3192 20704
rect 3256 20640 3262 20704
rect 2946 20639 3262 20640
rect 4546 20704 4862 20705
rect 4546 20640 4552 20704
rect 4616 20640 4632 20704
rect 4696 20640 4712 20704
rect 4776 20640 4792 20704
rect 4856 20640 4862 20704
rect 4546 20639 4862 20640
rect 6146 20704 6462 20705
rect 6146 20640 6152 20704
rect 6216 20640 6232 20704
rect 6296 20640 6312 20704
rect 6376 20640 6392 20704
rect 6456 20640 6462 20704
rect 6146 20639 6462 20640
rect 7746 20704 8062 20705
rect 7746 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8062 20704
rect 7746 20639 8062 20640
rect 9346 20704 9662 20705
rect 9346 20640 9352 20704
rect 9416 20640 9432 20704
rect 9496 20640 9512 20704
rect 9576 20640 9592 20704
rect 9656 20640 9662 20704
rect 108021 20660 108087 20663
rect 9346 20639 9662 20640
rect 107924 20658 108087 20660
rect 1393 20634 1459 20637
rect 0 20632 1459 20634
rect 0 20576 1398 20632
rect 1454 20576 1459 20632
rect 107924 20602 108026 20658
rect 108082 20602 108087 20658
rect 107924 20600 108087 20602
rect 108021 20597 108087 20600
rect 0 20574 1459 20576
rect 1393 20571 1459 20574
rect 3606 20160 3922 20161
rect 3606 20096 3612 20160
rect 3676 20096 3692 20160
rect 3756 20096 3772 20160
rect 3836 20096 3852 20160
rect 3916 20096 3922 20160
rect 3606 20095 3922 20096
rect 5206 20160 5522 20161
rect 5206 20096 5212 20160
rect 5276 20096 5292 20160
rect 5356 20096 5372 20160
rect 5436 20096 5452 20160
rect 5516 20096 5522 20160
rect 5206 20095 5522 20096
rect 6806 20160 7122 20161
rect 6806 20096 6812 20160
rect 6876 20096 6892 20160
rect 6956 20096 6972 20160
rect 7036 20096 7052 20160
rect 7116 20096 7122 20160
rect 6806 20095 7122 20096
rect 8406 20160 8722 20161
rect 8406 20096 8412 20160
rect 8476 20096 8492 20160
rect 8556 20096 8572 20160
rect 8636 20096 8652 20160
rect 8716 20096 8722 20160
rect 8406 20095 8722 20096
rect 933 19682 999 19685
rect 0 19680 999 19682
rect 0 19624 938 19680
rect 994 19624 999 19680
rect 0 19622 999 19624
rect 933 19619 999 19622
rect 2946 19616 3262 19617
rect 2946 19552 2952 19616
rect 3016 19552 3032 19616
rect 3096 19552 3112 19616
rect 3176 19552 3192 19616
rect 3256 19552 3262 19616
rect 2946 19551 3262 19552
rect 4546 19616 4862 19617
rect 4546 19552 4552 19616
rect 4616 19552 4632 19616
rect 4696 19552 4712 19616
rect 4776 19552 4792 19616
rect 4856 19552 4862 19616
rect 4546 19551 4862 19552
rect 6146 19616 6462 19617
rect 6146 19552 6152 19616
rect 6216 19552 6232 19616
rect 6296 19552 6312 19616
rect 6376 19552 6392 19616
rect 6456 19552 6462 19616
rect 6146 19551 6462 19552
rect 7746 19616 8062 19617
rect 7746 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8062 19616
rect 7746 19551 8062 19552
rect 9346 19616 9662 19617
rect 9346 19552 9352 19616
rect 9416 19552 9432 19616
rect 9496 19552 9512 19616
rect 9576 19552 9592 19616
rect 9656 19552 9662 19616
rect 9346 19551 9662 19552
rect 3606 19072 3922 19073
rect 3606 19008 3612 19072
rect 3676 19008 3692 19072
rect 3756 19008 3772 19072
rect 3836 19008 3852 19072
rect 3916 19008 3922 19072
rect 3606 19007 3922 19008
rect 5206 19072 5522 19073
rect 5206 19008 5212 19072
rect 5276 19008 5292 19072
rect 5356 19008 5372 19072
rect 5436 19008 5452 19072
rect 5516 19008 5522 19072
rect 5206 19007 5522 19008
rect 6806 19072 7122 19073
rect 6806 19008 6812 19072
rect 6876 19008 6892 19072
rect 6956 19008 6972 19072
rect 7036 19008 7052 19072
rect 7116 19008 7122 19072
rect 6806 19007 7122 19008
rect 8406 19072 8722 19073
rect 8406 19008 8412 19072
rect 8476 19008 8492 19072
rect 8556 19008 8572 19072
rect 8636 19008 8652 19072
rect 8716 19008 8722 19072
rect 8406 19007 8722 19008
rect 933 18730 999 18733
rect 0 18728 999 18730
rect 0 18672 938 18728
rect 994 18672 999 18728
rect 0 18670 999 18672
rect 933 18667 999 18670
rect 2946 18528 3262 18529
rect 2946 18464 2952 18528
rect 3016 18464 3032 18528
rect 3096 18464 3112 18528
rect 3176 18464 3192 18528
rect 3256 18464 3262 18528
rect 2946 18463 3262 18464
rect 4546 18528 4862 18529
rect 4546 18464 4552 18528
rect 4616 18464 4632 18528
rect 4696 18464 4712 18528
rect 4776 18464 4792 18528
rect 4856 18464 4862 18528
rect 4546 18463 4862 18464
rect 6146 18528 6462 18529
rect 6146 18464 6152 18528
rect 6216 18464 6232 18528
rect 6296 18464 6312 18528
rect 6376 18464 6392 18528
rect 6456 18464 6462 18528
rect 6146 18463 6462 18464
rect 7746 18528 8062 18529
rect 7746 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8062 18528
rect 7746 18463 8062 18464
rect 9346 18528 9662 18529
rect 9346 18464 9352 18528
rect 9416 18464 9432 18528
rect 9496 18464 9512 18528
rect 9576 18464 9592 18528
rect 9656 18464 9662 18528
rect 9346 18463 9662 18464
rect 107894 18461 107954 18998
rect 107894 18456 107995 18461
rect 107894 18400 107934 18456
rect 107990 18400 107995 18456
rect 107894 18398 107995 18400
rect 107929 18395 107995 18398
rect 3606 17984 3922 17985
rect 3606 17920 3612 17984
rect 3676 17920 3692 17984
rect 3756 17920 3772 17984
rect 3836 17920 3852 17984
rect 3916 17920 3922 17984
rect 3606 17919 3922 17920
rect 5206 17984 5522 17985
rect 5206 17920 5212 17984
rect 5276 17920 5292 17984
rect 5356 17920 5372 17984
rect 5436 17920 5452 17984
rect 5516 17920 5522 17984
rect 5206 17919 5522 17920
rect 6806 17984 7122 17985
rect 6806 17920 6812 17984
rect 6876 17920 6892 17984
rect 6956 17920 6972 17984
rect 7036 17920 7052 17984
rect 7116 17920 7122 17984
rect 6806 17919 7122 17920
rect 8406 17984 8722 17985
rect 8406 17920 8412 17984
rect 8476 17920 8492 17984
rect 8556 17920 8572 17984
rect 8636 17920 8652 17984
rect 8716 17920 8722 17984
rect 8406 17919 8722 17920
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 1577 17715 1643 17718
rect 108113 17668 108179 17671
rect 107924 17666 108179 17668
rect 107924 17610 108118 17666
rect 108174 17610 108179 17666
rect 107924 17608 108179 17610
rect 108113 17605 108179 17608
rect 2946 17440 3262 17441
rect 2946 17376 2952 17440
rect 3016 17376 3032 17440
rect 3096 17376 3112 17440
rect 3176 17376 3192 17440
rect 3256 17376 3262 17440
rect 2946 17375 3262 17376
rect 4546 17440 4862 17441
rect 4546 17376 4552 17440
rect 4616 17376 4632 17440
rect 4696 17376 4712 17440
rect 4776 17376 4792 17440
rect 4856 17376 4862 17440
rect 4546 17375 4862 17376
rect 6146 17440 6462 17441
rect 6146 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6392 17440
rect 6456 17376 6462 17440
rect 6146 17375 6462 17376
rect 7746 17440 8062 17441
rect 7746 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8062 17440
rect 7746 17375 8062 17376
rect 9346 17440 9662 17441
rect 9346 17376 9352 17440
rect 9416 17376 9432 17440
rect 9496 17376 9512 17440
rect 9576 17376 9592 17440
rect 9656 17376 9662 17440
rect 9346 17375 9662 17376
rect 3606 16896 3922 16897
rect 3606 16832 3612 16896
rect 3676 16832 3692 16896
rect 3756 16832 3772 16896
rect 3836 16832 3852 16896
rect 3916 16832 3922 16896
rect 3606 16831 3922 16832
rect 5206 16896 5522 16897
rect 5206 16832 5212 16896
rect 5276 16832 5292 16896
rect 5356 16832 5372 16896
rect 5436 16832 5452 16896
rect 5516 16832 5522 16896
rect 5206 16831 5522 16832
rect 6806 16896 7122 16897
rect 6806 16832 6812 16896
rect 6876 16832 6892 16896
rect 6956 16832 6972 16896
rect 7036 16832 7052 16896
rect 7116 16832 7122 16896
rect 6806 16831 7122 16832
rect 8406 16896 8722 16897
rect 8406 16832 8412 16896
rect 8476 16832 8492 16896
rect 8556 16832 8572 16896
rect 8636 16832 8652 16896
rect 8716 16832 8722 16896
rect 8406 16831 8722 16832
rect 933 16826 999 16829
rect 0 16824 999 16826
rect 0 16768 938 16824
rect 994 16768 999 16824
rect 0 16766 999 16768
rect 933 16763 999 16766
rect 2946 16352 3262 16353
rect 2946 16288 2952 16352
rect 3016 16288 3032 16352
rect 3096 16288 3112 16352
rect 3176 16288 3192 16352
rect 3256 16288 3262 16352
rect 2946 16287 3262 16288
rect 4546 16352 4862 16353
rect 4546 16288 4552 16352
rect 4616 16288 4632 16352
rect 4696 16288 4712 16352
rect 4776 16288 4792 16352
rect 4856 16288 4862 16352
rect 4546 16287 4862 16288
rect 6146 16352 6462 16353
rect 6146 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6392 16352
rect 6456 16288 6462 16352
rect 6146 16287 6462 16288
rect 7746 16352 8062 16353
rect 7746 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8062 16352
rect 7746 16287 8062 16288
rect 9346 16352 9662 16353
rect 9346 16288 9352 16352
rect 9416 16288 9432 16352
rect 9496 16288 9512 16352
rect 9576 16288 9592 16352
rect 9656 16288 9662 16352
rect 9346 16287 9662 16288
rect 933 15874 999 15877
rect 0 15872 999 15874
rect 0 15816 938 15872
rect 994 15816 999 15872
rect 0 15814 999 15816
rect 933 15811 999 15814
rect 3606 15808 3922 15809
rect 3606 15744 3612 15808
rect 3676 15744 3692 15808
rect 3756 15744 3772 15808
rect 3836 15744 3852 15808
rect 3916 15744 3922 15808
rect 3606 15743 3922 15744
rect 5206 15808 5522 15809
rect 5206 15744 5212 15808
rect 5276 15744 5292 15808
rect 5356 15744 5372 15808
rect 5436 15744 5452 15808
rect 5516 15744 5522 15808
rect 5206 15743 5522 15744
rect 6806 15808 7122 15809
rect 6806 15744 6812 15808
rect 6876 15744 6892 15808
rect 6956 15744 6972 15808
rect 7036 15744 7052 15808
rect 7116 15744 7122 15808
rect 6806 15743 7122 15744
rect 8406 15808 8722 15809
rect 8406 15744 8412 15808
rect 8476 15744 8492 15808
rect 8556 15744 8572 15808
rect 8636 15744 8652 15808
rect 8716 15744 8722 15808
rect 8406 15743 8722 15744
rect 2946 15264 3262 15265
rect 2946 15200 2952 15264
rect 3016 15200 3032 15264
rect 3096 15200 3112 15264
rect 3176 15200 3192 15264
rect 3256 15200 3262 15264
rect 2946 15199 3262 15200
rect 4546 15264 4862 15265
rect 4546 15200 4552 15264
rect 4616 15200 4632 15264
rect 4696 15200 4712 15264
rect 4776 15200 4792 15264
rect 4856 15200 4862 15264
rect 4546 15199 4862 15200
rect 6146 15264 6462 15265
rect 6146 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6392 15264
rect 6456 15200 6462 15264
rect 6146 15199 6462 15200
rect 7746 15264 8062 15265
rect 7746 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8062 15264
rect 7746 15199 8062 15200
rect 9346 15264 9662 15265
rect 9346 15200 9352 15264
rect 9416 15200 9432 15264
rect 9496 15200 9512 15264
rect 9576 15200 9592 15264
rect 9656 15200 9662 15264
rect 9346 15199 9662 15200
rect 933 14922 999 14925
rect 0 14920 999 14922
rect 0 14864 938 14920
rect 994 14864 999 14920
rect 0 14862 999 14864
rect 933 14859 999 14862
rect 3606 14720 3922 14721
rect 3606 14656 3612 14720
rect 3676 14656 3692 14720
rect 3756 14656 3772 14720
rect 3836 14656 3852 14720
rect 3916 14656 3922 14720
rect 3606 14655 3922 14656
rect 5206 14720 5522 14721
rect 5206 14656 5212 14720
rect 5276 14656 5292 14720
rect 5356 14656 5372 14720
rect 5436 14656 5452 14720
rect 5516 14656 5522 14720
rect 5206 14655 5522 14656
rect 6806 14720 7122 14721
rect 6806 14656 6812 14720
rect 6876 14656 6892 14720
rect 6956 14656 6972 14720
rect 7036 14656 7052 14720
rect 7116 14656 7122 14720
rect 6806 14655 7122 14656
rect 8406 14720 8722 14721
rect 8406 14656 8412 14720
rect 8476 14656 8492 14720
rect 8556 14656 8572 14720
rect 8636 14656 8652 14720
rect 8716 14656 8722 14720
rect 8406 14655 8722 14656
rect 2946 14176 3262 14177
rect 2946 14112 2952 14176
rect 3016 14112 3032 14176
rect 3096 14112 3112 14176
rect 3176 14112 3192 14176
rect 3256 14112 3262 14176
rect 2946 14111 3262 14112
rect 4546 14176 4862 14177
rect 4546 14112 4552 14176
rect 4616 14112 4632 14176
rect 4696 14112 4712 14176
rect 4776 14112 4792 14176
rect 4856 14112 4862 14176
rect 4546 14111 4862 14112
rect 6146 14176 6462 14177
rect 6146 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6392 14176
rect 6456 14112 6462 14176
rect 6146 14111 6462 14112
rect 7746 14176 8062 14177
rect 7746 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8062 14176
rect 7746 14111 8062 14112
rect 9346 14176 9662 14177
rect 9346 14112 9352 14176
rect 9416 14112 9432 14176
rect 9496 14112 9512 14176
rect 9576 14112 9592 14176
rect 9656 14112 9662 14176
rect 9346 14111 9662 14112
rect 933 13970 999 13973
rect 0 13968 999 13970
rect 0 13912 938 13968
rect 994 13912 999 13968
rect 0 13910 999 13912
rect 933 13907 999 13910
rect 3606 13632 3922 13633
rect 3606 13568 3612 13632
rect 3676 13568 3692 13632
rect 3756 13568 3772 13632
rect 3836 13568 3852 13632
rect 3916 13568 3922 13632
rect 3606 13567 3922 13568
rect 5206 13632 5522 13633
rect 5206 13568 5212 13632
rect 5276 13568 5292 13632
rect 5356 13568 5372 13632
rect 5436 13568 5452 13632
rect 5516 13568 5522 13632
rect 5206 13567 5522 13568
rect 6806 13632 7122 13633
rect 6806 13568 6812 13632
rect 6876 13568 6892 13632
rect 6956 13568 6972 13632
rect 7036 13568 7052 13632
rect 7116 13568 7122 13632
rect 6806 13567 7122 13568
rect 8406 13632 8722 13633
rect 8406 13568 8412 13632
rect 8476 13568 8492 13632
rect 8556 13568 8572 13632
rect 8636 13568 8652 13632
rect 8716 13568 8722 13632
rect 8406 13567 8722 13568
rect 2946 13088 3262 13089
rect 2946 13024 2952 13088
rect 3016 13024 3032 13088
rect 3096 13024 3112 13088
rect 3176 13024 3192 13088
rect 3256 13024 3262 13088
rect 2946 13023 3262 13024
rect 4546 13088 4862 13089
rect 4546 13024 4552 13088
rect 4616 13024 4632 13088
rect 4696 13024 4712 13088
rect 4776 13024 4792 13088
rect 4856 13024 4862 13088
rect 4546 13023 4862 13024
rect 6146 13088 6462 13089
rect 6146 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6392 13088
rect 6456 13024 6462 13088
rect 6146 13023 6462 13024
rect 7746 13088 8062 13089
rect 7746 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8062 13088
rect 7746 13023 8062 13024
rect 9346 13088 9662 13089
rect 9346 13024 9352 13088
rect 9416 13024 9432 13088
rect 9496 13024 9512 13088
rect 9576 13024 9592 13088
rect 9656 13024 9662 13088
rect 9346 13023 9662 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 933 12955 999 12958
rect 3606 12544 3922 12545
rect 3606 12480 3612 12544
rect 3676 12480 3692 12544
rect 3756 12480 3772 12544
rect 3836 12480 3852 12544
rect 3916 12480 3922 12544
rect 3606 12479 3922 12480
rect 5206 12544 5522 12545
rect 5206 12480 5212 12544
rect 5276 12480 5292 12544
rect 5356 12480 5372 12544
rect 5436 12480 5452 12544
rect 5516 12480 5522 12544
rect 5206 12479 5522 12480
rect 6806 12544 7122 12545
rect 6806 12480 6812 12544
rect 6876 12480 6892 12544
rect 6956 12480 6972 12544
rect 7036 12480 7052 12544
rect 7116 12480 7122 12544
rect 6806 12479 7122 12480
rect 8406 12544 8722 12545
rect 8406 12480 8412 12544
rect 8476 12480 8492 12544
rect 8556 12480 8572 12544
rect 8636 12480 8652 12544
rect 8716 12480 8722 12544
rect 8406 12479 8722 12480
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 933 12003 999 12006
rect 2946 12000 3262 12001
rect 2946 11936 2952 12000
rect 3016 11936 3032 12000
rect 3096 11936 3112 12000
rect 3176 11936 3192 12000
rect 3256 11936 3262 12000
rect 2946 11935 3262 11936
rect 4546 12000 4862 12001
rect 4546 11936 4552 12000
rect 4616 11936 4632 12000
rect 4696 11936 4712 12000
rect 4776 11936 4792 12000
rect 4856 11936 4862 12000
rect 4546 11935 4862 11936
rect 6146 12000 6462 12001
rect 6146 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6392 12000
rect 6456 11936 6462 12000
rect 6146 11935 6462 11936
rect 7746 12000 8062 12001
rect 7746 11936 7752 12000
rect 7816 11936 7832 12000
rect 7896 11936 7912 12000
rect 7976 11936 7992 12000
rect 8056 11936 8062 12000
rect 7746 11935 8062 11936
rect 9346 12000 9662 12001
rect 9346 11936 9352 12000
rect 9416 11936 9432 12000
rect 9496 11936 9512 12000
rect 9576 11936 9592 12000
rect 9656 11936 9662 12000
rect 9346 11935 9662 11936
rect 3606 11456 3922 11457
rect 3606 11392 3612 11456
rect 3676 11392 3692 11456
rect 3756 11392 3772 11456
rect 3836 11392 3852 11456
rect 3916 11392 3922 11456
rect 3606 11391 3922 11392
rect 5206 11456 5522 11457
rect 5206 11392 5212 11456
rect 5276 11392 5292 11456
rect 5356 11392 5372 11456
rect 5436 11392 5452 11456
rect 5516 11392 5522 11456
rect 5206 11391 5522 11392
rect 6806 11456 7122 11457
rect 6806 11392 6812 11456
rect 6876 11392 6892 11456
rect 6956 11392 6972 11456
rect 7036 11392 7052 11456
rect 7116 11392 7122 11456
rect 6806 11391 7122 11392
rect 8406 11456 8722 11457
rect 8406 11392 8412 11456
rect 8476 11392 8492 11456
rect 8556 11392 8572 11456
rect 8636 11392 8652 11456
rect 8716 11392 8722 11456
rect 8406 11391 8722 11392
rect 9581 11250 9647 11253
rect 11329 11250 11395 11253
rect 11470 11250 12052 11276
rect 9581 11248 12052 11250
rect 9581 11192 9586 11248
rect 9642 11192 11334 11248
rect 11390 11216 12052 11248
rect 11390 11192 11530 11216
rect 9581 11190 11530 11192
rect 9581 11187 9647 11190
rect 11329 11187 11395 11190
rect 933 11114 999 11117
rect 0 11112 999 11114
rect 0 11056 938 11112
rect 994 11056 999 11112
rect 0 11054 999 11056
rect 933 11051 999 11054
rect 2946 10912 3262 10913
rect 2946 10848 2952 10912
rect 3016 10848 3032 10912
rect 3096 10848 3112 10912
rect 3176 10848 3192 10912
rect 3256 10848 3262 10912
rect 2946 10847 3262 10848
rect 4546 10912 4862 10913
rect 4546 10848 4552 10912
rect 4616 10848 4632 10912
rect 4696 10848 4712 10912
rect 4776 10848 4792 10912
rect 4856 10848 4862 10912
rect 4546 10847 4862 10848
rect 6146 10912 6462 10913
rect 6146 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6392 10912
rect 6456 10848 6462 10912
rect 6146 10847 6462 10848
rect 7746 10912 8062 10913
rect 7746 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8062 10912
rect 7746 10847 8062 10848
rect 9346 10912 9662 10913
rect 9346 10848 9352 10912
rect 9416 10848 9432 10912
rect 9496 10848 9512 10912
rect 9576 10848 9592 10912
rect 9656 10848 9662 10912
rect 9346 10847 9662 10848
rect 3606 10368 3922 10369
rect 3606 10304 3612 10368
rect 3676 10304 3692 10368
rect 3756 10304 3772 10368
rect 3836 10304 3852 10368
rect 3916 10304 3922 10368
rect 3606 10303 3922 10304
rect 5206 10368 5522 10369
rect 5206 10304 5212 10368
rect 5276 10304 5292 10368
rect 5356 10304 5372 10368
rect 5436 10304 5452 10368
rect 5516 10304 5522 10368
rect 5206 10303 5522 10304
rect 6806 10368 7122 10369
rect 6806 10304 6812 10368
rect 6876 10304 6892 10368
rect 6956 10304 6972 10368
rect 7036 10304 7052 10368
rect 7116 10304 7122 10368
rect 6806 10303 7122 10304
rect 8406 10368 8722 10369
rect 8406 10304 8412 10368
rect 8476 10304 8492 10368
rect 8556 10304 8572 10368
rect 8636 10304 8652 10368
rect 8716 10304 8722 10368
rect 8406 10303 8722 10304
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 933 10099 999 10102
rect 2946 9824 3262 9825
rect 2946 9760 2952 9824
rect 3016 9760 3032 9824
rect 3096 9760 3112 9824
rect 3176 9760 3192 9824
rect 3256 9760 3262 9824
rect 2946 9759 3262 9760
rect 4546 9824 4862 9825
rect 4546 9760 4552 9824
rect 4616 9760 4632 9824
rect 4696 9760 4712 9824
rect 4776 9760 4792 9824
rect 4856 9760 4862 9824
rect 4546 9759 4862 9760
rect 6146 9824 6462 9825
rect 6146 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6392 9824
rect 6456 9760 6462 9824
rect 6146 9759 6462 9760
rect 7746 9824 8062 9825
rect 7746 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8062 9824
rect 7746 9759 8062 9760
rect 9346 9824 9662 9825
rect 9346 9760 9352 9824
rect 9416 9760 9432 9824
rect 9496 9760 9512 9824
rect 9576 9760 9592 9824
rect 9656 9760 9662 9824
rect 9346 9759 9662 9760
rect 11329 9618 11395 9621
rect 11470 9618 12052 9644
rect 11329 9616 12052 9618
rect 11329 9560 11334 9616
rect 11390 9584 12052 9616
rect 11390 9560 11530 9584
rect 11329 9558 11530 9560
rect 11329 9555 11395 9558
rect 3606 9280 3922 9281
rect 3606 9216 3612 9280
rect 3676 9216 3692 9280
rect 3756 9216 3772 9280
rect 3836 9216 3852 9280
rect 3916 9216 3922 9280
rect 3606 9215 3922 9216
rect 5206 9280 5522 9281
rect 5206 9216 5212 9280
rect 5276 9216 5292 9280
rect 5356 9216 5372 9280
rect 5436 9216 5452 9280
rect 5516 9216 5522 9280
rect 5206 9215 5522 9216
rect 6806 9280 7122 9281
rect 6806 9216 6812 9280
rect 6876 9216 6892 9280
rect 6956 9216 6972 9280
rect 7036 9216 7052 9280
rect 7116 9216 7122 9280
rect 6806 9215 7122 9216
rect 8406 9280 8722 9281
rect 8406 9216 8412 9280
rect 8476 9216 8492 9280
rect 8556 9216 8572 9280
rect 8636 9216 8652 9280
rect 8716 9216 8722 9280
rect 8406 9215 8722 9216
rect 933 9210 999 9213
rect 0 9208 999 9210
rect 0 9152 938 9208
rect 994 9152 999 9208
rect 0 9150 999 9152
rect 933 9147 999 9150
rect 2946 8736 3262 8737
rect 2946 8672 2952 8736
rect 3016 8672 3032 8736
rect 3096 8672 3112 8736
rect 3176 8672 3192 8736
rect 3256 8672 3262 8736
rect 2946 8671 3262 8672
rect 4546 8736 4862 8737
rect 4546 8672 4552 8736
rect 4616 8672 4632 8736
rect 4696 8672 4712 8736
rect 4776 8672 4792 8736
rect 4856 8672 4862 8736
rect 4546 8671 4862 8672
rect 6146 8736 6462 8737
rect 6146 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6392 8736
rect 6456 8672 6462 8736
rect 6146 8671 6462 8672
rect 7746 8736 8062 8737
rect 7746 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8062 8736
rect 7746 8671 8062 8672
rect 9346 8736 9662 8737
rect 9346 8672 9352 8736
rect 9416 8672 9432 8736
rect 9496 8672 9512 8736
rect 9576 8672 9592 8736
rect 9656 8672 9662 8736
rect 9346 8671 9662 8672
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 1393 8195 1459 8198
rect 3606 8192 3922 8193
rect 3606 8128 3612 8192
rect 3676 8128 3692 8192
rect 3756 8128 3772 8192
rect 3836 8128 3852 8192
rect 3916 8128 3922 8192
rect 3606 8127 3922 8128
rect 5206 8192 5522 8193
rect 5206 8128 5212 8192
rect 5276 8128 5292 8192
rect 5356 8128 5372 8192
rect 5436 8128 5452 8192
rect 5516 8128 5522 8192
rect 5206 8127 5522 8128
rect 6806 8192 7122 8193
rect 6806 8128 6812 8192
rect 6876 8128 6892 8192
rect 6956 8128 6972 8192
rect 7036 8128 7052 8192
rect 7116 8128 7122 8192
rect 6806 8127 7122 8128
rect 8406 8192 8722 8193
rect 8406 8128 8412 8192
rect 8476 8128 8492 8192
rect 8556 8128 8572 8192
rect 8636 8128 8652 8192
rect 8716 8128 8722 8192
rect 8406 8127 8722 8128
rect 2946 7648 3262 7649
rect 2946 7584 2952 7648
rect 3016 7584 3032 7648
rect 3096 7584 3112 7648
rect 3176 7584 3192 7648
rect 3256 7584 3262 7648
rect 2946 7583 3262 7584
rect 4546 7648 4862 7649
rect 4546 7584 4552 7648
rect 4616 7584 4632 7648
rect 4696 7584 4712 7648
rect 4776 7584 4792 7648
rect 4856 7584 4862 7648
rect 4546 7583 4862 7584
rect 6146 7648 6462 7649
rect 6146 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6392 7648
rect 6456 7584 6462 7648
rect 6146 7583 6462 7584
rect 7746 7648 8062 7649
rect 7746 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8062 7648
rect 7746 7583 8062 7584
rect 9346 7648 9662 7649
rect 9346 7584 9352 7648
rect 9416 7584 9432 7648
rect 9496 7584 9512 7648
rect 9576 7584 9592 7648
rect 9656 7584 9662 7648
rect 9346 7583 9662 7584
rect 933 7306 999 7309
rect 0 7304 999 7306
rect 0 7248 938 7304
rect 994 7248 999 7304
rect 0 7246 999 7248
rect 933 7243 999 7246
rect 3606 7104 3922 7105
rect 3606 7040 3612 7104
rect 3676 7040 3692 7104
rect 3756 7040 3772 7104
rect 3836 7040 3852 7104
rect 3916 7040 3922 7104
rect 3606 7039 3922 7040
rect 5206 7104 5522 7105
rect 5206 7040 5212 7104
rect 5276 7040 5292 7104
rect 5356 7040 5372 7104
rect 5436 7040 5452 7104
rect 5516 7040 5522 7104
rect 5206 7039 5522 7040
rect 6806 7104 7122 7105
rect 6806 7040 6812 7104
rect 6876 7040 6892 7104
rect 6956 7040 6972 7104
rect 7036 7040 7052 7104
rect 7116 7040 7122 7104
rect 6806 7039 7122 7040
rect 8406 7104 8722 7105
rect 8406 7040 8412 7104
rect 8476 7040 8492 7104
rect 8556 7040 8572 7104
rect 8636 7040 8652 7104
rect 8716 7040 8722 7104
rect 8406 7039 8722 7040
rect 2946 6560 3262 6561
rect 2946 6496 2952 6560
rect 3016 6496 3032 6560
rect 3096 6496 3112 6560
rect 3176 6496 3192 6560
rect 3256 6496 3262 6560
rect 2946 6495 3262 6496
rect 4546 6560 4862 6561
rect 4546 6496 4552 6560
rect 4616 6496 4632 6560
rect 4696 6496 4712 6560
rect 4776 6496 4792 6560
rect 4856 6496 4862 6560
rect 4546 6495 4862 6496
rect 6146 6560 6462 6561
rect 6146 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6392 6560
rect 6456 6496 6462 6560
rect 6146 6495 6462 6496
rect 7746 6560 8062 6561
rect 7746 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8062 6560
rect 7746 6495 8062 6496
rect 9346 6560 9662 6561
rect 9346 6496 9352 6560
rect 9416 6496 9432 6560
rect 9496 6496 9512 6560
rect 9576 6496 9592 6560
rect 9656 6496 9662 6560
rect 9346 6495 9662 6496
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 933 6291 999 6294
rect 3606 6016 3922 6017
rect 3606 5952 3612 6016
rect 3676 5952 3692 6016
rect 3756 5952 3772 6016
rect 3836 5952 3852 6016
rect 3916 5952 3922 6016
rect 3606 5951 3922 5952
rect 5206 6016 5522 6017
rect 5206 5952 5212 6016
rect 5276 5952 5292 6016
rect 5356 5952 5372 6016
rect 5436 5952 5452 6016
rect 5516 5952 5522 6016
rect 5206 5951 5522 5952
rect 6806 6016 7122 6017
rect 6806 5952 6812 6016
rect 6876 5952 6892 6016
rect 6956 5952 6972 6016
rect 7036 5952 7052 6016
rect 7116 5952 7122 6016
rect 6806 5951 7122 5952
rect 8406 6016 8722 6017
rect 8406 5952 8412 6016
rect 8476 5952 8492 6016
rect 8556 5952 8572 6016
rect 8636 5952 8652 6016
rect 8716 5952 8722 6016
rect 8406 5951 8722 5952
rect 1577 5538 1643 5541
rect 798 5536 1643 5538
rect 798 5480 1582 5536
rect 1638 5480 1643 5536
rect 798 5478 1643 5480
rect 798 5402 858 5478
rect 1577 5475 1643 5478
rect 2946 5472 3262 5473
rect 2946 5408 2952 5472
rect 3016 5408 3032 5472
rect 3096 5408 3112 5472
rect 3176 5408 3192 5472
rect 3256 5408 3262 5472
rect 2946 5407 3262 5408
rect 4546 5472 4862 5473
rect 4546 5408 4552 5472
rect 4616 5408 4632 5472
rect 4696 5408 4712 5472
rect 4776 5408 4792 5472
rect 4856 5408 4862 5472
rect 4546 5407 4862 5408
rect 6146 5472 6462 5473
rect 6146 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6392 5472
rect 6456 5408 6462 5472
rect 6146 5407 6462 5408
rect 7746 5472 8062 5473
rect 7746 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8062 5472
rect 7746 5407 8062 5408
rect 9346 5472 9662 5473
rect 9346 5408 9352 5472
rect 9416 5408 9432 5472
rect 9496 5408 9512 5472
rect 9576 5408 9592 5472
rect 9656 5408 9662 5472
rect 9346 5407 9662 5408
rect 0 5342 858 5402
rect 3606 4928 3922 4929
rect 3606 4864 3612 4928
rect 3676 4864 3692 4928
rect 3756 4864 3772 4928
rect 3836 4864 3852 4928
rect 3916 4864 3922 4928
rect 3606 4863 3922 4864
rect 5206 4928 5522 4929
rect 5206 4864 5212 4928
rect 5276 4864 5292 4928
rect 5356 4864 5372 4928
rect 5436 4864 5452 4928
rect 5516 4864 5522 4928
rect 5206 4863 5522 4864
rect 6806 4928 7122 4929
rect 6806 4864 6812 4928
rect 6876 4864 6892 4928
rect 6956 4864 6972 4928
rect 7036 4864 7052 4928
rect 7116 4864 7122 4928
rect 6806 4863 7122 4864
rect 8406 4928 8722 4929
rect 8406 4864 8412 4928
rect 8476 4864 8492 4928
rect 8556 4864 8572 4928
rect 8636 4864 8652 4928
rect 8716 4864 8722 4928
rect 8406 4863 8722 4864
rect 933 4450 999 4453
rect 0 4448 999 4450
rect 0 4392 938 4448
rect 994 4392 999 4448
rect 0 4390 999 4392
rect 933 4387 999 4390
rect 2946 4384 3262 4385
rect 2946 4320 2952 4384
rect 3016 4320 3032 4384
rect 3096 4320 3112 4384
rect 3176 4320 3192 4384
rect 3256 4320 3262 4384
rect 2946 4319 3262 4320
rect 4546 4384 4862 4385
rect 4546 4320 4552 4384
rect 4616 4320 4632 4384
rect 4696 4320 4712 4384
rect 4776 4320 4792 4384
rect 4856 4320 4862 4384
rect 4546 4319 4862 4320
rect 6146 4384 6462 4385
rect 6146 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6392 4384
rect 6456 4320 6462 4384
rect 6146 4319 6462 4320
rect 7746 4384 8062 4385
rect 7746 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8062 4384
rect 7746 4319 8062 4320
rect 9346 4384 9662 4385
rect 9346 4320 9352 4384
rect 9416 4320 9432 4384
rect 9496 4320 9512 4384
rect 9576 4320 9592 4384
rect 9656 4320 9662 4384
rect 9346 4319 9662 4320
rect 17861 3908 17927 3909
rect 39205 3908 39271 3909
rect 40309 3908 40375 3909
rect 17848 3844 17854 3908
rect 17918 3906 17927 3908
rect 39200 3906 39206 3908
rect 17918 3904 18010 3906
rect 17922 3848 18010 3904
rect 17918 3846 18010 3848
rect 39118 3846 39206 3906
rect 17918 3844 17927 3846
rect 39200 3844 39206 3846
rect 39270 3844 39276 3908
rect 40288 3844 40294 3908
rect 40358 3906 40375 3908
rect 45001 3908 45067 3909
rect 46105 3908 46171 3909
rect 50889 3908 50955 3909
rect 54385 3908 54451 3909
rect 45001 3906 45054 3908
rect 40358 3904 40450 3906
rect 40370 3848 40450 3904
rect 40358 3846 40450 3848
rect 44962 3904 45054 3906
rect 44962 3848 45006 3904
rect 44962 3846 45054 3848
rect 40358 3844 40375 3846
rect 17861 3843 17927 3844
rect 39205 3843 39271 3844
rect 40309 3843 40375 3844
rect 45001 3844 45054 3846
rect 45118 3844 45124 3908
rect 46105 3906 46142 3908
rect 46050 3904 46142 3906
rect 46050 3848 46110 3904
rect 46050 3846 46142 3848
rect 46105 3844 46142 3846
rect 46206 3844 46212 3908
rect 50889 3906 50902 3908
rect 50810 3904 50902 3906
rect 50810 3848 50894 3904
rect 50810 3846 50902 3848
rect 50889 3844 50902 3846
rect 50966 3844 50972 3908
rect 54385 3906 54438 3908
rect 54346 3904 54438 3906
rect 54346 3848 54390 3904
rect 54346 3846 54438 3848
rect 54385 3844 54438 3846
rect 54502 3844 54508 3908
rect 93894 3844 93900 3908
rect 93964 3906 93970 3908
rect 94960 3906 94966 3908
rect 93964 3846 94966 3906
rect 93964 3844 93970 3846
rect 94960 3844 94966 3846
rect 95030 3844 95036 3908
rect 45001 3843 45067 3844
rect 46105 3843 46171 3844
rect 50889 3843 50955 3844
rect 54385 3843 54451 3844
rect 3606 3840 3922 3841
rect 3606 3776 3612 3840
rect 3676 3776 3692 3840
rect 3756 3776 3772 3840
rect 3836 3776 3852 3840
rect 3916 3776 3922 3840
rect 3606 3775 3922 3776
rect 5206 3840 5522 3841
rect 5206 3776 5212 3840
rect 5276 3776 5292 3840
rect 5356 3776 5372 3840
rect 5436 3776 5452 3840
rect 5516 3776 5522 3840
rect 5206 3775 5522 3776
rect 6806 3840 7122 3841
rect 6806 3776 6812 3840
rect 6876 3776 6892 3840
rect 6956 3776 6972 3840
rect 7036 3776 7052 3840
rect 7116 3776 7122 3840
rect 6806 3775 7122 3776
rect 8406 3840 8722 3841
rect 8406 3776 8412 3840
rect 8476 3776 8492 3840
rect 8556 3776 8572 3840
rect 8636 3776 8652 3840
rect 8716 3776 8722 3840
rect 8406 3775 8722 3776
rect 28717 3772 28783 3773
rect 29821 3772 29887 3773
rect 47485 3772 47551 3773
rect 28717 3770 28734 3772
rect 28642 3768 28734 3770
rect 28642 3712 28722 3768
rect 28642 3710 28734 3712
rect 28717 3708 28734 3710
rect 28798 3708 28804 3772
rect 29816 3770 29822 3772
rect 29734 3710 29822 3770
rect 29816 3708 29822 3710
rect 29886 3708 29892 3772
rect 47485 3770 47502 3772
rect 47410 3768 47502 3770
rect 47410 3712 47490 3768
rect 47410 3710 47502 3712
rect 47485 3708 47502 3710
rect 47566 3708 47572 3772
rect 28717 3707 28783 3708
rect 29821 3707 29887 3708
rect 47485 3707 47551 3708
rect 5901 3634 5967 3637
rect 108113 3634 108179 3637
rect 5901 3632 108179 3634
rect 5901 3576 5906 3632
rect 5962 3576 108118 3632
rect 108174 3576 108179 3632
rect 5901 3574 108179 3576
rect 5901 3571 5967 3574
rect 108113 3571 108179 3574
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 933 3435 999 3438
rect 5717 3498 5783 3501
rect 108021 3498 108087 3501
rect 5717 3496 108087 3498
rect 5717 3440 5722 3496
rect 5778 3440 108026 3496
rect 108082 3440 108087 3496
rect 5717 3438 108087 3440
rect 5717 3435 5783 3438
rect 108021 3435 108087 3438
rect 10685 3362 10751 3365
rect 29637 3362 29703 3365
rect 10685 3360 29703 3362
rect 10685 3304 10690 3360
rect 10746 3304 29642 3360
rect 29698 3304 29703 3360
rect 10685 3302 29703 3304
rect 10685 3299 10751 3302
rect 29637 3299 29703 3302
rect 2946 3296 3262 3297
rect 2946 3232 2952 3296
rect 3016 3232 3032 3296
rect 3096 3232 3112 3296
rect 3176 3232 3192 3296
rect 3256 3232 3262 3296
rect 2946 3231 3262 3232
rect 4546 3296 4862 3297
rect 4546 3232 4552 3296
rect 4616 3232 4632 3296
rect 4696 3232 4712 3296
rect 4776 3232 4792 3296
rect 4856 3232 4862 3296
rect 4546 3231 4862 3232
rect 6146 3296 6462 3297
rect 6146 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6392 3296
rect 6456 3232 6462 3296
rect 6146 3231 6462 3232
rect 7746 3296 8062 3297
rect 7746 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8062 3296
rect 7746 3231 8062 3232
rect 9346 3296 9662 3297
rect 9346 3232 9352 3296
rect 9416 3232 9432 3296
rect 9496 3232 9512 3296
rect 9576 3232 9592 3296
rect 9656 3232 9662 3296
rect 9346 3231 9662 3232
rect 3606 2752 3922 2753
rect 3606 2688 3612 2752
rect 3676 2688 3692 2752
rect 3756 2688 3772 2752
rect 3836 2688 3852 2752
rect 3916 2688 3922 2752
rect 3606 2687 3922 2688
rect 5206 2752 5522 2753
rect 5206 2688 5212 2752
rect 5276 2688 5292 2752
rect 5356 2688 5372 2752
rect 5436 2688 5452 2752
rect 5516 2688 5522 2752
rect 5206 2687 5522 2688
rect 6806 2752 7122 2753
rect 6806 2688 6812 2752
rect 6876 2688 6892 2752
rect 6956 2688 6972 2752
rect 7036 2688 7052 2752
rect 7116 2688 7122 2752
rect 6806 2687 7122 2688
rect 8406 2752 8722 2753
rect 8406 2688 8412 2752
rect 8476 2688 8492 2752
rect 8556 2688 8572 2752
rect 8636 2688 8652 2752
rect 8716 2688 8722 2752
rect 8406 2687 8722 2688
rect 36997 2684 37063 2685
rect 49693 2684 49759 2685
rect 55397 2684 55463 2685
rect 57973 2684 58039 2685
rect 11830 2620 11836 2684
rect 11900 2682 11906 2684
rect 35566 2682 35572 2684
rect 11900 2622 35572 2682
rect 11900 2620 11906 2622
rect 35566 2620 35572 2622
rect 35636 2620 35642 2684
rect 36997 2682 37044 2684
rect 36952 2680 37044 2682
rect 36952 2624 37002 2680
rect 36952 2622 37044 2624
rect 36997 2620 37044 2622
rect 37108 2620 37114 2684
rect 49693 2682 49740 2684
rect 49648 2680 49740 2682
rect 49648 2624 49698 2680
rect 49648 2622 49740 2624
rect 49693 2620 49740 2622
rect 49804 2620 49810 2684
rect 55397 2682 55444 2684
rect 55352 2680 55444 2682
rect 55352 2624 55402 2680
rect 55352 2622 55444 2624
rect 55397 2620 55444 2622
rect 55508 2620 55514 2684
rect 57973 2682 58020 2684
rect 57928 2680 58020 2682
rect 57928 2624 57978 2680
rect 57928 2622 58020 2624
rect 57973 2620 58020 2622
rect 58084 2620 58090 2684
rect 36997 2619 37063 2620
rect 49693 2619 49759 2620
rect 55397 2619 55463 2620
rect 57973 2619 58039 2620
rect 1209 2546 1275 2549
rect 94957 2548 95023 2549
rect 94814 2546 94820 2548
rect 1209 2544 94820 2546
rect 1209 2488 1214 2544
rect 1270 2488 94820 2544
rect 1209 2486 94820 2488
rect 1209 2483 1275 2486
rect 94814 2484 94820 2486
rect 94884 2484 94890 2548
rect 94957 2544 95004 2548
rect 95068 2546 95074 2548
rect 94957 2488 94962 2544
rect 94957 2484 95004 2488
rect 95068 2486 95114 2546
rect 95068 2484 95074 2486
rect 94957 2483 95023 2484
rect 32029 2412 32095 2413
rect 42793 2412 42859 2413
rect 32029 2410 32076 2412
rect 31984 2408 32076 2410
rect 31984 2352 32034 2408
rect 31984 2350 32076 2352
rect 32029 2348 32076 2350
rect 32140 2348 32146 2412
rect 42742 2348 42748 2412
rect 42812 2410 42859 2412
rect 43805 2412 43871 2413
rect 48589 2412 48655 2413
rect 43805 2410 43852 2412
rect 42812 2408 42904 2410
rect 42854 2352 42904 2408
rect 42812 2350 42904 2352
rect 43760 2408 43852 2410
rect 43760 2352 43810 2408
rect 43760 2350 43852 2352
rect 42812 2348 42859 2350
rect 32029 2347 32095 2348
rect 42793 2347 42859 2348
rect 43805 2348 43852 2350
rect 43916 2348 43922 2412
rect 48589 2410 48636 2412
rect 48544 2408 48636 2410
rect 48544 2352 48594 2408
rect 48544 2350 48636 2352
rect 48589 2348 48636 2350
rect 48700 2348 48706 2412
rect 43805 2347 43871 2348
rect 48589 2347 48655 2348
rect 2946 2208 3262 2209
rect 2946 2144 2952 2208
rect 3016 2144 3032 2208
rect 3096 2144 3112 2208
rect 3176 2144 3192 2208
rect 3256 2144 3262 2208
rect 2946 2143 3262 2144
rect 4546 2208 4862 2209
rect 4546 2144 4552 2208
rect 4616 2144 4632 2208
rect 4696 2144 4712 2208
rect 4776 2144 4792 2208
rect 4856 2144 4862 2208
rect 4546 2143 4862 2144
rect 6146 2208 6462 2209
rect 6146 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6392 2208
rect 6456 2144 6462 2208
rect 6146 2143 6462 2144
rect 7746 2208 8062 2209
rect 7746 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8062 2208
rect 7746 2143 8062 2144
rect 9346 2208 9662 2209
rect 9346 2144 9352 2208
rect 9416 2144 9432 2208
rect 9496 2144 9512 2208
rect 9576 2144 9592 2208
rect 9656 2144 9662 2208
rect 9346 2143 9662 2144
rect 11646 2076 11652 2140
rect 11716 2138 11722 2140
rect 37457 2138 37523 2141
rect 11716 2136 37523 2138
rect 11716 2080 37462 2136
rect 37518 2080 37523 2136
rect 11716 2078 37523 2080
rect 11716 2076 11722 2078
rect 37457 2075 37523 2078
rect 1669 2002 1735 2005
rect 94630 2002 94636 2004
rect 1669 2000 94636 2002
rect 1669 1944 1674 2000
rect 1730 1944 94636 2000
rect 1669 1942 94636 1944
rect 1669 1939 1735 1942
rect 94630 1940 94636 1942
rect 94700 1940 94706 2004
rect 3606 1664 3922 1665
rect 3606 1600 3612 1664
rect 3676 1600 3692 1664
rect 3756 1600 3772 1664
rect 3836 1600 3852 1664
rect 3916 1600 3922 1664
rect 3606 1599 3922 1600
rect 5206 1664 5522 1665
rect 5206 1600 5212 1664
rect 5276 1600 5292 1664
rect 5356 1600 5372 1664
rect 5436 1600 5452 1664
rect 5516 1600 5522 1664
rect 5206 1599 5522 1600
rect 6806 1664 7122 1665
rect 6806 1600 6812 1664
rect 6876 1600 6892 1664
rect 6956 1600 6972 1664
rect 7036 1600 7052 1664
rect 7116 1600 7122 1664
rect 6806 1599 7122 1600
rect 8406 1664 8722 1665
rect 8406 1600 8412 1664
rect 8476 1600 8492 1664
rect 8556 1600 8572 1664
rect 8636 1600 8652 1664
rect 8716 1600 8722 1664
rect 8406 1599 8722 1600
rect 10006 1664 10322 1665
rect 10006 1600 10012 1664
rect 10076 1600 10092 1664
rect 10156 1600 10172 1664
rect 10236 1600 10252 1664
rect 10316 1600 10322 1664
rect 10006 1599 10322 1600
rect 11606 1664 11922 1665
rect 11606 1600 11612 1664
rect 11676 1600 11692 1664
rect 11756 1600 11772 1664
rect 11836 1600 11852 1664
rect 11916 1600 11922 1664
rect 11606 1599 11922 1600
rect 13206 1664 13522 1665
rect 13206 1600 13212 1664
rect 13276 1600 13292 1664
rect 13356 1600 13372 1664
rect 13436 1600 13452 1664
rect 13516 1600 13522 1664
rect 13206 1599 13522 1600
rect 14806 1664 15122 1665
rect 14806 1600 14812 1664
rect 14876 1600 14892 1664
rect 14956 1600 14972 1664
rect 15036 1600 15052 1664
rect 15116 1600 15122 1664
rect 14806 1599 15122 1600
rect 16406 1664 16722 1665
rect 16406 1600 16412 1664
rect 16476 1600 16492 1664
rect 16556 1600 16572 1664
rect 16636 1600 16652 1664
rect 16716 1600 16722 1664
rect 16406 1599 16722 1600
rect 18006 1664 18322 1665
rect 18006 1600 18012 1664
rect 18076 1600 18092 1664
rect 18156 1600 18172 1664
rect 18236 1600 18252 1664
rect 18316 1600 18322 1664
rect 18006 1599 18322 1600
rect 19606 1664 19922 1665
rect 19606 1600 19612 1664
rect 19676 1600 19692 1664
rect 19756 1600 19772 1664
rect 19836 1600 19852 1664
rect 19916 1600 19922 1664
rect 19606 1599 19922 1600
rect 21206 1664 21522 1665
rect 21206 1600 21212 1664
rect 21276 1600 21292 1664
rect 21356 1600 21372 1664
rect 21436 1600 21452 1664
rect 21516 1600 21522 1664
rect 21206 1599 21522 1600
rect 22806 1664 23122 1665
rect 22806 1600 22812 1664
rect 22876 1600 22892 1664
rect 22956 1600 22972 1664
rect 23036 1600 23052 1664
rect 23116 1600 23122 1664
rect 22806 1599 23122 1600
rect 24406 1664 24722 1665
rect 24406 1600 24412 1664
rect 24476 1600 24492 1664
rect 24556 1600 24572 1664
rect 24636 1600 24652 1664
rect 24716 1600 24722 1664
rect 24406 1599 24722 1600
rect 26006 1664 26322 1665
rect 26006 1600 26012 1664
rect 26076 1600 26092 1664
rect 26156 1600 26172 1664
rect 26236 1600 26252 1664
rect 26316 1600 26322 1664
rect 26006 1599 26322 1600
rect 27606 1664 27922 1665
rect 27606 1600 27612 1664
rect 27676 1600 27692 1664
rect 27756 1600 27772 1664
rect 27836 1600 27852 1664
rect 27916 1600 27922 1664
rect 27606 1599 27922 1600
rect 29206 1664 29522 1665
rect 29206 1600 29212 1664
rect 29276 1600 29292 1664
rect 29356 1600 29372 1664
rect 29436 1600 29452 1664
rect 29516 1600 29522 1664
rect 29206 1599 29522 1600
rect 30806 1664 31122 1665
rect 30806 1600 30812 1664
rect 30876 1600 30892 1664
rect 30956 1600 30972 1664
rect 31036 1600 31052 1664
rect 31116 1600 31122 1664
rect 30806 1599 31122 1600
rect 32406 1664 32722 1665
rect 32406 1600 32412 1664
rect 32476 1600 32492 1664
rect 32556 1600 32572 1664
rect 32636 1600 32652 1664
rect 32716 1600 32722 1664
rect 32406 1599 32722 1600
rect 34006 1664 34322 1665
rect 34006 1600 34012 1664
rect 34076 1600 34092 1664
rect 34156 1600 34172 1664
rect 34236 1600 34252 1664
rect 34316 1600 34322 1664
rect 34006 1599 34322 1600
rect 35606 1664 35922 1665
rect 35606 1600 35612 1664
rect 35676 1600 35692 1664
rect 35756 1600 35772 1664
rect 35836 1600 35852 1664
rect 35916 1600 35922 1664
rect 35606 1599 35922 1600
rect 37206 1664 37522 1665
rect 37206 1600 37212 1664
rect 37276 1600 37292 1664
rect 37356 1600 37372 1664
rect 37436 1600 37452 1664
rect 37516 1600 37522 1664
rect 37206 1599 37522 1600
rect 38806 1664 39122 1665
rect 38806 1600 38812 1664
rect 38876 1600 38892 1664
rect 38956 1600 38972 1664
rect 39036 1600 39052 1664
rect 39116 1600 39122 1664
rect 38806 1599 39122 1600
rect 40406 1664 40722 1665
rect 40406 1600 40412 1664
rect 40476 1600 40492 1664
rect 40556 1600 40572 1664
rect 40636 1600 40652 1664
rect 40716 1600 40722 1664
rect 40406 1599 40722 1600
rect 42006 1664 42322 1665
rect 42006 1600 42012 1664
rect 42076 1600 42092 1664
rect 42156 1600 42172 1664
rect 42236 1600 42252 1664
rect 42316 1600 42322 1664
rect 42006 1599 42322 1600
rect 43606 1664 43922 1665
rect 43606 1600 43612 1664
rect 43676 1600 43692 1664
rect 43756 1600 43772 1664
rect 43836 1600 43852 1664
rect 43916 1600 43922 1664
rect 43606 1599 43922 1600
rect 45206 1664 45522 1665
rect 45206 1600 45212 1664
rect 45276 1600 45292 1664
rect 45356 1600 45372 1664
rect 45436 1600 45452 1664
rect 45516 1600 45522 1664
rect 45206 1599 45522 1600
rect 46806 1664 47122 1665
rect 46806 1600 46812 1664
rect 46876 1600 46892 1664
rect 46956 1600 46972 1664
rect 47036 1600 47052 1664
rect 47116 1600 47122 1664
rect 46806 1599 47122 1600
rect 48406 1664 48722 1665
rect 48406 1600 48412 1664
rect 48476 1600 48492 1664
rect 48556 1600 48572 1664
rect 48636 1600 48652 1664
rect 48716 1600 48722 1664
rect 48406 1599 48722 1600
rect 50006 1664 50322 1665
rect 50006 1600 50012 1664
rect 50076 1600 50092 1664
rect 50156 1600 50172 1664
rect 50236 1600 50252 1664
rect 50316 1600 50322 1664
rect 50006 1599 50322 1600
rect 51606 1664 51922 1665
rect 51606 1600 51612 1664
rect 51676 1600 51692 1664
rect 51756 1600 51772 1664
rect 51836 1600 51852 1664
rect 51916 1600 51922 1664
rect 51606 1599 51922 1600
rect 53206 1664 53522 1665
rect 53206 1600 53212 1664
rect 53276 1600 53292 1664
rect 53356 1600 53372 1664
rect 53436 1600 53452 1664
rect 53516 1600 53522 1664
rect 53206 1599 53522 1600
rect 54806 1664 55122 1665
rect 54806 1600 54812 1664
rect 54876 1600 54892 1664
rect 54956 1600 54972 1664
rect 55036 1600 55052 1664
rect 55116 1600 55122 1664
rect 54806 1599 55122 1600
rect 56406 1664 56722 1665
rect 56406 1600 56412 1664
rect 56476 1600 56492 1664
rect 56556 1600 56572 1664
rect 56636 1600 56652 1664
rect 56716 1600 56722 1664
rect 56406 1599 56722 1600
rect 58006 1664 58322 1665
rect 58006 1600 58012 1664
rect 58076 1600 58092 1664
rect 58156 1600 58172 1664
rect 58236 1600 58252 1664
rect 58316 1600 58322 1664
rect 58006 1599 58322 1600
rect 59606 1664 59922 1665
rect 59606 1600 59612 1664
rect 59676 1600 59692 1664
rect 59756 1600 59772 1664
rect 59836 1600 59852 1664
rect 59916 1600 59922 1664
rect 59606 1599 59922 1600
rect 61206 1664 61522 1665
rect 61206 1600 61212 1664
rect 61276 1600 61292 1664
rect 61356 1600 61372 1664
rect 61436 1600 61452 1664
rect 61516 1600 61522 1664
rect 61206 1599 61522 1600
rect 62806 1664 63122 1665
rect 62806 1600 62812 1664
rect 62876 1600 62892 1664
rect 62956 1600 62972 1664
rect 63036 1600 63052 1664
rect 63116 1600 63122 1664
rect 62806 1599 63122 1600
rect 64406 1664 64722 1665
rect 64406 1600 64412 1664
rect 64476 1600 64492 1664
rect 64556 1600 64572 1664
rect 64636 1600 64652 1664
rect 64716 1600 64722 1664
rect 64406 1599 64722 1600
rect 66006 1664 66322 1665
rect 66006 1600 66012 1664
rect 66076 1600 66092 1664
rect 66156 1600 66172 1664
rect 66236 1600 66252 1664
rect 66316 1600 66322 1664
rect 66006 1599 66322 1600
rect 67606 1664 67922 1665
rect 67606 1600 67612 1664
rect 67676 1600 67692 1664
rect 67756 1600 67772 1664
rect 67836 1600 67852 1664
rect 67916 1600 67922 1664
rect 67606 1599 67922 1600
rect 69206 1664 69522 1665
rect 69206 1600 69212 1664
rect 69276 1600 69292 1664
rect 69356 1600 69372 1664
rect 69436 1600 69452 1664
rect 69516 1600 69522 1664
rect 69206 1599 69522 1600
rect 70806 1664 71122 1665
rect 70806 1600 70812 1664
rect 70876 1600 70892 1664
rect 70956 1600 70972 1664
rect 71036 1600 71052 1664
rect 71116 1600 71122 1664
rect 70806 1599 71122 1600
rect 72406 1664 72722 1665
rect 72406 1600 72412 1664
rect 72476 1600 72492 1664
rect 72556 1600 72572 1664
rect 72636 1600 72652 1664
rect 72716 1600 72722 1664
rect 72406 1599 72722 1600
rect 74006 1664 74322 1665
rect 74006 1600 74012 1664
rect 74076 1600 74092 1664
rect 74156 1600 74172 1664
rect 74236 1600 74252 1664
rect 74316 1600 74322 1664
rect 74006 1599 74322 1600
rect 75606 1664 75922 1665
rect 75606 1600 75612 1664
rect 75676 1600 75692 1664
rect 75756 1600 75772 1664
rect 75836 1600 75852 1664
rect 75916 1600 75922 1664
rect 75606 1599 75922 1600
rect 77206 1664 77522 1665
rect 77206 1600 77212 1664
rect 77276 1600 77292 1664
rect 77356 1600 77372 1664
rect 77436 1600 77452 1664
rect 77516 1600 77522 1664
rect 77206 1599 77522 1600
rect 78806 1664 79122 1665
rect 78806 1600 78812 1664
rect 78876 1600 78892 1664
rect 78956 1600 78972 1664
rect 79036 1600 79052 1664
rect 79116 1600 79122 1664
rect 78806 1599 79122 1600
rect 80406 1664 80722 1665
rect 80406 1600 80412 1664
rect 80476 1600 80492 1664
rect 80556 1600 80572 1664
rect 80636 1600 80652 1664
rect 80716 1600 80722 1664
rect 80406 1599 80722 1600
rect 82006 1664 82322 1665
rect 82006 1600 82012 1664
rect 82076 1600 82092 1664
rect 82156 1600 82172 1664
rect 82236 1600 82252 1664
rect 82316 1600 82322 1664
rect 82006 1599 82322 1600
rect 83606 1664 83922 1665
rect 83606 1600 83612 1664
rect 83676 1600 83692 1664
rect 83756 1600 83772 1664
rect 83836 1600 83852 1664
rect 83916 1600 83922 1664
rect 83606 1599 83922 1600
rect 85206 1664 85522 1665
rect 85206 1600 85212 1664
rect 85276 1600 85292 1664
rect 85356 1600 85372 1664
rect 85436 1600 85452 1664
rect 85516 1600 85522 1664
rect 85206 1599 85522 1600
rect 86806 1664 87122 1665
rect 86806 1600 86812 1664
rect 86876 1600 86892 1664
rect 86956 1600 86972 1664
rect 87036 1600 87052 1664
rect 87116 1600 87122 1664
rect 86806 1599 87122 1600
rect 88406 1664 88722 1665
rect 88406 1600 88412 1664
rect 88476 1600 88492 1664
rect 88556 1600 88572 1664
rect 88636 1600 88652 1664
rect 88716 1600 88722 1664
rect 88406 1599 88722 1600
rect 90006 1664 90322 1665
rect 90006 1600 90012 1664
rect 90076 1600 90092 1664
rect 90156 1600 90172 1664
rect 90236 1600 90252 1664
rect 90316 1600 90322 1664
rect 90006 1599 90322 1600
rect 91606 1664 91922 1665
rect 91606 1600 91612 1664
rect 91676 1600 91692 1664
rect 91756 1600 91772 1664
rect 91836 1600 91852 1664
rect 91916 1600 91922 1664
rect 91606 1599 91922 1600
rect 93206 1664 93522 1665
rect 93206 1600 93212 1664
rect 93276 1600 93292 1664
rect 93356 1600 93372 1664
rect 93436 1600 93452 1664
rect 93516 1600 93522 1664
rect 93206 1599 93522 1600
rect 94806 1664 95122 1665
rect 94806 1600 94812 1664
rect 94876 1600 94892 1664
rect 94956 1600 94972 1664
rect 95036 1600 95052 1664
rect 95116 1600 95122 1664
rect 94806 1599 95122 1600
rect 96406 1664 96722 1665
rect 96406 1600 96412 1664
rect 96476 1600 96492 1664
rect 96556 1600 96572 1664
rect 96636 1600 96652 1664
rect 96716 1600 96722 1664
rect 96406 1599 96722 1600
rect 98006 1664 98322 1665
rect 98006 1600 98012 1664
rect 98076 1600 98092 1664
rect 98156 1600 98172 1664
rect 98236 1600 98252 1664
rect 98316 1600 98322 1664
rect 98006 1599 98322 1600
rect 99606 1664 99922 1665
rect 99606 1600 99612 1664
rect 99676 1600 99692 1664
rect 99756 1600 99772 1664
rect 99836 1600 99852 1664
rect 99916 1600 99922 1664
rect 99606 1599 99922 1600
rect 101206 1664 101522 1665
rect 101206 1600 101212 1664
rect 101276 1600 101292 1664
rect 101356 1600 101372 1664
rect 101436 1600 101452 1664
rect 101516 1600 101522 1664
rect 101206 1599 101522 1600
rect 102806 1664 103122 1665
rect 102806 1600 102812 1664
rect 102876 1600 102892 1664
rect 102956 1600 102972 1664
rect 103036 1600 103052 1664
rect 103116 1600 103122 1664
rect 102806 1599 103122 1600
rect 104406 1664 104722 1665
rect 104406 1600 104412 1664
rect 104476 1600 104492 1664
rect 104556 1600 104572 1664
rect 104636 1600 104652 1664
rect 104716 1600 104722 1664
rect 104406 1599 104722 1600
rect 106006 1664 106322 1665
rect 106006 1600 106012 1664
rect 106076 1600 106092 1664
rect 106156 1600 106172 1664
rect 106236 1600 106252 1664
rect 106316 1600 106322 1664
rect 106006 1599 106322 1600
rect 107606 1664 107922 1665
rect 107606 1600 107612 1664
rect 107676 1600 107692 1664
rect 107756 1600 107772 1664
rect 107836 1600 107852 1664
rect 107916 1600 107922 1664
rect 107606 1599 107922 1600
rect 30557 1322 30623 1325
rect 33225 1324 33291 1325
rect 34513 1324 34579 1325
rect 31334 1322 31340 1324
rect 30557 1320 31340 1322
rect 30557 1264 30562 1320
rect 30618 1264 31340 1320
rect 30557 1262 31340 1264
rect 30557 1259 30623 1262
rect 31334 1260 31340 1262
rect 31404 1260 31410 1324
rect 33174 1260 33180 1324
rect 33244 1322 33291 1324
rect 33244 1320 33336 1322
rect 33286 1264 33336 1320
rect 33244 1262 33336 1264
rect 33244 1260 33291 1262
rect 34462 1260 34468 1324
rect 34532 1322 34579 1324
rect 37273 1322 37339 1325
rect 37958 1322 37964 1324
rect 34532 1320 34624 1322
rect 34574 1264 34624 1320
rect 34532 1262 34624 1264
rect 37273 1320 37964 1322
rect 37273 1264 37278 1320
rect 37334 1264 37964 1320
rect 37273 1262 37964 1264
rect 34532 1260 34579 1262
rect 33225 1259 33291 1260
rect 34513 1259 34579 1260
rect 37273 1259 37339 1262
rect 37958 1260 37964 1262
rect 38028 1260 38034 1324
rect 56593 1322 56659 1325
rect 56910 1322 56916 1324
rect 56593 1320 56916 1322
rect 56593 1264 56598 1320
rect 56654 1264 56916 1320
rect 56593 1262 56916 1264
rect 56593 1259 56659 1262
rect 56910 1260 56916 1262
rect 56980 1260 56986 1324
rect 57973 1322 58039 1325
rect 58750 1322 58756 1324
rect 57973 1320 58756 1322
rect 57973 1264 57978 1320
rect 58034 1264 58756 1320
rect 57973 1262 58756 1264
rect 57973 1259 58039 1262
rect 58750 1260 58756 1262
rect 58820 1260 58826 1324
rect 59353 1322 59419 1325
rect 60917 1324 60983 1325
rect 60222 1322 60228 1324
rect 59353 1320 60228 1322
rect 59353 1264 59358 1320
rect 59414 1264 60228 1320
rect 59353 1262 60228 1264
rect 59353 1259 59419 1262
rect 60222 1260 60228 1262
rect 60292 1260 60298 1324
rect 60917 1322 60964 1324
rect 60872 1320 60964 1322
rect 60872 1264 60922 1320
rect 60872 1262 60964 1264
rect 60917 1260 60964 1262
rect 61028 1260 61034 1324
rect 62481 1322 62547 1325
rect 63493 1324 63559 1325
rect 62614 1322 62620 1324
rect 62481 1320 62620 1322
rect 62481 1264 62486 1320
rect 62542 1264 62620 1320
rect 62481 1262 62620 1264
rect 60917 1259 60983 1260
rect 62481 1259 62547 1262
rect 62614 1260 62620 1262
rect 62684 1260 62690 1324
rect 63493 1322 63540 1324
rect 63448 1320 63540 1322
rect 63448 1264 63498 1320
rect 63448 1262 63540 1264
rect 63493 1260 63540 1262
rect 63604 1260 63610 1324
rect 64873 1322 64939 1325
rect 65006 1322 65012 1324
rect 64873 1320 65012 1322
rect 64873 1264 64878 1320
rect 64934 1264 65012 1320
rect 64873 1262 65012 1264
rect 63493 1259 63559 1260
rect 64873 1259 64939 1262
rect 65006 1260 65012 1262
rect 65076 1260 65082 1324
rect 65149 1322 65215 1325
rect 65742 1322 65748 1324
rect 65149 1320 65748 1322
rect 65149 1264 65154 1320
rect 65210 1264 65748 1320
rect 65149 1262 65748 1264
rect 65149 1259 65215 1262
rect 65742 1260 65748 1262
rect 65812 1260 65818 1324
rect 66253 1322 66319 1325
rect 67398 1322 67404 1324
rect 66253 1320 67404 1322
rect 66253 1264 66258 1320
rect 66314 1264 67404 1320
rect 66253 1262 67404 1264
rect 66253 1259 66319 1262
rect 67398 1260 67404 1262
rect 67468 1260 67474 1324
rect 67633 1322 67699 1325
rect 68318 1322 68324 1324
rect 67633 1320 68324 1322
rect 67633 1264 67638 1320
rect 67694 1264 68324 1320
rect 67633 1262 68324 1264
rect 67633 1259 67699 1262
rect 68318 1260 68324 1262
rect 68388 1260 68394 1324
rect 69013 1322 69079 1325
rect 69606 1322 69612 1324
rect 69013 1320 69612 1322
rect 69013 1264 69018 1320
rect 69074 1264 69612 1320
rect 69013 1262 69612 1264
rect 69013 1259 69079 1262
rect 69606 1260 69612 1262
rect 69676 1260 69682 1324
rect 2946 1120 3262 1121
rect 2946 1056 2952 1120
rect 3016 1056 3032 1120
rect 3096 1056 3112 1120
rect 3176 1056 3192 1120
rect 3256 1056 3262 1120
rect 2946 1055 3262 1056
rect 4546 1120 4862 1121
rect 4546 1056 4552 1120
rect 4616 1056 4632 1120
rect 4696 1056 4712 1120
rect 4776 1056 4792 1120
rect 4856 1056 4862 1120
rect 4546 1055 4862 1056
rect 6146 1120 6462 1121
rect 6146 1056 6152 1120
rect 6216 1056 6232 1120
rect 6296 1056 6312 1120
rect 6376 1056 6392 1120
rect 6456 1056 6462 1120
rect 6146 1055 6462 1056
rect 7746 1120 8062 1121
rect 7746 1056 7752 1120
rect 7816 1056 7832 1120
rect 7896 1056 7912 1120
rect 7976 1056 7992 1120
rect 8056 1056 8062 1120
rect 7746 1055 8062 1056
rect 9346 1120 9662 1121
rect 9346 1056 9352 1120
rect 9416 1056 9432 1120
rect 9496 1056 9512 1120
rect 9576 1056 9592 1120
rect 9656 1056 9662 1120
rect 9346 1055 9662 1056
rect 10946 1120 11262 1121
rect 10946 1056 10952 1120
rect 11016 1056 11032 1120
rect 11096 1056 11112 1120
rect 11176 1056 11192 1120
rect 11256 1056 11262 1120
rect 10946 1055 11262 1056
rect 12546 1120 12862 1121
rect 12546 1056 12552 1120
rect 12616 1056 12632 1120
rect 12696 1056 12712 1120
rect 12776 1056 12792 1120
rect 12856 1056 12862 1120
rect 12546 1055 12862 1056
rect 14146 1120 14462 1121
rect 14146 1056 14152 1120
rect 14216 1056 14232 1120
rect 14296 1056 14312 1120
rect 14376 1056 14392 1120
rect 14456 1056 14462 1120
rect 14146 1055 14462 1056
rect 15746 1120 16062 1121
rect 15746 1056 15752 1120
rect 15816 1056 15832 1120
rect 15896 1056 15912 1120
rect 15976 1056 15992 1120
rect 16056 1056 16062 1120
rect 15746 1055 16062 1056
rect 17346 1120 17662 1121
rect 17346 1056 17352 1120
rect 17416 1056 17432 1120
rect 17496 1056 17512 1120
rect 17576 1056 17592 1120
rect 17656 1056 17662 1120
rect 17346 1055 17662 1056
rect 18946 1120 19262 1121
rect 18946 1056 18952 1120
rect 19016 1056 19032 1120
rect 19096 1056 19112 1120
rect 19176 1056 19192 1120
rect 19256 1056 19262 1120
rect 18946 1055 19262 1056
rect 20546 1120 20862 1121
rect 20546 1056 20552 1120
rect 20616 1056 20632 1120
rect 20696 1056 20712 1120
rect 20776 1056 20792 1120
rect 20856 1056 20862 1120
rect 20546 1055 20862 1056
rect 22146 1120 22462 1121
rect 22146 1056 22152 1120
rect 22216 1056 22232 1120
rect 22296 1056 22312 1120
rect 22376 1056 22392 1120
rect 22456 1056 22462 1120
rect 22146 1055 22462 1056
rect 23746 1120 24062 1121
rect 23746 1056 23752 1120
rect 23816 1056 23832 1120
rect 23896 1056 23912 1120
rect 23976 1056 23992 1120
rect 24056 1056 24062 1120
rect 23746 1055 24062 1056
rect 25346 1120 25662 1121
rect 25346 1056 25352 1120
rect 25416 1056 25432 1120
rect 25496 1056 25512 1120
rect 25576 1056 25592 1120
rect 25656 1056 25662 1120
rect 25346 1055 25662 1056
rect 26946 1120 27262 1121
rect 26946 1056 26952 1120
rect 27016 1056 27032 1120
rect 27096 1056 27112 1120
rect 27176 1056 27192 1120
rect 27256 1056 27262 1120
rect 26946 1055 27262 1056
rect 28546 1120 28862 1121
rect 28546 1056 28552 1120
rect 28616 1056 28632 1120
rect 28696 1056 28712 1120
rect 28776 1056 28792 1120
rect 28856 1056 28862 1120
rect 28546 1055 28862 1056
rect 30146 1120 30462 1121
rect 30146 1056 30152 1120
rect 30216 1056 30232 1120
rect 30296 1056 30312 1120
rect 30376 1056 30392 1120
rect 30456 1056 30462 1120
rect 30146 1055 30462 1056
rect 31746 1120 32062 1121
rect 31746 1056 31752 1120
rect 31816 1056 31832 1120
rect 31896 1056 31912 1120
rect 31976 1056 31992 1120
rect 32056 1056 32062 1120
rect 31746 1055 32062 1056
rect 33346 1120 33662 1121
rect 33346 1056 33352 1120
rect 33416 1056 33432 1120
rect 33496 1056 33512 1120
rect 33576 1056 33592 1120
rect 33656 1056 33662 1120
rect 33346 1055 33662 1056
rect 34946 1120 35262 1121
rect 34946 1056 34952 1120
rect 35016 1056 35032 1120
rect 35096 1056 35112 1120
rect 35176 1056 35192 1120
rect 35256 1056 35262 1120
rect 34946 1055 35262 1056
rect 36546 1120 36862 1121
rect 36546 1056 36552 1120
rect 36616 1056 36632 1120
rect 36696 1056 36712 1120
rect 36776 1056 36792 1120
rect 36856 1056 36862 1120
rect 36546 1055 36862 1056
rect 38146 1120 38462 1121
rect 38146 1056 38152 1120
rect 38216 1056 38232 1120
rect 38296 1056 38312 1120
rect 38376 1056 38392 1120
rect 38456 1056 38462 1120
rect 38146 1055 38462 1056
rect 39746 1120 40062 1121
rect 39746 1056 39752 1120
rect 39816 1056 39832 1120
rect 39896 1056 39912 1120
rect 39976 1056 39992 1120
rect 40056 1056 40062 1120
rect 39746 1055 40062 1056
rect 41346 1120 41662 1121
rect 41346 1056 41352 1120
rect 41416 1056 41432 1120
rect 41496 1056 41512 1120
rect 41576 1056 41592 1120
rect 41656 1056 41662 1120
rect 41346 1055 41662 1056
rect 42946 1120 43262 1121
rect 42946 1056 42952 1120
rect 43016 1056 43032 1120
rect 43096 1056 43112 1120
rect 43176 1056 43192 1120
rect 43256 1056 43262 1120
rect 42946 1055 43262 1056
rect 44546 1120 44862 1121
rect 44546 1056 44552 1120
rect 44616 1056 44632 1120
rect 44696 1056 44712 1120
rect 44776 1056 44792 1120
rect 44856 1056 44862 1120
rect 44546 1055 44862 1056
rect 46146 1120 46462 1121
rect 46146 1056 46152 1120
rect 46216 1056 46232 1120
rect 46296 1056 46312 1120
rect 46376 1056 46392 1120
rect 46456 1056 46462 1120
rect 46146 1055 46462 1056
rect 47746 1120 48062 1121
rect 47746 1056 47752 1120
rect 47816 1056 47832 1120
rect 47896 1056 47912 1120
rect 47976 1056 47992 1120
rect 48056 1056 48062 1120
rect 47746 1055 48062 1056
rect 49346 1120 49662 1121
rect 49346 1056 49352 1120
rect 49416 1056 49432 1120
rect 49496 1056 49512 1120
rect 49576 1056 49592 1120
rect 49656 1056 49662 1120
rect 49346 1055 49662 1056
rect 50946 1120 51262 1121
rect 50946 1056 50952 1120
rect 51016 1056 51032 1120
rect 51096 1056 51112 1120
rect 51176 1056 51192 1120
rect 51256 1056 51262 1120
rect 50946 1055 51262 1056
rect 52546 1120 52862 1121
rect 52546 1056 52552 1120
rect 52616 1056 52632 1120
rect 52696 1056 52712 1120
rect 52776 1056 52792 1120
rect 52856 1056 52862 1120
rect 52546 1055 52862 1056
rect 54146 1120 54462 1121
rect 54146 1056 54152 1120
rect 54216 1056 54232 1120
rect 54296 1056 54312 1120
rect 54376 1056 54392 1120
rect 54456 1056 54462 1120
rect 54146 1055 54462 1056
rect 55746 1120 56062 1121
rect 55746 1056 55752 1120
rect 55816 1056 55832 1120
rect 55896 1056 55912 1120
rect 55976 1056 55992 1120
rect 56056 1056 56062 1120
rect 55746 1055 56062 1056
rect 57346 1120 57662 1121
rect 57346 1056 57352 1120
rect 57416 1056 57432 1120
rect 57496 1056 57512 1120
rect 57576 1056 57592 1120
rect 57656 1056 57662 1120
rect 57346 1055 57662 1056
rect 58946 1120 59262 1121
rect 58946 1056 58952 1120
rect 59016 1056 59032 1120
rect 59096 1056 59112 1120
rect 59176 1056 59192 1120
rect 59256 1056 59262 1120
rect 58946 1055 59262 1056
rect 60546 1120 60862 1121
rect 60546 1056 60552 1120
rect 60616 1056 60632 1120
rect 60696 1056 60712 1120
rect 60776 1056 60792 1120
rect 60856 1056 60862 1120
rect 60546 1055 60862 1056
rect 62146 1120 62462 1121
rect 62146 1056 62152 1120
rect 62216 1056 62232 1120
rect 62296 1056 62312 1120
rect 62376 1056 62392 1120
rect 62456 1056 62462 1120
rect 62146 1055 62462 1056
rect 63746 1120 64062 1121
rect 63746 1056 63752 1120
rect 63816 1056 63832 1120
rect 63896 1056 63912 1120
rect 63976 1056 63992 1120
rect 64056 1056 64062 1120
rect 63746 1055 64062 1056
rect 65346 1120 65662 1121
rect 65346 1056 65352 1120
rect 65416 1056 65432 1120
rect 65496 1056 65512 1120
rect 65576 1056 65592 1120
rect 65656 1056 65662 1120
rect 65346 1055 65662 1056
rect 66946 1120 67262 1121
rect 66946 1056 66952 1120
rect 67016 1056 67032 1120
rect 67096 1056 67112 1120
rect 67176 1056 67192 1120
rect 67256 1056 67262 1120
rect 66946 1055 67262 1056
rect 68546 1120 68862 1121
rect 68546 1056 68552 1120
rect 68616 1056 68632 1120
rect 68696 1056 68712 1120
rect 68776 1056 68792 1120
rect 68856 1056 68862 1120
rect 68546 1055 68862 1056
rect 70146 1120 70462 1121
rect 70146 1056 70152 1120
rect 70216 1056 70232 1120
rect 70296 1056 70312 1120
rect 70376 1056 70392 1120
rect 70456 1056 70462 1120
rect 70146 1055 70462 1056
rect 71746 1120 72062 1121
rect 71746 1056 71752 1120
rect 71816 1056 71832 1120
rect 71896 1056 71912 1120
rect 71976 1056 71992 1120
rect 72056 1056 72062 1120
rect 71746 1055 72062 1056
rect 73346 1120 73662 1121
rect 73346 1056 73352 1120
rect 73416 1056 73432 1120
rect 73496 1056 73512 1120
rect 73576 1056 73592 1120
rect 73656 1056 73662 1120
rect 73346 1055 73662 1056
rect 74946 1120 75262 1121
rect 74946 1056 74952 1120
rect 75016 1056 75032 1120
rect 75096 1056 75112 1120
rect 75176 1056 75192 1120
rect 75256 1056 75262 1120
rect 74946 1055 75262 1056
rect 76546 1120 76862 1121
rect 76546 1056 76552 1120
rect 76616 1056 76632 1120
rect 76696 1056 76712 1120
rect 76776 1056 76792 1120
rect 76856 1056 76862 1120
rect 76546 1055 76862 1056
rect 78146 1120 78462 1121
rect 78146 1056 78152 1120
rect 78216 1056 78232 1120
rect 78296 1056 78312 1120
rect 78376 1056 78392 1120
rect 78456 1056 78462 1120
rect 78146 1055 78462 1056
rect 79746 1120 80062 1121
rect 79746 1056 79752 1120
rect 79816 1056 79832 1120
rect 79896 1056 79912 1120
rect 79976 1056 79992 1120
rect 80056 1056 80062 1120
rect 79746 1055 80062 1056
rect 81346 1120 81662 1121
rect 81346 1056 81352 1120
rect 81416 1056 81432 1120
rect 81496 1056 81512 1120
rect 81576 1056 81592 1120
rect 81656 1056 81662 1120
rect 81346 1055 81662 1056
rect 82946 1120 83262 1121
rect 82946 1056 82952 1120
rect 83016 1056 83032 1120
rect 83096 1056 83112 1120
rect 83176 1056 83192 1120
rect 83256 1056 83262 1120
rect 82946 1055 83262 1056
rect 84546 1120 84862 1121
rect 84546 1056 84552 1120
rect 84616 1056 84632 1120
rect 84696 1056 84712 1120
rect 84776 1056 84792 1120
rect 84856 1056 84862 1120
rect 84546 1055 84862 1056
rect 86146 1120 86462 1121
rect 86146 1056 86152 1120
rect 86216 1056 86232 1120
rect 86296 1056 86312 1120
rect 86376 1056 86392 1120
rect 86456 1056 86462 1120
rect 86146 1055 86462 1056
rect 87746 1120 88062 1121
rect 87746 1056 87752 1120
rect 87816 1056 87832 1120
rect 87896 1056 87912 1120
rect 87976 1056 87992 1120
rect 88056 1056 88062 1120
rect 87746 1055 88062 1056
rect 89346 1120 89662 1121
rect 89346 1056 89352 1120
rect 89416 1056 89432 1120
rect 89496 1056 89512 1120
rect 89576 1056 89592 1120
rect 89656 1056 89662 1120
rect 89346 1055 89662 1056
rect 90946 1120 91262 1121
rect 90946 1056 90952 1120
rect 91016 1056 91032 1120
rect 91096 1056 91112 1120
rect 91176 1056 91192 1120
rect 91256 1056 91262 1120
rect 90946 1055 91262 1056
rect 92546 1120 92862 1121
rect 92546 1056 92552 1120
rect 92616 1056 92632 1120
rect 92696 1056 92712 1120
rect 92776 1056 92792 1120
rect 92856 1056 92862 1120
rect 92546 1055 92862 1056
rect 94146 1120 94462 1121
rect 94146 1056 94152 1120
rect 94216 1056 94232 1120
rect 94296 1056 94312 1120
rect 94376 1056 94392 1120
rect 94456 1056 94462 1120
rect 94146 1055 94462 1056
rect 95746 1120 96062 1121
rect 95746 1056 95752 1120
rect 95816 1056 95832 1120
rect 95896 1056 95912 1120
rect 95976 1056 95992 1120
rect 96056 1056 96062 1120
rect 95746 1055 96062 1056
rect 97346 1120 97662 1121
rect 97346 1056 97352 1120
rect 97416 1056 97432 1120
rect 97496 1056 97512 1120
rect 97576 1056 97592 1120
rect 97656 1056 97662 1120
rect 97346 1055 97662 1056
rect 98946 1120 99262 1121
rect 98946 1056 98952 1120
rect 99016 1056 99032 1120
rect 99096 1056 99112 1120
rect 99176 1056 99192 1120
rect 99256 1056 99262 1120
rect 98946 1055 99262 1056
rect 100546 1120 100862 1121
rect 100546 1056 100552 1120
rect 100616 1056 100632 1120
rect 100696 1056 100712 1120
rect 100776 1056 100792 1120
rect 100856 1056 100862 1120
rect 100546 1055 100862 1056
rect 102146 1120 102462 1121
rect 102146 1056 102152 1120
rect 102216 1056 102232 1120
rect 102296 1056 102312 1120
rect 102376 1056 102392 1120
rect 102456 1056 102462 1120
rect 102146 1055 102462 1056
rect 103746 1120 104062 1121
rect 103746 1056 103752 1120
rect 103816 1056 103832 1120
rect 103896 1056 103912 1120
rect 103976 1056 103992 1120
rect 104056 1056 104062 1120
rect 103746 1055 104062 1056
rect 105346 1120 105662 1121
rect 105346 1056 105352 1120
rect 105416 1056 105432 1120
rect 105496 1056 105512 1120
rect 105576 1056 105592 1120
rect 105656 1056 105662 1120
rect 105346 1055 105662 1056
rect 106946 1120 107262 1121
rect 106946 1056 106952 1120
rect 107016 1056 107032 1120
rect 107096 1056 107112 1120
rect 107176 1056 107192 1120
rect 107256 1056 107262 1120
rect 106946 1055 107262 1056
rect 108546 1120 108862 1121
rect 108546 1056 108552 1120
rect 108616 1056 108632 1120
rect 108696 1056 108712 1120
rect 108776 1056 108792 1120
rect 108856 1056 108862 1120
rect 108546 1055 108862 1056
rect 26325 914 26391 917
rect 53046 914 53052 916
rect 26325 912 53052 914
rect 26325 856 26330 912
rect 26386 856 53052 912
rect 26325 854 53052 856
rect 26325 851 26391 854
rect 53046 852 53052 854
rect 53116 852 53122 916
rect 4981 778 5047 781
rect 93894 778 93900 780
rect 4981 776 93900 778
rect 4981 720 4986 776
rect 5042 720 93900 776
rect 4981 718 93900 720
rect 4981 715 5047 718
rect 93894 716 93900 718
rect 93964 716 93970 780
rect 10726 580 10732 644
rect 10796 642 10802 644
rect 27470 642 27476 644
rect 10796 582 27476 642
rect 10796 580 10802 582
rect 27470 580 27476 582
rect 27540 580 27546 644
rect 32213 642 32279 645
rect 52310 642 52316 644
rect 32213 640 52316 642
rect 32213 584 32218 640
rect 32274 584 52316 640
rect 32213 582 52316 584
rect 32213 579 32279 582
rect 52310 580 52316 582
rect 52380 580 52386 644
rect 10593 506 10659 509
rect 41822 506 41828 508
rect 10593 504 41828 506
rect 10593 448 10598 504
rect 10654 448 41828 504
rect 10593 446 41828 448
rect 10593 443 10659 446
rect 41822 444 41828 446
rect 41892 444 41898 508
rect 1301 370 1367 373
rect 33133 370 33199 373
rect 1301 368 33199 370
rect 1301 312 1306 368
rect 1362 312 33138 368
rect 33194 312 33199 368
rect 1301 310 33199 312
rect 1301 307 1367 310
rect 33133 307 33199 310
<< via3 >>
rect 3612 86524 3676 86528
rect 3612 86468 3616 86524
rect 3616 86468 3672 86524
rect 3672 86468 3676 86524
rect 3612 86464 3676 86468
rect 3692 86524 3756 86528
rect 3692 86468 3696 86524
rect 3696 86468 3752 86524
rect 3752 86468 3756 86524
rect 3692 86464 3756 86468
rect 3772 86524 3836 86528
rect 3772 86468 3776 86524
rect 3776 86468 3832 86524
rect 3832 86468 3836 86524
rect 3772 86464 3836 86468
rect 3852 86524 3916 86528
rect 3852 86468 3856 86524
rect 3856 86468 3912 86524
rect 3912 86468 3916 86524
rect 3852 86464 3916 86468
rect 5212 86524 5276 86528
rect 5212 86468 5216 86524
rect 5216 86468 5272 86524
rect 5272 86468 5276 86524
rect 5212 86464 5276 86468
rect 5292 86524 5356 86528
rect 5292 86468 5296 86524
rect 5296 86468 5352 86524
rect 5352 86468 5356 86524
rect 5292 86464 5356 86468
rect 5372 86524 5436 86528
rect 5372 86468 5376 86524
rect 5376 86468 5432 86524
rect 5432 86468 5436 86524
rect 5372 86464 5436 86468
rect 5452 86524 5516 86528
rect 5452 86468 5456 86524
rect 5456 86468 5512 86524
rect 5512 86468 5516 86524
rect 5452 86464 5516 86468
rect 6812 86524 6876 86528
rect 6812 86468 6816 86524
rect 6816 86468 6872 86524
rect 6872 86468 6876 86524
rect 6812 86464 6876 86468
rect 6892 86524 6956 86528
rect 6892 86468 6896 86524
rect 6896 86468 6952 86524
rect 6952 86468 6956 86524
rect 6892 86464 6956 86468
rect 6972 86524 7036 86528
rect 6972 86468 6976 86524
rect 6976 86468 7032 86524
rect 7032 86468 7036 86524
rect 6972 86464 7036 86468
rect 7052 86524 7116 86528
rect 7052 86468 7056 86524
rect 7056 86468 7112 86524
rect 7112 86468 7116 86524
rect 7052 86464 7116 86468
rect 8412 86524 8476 86528
rect 8412 86468 8416 86524
rect 8416 86468 8472 86524
rect 8472 86468 8476 86524
rect 8412 86464 8476 86468
rect 8492 86524 8556 86528
rect 8492 86468 8496 86524
rect 8496 86468 8552 86524
rect 8552 86468 8556 86524
rect 8492 86464 8556 86468
rect 8572 86524 8636 86528
rect 8572 86468 8576 86524
rect 8576 86468 8632 86524
rect 8632 86468 8636 86524
rect 8572 86464 8636 86468
rect 8652 86524 8716 86528
rect 8652 86468 8656 86524
rect 8656 86468 8712 86524
rect 8712 86468 8716 86524
rect 8652 86464 8716 86468
rect 10012 86524 10076 86528
rect 10012 86468 10016 86524
rect 10016 86468 10072 86524
rect 10072 86468 10076 86524
rect 10012 86464 10076 86468
rect 10092 86524 10156 86528
rect 10092 86468 10096 86524
rect 10096 86468 10152 86524
rect 10152 86468 10156 86524
rect 10092 86464 10156 86468
rect 10172 86524 10236 86528
rect 10172 86468 10176 86524
rect 10176 86468 10232 86524
rect 10232 86468 10236 86524
rect 10172 86464 10236 86468
rect 10252 86524 10316 86528
rect 10252 86468 10256 86524
rect 10256 86468 10312 86524
rect 10312 86468 10316 86524
rect 10252 86464 10316 86468
rect 11612 86524 11676 86528
rect 11612 86468 11616 86524
rect 11616 86468 11672 86524
rect 11672 86468 11676 86524
rect 11612 86464 11676 86468
rect 11692 86524 11756 86528
rect 11692 86468 11696 86524
rect 11696 86468 11752 86524
rect 11752 86468 11756 86524
rect 11692 86464 11756 86468
rect 11772 86524 11836 86528
rect 11772 86468 11776 86524
rect 11776 86468 11832 86524
rect 11832 86468 11836 86524
rect 11772 86464 11836 86468
rect 11852 86524 11916 86528
rect 11852 86468 11856 86524
rect 11856 86468 11912 86524
rect 11912 86468 11916 86524
rect 11852 86464 11916 86468
rect 13212 86524 13276 86528
rect 13212 86468 13216 86524
rect 13216 86468 13272 86524
rect 13272 86468 13276 86524
rect 13212 86464 13276 86468
rect 13292 86524 13356 86528
rect 13292 86468 13296 86524
rect 13296 86468 13352 86524
rect 13352 86468 13356 86524
rect 13292 86464 13356 86468
rect 13372 86524 13436 86528
rect 13372 86468 13376 86524
rect 13376 86468 13432 86524
rect 13432 86468 13436 86524
rect 13372 86464 13436 86468
rect 13452 86524 13516 86528
rect 13452 86468 13456 86524
rect 13456 86468 13512 86524
rect 13512 86468 13516 86524
rect 13452 86464 13516 86468
rect 14812 86524 14876 86528
rect 14812 86468 14816 86524
rect 14816 86468 14872 86524
rect 14872 86468 14876 86524
rect 14812 86464 14876 86468
rect 14892 86524 14956 86528
rect 14892 86468 14896 86524
rect 14896 86468 14952 86524
rect 14952 86468 14956 86524
rect 14892 86464 14956 86468
rect 14972 86524 15036 86528
rect 14972 86468 14976 86524
rect 14976 86468 15032 86524
rect 15032 86468 15036 86524
rect 14972 86464 15036 86468
rect 15052 86524 15116 86528
rect 15052 86468 15056 86524
rect 15056 86468 15112 86524
rect 15112 86468 15116 86524
rect 15052 86464 15116 86468
rect 16412 86524 16476 86528
rect 16412 86468 16416 86524
rect 16416 86468 16472 86524
rect 16472 86468 16476 86524
rect 16412 86464 16476 86468
rect 16492 86524 16556 86528
rect 16492 86468 16496 86524
rect 16496 86468 16552 86524
rect 16552 86468 16556 86524
rect 16492 86464 16556 86468
rect 16572 86524 16636 86528
rect 16572 86468 16576 86524
rect 16576 86468 16632 86524
rect 16632 86468 16636 86524
rect 16572 86464 16636 86468
rect 16652 86524 16716 86528
rect 16652 86468 16656 86524
rect 16656 86468 16712 86524
rect 16712 86468 16716 86524
rect 16652 86464 16716 86468
rect 18012 86524 18076 86528
rect 18012 86468 18016 86524
rect 18016 86468 18072 86524
rect 18072 86468 18076 86524
rect 18012 86464 18076 86468
rect 18092 86524 18156 86528
rect 18092 86468 18096 86524
rect 18096 86468 18152 86524
rect 18152 86468 18156 86524
rect 18092 86464 18156 86468
rect 18172 86524 18236 86528
rect 18172 86468 18176 86524
rect 18176 86468 18232 86524
rect 18232 86468 18236 86524
rect 18172 86464 18236 86468
rect 18252 86524 18316 86528
rect 18252 86468 18256 86524
rect 18256 86468 18312 86524
rect 18312 86468 18316 86524
rect 18252 86464 18316 86468
rect 19612 86524 19676 86528
rect 19612 86468 19616 86524
rect 19616 86468 19672 86524
rect 19672 86468 19676 86524
rect 19612 86464 19676 86468
rect 19692 86524 19756 86528
rect 19692 86468 19696 86524
rect 19696 86468 19752 86524
rect 19752 86468 19756 86524
rect 19692 86464 19756 86468
rect 19772 86524 19836 86528
rect 19772 86468 19776 86524
rect 19776 86468 19832 86524
rect 19832 86468 19836 86524
rect 19772 86464 19836 86468
rect 19852 86524 19916 86528
rect 19852 86468 19856 86524
rect 19856 86468 19912 86524
rect 19912 86468 19916 86524
rect 19852 86464 19916 86468
rect 21212 86524 21276 86528
rect 21212 86468 21216 86524
rect 21216 86468 21272 86524
rect 21272 86468 21276 86524
rect 21212 86464 21276 86468
rect 21292 86524 21356 86528
rect 21292 86468 21296 86524
rect 21296 86468 21352 86524
rect 21352 86468 21356 86524
rect 21292 86464 21356 86468
rect 21372 86524 21436 86528
rect 21372 86468 21376 86524
rect 21376 86468 21432 86524
rect 21432 86468 21436 86524
rect 21372 86464 21436 86468
rect 21452 86524 21516 86528
rect 21452 86468 21456 86524
rect 21456 86468 21512 86524
rect 21512 86468 21516 86524
rect 21452 86464 21516 86468
rect 22812 86524 22876 86528
rect 22812 86468 22816 86524
rect 22816 86468 22872 86524
rect 22872 86468 22876 86524
rect 22812 86464 22876 86468
rect 22892 86524 22956 86528
rect 22892 86468 22896 86524
rect 22896 86468 22952 86524
rect 22952 86468 22956 86524
rect 22892 86464 22956 86468
rect 22972 86524 23036 86528
rect 22972 86468 22976 86524
rect 22976 86468 23032 86524
rect 23032 86468 23036 86524
rect 22972 86464 23036 86468
rect 23052 86524 23116 86528
rect 23052 86468 23056 86524
rect 23056 86468 23112 86524
rect 23112 86468 23116 86524
rect 23052 86464 23116 86468
rect 24412 86524 24476 86528
rect 24412 86468 24416 86524
rect 24416 86468 24472 86524
rect 24472 86468 24476 86524
rect 24412 86464 24476 86468
rect 24492 86524 24556 86528
rect 24492 86468 24496 86524
rect 24496 86468 24552 86524
rect 24552 86468 24556 86524
rect 24492 86464 24556 86468
rect 24572 86524 24636 86528
rect 24572 86468 24576 86524
rect 24576 86468 24632 86524
rect 24632 86468 24636 86524
rect 24572 86464 24636 86468
rect 24652 86524 24716 86528
rect 24652 86468 24656 86524
rect 24656 86468 24712 86524
rect 24712 86468 24716 86524
rect 24652 86464 24716 86468
rect 26012 86524 26076 86528
rect 26012 86468 26016 86524
rect 26016 86468 26072 86524
rect 26072 86468 26076 86524
rect 26012 86464 26076 86468
rect 26092 86524 26156 86528
rect 26092 86468 26096 86524
rect 26096 86468 26152 86524
rect 26152 86468 26156 86524
rect 26092 86464 26156 86468
rect 26172 86524 26236 86528
rect 26172 86468 26176 86524
rect 26176 86468 26232 86524
rect 26232 86468 26236 86524
rect 26172 86464 26236 86468
rect 26252 86524 26316 86528
rect 26252 86468 26256 86524
rect 26256 86468 26312 86524
rect 26312 86468 26316 86524
rect 26252 86464 26316 86468
rect 27612 86524 27676 86528
rect 27612 86468 27616 86524
rect 27616 86468 27672 86524
rect 27672 86468 27676 86524
rect 27612 86464 27676 86468
rect 27692 86524 27756 86528
rect 27692 86468 27696 86524
rect 27696 86468 27752 86524
rect 27752 86468 27756 86524
rect 27692 86464 27756 86468
rect 27772 86524 27836 86528
rect 27772 86468 27776 86524
rect 27776 86468 27832 86524
rect 27832 86468 27836 86524
rect 27772 86464 27836 86468
rect 27852 86524 27916 86528
rect 27852 86468 27856 86524
rect 27856 86468 27912 86524
rect 27912 86468 27916 86524
rect 27852 86464 27916 86468
rect 29212 86524 29276 86528
rect 29212 86468 29216 86524
rect 29216 86468 29272 86524
rect 29272 86468 29276 86524
rect 29212 86464 29276 86468
rect 29292 86524 29356 86528
rect 29292 86468 29296 86524
rect 29296 86468 29352 86524
rect 29352 86468 29356 86524
rect 29292 86464 29356 86468
rect 29372 86524 29436 86528
rect 29372 86468 29376 86524
rect 29376 86468 29432 86524
rect 29432 86468 29436 86524
rect 29372 86464 29436 86468
rect 29452 86524 29516 86528
rect 29452 86468 29456 86524
rect 29456 86468 29512 86524
rect 29512 86468 29516 86524
rect 29452 86464 29516 86468
rect 30812 86524 30876 86528
rect 30812 86468 30816 86524
rect 30816 86468 30872 86524
rect 30872 86468 30876 86524
rect 30812 86464 30876 86468
rect 30892 86524 30956 86528
rect 30892 86468 30896 86524
rect 30896 86468 30952 86524
rect 30952 86468 30956 86524
rect 30892 86464 30956 86468
rect 30972 86524 31036 86528
rect 30972 86468 30976 86524
rect 30976 86468 31032 86524
rect 31032 86468 31036 86524
rect 30972 86464 31036 86468
rect 31052 86524 31116 86528
rect 31052 86468 31056 86524
rect 31056 86468 31112 86524
rect 31112 86468 31116 86524
rect 31052 86464 31116 86468
rect 32412 86524 32476 86528
rect 32412 86468 32416 86524
rect 32416 86468 32472 86524
rect 32472 86468 32476 86524
rect 32412 86464 32476 86468
rect 32492 86524 32556 86528
rect 32492 86468 32496 86524
rect 32496 86468 32552 86524
rect 32552 86468 32556 86524
rect 32492 86464 32556 86468
rect 32572 86524 32636 86528
rect 32572 86468 32576 86524
rect 32576 86468 32632 86524
rect 32632 86468 32636 86524
rect 32572 86464 32636 86468
rect 32652 86524 32716 86528
rect 32652 86468 32656 86524
rect 32656 86468 32712 86524
rect 32712 86468 32716 86524
rect 32652 86464 32716 86468
rect 34012 86524 34076 86528
rect 34012 86468 34016 86524
rect 34016 86468 34072 86524
rect 34072 86468 34076 86524
rect 34012 86464 34076 86468
rect 34092 86524 34156 86528
rect 34092 86468 34096 86524
rect 34096 86468 34152 86524
rect 34152 86468 34156 86524
rect 34092 86464 34156 86468
rect 34172 86524 34236 86528
rect 34172 86468 34176 86524
rect 34176 86468 34232 86524
rect 34232 86468 34236 86524
rect 34172 86464 34236 86468
rect 34252 86524 34316 86528
rect 34252 86468 34256 86524
rect 34256 86468 34312 86524
rect 34312 86468 34316 86524
rect 34252 86464 34316 86468
rect 35612 86524 35676 86528
rect 35612 86468 35616 86524
rect 35616 86468 35672 86524
rect 35672 86468 35676 86524
rect 35612 86464 35676 86468
rect 35692 86524 35756 86528
rect 35692 86468 35696 86524
rect 35696 86468 35752 86524
rect 35752 86468 35756 86524
rect 35692 86464 35756 86468
rect 35772 86524 35836 86528
rect 35772 86468 35776 86524
rect 35776 86468 35832 86524
rect 35832 86468 35836 86524
rect 35772 86464 35836 86468
rect 35852 86524 35916 86528
rect 35852 86468 35856 86524
rect 35856 86468 35912 86524
rect 35912 86468 35916 86524
rect 35852 86464 35916 86468
rect 37212 86524 37276 86528
rect 37212 86468 37216 86524
rect 37216 86468 37272 86524
rect 37272 86468 37276 86524
rect 37212 86464 37276 86468
rect 37292 86524 37356 86528
rect 37292 86468 37296 86524
rect 37296 86468 37352 86524
rect 37352 86468 37356 86524
rect 37292 86464 37356 86468
rect 37372 86524 37436 86528
rect 37372 86468 37376 86524
rect 37376 86468 37432 86524
rect 37432 86468 37436 86524
rect 37372 86464 37436 86468
rect 37452 86524 37516 86528
rect 37452 86468 37456 86524
rect 37456 86468 37512 86524
rect 37512 86468 37516 86524
rect 37452 86464 37516 86468
rect 38812 86524 38876 86528
rect 38812 86468 38816 86524
rect 38816 86468 38872 86524
rect 38872 86468 38876 86524
rect 38812 86464 38876 86468
rect 38892 86524 38956 86528
rect 38892 86468 38896 86524
rect 38896 86468 38952 86524
rect 38952 86468 38956 86524
rect 38892 86464 38956 86468
rect 38972 86524 39036 86528
rect 38972 86468 38976 86524
rect 38976 86468 39032 86524
rect 39032 86468 39036 86524
rect 38972 86464 39036 86468
rect 39052 86524 39116 86528
rect 39052 86468 39056 86524
rect 39056 86468 39112 86524
rect 39112 86468 39116 86524
rect 39052 86464 39116 86468
rect 40412 86524 40476 86528
rect 40412 86468 40416 86524
rect 40416 86468 40472 86524
rect 40472 86468 40476 86524
rect 40412 86464 40476 86468
rect 40492 86524 40556 86528
rect 40492 86468 40496 86524
rect 40496 86468 40552 86524
rect 40552 86468 40556 86524
rect 40492 86464 40556 86468
rect 40572 86524 40636 86528
rect 40572 86468 40576 86524
rect 40576 86468 40632 86524
rect 40632 86468 40636 86524
rect 40572 86464 40636 86468
rect 40652 86524 40716 86528
rect 40652 86468 40656 86524
rect 40656 86468 40712 86524
rect 40712 86468 40716 86524
rect 40652 86464 40716 86468
rect 42012 86524 42076 86528
rect 42012 86468 42016 86524
rect 42016 86468 42072 86524
rect 42072 86468 42076 86524
rect 42012 86464 42076 86468
rect 42092 86524 42156 86528
rect 42092 86468 42096 86524
rect 42096 86468 42152 86524
rect 42152 86468 42156 86524
rect 42092 86464 42156 86468
rect 42172 86524 42236 86528
rect 42172 86468 42176 86524
rect 42176 86468 42232 86524
rect 42232 86468 42236 86524
rect 42172 86464 42236 86468
rect 42252 86524 42316 86528
rect 42252 86468 42256 86524
rect 42256 86468 42312 86524
rect 42312 86468 42316 86524
rect 42252 86464 42316 86468
rect 43612 86524 43676 86528
rect 43612 86468 43616 86524
rect 43616 86468 43672 86524
rect 43672 86468 43676 86524
rect 43612 86464 43676 86468
rect 43692 86524 43756 86528
rect 43692 86468 43696 86524
rect 43696 86468 43752 86524
rect 43752 86468 43756 86524
rect 43692 86464 43756 86468
rect 43772 86524 43836 86528
rect 43772 86468 43776 86524
rect 43776 86468 43832 86524
rect 43832 86468 43836 86524
rect 43772 86464 43836 86468
rect 43852 86524 43916 86528
rect 43852 86468 43856 86524
rect 43856 86468 43912 86524
rect 43912 86468 43916 86524
rect 43852 86464 43916 86468
rect 45212 86524 45276 86528
rect 45212 86468 45216 86524
rect 45216 86468 45272 86524
rect 45272 86468 45276 86524
rect 45212 86464 45276 86468
rect 45292 86524 45356 86528
rect 45292 86468 45296 86524
rect 45296 86468 45352 86524
rect 45352 86468 45356 86524
rect 45292 86464 45356 86468
rect 45372 86524 45436 86528
rect 45372 86468 45376 86524
rect 45376 86468 45432 86524
rect 45432 86468 45436 86524
rect 45372 86464 45436 86468
rect 45452 86524 45516 86528
rect 45452 86468 45456 86524
rect 45456 86468 45512 86524
rect 45512 86468 45516 86524
rect 45452 86464 45516 86468
rect 46812 86524 46876 86528
rect 46812 86468 46816 86524
rect 46816 86468 46872 86524
rect 46872 86468 46876 86524
rect 46812 86464 46876 86468
rect 46892 86524 46956 86528
rect 46892 86468 46896 86524
rect 46896 86468 46952 86524
rect 46952 86468 46956 86524
rect 46892 86464 46956 86468
rect 46972 86524 47036 86528
rect 46972 86468 46976 86524
rect 46976 86468 47032 86524
rect 47032 86468 47036 86524
rect 46972 86464 47036 86468
rect 47052 86524 47116 86528
rect 47052 86468 47056 86524
rect 47056 86468 47112 86524
rect 47112 86468 47116 86524
rect 47052 86464 47116 86468
rect 48412 86524 48476 86528
rect 48412 86468 48416 86524
rect 48416 86468 48472 86524
rect 48472 86468 48476 86524
rect 48412 86464 48476 86468
rect 48492 86524 48556 86528
rect 48492 86468 48496 86524
rect 48496 86468 48552 86524
rect 48552 86468 48556 86524
rect 48492 86464 48556 86468
rect 48572 86524 48636 86528
rect 48572 86468 48576 86524
rect 48576 86468 48632 86524
rect 48632 86468 48636 86524
rect 48572 86464 48636 86468
rect 48652 86524 48716 86528
rect 48652 86468 48656 86524
rect 48656 86468 48712 86524
rect 48712 86468 48716 86524
rect 48652 86464 48716 86468
rect 50012 86524 50076 86528
rect 50012 86468 50016 86524
rect 50016 86468 50072 86524
rect 50072 86468 50076 86524
rect 50012 86464 50076 86468
rect 50092 86524 50156 86528
rect 50092 86468 50096 86524
rect 50096 86468 50152 86524
rect 50152 86468 50156 86524
rect 50092 86464 50156 86468
rect 50172 86524 50236 86528
rect 50172 86468 50176 86524
rect 50176 86468 50232 86524
rect 50232 86468 50236 86524
rect 50172 86464 50236 86468
rect 50252 86524 50316 86528
rect 50252 86468 50256 86524
rect 50256 86468 50312 86524
rect 50312 86468 50316 86524
rect 50252 86464 50316 86468
rect 51612 86524 51676 86528
rect 51612 86468 51616 86524
rect 51616 86468 51672 86524
rect 51672 86468 51676 86524
rect 51612 86464 51676 86468
rect 51692 86524 51756 86528
rect 51692 86468 51696 86524
rect 51696 86468 51752 86524
rect 51752 86468 51756 86524
rect 51692 86464 51756 86468
rect 51772 86524 51836 86528
rect 51772 86468 51776 86524
rect 51776 86468 51832 86524
rect 51832 86468 51836 86524
rect 51772 86464 51836 86468
rect 51852 86524 51916 86528
rect 51852 86468 51856 86524
rect 51856 86468 51912 86524
rect 51912 86468 51916 86524
rect 51852 86464 51916 86468
rect 53212 86524 53276 86528
rect 53212 86468 53216 86524
rect 53216 86468 53272 86524
rect 53272 86468 53276 86524
rect 53212 86464 53276 86468
rect 53292 86524 53356 86528
rect 53292 86468 53296 86524
rect 53296 86468 53352 86524
rect 53352 86468 53356 86524
rect 53292 86464 53356 86468
rect 53372 86524 53436 86528
rect 53372 86468 53376 86524
rect 53376 86468 53432 86524
rect 53432 86468 53436 86524
rect 53372 86464 53436 86468
rect 53452 86524 53516 86528
rect 53452 86468 53456 86524
rect 53456 86468 53512 86524
rect 53512 86468 53516 86524
rect 53452 86464 53516 86468
rect 54812 86524 54876 86528
rect 54812 86468 54816 86524
rect 54816 86468 54872 86524
rect 54872 86468 54876 86524
rect 54812 86464 54876 86468
rect 54892 86524 54956 86528
rect 54892 86468 54896 86524
rect 54896 86468 54952 86524
rect 54952 86468 54956 86524
rect 54892 86464 54956 86468
rect 54972 86524 55036 86528
rect 54972 86468 54976 86524
rect 54976 86468 55032 86524
rect 55032 86468 55036 86524
rect 54972 86464 55036 86468
rect 55052 86524 55116 86528
rect 55052 86468 55056 86524
rect 55056 86468 55112 86524
rect 55112 86468 55116 86524
rect 55052 86464 55116 86468
rect 56412 86524 56476 86528
rect 56412 86468 56416 86524
rect 56416 86468 56472 86524
rect 56472 86468 56476 86524
rect 56412 86464 56476 86468
rect 56492 86524 56556 86528
rect 56492 86468 56496 86524
rect 56496 86468 56552 86524
rect 56552 86468 56556 86524
rect 56492 86464 56556 86468
rect 56572 86524 56636 86528
rect 56572 86468 56576 86524
rect 56576 86468 56632 86524
rect 56632 86468 56636 86524
rect 56572 86464 56636 86468
rect 56652 86524 56716 86528
rect 56652 86468 56656 86524
rect 56656 86468 56712 86524
rect 56712 86468 56716 86524
rect 56652 86464 56716 86468
rect 58012 86524 58076 86528
rect 58012 86468 58016 86524
rect 58016 86468 58072 86524
rect 58072 86468 58076 86524
rect 58012 86464 58076 86468
rect 58092 86524 58156 86528
rect 58092 86468 58096 86524
rect 58096 86468 58152 86524
rect 58152 86468 58156 86524
rect 58092 86464 58156 86468
rect 58172 86524 58236 86528
rect 58172 86468 58176 86524
rect 58176 86468 58232 86524
rect 58232 86468 58236 86524
rect 58172 86464 58236 86468
rect 58252 86524 58316 86528
rect 58252 86468 58256 86524
rect 58256 86468 58312 86524
rect 58312 86468 58316 86524
rect 58252 86464 58316 86468
rect 59612 86524 59676 86528
rect 59612 86468 59616 86524
rect 59616 86468 59672 86524
rect 59672 86468 59676 86524
rect 59612 86464 59676 86468
rect 59692 86524 59756 86528
rect 59692 86468 59696 86524
rect 59696 86468 59752 86524
rect 59752 86468 59756 86524
rect 59692 86464 59756 86468
rect 59772 86524 59836 86528
rect 59772 86468 59776 86524
rect 59776 86468 59832 86524
rect 59832 86468 59836 86524
rect 59772 86464 59836 86468
rect 59852 86524 59916 86528
rect 59852 86468 59856 86524
rect 59856 86468 59912 86524
rect 59912 86468 59916 86524
rect 59852 86464 59916 86468
rect 61212 86524 61276 86528
rect 61212 86468 61216 86524
rect 61216 86468 61272 86524
rect 61272 86468 61276 86524
rect 61212 86464 61276 86468
rect 61292 86524 61356 86528
rect 61292 86468 61296 86524
rect 61296 86468 61352 86524
rect 61352 86468 61356 86524
rect 61292 86464 61356 86468
rect 61372 86524 61436 86528
rect 61372 86468 61376 86524
rect 61376 86468 61432 86524
rect 61432 86468 61436 86524
rect 61372 86464 61436 86468
rect 61452 86524 61516 86528
rect 61452 86468 61456 86524
rect 61456 86468 61512 86524
rect 61512 86468 61516 86524
rect 61452 86464 61516 86468
rect 62812 86524 62876 86528
rect 62812 86468 62816 86524
rect 62816 86468 62872 86524
rect 62872 86468 62876 86524
rect 62812 86464 62876 86468
rect 62892 86524 62956 86528
rect 62892 86468 62896 86524
rect 62896 86468 62952 86524
rect 62952 86468 62956 86524
rect 62892 86464 62956 86468
rect 62972 86524 63036 86528
rect 62972 86468 62976 86524
rect 62976 86468 63032 86524
rect 63032 86468 63036 86524
rect 62972 86464 63036 86468
rect 63052 86524 63116 86528
rect 63052 86468 63056 86524
rect 63056 86468 63112 86524
rect 63112 86468 63116 86524
rect 63052 86464 63116 86468
rect 64412 86524 64476 86528
rect 64412 86468 64416 86524
rect 64416 86468 64472 86524
rect 64472 86468 64476 86524
rect 64412 86464 64476 86468
rect 64492 86524 64556 86528
rect 64492 86468 64496 86524
rect 64496 86468 64552 86524
rect 64552 86468 64556 86524
rect 64492 86464 64556 86468
rect 64572 86524 64636 86528
rect 64572 86468 64576 86524
rect 64576 86468 64632 86524
rect 64632 86468 64636 86524
rect 64572 86464 64636 86468
rect 64652 86524 64716 86528
rect 64652 86468 64656 86524
rect 64656 86468 64712 86524
rect 64712 86468 64716 86524
rect 64652 86464 64716 86468
rect 66012 86524 66076 86528
rect 66012 86468 66016 86524
rect 66016 86468 66072 86524
rect 66072 86468 66076 86524
rect 66012 86464 66076 86468
rect 66092 86524 66156 86528
rect 66092 86468 66096 86524
rect 66096 86468 66152 86524
rect 66152 86468 66156 86524
rect 66092 86464 66156 86468
rect 66172 86524 66236 86528
rect 66172 86468 66176 86524
rect 66176 86468 66232 86524
rect 66232 86468 66236 86524
rect 66172 86464 66236 86468
rect 66252 86524 66316 86528
rect 66252 86468 66256 86524
rect 66256 86468 66312 86524
rect 66312 86468 66316 86524
rect 66252 86464 66316 86468
rect 67612 86524 67676 86528
rect 67612 86468 67616 86524
rect 67616 86468 67672 86524
rect 67672 86468 67676 86524
rect 67612 86464 67676 86468
rect 67692 86524 67756 86528
rect 67692 86468 67696 86524
rect 67696 86468 67752 86524
rect 67752 86468 67756 86524
rect 67692 86464 67756 86468
rect 67772 86524 67836 86528
rect 67772 86468 67776 86524
rect 67776 86468 67832 86524
rect 67832 86468 67836 86524
rect 67772 86464 67836 86468
rect 67852 86524 67916 86528
rect 67852 86468 67856 86524
rect 67856 86468 67912 86524
rect 67912 86468 67916 86524
rect 67852 86464 67916 86468
rect 69212 86524 69276 86528
rect 69212 86468 69216 86524
rect 69216 86468 69272 86524
rect 69272 86468 69276 86524
rect 69212 86464 69276 86468
rect 69292 86524 69356 86528
rect 69292 86468 69296 86524
rect 69296 86468 69352 86524
rect 69352 86468 69356 86524
rect 69292 86464 69356 86468
rect 69372 86524 69436 86528
rect 69372 86468 69376 86524
rect 69376 86468 69432 86524
rect 69432 86468 69436 86524
rect 69372 86464 69436 86468
rect 69452 86524 69516 86528
rect 69452 86468 69456 86524
rect 69456 86468 69512 86524
rect 69512 86468 69516 86524
rect 69452 86464 69516 86468
rect 70812 86524 70876 86528
rect 70812 86468 70816 86524
rect 70816 86468 70872 86524
rect 70872 86468 70876 86524
rect 70812 86464 70876 86468
rect 70892 86524 70956 86528
rect 70892 86468 70896 86524
rect 70896 86468 70952 86524
rect 70952 86468 70956 86524
rect 70892 86464 70956 86468
rect 70972 86524 71036 86528
rect 70972 86468 70976 86524
rect 70976 86468 71032 86524
rect 71032 86468 71036 86524
rect 70972 86464 71036 86468
rect 71052 86524 71116 86528
rect 71052 86468 71056 86524
rect 71056 86468 71112 86524
rect 71112 86468 71116 86524
rect 71052 86464 71116 86468
rect 72412 86524 72476 86528
rect 72412 86468 72416 86524
rect 72416 86468 72472 86524
rect 72472 86468 72476 86524
rect 72412 86464 72476 86468
rect 72492 86524 72556 86528
rect 72492 86468 72496 86524
rect 72496 86468 72552 86524
rect 72552 86468 72556 86524
rect 72492 86464 72556 86468
rect 72572 86524 72636 86528
rect 72572 86468 72576 86524
rect 72576 86468 72632 86524
rect 72632 86468 72636 86524
rect 72572 86464 72636 86468
rect 72652 86524 72716 86528
rect 72652 86468 72656 86524
rect 72656 86468 72712 86524
rect 72712 86468 72716 86524
rect 72652 86464 72716 86468
rect 74012 86524 74076 86528
rect 74012 86468 74016 86524
rect 74016 86468 74072 86524
rect 74072 86468 74076 86524
rect 74012 86464 74076 86468
rect 74092 86524 74156 86528
rect 74092 86468 74096 86524
rect 74096 86468 74152 86524
rect 74152 86468 74156 86524
rect 74092 86464 74156 86468
rect 74172 86524 74236 86528
rect 74172 86468 74176 86524
rect 74176 86468 74232 86524
rect 74232 86468 74236 86524
rect 74172 86464 74236 86468
rect 74252 86524 74316 86528
rect 74252 86468 74256 86524
rect 74256 86468 74312 86524
rect 74312 86468 74316 86524
rect 74252 86464 74316 86468
rect 75612 86524 75676 86528
rect 75612 86468 75616 86524
rect 75616 86468 75672 86524
rect 75672 86468 75676 86524
rect 75612 86464 75676 86468
rect 75692 86524 75756 86528
rect 75692 86468 75696 86524
rect 75696 86468 75752 86524
rect 75752 86468 75756 86524
rect 75692 86464 75756 86468
rect 75772 86524 75836 86528
rect 75772 86468 75776 86524
rect 75776 86468 75832 86524
rect 75832 86468 75836 86524
rect 75772 86464 75836 86468
rect 75852 86524 75916 86528
rect 75852 86468 75856 86524
rect 75856 86468 75912 86524
rect 75912 86468 75916 86524
rect 75852 86464 75916 86468
rect 77212 86524 77276 86528
rect 77212 86468 77216 86524
rect 77216 86468 77272 86524
rect 77272 86468 77276 86524
rect 77212 86464 77276 86468
rect 77292 86524 77356 86528
rect 77292 86468 77296 86524
rect 77296 86468 77352 86524
rect 77352 86468 77356 86524
rect 77292 86464 77356 86468
rect 77372 86524 77436 86528
rect 77372 86468 77376 86524
rect 77376 86468 77432 86524
rect 77432 86468 77436 86524
rect 77372 86464 77436 86468
rect 77452 86524 77516 86528
rect 77452 86468 77456 86524
rect 77456 86468 77512 86524
rect 77512 86468 77516 86524
rect 77452 86464 77516 86468
rect 78812 86524 78876 86528
rect 78812 86468 78816 86524
rect 78816 86468 78872 86524
rect 78872 86468 78876 86524
rect 78812 86464 78876 86468
rect 78892 86524 78956 86528
rect 78892 86468 78896 86524
rect 78896 86468 78952 86524
rect 78952 86468 78956 86524
rect 78892 86464 78956 86468
rect 78972 86524 79036 86528
rect 78972 86468 78976 86524
rect 78976 86468 79032 86524
rect 79032 86468 79036 86524
rect 78972 86464 79036 86468
rect 79052 86524 79116 86528
rect 79052 86468 79056 86524
rect 79056 86468 79112 86524
rect 79112 86468 79116 86524
rect 79052 86464 79116 86468
rect 80412 86524 80476 86528
rect 80412 86468 80416 86524
rect 80416 86468 80472 86524
rect 80472 86468 80476 86524
rect 80412 86464 80476 86468
rect 80492 86524 80556 86528
rect 80492 86468 80496 86524
rect 80496 86468 80552 86524
rect 80552 86468 80556 86524
rect 80492 86464 80556 86468
rect 80572 86524 80636 86528
rect 80572 86468 80576 86524
rect 80576 86468 80632 86524
rect 80632 86468 80636 86524
rect 80572 86464 80636 86468
rect 80652 86524 80716 86528
rect 80652 86468 80656 86524
rect 80656 86468 80712 86524
rect 80712 86468 80716 86524
rect 80652 86464 80716 86468
rect 82012 86524 82076 86528
rect 82012 86468 82016 86524
rect 82016 86468 82072 86524
rect 82072 86468 82076 86524
rect 82012 86464 82076 86468
rect 82092 86524 82156 86528
rect 82092 86468 82096 86524
rect 82096 86468 82152 86524
rect 82152 86468 82156 86524
rect 82092 86464 82156 86468
rect 82172 86524 82236 86528
rect 82172 86468 82176 86524
rect 82176 86468 82232 86524
rect 82232 86468 82236 86524
rect 82172 86464 82236 86468
rect 82252 86524 82316 86528
rect 82252 86468 82256 86524
rect 82256 86468 82312 86524
rect 82312 86468 82316 86524
rect 82252 86464 82316 86468
rect 83612 86524 83676 86528
rect 83612 86468 83616 86524
rect 83616 86468 83672 86524
rect 83672 86468 83676 86524
rect 83612 86464 83676 86468
rect 83692 86524 83756 86528
rect 83692 86468 83696 86524
rect 83696 86468 83752 86524
rect 83752 86468 83756 86524
rect 83692 86464 83756 86468
rect 83772 86524 83836 86528
rect 83772 86468 83776 86524
rect 83776 86468 83832 86524
rect 83832 86468 83836 86524
rect 83772 86464 83836 86468
rect 83852 86524 83916 86528
rect 83852 86468 83856 86524
rect 83856 86468 83912 86524
rect 83912 86468 83916 86524
rect 83852 86464 83916 86468
rect 85212 86524 85276 86528
rect 85212 86468 85216 86524
rect 85216 86468 85272 86524
rect 85272 86468 85276 86524
rect 85212 86464 85276 86468
rect 85292 86524 85356 86528
rect 85292 86468 85296 86524
rect 85296 86468 85352 86524
rect 85352 86468 85356 86524
rect 85292 86464 85356 86468
rect 85372 86524 85436 86528
rect 85372 86468 85376 86524
rect 85376 86468 85432 86524
rect 85432 86468 85436 86524
rect 85372 86464 85436 86468
rect 85452 86524 85516 86528
rect 85452 86468 85456 86524
rect 85456 86468 85512 86524
rect 85512 86468 85516 86524
rect 85452 86464 85516 86468
rect 86812 86524 86876 86528
rect 86812 86468 86816 86524
rect 86816 86468 86872 86524
rect 86872 86468 86876 86524
rect 86812 86464 86876 86468
rect 86892 86524 86956 86528
rect 86892 86468 86896 86524
rect 86896 86468 86952 86524
rect 86952 86468 86956 86524
rect 86892 86464 86956 86468
rect 86972 86524 87036 86528
rect 86972 86468 86976 86524
rect 86976 86468 87032 86524
rect 87032 86468 87036 86524
rect 86972 86464 87036 86468
rect 87052 86524 87116 86528
rect 87052 86468 87056 86524
rect 87056 86468 87112 86524
rect 87112 86468 87116 86524
rect 87052 86464 87116 86468
rect 88412 86524 88476 86528
rect 88412 86468 88416 86524
rect 88416 86468 88472 86524
rect 88472 86468 88476 86524
rect 88412 86464 88476 86468
rect 88492 86524 88556 86528
rect 88492 86468 88496 86524
rect 88496 86468 88552 86524
rect 88552 86468 88556 86524
rect 88492 86464 88556 86468
rect 88572 86524 88636 86528
rect 88572 86468 88576 86524
rect 88576 86468 88632 86524
rect 88632 86468 88636 86524
rect 88572 86464 88636 86468
rect 88652 86524 88716 86528
rect 88652 86468 88656 86524
rect 88656 86468 88712 86524
rect 88712 86468 88716 86524
rect 88652 86464 88716 86468
rect 90012 86524 90076 86528
rect 90012 86468 90016 86524
rect 90016 86468 90072 86524
rect 90072 86468 90076 86524
rect 90012 86464 90076 86468
rect 90092 86524 90156 86528
rect 90092 86468 90096 86524
rect 90096 86468 90152 86524
rect 90152 86468 90156 86524
rect 90092 86464 90156 86468
rect 90172 86524 90236 86528
rect 90172 86468 90176 86524
rect 90176 86468 90232 86524
rect 90232 86468 90236 86524
rect 90172 86464 90236 86468
rect 90252 86524 90316 86528
rect 90252 86468 90256 86524
rect 90256 86468 90312 86524
rect 90312 86468 90316 86524
rect 90252 86464 90316 86468
rect 91612 86524 91676 86528
rect 91612 86468 91616 86524
rect 91616 86468 91672 86524
rect 91672 86468 91676 86524
rect 91612 86464 91676 86468
rect 91692 86524 91756 86528
rect 91692 86468 91696 86524
rect 91696 86468 91752 86524
rect 91752 86468 91756 86524
rect 91692 86464 91756 86468
rect 91772 86524 91836 86528
rect 91772 86468 91776 86524
rect 91776 86468 91832 86524
rect 91832 86468 91836 86524
rect 91772 86464 91836 86468
rect 91852 86524 91916 86528
rect 91852 86468 91856 86524
rect 91856 86468 91912 86524
rect 91912 86468 91916 86524
rect 91852 86464 91916 86468
rect 93212 86524 93276 86528
rect 93212 86468 93216 86524
rect 93216 86468 93272 86524
rect 93272 86468 93276 86524
rect 93212 86464 93276 86468
rect 93292 86524 93356 86528
rect 93292 86468 93296 86524
rect 93296 86468 93352 86524
rect 93352 86468 93356 86524
rect 93292 86464 93356 86468
rect 93372 86524 93436 86528
rect 93372 86468 93376 86524
rect 93376 86468 93432 86524
rect 93432 86468 93436 86524
rect 93372 86464 93436 86468
rect 93452 86524 93516 86528
rect 93452 86468 93456 86524
rect 93456 86468 93512 86524
rect 93512 86468 93516 86524
rect 93452 86464 93516 86468
rect 94812 86524 94876 86528
rect 94812 86468 94816 86524
rect 94816 86468 94872 86524
rect 94872 86468 94876 86524
rect 94812 86464 94876 86468
rect 94892 86524 94956 86528
rect 94892 86468 94896 86524
rect 94896 86468 94952 86524
rect 94952 86468 94956 86524
rect 94892 86464 94956 86468
rect 94972 86524 95036 86528
rect 94972 86468 94976 86524
rect 94976 86468 95032 86524
rect 95032 86468 95036 86524
rect 94972 86464 95036 86468
rect 95052 86524 95116 86528
rect 95052 86468 95056 86524
rect 95056 86468 95112 86524
rect 95112 86468 95116 86524
rect 95052 86464 95116 86468
rect 96412 86524 96476 86528
rect 96412 86468 96416 86524
rect 96416 86468 96472 86524
rect 96472 86468 96476 86524
rect 96412 86464 96476 86468
rect 96492 86524 96556 86528
rect 96492 86468 96496 86524
rect 96496 86468 96552 86524
rect 96552 86468 96556 86524
rect 96492 86464 96556 86468
rect 96572 86524 96636 86528
rect 96572 86468 96576 86524
rect 96576 86468 96632 86524
rect 96632 86468 96636 86524
rect 96572 86464 96636 86468
rect 96652 86524 96716 86528
rect 96652 86468 96656 86524
rect 96656 86468 96712 86524
rect 96712 86468 96716 86524
rect 96652 86464 96716 86468
rect 98012 86524 98076 86528
rect 98012 86468 98016 86524
rect 98016 86468 98072 86524
rect 98072 86468 98076 86524
rect 98012 86464 98076 86468
rect 98092 86524 98156 86528
rect 98092 86468 98096 86524
rect 98096 86468 98152 86524
rect 98152 86468 98156 86524
rect 98092 86464 98156 86468
rect 98172 86524 98236 86528
rect 98172 86468 98176 86524
rect 98176 86468 98232 86524
rect 98232 86468 98236 86524
rect 98172 86464 98236 86468
rect 98252 86524 98316 86528
rect 98252 86468 98256 86524
rect 98256 86468 98312 86524
rect 98312 86468 98316 86524
rect 98252 86464 98316 86468
rect 99612 86524 99676 86528
rect 99612 86468 99616 86524
rect 99616 86468 99672 86524
rect 99672 86468 99676 86524
rect 99612 86464 99676 86468
rect 99692 86524 99756 86528
rect 99692 86468 99696 86524
rect 99696 86468 99752 86524
rect 99752 86468 99756 86524
rect 99692 86464 99756 86468
rect 99772 86524 99836 86528
rect 99772 86468 99776 86524
rect 99776 86468 99832 86524
rect 99832 86468 99836 86524
rect 99772 86464 99836 86468
rect 99852 86524 99916 86528
rect 99852 86468 99856 86524
rect 99856 86468 99912 86524
rect 99912 86468 99916 86524
rect 99852 86464 99916 86468
rect 101212 86524 101276 86528
rect 101212 86468 101216 86524
rect 101216 86468 101272 86524
rect 101272 86468 101276 86524
rect 101212 86464 101276 86468
rect 101292 86524 101356 86528
rect 101292 86468 101296 86524
rect 101296 86468 101352 86524
rect 101352 86468 101356 86524
rect 101292 86464 101356 86468
rect 101372 86524 101436 86528
rect 101372 86468 101376 86524
rect 101376 86468 101432 86524
rect 101432 86468 101436 86524
rect 101372 86464 101436 86468
rect 101452 86524 101516 86528
rect 101452 86468 101456 86524
rect 101456 86468 101512 86524
rect 101512 86468 101516 86524
rect 101452 86464 101516 86468
rect 102812 86524 102876 86528
rect 102812 86468 102816 86524
rect 102816 86468 102872 86524
rect 102872 86468 102876 86524
rect 102812 86464 102876 86468
rect 102892 86524 102956 86528
rect 102892 86468 102896 86524
rect 102896 86468 102952 86524
rect 102952 86468 102956 86524
rect 102892 86464 102956 86468
rect 102972 86524 103036 86528
rect 102972 86468 102976 86524
rect 102976 86468 103032 86524
rect 103032 86468 103036 86524
rect 102972 86464 103036 86468
rect 103052 86524 103116 86528
rect 103052 86468 103056 86524
rect 103056 86468 103112 86524
rect 103112 86468 103116 86524
rect 103052 86464 103116 86468
rect 104412 86524 104476 86528
rect 104412 86468 104416 86524
rect 104416 86468 104472 86524
rect 104472 86468 104476 86524
rect 104412 86464 104476 86468
rect 104492 86524 104556 86528
rect 104492 86468 104496 86524
rect 104496 86468 104552 86524
rect 104552 86468 104556 86524
rect 104492 86464 104556 86468
rect 104572 86524 104636 86528
rect 104572 86468 104576 86524
rect 104576 86468 104632 86524
rect 104632 86468 104636 86524
rect 104572 86464 104636 86468
rect 104652 86524 104716 86528
rect 104652 86468 104656 86524
rect 104656 86468 104712 86524
rect 104712 86468 104716 86524
rect 104652 86464 104716 86468
rect 106012 86524 106076 86528
rect 106012 86468 106016 86524
rect 106016 86468 106072 86524
rect 106072 86468 106076 86524
rect 106012 86464 106076 86468
rect 106092 86524 106156 86528
rect 106092 86468 106096 86524
rect 106096 86468 106152 86524
rect 106152 86468 106156 86524
rect 106092 86464 106156 86468
rect 106172 86524 106236 86528
rect 106172 86468 106176 86524
rect 106176 86468 106232 86524
rect 106232 86468 106236 86524
rect 106172 86464 106236 86468
rect 106252 86524 106316 86528
rect 106252 86468 106256 86524
rect 106256 86468 106312 86524
rect 106312 86468 106316 86524
rect 106252 86464 106316 86468
rect 107612 86524 107676 86528
rect 107612 86468 107616 86524
rect 107616 86468 107672 86524
rect 107672 86468 107676 86524
rect 107612 86464 107676 86468
rect 107692 86524 107756 86528
rect 107692 86468 107696 86524
rect 107696 86468 107752 86524
rect 107752 86468 107756 86524
rect 107692 86464 107756 86468
rect 107772 86524 107836 86528
rect 107772 86468 107776 86524
rect 107776 86468 107832 86524
rect 107832 86468 107836 86524
rect 107772 86464 107836 86468
rect 107852 86524 107916 86528
rect 107852 86468 107856 86524
rect 107856 86468 107912 86524
rect 107912 86468 107916 86524
rect 107852 86464 107916 86468
rect 11468 86124 11532 86188
rect 2952 85980 3016 85984
rect 2952 85924 2956 85980
rect 2956 85924 3012 85980
rect 3012 85924 3016 85980
rect 2952 85920 3016 85924
rect 3032 85980 3096 85984
rect 3032 85924 3036 85980
rect 3036 85924 3092 85980
rect 3092 85924 3096 85980
rect 3032 85920 3096 85924
rect 3112 85980 3176 85984
rect 3112 85924 3116 85980
rect 3116 85924 3172 85980
rect 3172 85924 3176 85980
rect 3112 85920 3176 85924
rect 3192 85980 3256 85984
rect 3192 85924 3196 85980
rect 3196 85924 3252 85980
rect 3252 85924 3256 85980
rect 3192 85920 3256 85924
rect 4552 85980 4616 85984
rect 4552 85924 4556 85980
rect 4556 85924 4612 85980
rect 4612 85924 4616 85980
rect 4552 85920 4616 85924
rect 4632 85980 4696 85984
rect 4632 85924 4636 85980
rect 4636 85924 4692 85980
rect 4692 85924 4696 85980
rect 4632 85920 4696 85924
rect 4712 85980 4776 85984
rect 4712 85924 4716 85980
rect 4716 85924 4772 85980
rect 4772 85924 4776 85980
rect 4712 85920 4776 85924
rect 4792 85980 4856 85984
rect 4792 85924 4796 85980
rect 4796 85924 4852 85980
rect 4852 85924 4856 85980
rect 4792 85920 4856 85924
rect 6152 85980 6216 85984
rect 6152 85924 6156 85980
rect 6156 85924 6212 85980
rect 6212 85924 6216 85980
rect 6152 85920 6216 85924
rect 6232 85980 6296 85984
rect 6232 85924 6236 85980
rect 6236 85924 6292 85980
rect 6292 85924 6296 85980
rect 6232 85920 6296 85924
rect 6312 85980 6376 85984
rect 6312 85924 6316 85980
rect 6316 85924 6372 85980
rect 6372 85924 6376 85980
rect 6312 85920 6376 85924
rect 6392 85980 6456 85984
rect 6392 85924 6396 85980
rect 6396 85924 6452 85980
rect 6452 85924 6456 85980
rect 6392 85920 6456 85924
rect 7752 85980 7816 85984
rect 7752 85924 7756 85980
rect 7756 85924 7812 85980
rect 7812 85924 7816 85980
rect 7752 85920 7816 85924
rect 7832 85980 7896 85984
rect 7832 85924 7836 85980
rect 7836 85924 7892 85980
rect 7892 85924 7896 85980
rect 7832 85920 7896 85924
rect 7912 85980 7976 85984
rect 7912 85924 7916 85980
rect 7916 85924 7972 85980
rect 7972 85924 7976 85980
rect 7912 85920 7976 85924
rect 7992 85980 8056 85984
rect 7992 85924 7996 85980
rect 7996 85924 8052 85980
rect 8052 85924 8056 85980
rect 7992 85920 8056 85924
rect 9352 85980 9416 85984
rect 9352 85924 9356 85980
rect 9356 85924 9412 85980
rect 9412 85924 9416 85980
rect 9352 85920 9416 85924
rect 9432 85980 9496 85984
rect 9432 85924 9436 85980
rect 9436 85924 9492 85980
rect 9492 85924 9496 85980
rect 9432 85920 9496 85924
rect 9512 85980 9576 85984
rect 9512 85924 9516 85980
rect 9516 85924 9572 85980
rect 9572 85924 9576 85980
rect 9512 85920 9576 85924
rect 9592 85980 9656 85984
rect 9592 85924 9596 85980
rect 9596 85924 9652 85980
rect 9652 85924 9656 85980
rect 9592 85920 9656 85924
rect 10952 85980 11016 85984
rect 10952 85924 10956 85980
rect 10956 85924 11012 85980
rect 11012 85924 11016 85980
rect 10952 85920 11016 85924
rect 11032 85980 11096 85984
rect 11032 85924 11036 85980
rect 11036 85924 11092 85980
rect 11092 85924 11096 85980
rect 11032 85920 11096 85924
rect 11112 85980 11176 85984
rect 11112 85924 11116 85980
rect 11116 85924 11172 85980
rect 11172 85924 11176 85980
rect 11112 85920 11176 85924
rect 11192 85980 11256 85984
rect 11192 85924 11196 85980
rect 11196 85924 11252 85980
rect 11252 85924 11256 85980
rect 11192 85920 11256 85924
rect 12552 85980 12616 85984
rect 12552 85924 12556 85980
rect 12556 85924 12612 85980
rect 12612 85924 12616 85980
rect 12552 85920 12616 85924
rect 12632 85980 12696 85984
rect 12632 85924 12636 85980
rect 12636 85924 12692 85980
rect 12692 85924 12696 85980
rect 12632 85920 12696 85924
rect 12712 85980 12776 85984
rect 12712 85924 12716 85980
rect 12716 85924 12772 85980
rect 12772 85924 12776 85980
rect 12712 85920 12776 85924
rect 12792 85980 12856 85984
rect 12792 85924 12796 85980
rect 12796 85924 12852 85980
rect 12852 85924 12856 85980
rect 12792 85920 12856 85924
rect 14152 85980 14216 85984
rect 14152 85924 14156 85980
rect 14156 85924 14212 85980
rect 14212 85924 14216 85980
rect 14152 85920 14216 85924
rect 14232 85980 14296 85984
rect 14232 85924 14236 85980
rect 14236 85924 14292 85980
rect 14292 85924 14296 85980
rect 14232 85920 14296 85924
rect 14312 85980 14376 85984
rect 14312 85924 14316 85980
rect 14316 85924 14372 85980
rect 14372 85924 14376 85980
rect 14312 85920 14376 85924
rect 14392 85980 14456 85984
rect 14392 85924 14396 85980
rect 14396 85924 14452 85980
rect 14452 85924 14456 85980
rect 14392 85920 14456 85924
rect 15752 85980 15816 85984
rect 15752 85924 15756 85980
rect 15756 85924 15812 85980
rect 15812 85924 15816 85980
rect 15752 85920 15816 85924
rect 15832 85980 15896 85984
rect 15832 85924 15836 85980
rect 15836 85924 15892 85980
rect 15892 85924 15896 85980
rect 15832 85920 15896 85924
rect 15912 85980 15976 85984
rect 15912 85924 15916 85980
rect 15916 85924 15972 85980
rect 15972 85924 15976 85980
rect 15912 85920 15976 85924
rect 15992 85980 16056 85984
rect 15992 85924 15996 85980
rect 15996 85924 16052 85980
rect 16052 85924 16056 85980
rect 15992 85920 16056 85924
rect 17352 85980 17416 85984
rect 17352 85924 17356 85980
rect 17356 85924 17412 85980
rect 17412 85924 17416 85980
rect 17352 85920 17416 85924
rect 17432 85980 17496 85984
rect 17432 85924 17436 85980
rect 17436 85924 17492 85980
rect 17492 85924 17496 85980
rect 17432 85920 17496 85924
rect 17512 85980 17576 85984
rect 17512 85924 17516 85980
rect 17516 85924 17572 85980
rect 17572 85924 17576 85980
rect 17512 85920 17576 85924
rect 17592 85980 17656 85984
rect 17592 85924 17596 85980
rect 17596 85924 17652 85980
rect 17652 85924 17656 85980
rect 17592 85920 17656 85924
rect 18952 85980 19016 85984
rect 18952 85924 18956 85980
rect 18956 85924 19012 85980
rect 19012 85924 19016 85980
rect 18952 85920 19016 85924
rect 19032 85980 19096 85984
rect 19032 85924 19036 85980
rect 19036 85924 19092 85980
rect 19092 85924 19096 85980
rect 19032 85920 19096 85924
rect 19112 85980 19176 85984
rect 19112 85924 19116 85980
rect 19116 85924 19172 85980
rect 19172 85924 19176 85980
rect 19112 85920 19176 85924
rect 19192 85980 19256 85984
rect 19192 85924 19196 85980
rect 19196 85924 19252 85980
rect 19252 85924 19256 85980
rect 19192 85920 19256 85924
rect 20552 85980 20616 85984
rect 20552 85924 20556 85980
rect 20556 85924 20612 85980
rect 20612 85924 20616 85980
rect 20552 85920 20616 85924
rect 20632 85980 20696 85984
rect 20632 85924 20636 85980
rect 20636 85924 20692 85980
rect 20692 85924 20696 85980
rect 20632 85920 20696 85924
rect 20712 85980 20776 85984
rect 20712 85924 20716 85980
rect 20716 85924 20772 85980
rect 20772 85924 20776 85980
rect 20712 85920 20776 85924
rect 20792 85980 20856 85984
rect 20792 85924 20796 85980
rect 20796 85924 20852 85980
rect 20852 85924 20856 85980
rect 20792 85920 20856 85924
rect 22152 85980 22216 85984
rect 22152 85924 22156 85980
rect 22156 85924 22212 85980
rect 22212 85924 22216 85980
rect 22152 85920 22216 85924
rect 22232 85980 22296 85984
rect 22232 85924 22236 85980
rect 22236 85924 22292 85980
rect 22292 85924 22296 85980
rect 22232 85920 22296 85924
rect 22312 85980 22376 85984
rect 22312 85924 22316 85980
rect 22316 85924 22372 85980
rect 22372 85924 22376 85980
rect 22312 85920 22376 85924
rect 22392 85980 22456 85984
rect 22392 85924 22396 85980
rect 22396 85924 22452 85980
rect 22452 85924 22456 85980
rect 22392 85920 22456 85924
rect 23752 85980 23816 85984
rect 23752 85924 23756 85980
rect 23756 85924 23812 85980
rect 23812 85924 23816 85980
rect 23752 85920 23816 85924
rect 23832 85980 23896 85984
rect 23832 85924 23836 85980
rect 23836 85924 23892 85980
rect 23892 85924 23896 85980
rect 23832 85920 23896 85924
rect 23912 85980 23976 85984
rect 23912 85924 23916 85980
rect 23916 85924 23972 85980
rect 23972 85924 23976 85980
rect 23912 85920 23976 85924
rect 23992 85980 24056 85984
rect 23992 85924 23996 85980
rect 23996 85924 24052 85980
rect 24052 85924 24056 85980
rect 23992 85920 24056 85924
rect 25352 85980 25416 85984
rect 25352 85924 25356 85980
rect 25356 85924 25412 85980
rect 25412 85924 25416 85980
rect 25352 85920 25416 85924
rect 25432 85980 25496 85984
rect 25432 85924 25436 85980
rect 25436 85924 25492 85980
rect 25492 85924 25496 85980
rect 25432 85920 25496 85924
rect 25512 85980 25576 85984
rect 25512 85924 25516 85980
rect 25516 85924 25572 85980
rect 25572 85924 25576 85980
rect 25512 85920 25576 85924
rect 25592 85980 25656 85984
rect 25592 85924 25596 85980
rect 25596 85924 25652 85980
rect 25652 85924 25656 85980
rect 25592 85920 25656 85924
rect 26952 85980 27016 85984
rect 26952 85924 26956 85980
rect 26956 85924 27012 85980
rect 27012 85924 27016 85980
rect 26952 85920 27016 85924
rect 27032 85980 27096 85984
rect 27032 85924 27036 85980
rect 27036 85924 27092 85980
rect 27092 85924 27096 85980
rect 27032 85920 27096 85924
rect 27112 85980 27176 85984
rect 27112 85924 27116 85980
rect 27116 85924 27172 85980
rect 27172 85924 27176 85980
rect 27112 85920 27176 85924
rect 27192 85980 27256 85984
rect 27192 85924 27196 85980
rect 27196 85924 27252 85980
rect 27252 85924 27256 85980
rect 27192 85920 27256 85924
rect 28552 85980 28616 85984
rect 28552 85924 28556 85980
rect 28556 85924 28612 85980
rect 28612 85924 28616 85980
rect 28552 85920 28616 85924
rect 28632 85980 28696 85984
rect 28632 85924 28636 85980
rect 28636 85924 28692 85980
rect 28692 85924 28696 85980
rect 28632 85920 28696 85924
rect 28712 85980 28776 85984
rect 28712 85924 28716 85980
rect 28716 85924 28772 85980
rect 28772 85924 28776 85980
rect 28712 85920 28776 85924
rect 28792 85980 28856 85984
rect 28792 85924 28796 85980
rect 28796 85924 28852 85980
rect 28852 85924 28856 85980
rect 28792 85920 28856 85924
rect 30152 85980 30216 85984
rect 30152 85924 30156 85980
rect 30156 85924 30212 85980
rect 30212 85924 30216 85980
rect 30152 85920 30216 85924
rect 30232 85980 30296 85984
rect 30232 85924 30236 85980
rect 30236 85924 30292 85980
rect 30292 85924 30296 85980
rect 30232 85920 30296 85924
rect 30312 85980 30376 85984
rect 30312 85924 30316 85980
rect 30316 85924 30372 85980
rect 30372 85924 30376 85980
rect 30312 85920 30376 85924
rect 30392 85980 30456 85984
rect 30392 85924 30396 85980
rect 30396 85924 30452 85980
rect 30452 85924 30456 85980
rect 30392 85920 30456 85924
rect 31752 85980 31816 85984
rect 31752 85924 31756 85980
rect 31756 85924 31812 85980
rect 31812 85924 31816 85980
rect 31752 85920 31816 85924
rect 31832 85980 31896 85984
rect 31832 85924 31836 85980
rect 31836 85924 31892 85980
rect 31892 85924 31896 85980
rect 31832 85920 31896 85924
rect 31912 85980 31976 85984
rect 31912 85924 31916 85980
rect 31916 85924 31972 85980
rect 31972 85924 31976 85980
rect 31912 85920 31976 85924
rect 31992 85980 32056 85984
rect 31992 85924 31996 85980
rect 31996 85924 32052 85980
rect 32052 85924 32056 85980
rect 31992 85920 32056 85924
rect 33352 85980 33416 85984
rect 33352 85924 33356 85980
rect 33356 85924 33412 85980
rect 33412 85924 33416 85980
rect 33352 85920 33416 85924
rect 33432 85980 33496 85984
rect 33432 85924 33436 85980
rect 33436 85924 33492 85980
rect 33492 85924 33496 85980
rect 33432 85920 33496 85924
rect 33512 85980 33576 85984
rect 33512 85924 33516 85980
rect 33516 85924 33572 85980
rect 33572 85924 33576 85980
rect 33512 85920 33576 85924
rect 33592 85980 33656 85984
rect 33592 85924 33596 85980
rect 33596 85924 33652 85980
rect 33652 85924 33656 85980
rect 33592 85920 33656 85924
rect 34952 85980 35016 85984
rect 34952 85924 34956 85980
rect 34956 85924 35012 85980
rect 35012 85924 35016 85980
rect 34952 85920 35016 85924
rect 35032 85980 35096 85984
rect 35032 85924 35036 85980
rect 35036 85924 35092 85980
rect 35092 85924 35096 85980
rect 35032 85920 35096 85924
rect 35112 85980 35176 85984
rect 35112 85924 35116 85980
rect 35116 85924 35172 85980
rect 35172 85924 35176 85980
rect 35112 85920 35176 85924
rect 35192 85980 35256 85984
rect 35192 85924 35196 85980
rect 35196 85924 35252 85980
rect 35252 85924 35256 85980
rect 35192 85920 35256 85924
rect 36552 85980 36616 85984
rect 36552 85924 36556 85980
rect 36556 85924 36612 85980
rect 36612 85924 36616 85980
rect 36552 85920 36616 85924
rect 36632 85980 36696 85984
rect 36632 85924 36636 85980
rect 36636 85924 36692 85980
rect 36692 85924 36696 85980
rect 36632 85920 36696 85924
rect 36712 85980 36776 85984
rect 36712 85924 36716 85980
rect 36716 85924 36772 85980
rect 36772 85924 36776 85980
rect 36712 85920 36776 85924
rect 36792 85980 36856 85984
rect 36792 85924 36796 85980
rect 36796 85924 36852 85980
rect 36852 85924 36856 85980
rect 36792 85920 36856 85924
rect 38152 85980 38216 85984
rect 38152 85924 38156 85980
rect 38156 85924 38212 85980
rect 38212 85924 38216 85980
rect 38152 85920 38216 85924
rect 38232 85980 38296 85984
rect 38232 85924 38236 85980
rect 38236 85924 38292 85980
rect 38292 85924 38296 85980
rect 38232 85920 38296 85924
rect 38312 85980 38376 85984
rect 38312 85924 38316 85980
rect 38316 85924 38372 85980
rect 38372 85924 38376 85980
rect 38312 85920 38376 85924
rect 38392 85980 38456 85984
rect 38392 85924 38396 85980
rect 38396 85924 38452 85980
rect 38452 85924 38456 85980
rect 38392 85920 38456 85924
rect 39752 85980 39816 85984
rect 39752 85924 39756 85980
rect 39756 85924 39812 85980
rect 39812 85924 39816 85980
rect 39752 85920 39816 85924
rect 39832 85980 39896 85984
rect 39832 85924 39836 85980
rect 39836 85924 39892 85980
rect 39892 85924 39896 85980
rect 39832 85920 39896 85924
rect 39912 85980 39976 85984
rect 39912 85924 39916 85980
rect 39916 85924 39972 85980
rect 39972 85924 39976 85980
rect 39912 85920 39976 85924
rect 39992 85980 40056 85984
rect 39992 85924 39996 85980
rect 39996 85924 40052 85980
rect 40052 85924 40056 85980
rect 39992 85920 40056 85924
rect 41352 85980 41416 85984
rect 41352 85924 41356 85980
rect 41356 85924 41412 85980
rect 41412 85924 41416 85980
rect 41352 85920 41416 85924
rect 41432 85980 41496 85984
rect 41432 85924 41436 85980
rect 41436 85924 41492 85980
rect 41492 85924 41496 85980
rect 41432 85920 41496 85924
rect 41512 85980 41576 85984
rect 41512 85924 41516 85980
rect 41516 85924 41572 85980
rect 41572 85924 41576 85980
rect 41512 85920 41576 85924
rect 41592 85980 41656 85984
rect 41592 85924 41596 85980
rect 41596 85924 41652 85980
rect 41652 85924 41656 85980
rect 41592 85920 41656 85924
rect 42952 85980 43016 85984
rect 42952 85924 42956 85980
rect 42956 85924 43012 85980
rect 43012 85924 43016 85980
rect 42952 85920 43016 85924
rect 43032 85980 43096 85984
rect 43032 85924 43036 85980
rect 43036 85924 43092 85980
rect 43092 85924 43096 85980
rect 43032 85920 43096 85924
rect 43112 85980 43176 85984
rect 43112 85924 43116 85980
rect 43116 85924 43172 85980
rect 43172 85924 43176 85980
rect 43112 85920 43176 85924
rect 43192 85980 43256 85984
rect 43192 85924 43196 85980
rect 43196 85924 43252 85980
rect 43252 85924 43256 85980
rect 43192 85920 43256 85924
rect 44552 85980 44616 85984
rect 44552 85924 44556 85980
rect 44556 85924 44612 85980
rect 44612 85924 44616 85980
rect 44552 85920 44616 85924
rect 44632 85980 44696 85984
rect 44632 85924 44636 85980
rect 44636 85924 44692 85980
rect 44692 85924 44696 85980
rect 44632 85920 44696 85924
rect 44712 85980 44776 85984
rect 44712 85924 44716 85980
rect 44716 85924 44772 85980
rect 44772 85924 44776 85980
rect 44712 85920 44776 85924
rect 44792 85980 44856 85984
rect 44792 85924 44796 85980
rect 44796 85924 44852 85980
rect 44852 85924 44856 85980
rect 44792 85920 44856 85924
rect 46152 85980 46216 85984
rect 46152 85924 46156 85980
rect 46156 85924 46212 85980
rect 46212 85924 46216 85980
rect 46152 85920 46216 85924
rect 46232 85980 46296 85984
rect 46232 85924 46236 85980
rect 46236 85924 46292 85980
rect 46292 85924 46296 85980
rect 46232 85920 46296 85924
rect 46312 85980 46376 85984
rect 46312 85924 46316 85980
rect 46316 85924 46372 85980
rect 46372 85924 46376 85980
rect 46312 85920 46376 85924
rect 46392 85980 46456 85984
rect 46392 85924 46396 85980
rect 46396 85924 46452 85980
rect 46452 85924 46456 85980
rect 46392 85920 46456 85924
rect 47752 85980 47816 85984
rect 47752 85924 47756 85980
rect 47756 85924 47812 85980
rect 47812 85924 47816 85980
rect 47752 85920 47816 85924
rect 47832 85980 47896 85984
rect 47832 85924 47836 85980
rect 47836 85924 47892 85980
rect 47892 85924 47896 85980
rect 47832 85920 47896 85924
rect 47912 85980 47976 85984
rect 47912 85924 47916 85980
rect 47916 85924 47972 85980
rect 47972 85924 47976 85980
rect 47912 85920 47976 85924
rect 47992 85980 48056 85984
rect 47992 85924 47996 85980
rect 47996 85924 48052 85980
rect 48052 85924 48056 85980
rect 47992 85920 48056 85924
rect 49352 85980 49416 85984
rect 49352 85924 49356 85980
rect 49356 85924 49412 85980
rect 49412 85924 49416 85980
rect 49352 85920 49416 85924
rect 49432 85980 49496 85984
rect 49432 85924 49436 85980
rect 49436 85924 49492 85980
rect 49492 85924 49496 85980
rect 49432 85920 49496 85924
rect 49512 85980 49576 85984
rect 49512 85924 49516 85980
rect 49516 85924 49572 85980
rect 49572 85924 49576 85980
rect 49512 85920 49576 85924
rect 49592 85980 49656 85984
rect 49592 85924 49596 85980
rect 49596 85924 49652 85980
rect 49652 85924 49656 85980
rect 49592 85920 49656 85924
rect 50952 85980 51016 85984
rect 50952 85924 50956 85980
rect 50956 85924 51012 85980
rect 51012 85924 51016 85980
rect 50952 85920 51016 85924
rect 51032 85980 51096 85984
rect 51032 85924 51036 85980
rect 51036 85924 51092 85980
rect 51092 85924 51096 85980
rect 51032 85920 51096 85924
rect 51112 85980 51176 85984
rect 51112 85924 51116 85980
rect 51116 85924 51172 85980
rect 51172 85924 51176 85980
rect 51112 85920 51176 85924
rect 51192 85980 51256 85984
rect 51192 85924 51196 85980
rect 51196 85924 51252 85980
rect 51252 85924 51256 85980
rect 51192 85920 51256 85924
rect 52552 85980 52616 85984
rect 52552 85924 52556 85980
rect 52556 85924 52612 85980
rect 52612 85924 52616 85980
rect 52552 85920 52616 85924
rect 52632 85980 52696 85984
rect 52632 85924 52636 85980
rect 52636 85924 52692 85980
rect 52692 85924 52696 85980
rect 52632 85920 52696 85924
rect 52712 85980 52776 85984
rect 52712 85924 52716 85980
rect 52716 85924 52772 85980
rect 52772 85924 52776 85980
rect 52712 85920 52776 85924
rect 52792 85980 52856 85984
rect 52792 85924 52796 85980
rect 52796 85924 52852 85980
rect 52852 85924 52856 85980
rect 52792 85920 52856 85924
rect 54152 85980 54216 85984
rect 54152 85924 54156 85980
rect 54156 85924 54212 85980
rect 54212 85924 54216 85980
rect 54152 85920 54216 85924
rect 54232 85980 54296 85984
rect 54232 85924 54236 85980
rect 54236 85924 54292 85980
rect 54292 85924 54296 85980
rect 54232 85920 54296 85924
rect 54312 85980 54376 85984
rect 54312 85924 54316 85980
rect 54316 85924 54372 85980
rect 54372 85924 54376 85980
rect 54312 85920 54376 85924
rect 54392 85980 54456 85984
rect 54392 85924 54396 85980
rect 54396 85924 54452 85980
rect 54452 85924 54456 85980
rect 54392 85920 54456 85924
rect 55752 85980 55816 85984
rect 55752 85924 55756 85980
rect 55756 85924 55812 85980
rect 55812 85924 55816 85980
rect 55752 85920 55816 85924
rect 55832 85980 55896 85984
rect 55832 85924 55836 85980
rect 55836 85924 55892 85980
rect 55892 85924 55896 85980
rect 55832 85920 55896 85924
rect 55912 85980 55976 85984
rect 55912 85924 55916 85980
rect 55916 85924 55972 85980
rect 55972 85924 55976 85980
rect 55912 85920 55976 85924
rect 55992 85980 56056 85984
rect 55992 85924 55996 85980
rect 55996 85924 56052 85980
rect 56052 85924 56056 85980
rect 55992 85920 56056 85924
rect 57352 85980 57416 85984
rect 57352 85924 57356 85980
rect 57356 85924 57412 85980
rect 57412 85924 57416 85980
rect 57352 85920 57416 85924
rect 57432 85980 57496 85984
rect 57432 85924 57436 85980
rect 57436 85924 57492 85980
rect 57492 85924 57496 85980
rect 57432 85920 57496 85924
rect 57512 85980 57576 85984
rect 57512 85924 57516 85980
rect 57516 85924 57572 85980
rect 57572 85924 57576 85980
rect 57512 85920 57576 85924
rect 57592 85980 57656 85984
rect 57592 85924 57596 85980
rect 57596 85924 57652 85980
rect 57652 85924 57656 85980
rect 57592 85920 57656 85924
rect 58952 85980 59016 85984
rect 58952 85924 58956 85980
rect 58956 85924 59012 85980
rect 59012 85924 59016 85980
rect 58952 85920 59016 85924
rect 59032 85980 59096 85984
rect 59032 85924 59036 85980
rect 59036 85924 59092 85980
rect 59092 85924 59096 85980
rect 59032 85920 59096 85924
rect 59112 85980 59176 85984
rect 59112 85924 59116 85980
rect 59116 85924 59172 85980
rect 59172 85924 59176 85980
rect 59112 85920 59176 85924
rect 59192 85980 59256 85984
rect 59192 85924 59196 85980
rect 59196 85924 59252 85980
rect 59252 85924 59256 85980
rect 59192 85920 59256 85924
rect 60552 85980 60616 85984
rect 60552 85924 60556 85980
rect 60556 85924 60612 85980
rect 60612 85924 60616 85980
rect 60552 85920 60616 85924
rect 60632 85980 60696 85984
rect 60632 85924 60636 85980
rect 60636 85924 60692 85980
rect 60692 85924 60696 85980
rect 60632 85920 60696 85924
rect 60712 85980 60776 85984
rect 60712 85924 60716 85980
rect 60716 85924 60772 85980
rect 60772 85924 60776 85980
rect 60712 85920 60776 85924
rect 60792 85980 60856 85984
rect 60792 85924 60796 85980
rect 60796 85924 60852 85980
rect 60852 85924 60856 85980
rect 60792 85920 60856 85924
rect 62152 85980 62216 85984
rect 62152 85924 62156 85980
rect 62156 85924 62212 85980
rect 62212 85924 62216 85980
rect 62152 85920 62216 85924
rect 62232 85980 62296 85984
rect 62232 85924 62236 85980
rect 62236 85924 62292 85980
rect 62292 85924 62296 85980
rect 62232 85920 62296 85924
rect 62312 85980 62376 85984
rect 62312 85924 62316 85980
rect 62316 85924 62372 85980
rect 62372 85924 62376 85980
rect 62312 85920 62376 85924
rect 62392 85980 62456 85984
rect 62392 85924 62396 85980
rect 62396 85924 62452 85980
rect 62452 85924 62456 85980
rect 62392 85920 62456 85924
rect 63752 85980 63816 85984
rect 63752 85924 63756 85980
rect 63756 85924 63812 85980
rect 63812 85924 63816 85980
rect 63752 85920 63816 85924
rect 63832 85980 63896 85984
rect 63832 85924 63836 85980
rect 63836 85924 63892 85980
rect 63892 85924 63896 85980
rect 63832 85920 63896 85924
rect 63912 85980 63976 85984
rect 63912 85924 63916 85980
rect 63916 85924 63972 85980
rect 63972 85924 63976 85980
rect 63912 85920 63976 85924
rect 63992 85980 64056 85984
rect 63992 85924 63996 85980
rect 63996 85924 64052 85980
rect 64052 85924 64056 85980
rect 63992 85920 64056 85924
rect 65352 85980 65416 85984
rect 65352 85924 65356 85980
rect 65356 85924 65412 85980
rect 65412 85924 65416 85980
rect 65352 85920 65416 85924
rect 65432 85980 65496 85984
rect 65432 85924 65436 85980
rect 65436 85924 65492 85980
rect 65492 85924 65496 85980
rect 65432 85920 65496 85924
rect 65512 85980 65576 85984
rect 65512 85924 65516 85980
rect 65516 85924 65572 85980
rect 65572 85924 65576 85980
rect 65512 85920 65576 85924
rect 65592 85980 65656 85984
rect 65592 85924 65596 85980
rect 65596 85924 65652 85980
rect 65652 85924 65656 85980
rect 65592 85920 65656 85924
rect 66952 85980 67016 85984
rect 66952 85924 66956 85980
rect 66956 85924 67012 85980
rect 67012 85924 67016 85980
rect 66952 85920 67016 85924
rect 67032 85980 67096 85984
rect 67032 85924 67036 85980
rect 67036 85924 67092 85980
rect 67092 85924 67096 85980
rect 67032 85920 67096 85924
rect 67112 85980 67176 85984
rect 67112 85924 67116 85980
rect 67116 85924 67172 85980
rect 67172 85924 67176 85980
rect 67112 85920 67176 85924
rect 67192 85980 67256 85984
rect 67192 85924 67196 85980
rect 67196 85924 67252 85980
rect 67252 85924 67256 85980
rect 67192 85920 67256 85924
rect 68552 85980 68616 85984
rect 68552 85924 68556 85980
rect 68556 85924 68612 85980
rect 68612 85924 68616 85980
rect 68552 85920 68616 85924
rect 68632 85980 68696 85984
rect 68632 85924 68636 85980
rect 68636 85924 68692 85980
rect 68692 85924 68696 85980
rect 68632 85920 68696 85924
rect 68712 85980 68776 85984
rect 68712 85924 68716 85980
rect 68716 85924 68772 85980
rect 68772 85924 68776 85980
rect 68712 85920 68776 85924
rect 68792 85980 68856 85984
rect 68792 85924 68796 85980
rect 68796 85924 68852 85980
rect 68852 85924 68856 85980
rect 68792 85920 68856 85924
rect 70152 85980 70216 85984
rect 70152 85924 70156 85980
rect 70156 85924 70212 85980
rect 70212 85924 70216 85980
rect 70152 85920 70216 85924
rect 70232 85980 70296 85984
rect 70232 85924 70236 85980
rect 70236 85924 70292 85980
rect 70292 85924 70296 85980
rect 70232 85920 70296 85924
rect 70312 85980 70376 85984
rect 70312 85924 70316 85980
rect 70316 85924 70372 85980
rect 70372 85924 70376 85980
rect 70312 85920 70376 85924
rect 70392 85980 70456 85984
rect 70392 85924 70396 85980
rect 70396 85924 70452 85980
rect 70452 85924 70456 85980
rect 70392 85920 70456 85924
rect 71752 85980 71816 85984
rect 71752 85924 71756 85980
rect 71756 85924 71812 85980
rect 71812 85924 71816 85980
rect 71752 85920 71816 85924
rect 71832 85980 71896 85984
rect 71832 85924 71836 85980
rect 71836 85924 71892 85980
rect 71892 85924 71896 85980
rect 71832 85920 71896 85924
rect 71912 85980 71976 85984
rect 71912 85924 71916 85980
rect 71916 85924 71972 85980
rect 71972 85924 71976 85980
rect 71912 85920 71976 85924
rect 71992 85980 72056 85984
rect 71992 85924 71996 85980
rect 71996 85924 72052 85980
rect 72052 85924 72056 85980
rect 71992 85920 72056 85924
rect 73352 85980 73416 85984
rect 73352 85924 73356 85980
rect 73356 85924 73412 85980
rect 73412 85924 73416 85980
rect 73352 85920 73416 85924
rect 73432 85980 73496 85984
rect 73432 85924 73436 85980
rect 73436 85924 73492 85980
rect 73492 85924 73496 85980
rect 73432 85920 73496 85924
rect 73512 85980 73576 85984
rect 73512 85924 73516 85980
rect 73516 85924 73572 85980
rect 73572 85924 73576 85980
rect 73512 85920 73576 85924
rect 73592 85980 73656 85984
rect 73592 85924 73596 85980
rect 73596 85924 73652 85980
rect 73652 85924 73656 85980
rect 73592 85920 73656 85924
rect 74952 85980 75016 85984
rect 74952 85924 74956 85980
rect 74956 85924 75012 85980
rect 75012 85924 75016 85980
rect 74952 85920 75016 85924
rect 75032 85980 75096 85984
rect 75032 85924 75036 85980
rect 75036 85924 75092 85980
rect 75092 85924 75096 85980
rect 75032 85920 75096 85924
rect 75112 85980 75176 85984
rect 75112 85924 75116 85980
rect 75116 85924 75172 85980
rect 75172 85924 75176 85980
rect 75112 85920 75176 85924
rect 75192 85980 75256 85984
rect 75192 85924 75196 85980
rect 75196 85924 75252 85980
rect 75252 85924 75256 85980
rect 75192 85920 75256 85924
rect 76552 85980 76616 85984
rect 76552 85924 76556 85980
rect 76556 85924 76612 85980
rect 76612 85924 76616 85980
rect 76552 85920 76616 85924
rect 76632 85980 76696 85984
rect 76632 85924 76636 85980
rect 76636 85924 76692 85980
rect 76692 85924 76696 85980
rect 76632 85920 76696 85924
rect 76712 85980 76776 85984
rect 76712 85924 76716 85980
rect 76716 85924 76772 85980
rect 76772 85924 76776 85980
rect 76712 85920 76776 85924
rect 76792 85980 76856 85984
rect 76792 85924 76796 85980
rect 76796 85924 76852 85980
rect 76852 85924 76856 85980
rect 76792 85920 76856 85924
rect 78152 85980 78216 85984
rect 78152 85924 78156 85980
rect 78156 85924 78212 85980
rect 78212 85924 78216 85980
rect 78152 85920 78216 85924
rect 78232 85980 78296 85984
rect 78232 85924 78236 85980
rect 78236 85924 78292 85980
rect 78292 85924 78296 85980
rect 78232 85920 78296 85924
rect 78312 85980 78376 85984
rect 78312 85924 78316 85980
rect 78316 85924 78372 85980
rect 78372 85924 78376 85980
rect 78312 85920 78376 85924
rect 78392 85980 78456 85984
rect 78392 85924 78396 85980
rect 78396 85924 78452 85980
rect 78452 85924 78456 85980
rect 78392 85920 78456 85924
rect 79752 85980 79816 85984
rect 79752 85924 79756 85980
rect 79756 85924 79812 85980
rect 79812 85924 79816 85980
rect 79752 85920 79816 85924
rect 79832 85980 79896 85984
rect 79832 85924 79836 85980
rect 79836 85924 79892 85980
rect 79892 85924 79896 85980
rect 79832 85920 79896 85924
rect 79912 85980 79976 85984
rect 79912 85924 79916 85980
rect 79916 85924 79972 85980
rect 79972 85924 79976 85980
rect 79912 85920 79976 85924
rect 79992 85980 80056 85984
rect 79992 85924 79996 85980
rect 79996 85924 80052 85980
rect 80052 85924 80056 85980
rect 79992 85920 80056 85924
rect 81352 85980 81416 85984
rect 81352 85924 81356 85980
rect 81356 85924 81412 85980
rect 81412 85924 81416 85980
rect 81352 85920 81416 85924
rect 81432 85980 81496 85984
rect 81432 85924 81436 85980
rect 81436 85924 81492 85980
rect 81492 85924 81496 85980
rect 81432 85920 81496 85924
rect 81512 85980 81576 85984
rect 81512 85924 81516 85980
rect 81516 85924 81572 85980
rect 81572 85924 81576 85980
rect 81512 85920 81576 85924
rect 81592 85980 81656 85984
rect 81592 85924 81596 85980
rect 81596 85924 81652 85980
rect 81652 85924 81656 85980
rect 81592 85920 81656 85924
rect 82952 85980 83016 85984
rect 82952 85924 82956 85980
rect 82956 85924 83012 85980
rect 83012 85924 83016 85980
rect 82952 85920 83016 85924
rect 83032 85980 83096 85984
rect 83032 85924 83036 85980
rect 83036 85924 83092 85980
rect 83092 85924 83096 85980
rect 83032 85920 83096 85924
rect 83112 85980 83176 85984
rect 83112 85924 83116 85980
rect 83116 85924 83172 85980
rect 83172 85924 83176 85980
rect 83112 85920 83176 85924
rect 83192 85980 83256 85984
rect 83192 85924 83196 85980
rect 83196 85924 83252 85980
rect 83252 85924 83256 85980
rect 83192 85920 83256 85924
rect 84552 85980 84616 85984
rect 84552 85924 84556 85980
rect 84556 85924 84612 85980
rect 84612 85924 84616 85980
rect 84552 85920 84616 85924
rect 84632 85980 84696 85984
rect 84632 85924 84636 85980
rect 84636 85924 84692 85980
rect 84692 85924 84696 85980
rect 84632 85920 84696 85924
rect 84712 85980 84776 85984
rect 84712 85924 84716 85980
rect 84716 85924 84772 85980
rect 84772 85924 84776 85980
rect 84712 85920 84776 85924
rect 84792 85980 84856 85984
rect 84792 85924 84796 85980
rect 84796 85924 84852 85980
rect 84852 85924 84856 85980
rect 84792 85920 84856 85924
rect 86152 85980 86216 85984
rect 86152 85924 86156 85980
rect 86156 85924 86212 85980
rect 86212 85924 86216 85980
rect 86152 85920 86216 85924
rect 86232 85980 86296 85984
rect 86232 85924 86236 85980
rect 86236 85924 86292 85980
rect 86292 85924 86296 85980
rect 86232 85920 86296 85924
rect 86312 85980 86376 85984
rect 86312 85924 86316 85980
rect 86316 85924 86372 85980
rect 86372 85924 86376 85980
rect 86312 85920 86376 85924
rect 86392 85980 86456 85984
rect 86392 85924 86396 85980
rect 86396 85924 86452 85980
rect 86452 85924 86456 85980
rect 86392 85920 86456 85924
rect 87752 85980 87816 85984
rect 87752 85924 87756 85980
rect 87756 85924 87812 85980
rect 87812 85924 87816 85980
rect 87752 85920 87816 85924
rect 87832 85980 87896 85984
rect 87832 85924 87836 85980
rect 87836 85924 87892 85980
rect 87892 85924 87896 85980
rect 87832 85920 87896 85924
rect 87912 85980 87976 85984
rect 87912 85924 87916 85980
rect 87916 85924 87972 85980
rect 87972 85924 87976 85980
rect 87912 85920 87976 85924
rect 87992 85980 88056 85984
rect 87992 85924 87996 85980
rect 87996 85924 88052 85980
rect 88052 85924 88056 85980
rect 87992 85920 88056 85924
rect 89352 85980 89416 85984
rect 89352 85924 89356 85980
rect 89356 85924 89412 85980
rect 89412 85924 89416 85980
rect 89352 85920 89416 85924
rect 89432 85980 89496 85984
rect 89432 85924 89436 85980
rect 89436 85924 89492 85980
rect 89492 85924 89496 85980
rect 89432 85920 89496 85924
rect 89512 85980 89576 85984
rect 89512 85924 89516 85980
rect 89516 85924 89572 85980
rect 89572 85924 89576 85980
rect 89512 85920 89576 85924
rect 89592 85980 89656 85984
rect 89592 85924 89596 85980
rect 89596 85924 89652 85980
rect 89652 85924 89656 85980
rect 89592 85920 89656 85924
rect 90952 85980 91016 85984
rect 90952 85924 90956 85980
rect 90956 85924 91012 85980
rect 91012 85924 91016 85980
rect 90952 85920 91016 85924
rect 91032 85980 91096 85984
rect 91032 85924 91036 85980
rect 91036 85924 91092 85980
rect 91092 85924 91096 85980
rect 91032 85920 91096 85924
rect 91112 85980 91176 85984
rect 91112 85924 91116 85980
rect 91116 85924 91172 85980
rect 91172 85924 91176 85980
rect 91112 85920 91176 85924
rect 91192 85980 91256 85984
rect 91192 85924 91196 85980
rect 91196 85924 91252 85980
rect 91252 85924 91256 85980
rect 91192 85920 91256 85924
rect 92552 85980 92616 85984
rect 92552 85924 92556 85980
rect 92556 85924 92612 85980
rect 92612 85924 92616 85980
rect 92552 85920 92616 85924
rect 92632 85980 92696 85984
rect 92632 85924 92636 85980
rect 92636 85924 92692 85980
rect 92692 85924 92696 85980
rect 92632 85920 92696 85924
rect 92712 85980 92776 85984
rect 92712 85924 92716 85980
rect 92716 85924 92772 85980
rect 92772 85924 92776 85980
rect 92712 85920 92776 85924
rect 92792 85980 92856 85984
rect 92792 85924 92796 85980
rect 92796 85924 92852 85980
rect 92852 85924 92856 85980
rect 92792 85920 92856 85924
rect 94152 85980 94216 85984
rect 94152 85924 94156 85980
rect 94156 85924 94212 85980
rect 94212 85924 94216 85980
rect 94152 85920 94216 85924
rect 94232 85980 94296 85984
rect 94232 85924 94236 85980
rect 94236 85924 94292 85980
rect 94292 85924 94296 85980
rect 94232 85920 94296 85924
rect 94312 85980 94376 85984
rect 94312 85924 94316 85980
rect 94316 85924 94372 85980
rect 94372 85924 94376 85980
rect 94312 85920 94376 85924
rect 94392 85980 94456 85984
rect 94392 85924 94396 85980
rect 94396 85924 94452 85980
rect 94452 85924 94456 85980
rect 94392 85920 94456 85924
rect 95752 85980 95816 85984
rect 95752 85924 95756 85980
rect 95756 85924 95812 85980
rect 95812 85924 95816 85980
rect 95752 85920 95816 85924
rect 95832 85980 95896 85984
rect 95832 85924 95836 85980
rect 95836 85924 95892 85980
rect 95892 85924 95896 85980
rect 95832 85920 95896 85924
rect 95912 85980 95976 85984
rect 95912 85924 95916 85980
rect 95916 85924 95972 85980
rect 95972 85924 95976 85980
rect 95912 85920 95976 85924
rect 95992 85980 96056 85984
rect 95992 85924 95996 85980
rect 95996 85924 96052 85980
rect 96052 85924 96056 85980
rect 95992 85920 96056 85924
rect 97352 85980 97416 85984
rect 97352 85924 97356 85980
rect 97356 85924 97412 85980
rect 97412 85924 97416 85980
rect 97352 85920 97416 85924
rect 97432 85980 97496 85984
rect 97432 85924 97436 85980
rect 97436 85924 97492 85980
rect 97492 85924 97496 85980
rect 97432 85920 97496 85924
rect 97512 85980 97576 85984
rect 97512 85924 97516 85980
rect 97516 85924 97572 85980
rect 97572 85924 97576 85980
rect 97512 85920 97576 85924
rect 97592 85980 97656 85984
rect 97592 85924 97596 85980
rect 97596 85924 97652 85980
rect 97652 85924 97656 85980
rect 97592 85920 97656 85924
rect 98952 85980 99016 85984
rect 98952 85924 98956 85980
rect 98956 85924 99012 85980
rect 99012 85924 99016 85980
rect 98952 85920 99016 85924
rect 99032 85980 99096 85984
rect 99032 85924 99036 85980
rect 99036 85924 99092 85980
rect 99092 85924 99096 85980
rect 99032 85920 99096 85924
rect 99112 85980 99176 85984
rect 99112 85924 99116 85980
rect 99116 85924 99172 85980
rect 99172 85924 99176 85980
rect 99112 85920 99176 85924
rect 99192 85980 99256 85984
rect 99192 85924 99196 85980
rect 99196 85924 99252 85980
rect 99252 85924 99256 85980
rect 99192 85920 99256 85924
rect 100552 85980 100616 85984
rect 100552 85924 100556 85980
rect 100556 85924 100612 85980
rect 100612 85924 100616 85980
rect 100552 85920 100616 85924
rect 100632 85980 100696 85984
rect 100632 85924 100636 85980
rect 100636 85924 100692 85980
rect 100692 85924 100696 85980
rect 100632 85920 100696 85924
rect 100712 85980 100776 85984
rect 100712 85924 100716 85980
rect 100716 85924 100772 85980
rect 100772 85924 100776 85980
rect 100712 85920 100776 85924
rect 100792 85980 100856 85984
rect 100792 85924 100796 85980
rect 100796 85924 100852 85980
rect 100852 85924 100856 85980
rect 100792 85920 100856 85924
rect 102152 85980 102216 85984
rect 102152 85924 102156 85980
rect 102156 85924 102212 85980
rect 102212 85924 102216 85980
rect 102152 85920 102216 85924
rect 102232 85980 102296 85984
rect 102232 85924 102236 85980
rect 102236 85924 102292 85980
rect 102292 85924 102296 85980
rect 102232 85920 102296 85924
rect 102312 85980 102376 85984
rect 102312 85924 102316 85980
rect 102316 85924 102372 85980
rect 102372 85924 102376 85980
rect 102312 85920 102376 85924
rect 102392 85980 102456 85984
rect 102392 85924 102396 85980
rect 102396 85924 102452 85980
rect 102452 85924 102456 85980
rect 102392 85920 102456 85924
rect 103752 85980 103816 85984
rect 103752 85924 103756 85980
rect 103756 85924 103812 85980
rect 103812 85924 103816 85980
rect 103752 85920 103816 85924
rect 103832 85980 103896 85984
rect 103832 85924 103836 85980
rect 103836 85924 103892 85980
rect 103892 85924 103896 85980
rect 103832 85920 103896 85924
rect 103912 85980 103976 85984
rect 103912 85924 103916 85980
rect 103916 85924 103972 85980
rect 103972 85924 103976 85980
rect 103912 85920 103976 85924
rect 103992 85980 104056 85984
rect 103992 85924 103996 85980
rect 103996 85924 104052 85980
rect 104052 85924 104056 85980
rect 103992 85920 104056 85924
rect 105352 85980 105416 85984
rect 105352 85924 105356 85980
rect 105356 85924 105412 85980
rect 105412 85924 105416 85980
rect 105352 85920 105416 85924
rect 105432 85980 105496 85984
rect 105432 85924 105436 85980
rect 105436 85924 105492 85980
rect 105492 85924 105496 85980
rect 105432 85920 105496 85924
rect 105512 85980 105576 85984
rect 105512 85924 105516 85980
rect 105516 85924 105572 85980
rect 105572 85924 105576 85980
rect 105512 85920 105576 85924
rect 105592 85980 105656 85984
rect 105592 85924 105596 85980
rect 105596 85924 105652 85980
rect 105652 85924 105656 85980
rect 105592 85920 105656 85924
rect 106952 85980 107016 85984
rect 106952 85924 106956 85980
rect 106956 85924 107012 85980
rect 107012 85924 107016 85980
rect 106952 85920 107016 85924
rect 107032 85980 107096 85984
rect 107032 85924 107036 85980
rect 107036 85924 107092 85980
rect 107092 85924 107096 85980
rect 107032 85920 107096 85924
rect 107112 85980 107176 85984
rect 107112 85924 107116 85980
rect 107116 85924 107172 85980
rect 107172 85924 107176 85980
rect 107112 85920 107176 85924
rect 107192 85980 107256 85984
rect 107192 85924 107196 85980
rect 107196 85924 107252 85980
rect 107252 85924 107256 85980
rect 107192 85920 107256 85924
rect 108552 85980 108616 85984
rect 108552 85924 108556 85980
rect 108556 85924 108612 85980
rect 108612 85924 108616 85980
rect 108552 85920 108616 85924
rect 108632 85980 108696 85984
rect 108632 85924 108636 85980
rect 108636 85924 108692 85980
rect 108692 85924 108696 85980
rect 108632 85920 108696 85924
rect 108712 85980 108776 85984
rect 108712 85924 108716 85980
rect 108716 85924 108772 85980
rect 108772 85924 108776 85980
rect 108712 85920 108776 85924
rect 108792 85980 108856 85984
rect 108792 85924 108796 85980
rect 108796 85924 108852 85980
rect 108852 85924 108856 85980
rect 108792 85920 108856 85924
rect 60964 85912 61028 85916
rect 60964 85856 61014 85912
rect 61014 85856 61028 85912
rect 60964 85852 61028 85856
rect 63540 85912 63604 85916
rect 63540 85856 63554 85912
rect 63554 85856 63604 85912
rect 63540 85852 63604 85856
rect 68140 85912 68204 85916
rect 68140 85856 68154 85912
rect 68154 85856 68204 85912
rect 68140 85852 68204 85856
rect 72188 85912 72252 85916
rect 72188 85856 72202 85912
rect 72202 85856 72252 85912
rect 72188 85852 72252 85856
rect 68324 85716 68388 85780
rect 40172 85580 40236 85644
rect 41828 85640 41892 85644
rect 41828 85584 41842 85640
rect 41842 85584 41892 85640
rect 41828 85580 41892 85584
rect 44036 85580 44100 85644
rect 46612 85640 46676 85644
rect 46612 85584 46626 85640
rect 46626 85584 46676 85640
rect 46612 85580 46676 85584
rect 47348 85640 47412 85644
rect 47348 85584 47362 85640
rect 47362 85584 47412 85640
rect 47348 85580 47412 85584
rect 49004 85580 49068 85644
rect 50476 85580 50540 85644
rect 55260 85640 55324 85644
rect 55260 85584 55274 85640
rect 55274 85584 55324 85640
rect 55260 85580 55324 85584
rect 56180 85580 56244 85644
rect 58756 85580 58820 85644
rect 62620 85580 62684 85644
rect 73844 85580 73908 85644
rect 76236 85580 76300 85644
rect 77708 85640 77772 85644
rect 77708 85584 77722 85640
rect 77722 85584 77772 85640
rect 77708 85580 77772 85584
rect 101996 85580 102060 85644
rect 75316 85444 75380 85508
rect 91508 85444 91572 85508
rect 3612 85436 3676 85440
rect 3612 85380 3616 85436
rect 3616 85380 3672 85436
rect 3672 85380 3676 85436
rect 3612 85376 3676 85380
rect 3692 85436 3756 85440
rect 3692 85380 3696 85436
rect 3696 85380 3752 85436
rect 3752 85380 3756 85436
rect 3692 85376 3756 85380
rect 3772 85436 3836 85440
rect 3772 85380 3776 85436
rect 3776 85380 3832 85436
rect 3832 85380 3836 85436
rect 3772 85376 3836 85380
rect 3852 85436 3916 85440
rect 3852 85380 3856 85436
rect 3856 85380 3912 85436
rect 3912 85380 3916 85436
rect 3852 85376 3916 85380
rect 5212 85436 5276 85440
rect 5212 85380 5216 85436
rect 5216 85380 5272 85436
rect 5272 85380 5276 85436
rect 5212 85376 5276 85380
rect 5292 85436 5356 85440
rect 5292 85380 5296 85436
rect 5296 85380 5352 85436
rect 5352 85380 5356 85436
rect 5292 85376 5356 85380
rect 5372 85436 5436 85440
rect 5372 85380 5376 85436
rect 5376 85380 5432 85436
rect 5432 85380 5436 85436
rect 5372 85376 5436 85380
rect 5452 85436 5516 85440
rect 5452 85380 5456 85436
rect 5456 85380 5512 85436
rect 5512 85380 5516 85436
rect 5452 85376 5516 85380
rect 6812 85436 6876 85440
rect 6812 85380 6816 85436
rect 6816 85380 6872 85436
rect 6872 85380 6876 85436
rect 6812 85376 6876 85380
rect 6892 85436 6956 85440
rect 6892 85380 6896 85436
rect 6896 85380 6952 85436
rect 6952 85380 6956 85436
rect 6892 85376 6956 85380
rect 6972 85436 7036 85440
rect 6972 85380 6976 85436
rect 6976 85380 7032 85436
rect 7032 85380 7036 85436
rect 6972 85376 7036 85380
rect 7052 85436 7116 85440
rect 7052 85380 7056 85436
rect 7056 85380 7112 85436
rect 7112 85380 7116 85436
rect 7052 85376 7116 85380
rect 8412 85436 8476 85440
rect 8412 85380 8416 85436
rect 8416 85380 8472 85436
rect 8472 85380 8476 85436
rect 8412 85376 8476 85380
rect 8492 85436 8556 85440
rect 8492 85380 8496 85436
rect 8496 85380 8552 85436
rect 8552 85380 8556 85436
rect 8492 85376 8556 85380
rect 8572 85436 8636 85440
rect 8572 85380 8576 85436
rect 8576 85380 8632 85436
rect 8632 85380 8636 85436
rect 8572 85376 8636 85380
rect 8652 85436 8716 85440
rect 8652 85380 8656 85436
rect 8656 85380 8712 85436
rect 8712 85380 8716 85436
rect 8652 85376 8716 85380
rect 2952 84892 3016 84896
rect 2952 84836 2956 84892
rect 2956 84836 3012 84892
rect 3012 84836 3016 84892
rect 2952 84832 3016 84836
rect 3032 84892 3096 84896
rect 3032 84836 3036 84892
rect 3036 84836 3092 84892
rect 3092 84836 3096 84892
rect 3032 84832 3096 84836
rect 3112 84892 3176 84896
rect 3112 84836 3116 84892
rect 3116 84836 3172 84892
rect 3172 84836 3176 84892
rect 3112 84832 3176 84836
rect 3192 84892 3256 84896
rect 3192 84836 3196 84892
rect 3196 84836 3252 84892
rect 3252 84836 3256 84892
rect 3192 84832 3256 84836
rect 4552 84892 4616 84896
rect 4552 84836 4556 84892
rect 4556 84836 4612 84892
rect 4612 84836 4616 84892
rect 4552 84832 4616 84836
rect 4632 84892 4696 84896
rect 4632 84836 4636 84892
rect 4636 84836 4692 84892
rect 4692 84836 4696 84892
rect 4632 84832 4696 84836
rect 4712 84892 4776 84896
rect 4712 84836 4716 84892
rect 4716 84836 4772 84892
rect 4772 84836 4776 84892
rect 4712 84832 4776 84836
rect 4792 84892 4856 84896
rect 4792 84836 4796 84892
rect 4796 84836 4852 84892
rect 4852 84836 4856 84892
rect 4792 84832 4856 84836
rect 6152 84892 6216 84896
rect 6152 84836 6156 84892
rect 6156 84836 6212 84892
rect 6212 84836 6216 84892
rect 6152 84832 6216 84836
rect 6232 84892 6296 84896
rect 6232 84836 6236 84892
rect 6236 84836 6292 84892
rect 6292 84836 6296 84892
rect 6232 84832 6296 84836
rect 6312 84892 6376 84896
rect 6312 84836 6316 84892
rect 6316 84836 6372 84892
rect 6372 84836 6376 84892
rect 6312 84832 6376 84836
rect 6392 84892 6456 84896
rect 6392 84836 6396 84892
rect 6396 84836 6452 84892
rect 6452 84836 6456 84892
rect 6392 84832 6456 84836
rect 7752 84892 7816 84896
rect 7752 84836 7756 84892
rect 7756 84836 7812 84892
rect 7812 84836 7816 84892
rect 7752 84832 7816 84836
rect 7832 84892 7896 84896
rect 7832 84836 7836 84892
rect 7836 84836 7892 84892
rect 7892 84836 7896 84892
rect 7832 84832 7896 84836
rect 7912 84892 7976 84896
rect 7912 84836 7916 84892
rect 7916 84836 7972 84892
rect 7972 84836 7976 84892
rect 7912 84832 7976 84836
rect 7992 84892 8056 84896
rect 7992 84836 7996 84892
rect 7996 84836 8052 84892
rect 8052 84836 8056 84892
rect 7992 84832 8056 84836
rect 9352 84892 9416 84896
rect 9352 84836 9356 84892
rect 9356 84836 9412 84892
rect 9412 84836 9416 84892
rect 9352 84832 9416 84836
rect 9432 84892 9496 84896
rect 9432 84836 9436 84892
rect 9436 84836 9492 84892
rect 9492 84836 9496 84892
rect 9432 84832 9496 84836
rect 9512 84892 9576 84896
rect 9512 84836 9516 84892
rect 9516 84836 9572 84892
rect 9572 84836 9576 84892
rect 9512 84832 9576 84836
rect 9592 84892 9656 84896
rect 9592 84836 9596 84892
rect 9596 84836 9652 84892
rect 9652 84836 9656 84892
rect 9592 84832 9656 84836
rect 52500 84824 52564 84828
rect 52500 84768 52514 84824
rect 52514 84768 52564 84824
rect 52500 84764 52564 84768
rect 51212 84688 51276 84692
rect 51212 84632 51226 84688
rect 51226 84632 51276 84688
rect 51212 84628 51276 84632
rect 53788 84688 53852 84692
rect 53788 84632 53838 84688
rect 53838 84632 53852 84688
rect 53788 84628 53852 84632
rect 66300 84688 66364 84692
rect 66300 84632 66314 84688
rect 66314 84632 66364 84688
rect 66300 84628 66364 84632
rect 71268 84688 71332 84692
rect 71268 84632 71282 84688
rect 71282 84632 71332 84688
rect 71268 84628 71332 84632
rect 57652 84552 57716 84556
rect 57652 84496 57666 84552
rect 57666 84496 57716 84552
rect 57652 84492 57716 84496
rect 78628 84552 78692 84556
rect 78628 84496 78678 84552
rect 78678 84496 78692 84552
rect 78628 84492 78692 84496
rect 42564 84416 42628 84420
rect 42564 84360 42578 84416
rect 42578 84360 42628 84416
rect 42564 84356 42628 84360
rect 44772 84416 44836 84420
rect 44772 84360 44786 84416
rect 44786 84360 44836 84416
rect 44772 84356 44836 84360
rect 3612 84348 3676 84352
rect 3612 84292 3616 84348
rect 3616 84292 3672 84348
rect 3672 84292 3676 84348
rect 3612 84288 3676 84292
rect 3692 84348 3756 84352
rect 3692 84292 3696 84348
rect 3696 84292 3752 84348
rect 3752 84292 3756 84348
rect 3692 84288 3756 84292
rect 3772 84348 3836 84352
rect 3772 84292 3776 84348
rect 3776 84292 3832 84348
rect 3832 84292 3836 84348
rect 3772 84288 3836 84292
rect 3852 84348 3916 84352
rect 3852 84292 3856 84348
rect 3856 84292 3912 84348
rect 3912 84292 3916 84348
rect 3852 84288 3916 84292
rect 5212 84348 5276 84352
rect 5212 84292 5216 84348
rect 5216 84292 5272 84348
rect 5272 84292 5276 84348
rect 5212 84288 5276 84292
rect 5292 84348 5356 84352
rect 5292 84292 5296 84348
rect 5296 84292 5352 84348
rect 5352 84292 5356 84348
rect 5292 84288 5356 84292
rect 5372 84348 5436 84352
rect 5372 84292 5376 84348
rect 5376 84292 5432 84348
rect 5432 84292 5436 84348
rect 5372 84288 5436 84292
rect 5452 84348 5516 84352
rect 5452 84292 5456 84348
rect 5456 84292 5512 84348
rect 5512 84292 5516 84348
rect 5452 84288 5516 84292
rect 6812 84348 6876 84352
rect 6812 84292 6816 84348
rect 6816 84292 6872 84348
rect 6872 84292 6876 84348
rect 6812 84288 6876 84292
rect 6892 84348 6956 84352
rect 6892 84292 6896 84348
rect 6896 84292 6952 84348
rect 6952 84292 6956 84348
rect 6892 84288 6956 84292
rect 6972 84348 7036 84352
rect 6972 84292 6976 84348
rect 6976 84292 7032 84348
rect 7032 84292 7036 84348
rect 6972 84288 7036 84292
rect 7052 84348 7116 84352
rect 7052 84292 7056 84348
rect 7056 84292 7112 84348
rect 7112 84292 7116 84348
rect 7052 84288 7116 84292
rect 8412 84348 8476 84352
rect 8412 84292 8416 84348
rect 8416 84292 8472 84348
rect 8472 84292 8476 84348
rect 8412 84288 8476 84292
rect 8492 84348 8556 84352
rect 8492 84292 8496 84348
rect 8496 84292 8552 84348
rect 8552 84292 8556 84348
rect 8492 84288 8556 84292
rect 8572 84348 8636 84352
rect 8572 84292 8576 84348
rect 8576 84292 8632 84348
rect 8632 84292 8636 84348
rect 8572 84288 8636 84292
rect 8652 84348 8716 84352
rect 8652 84292 8656 84348
rect 8656 84292 8712 84348
rect 8712 84292 8716 84348
rect 8652 84288 8716 84292
rect 10916 84220 10980 84284
rect 65012 84220 65076 84284
rect 2952 83804 3016 83808
rect 2952 83748 2956 83804
rect 2956 83748 3012 83804
rect 3012 83748 3016 83804
rect 2952 83744 3016 83748
rect 3032 83804 3096 83808
rect 3032 83748 3036 83804
rect 3036 83748 3092 83804
rect 3092 83748 3096 83804
rect 3032 83744 3096 83748
rect 3112 83804 3176 83808
rect 3112 83748 3116 83804
rect 3116 83748 3172 83804
rect 3172 83748 3176 83804
rect 3112 83744 3176 83748
rect 3192 83804 3256 83808
rect 3192 83748 3196 83804
rect 3196 83748 3252 83804
rect 3252 83748 3256 83804
rect 3192 83744 3256 83748
rect 4552 83804 4616 83808
rect 4552 83748 4556 83804
rect 4556 83748 4612 83804
rect 4612 83748 4616 83804
rect 4552 83744 4616 83748
rect 4632 83804 4696 83808
rect 4632 83748 4636 83804
rect 4636 83748 4692 83804
rect 4692 83748 4696 83804
rect 4632 83744 4696 83748
rect 4712 83804 4776 83808
rect 4712 83748 4716 83804
rect 4716 83748 4772 83804
rect 4772 83748 4776 83804
rect 4712 83744 4776 83748
rect 4792 83804 4856 83808
rect 4792 83748 4796 83804
rect 4796 83748 4852 83804
rect 4852 83748 4856 83804
rect 4792 83744 4856 83748
rect 6152 83804 6216 83808
rect 6152 83748 6156 83804
rect 6156 83748 6212 83804
rect 6212 83748 6216 83804
rect 6152 83744 6216 83748
rect 6232 83804 6296 83808
rect 6232 83748 6236 83804
rect 6236 83748 6292 83804
rect 6292 83748 6296 83804
rect 6232 83744 6296 83748
rect 6312 83804 6376 83808
rect 6312 83748 6316 83804
rect 6316 83748 6372 83804
rect 6372 83748 6376 83804
rect 6312 83744 6376 83748
rect 6392 83804 6456 83808
rect 6392 83748 6396 83804
rect 6396 83748 6452 83804
rect 6452 83748 6456 83804
rect 6392 83744 6456 83748
rect 7752 83804 7816 83808
rect 7752 83748 7756 83804
rect 7756 83748 7812 83804
rect 7812 83748 7816 83804
rect 7752 83744 7816 83748
rect 7832 83804 7896 83808
rect 7832 83748 7836 83804
rect 7836 83748 7892 83804
rect 7892 83748 7896 83804
rect 7832 83744 7896 83748
rect 7912 83804 7976 83808
rect 7912 83748 7916 83804
rect 7916 83748 7972 83804
rect 7972 83748 7976 83804
rect 7912 83744 7976 83748
rect 7992 83804 8056 83808
rect 7992 83748 7996 83804
rect 7996 83748 8052 83804
rect 8052 83748 8056 83804
rect 7992 83744 8056 83748
rect 9352 83804 9416 83808
rect 9352 83748 9356 83804
rect 9356 83748 9412 83804
rect 9412 83748 9416 83804
rect 9352 83744 9416 83748
rect 9432 83804 9496 83808
rect 9432 83748 9436 83804
rect 9436 83748 9492 83804
rect 9492 83748 9496 83804
rect 9432 83744 9496 83748
rect 9512 83804 9576 83808
rect 9512 83748 9516 83804
rect 9516 83748 9572 83804
rect 9572 83748 9576 83804
rect 9512 83744 9576 83748
rect 9592 83804 9656 83808
rect 9592 83748 9596 83804
rect 9596 83748 9652 83804
rect 9652 83748 9656 83804
rect 9592 83744 9656 83748
rect 60150 83676 60214 83740
rect 70214 83736 70278 83740
rect 70214 83680 70270 83736
rect 70270 83680 70278 83736
rect 70214 83676 70278 83680
rect 3612 83260 3676 83264
rect 3612 83204 3616 83260
rect 3616 83204 3672 83260
rect 3672 83204 3676 83260
rect 3612 83200 3676 83204
rect 3692 83260 3756 83264
rect 3692 83204 3696 83260
rect 3696 83204 3752 83260
rect 3752 83204 3756 83260
rect 3692 83200 3756 83204
rect 3772 83260 3836 83264
rect 3772 83204 3776 83260
rect 3776 83204 3832 83260
rect 3832 83204 3836 83260
rect 3772 83200 3836 83204
rect 3852 83260 3916 83264
rect 3852 83204 3856 83260
rect 3856 83204 3912 83260
rect 3912 83204 3916 83260
rect 3852 83200 3916 83204
rect 5212 83260 5276 83264
rect 5212 83204 5216 83260
rect 5216 83204 5272 83260
rect 5272 83204 5276 83260
rect 5212 83200 5276 83204
rect 5292 83260 5356 83264
rect 5292 83204 5296 83260
rect 5296 83204 5352 83260
rect 5352 83204 5356 83260
rect 5292 83200 5356 83204
rect 5372 83260 5436 83264
rect 5372 83204 5376 83260
rect 5376 83204 5432 83260
rect 5432 83204 5436 83260
rect 5372 83200 5436 83204
rect 5452 83260 5516 83264
rect 5452 83204 5456 83260
rect 5456 83204 5512 83260
rect 5512 83204 5516 83260
rect 5452 83200 5516 83204
rect 6812 83260 6876 83264
rect 6812 83204 6816 83260
rect 6816 83204 6872 83260
rect 6872 83204 6876 83260
rect 6812 83200 6876 83204
rect 6892 83260 6956 83264
rect 6892 83204 6896 83260
rect 6896 83204 6952 83260
rect 6952 83204 6956 83260
rect 6892 83200 6956 83204
rect 6972 83260 7036 83264
rect 6972 83204 6976 83260
rect 6976 83204 7032 83260
rect 7032 83204 7036 83260
rect 6972 83200 7036 83204
rect 7052 83260 7116 83264
rect 7052 83204 7056 83260
rect 7056 83204 7112 83260
rect 7112 83204 7116 83260
rect 7052 83200 7116 83204
rect 8412 83260 8476 83264
rect 8412 83204 8416 83260
rect 8416 83204 8472 83260
rect 8472 83204 8476 83260
rect 8412 83200 8476 83204
rect 8492 83260 8556 83264
rect 8492 83204 8496 83260
rect 8496 83204 8552 83260
rect 8552 83204 8556 83260
rect 8492 83200 8556 83204
rect 8572 83260 8636 83264
rect 8572 83204 8576 83260
rect 8576 83204 8632 83260
rect 8632 83204 8636 83260
rect 8572 83200 8636 83204
rect 8652 83260 8716 83264
rect 8652 83204 8656 83260
rect 8656 83204 8712 83260
rect 8712 83204 8716 83260
rect 8652 83200 8716 83204
rect 2952 82716 3016 82720
rect 2952 82660 2956 82716
rect 2956 82660 3012 82716
rect 3012 82660 3016 82716
rect 2952 82656 3016 82660
rect 3032 82716 3096 82720
rect 3032 82660 3036 82716
rect 3036 82660 3092 82716
rect 3092 82660 3096 82716
rect 3032 82656 3096 82660
rect 3112 82716 3176 82720
rect 3112 82660 3116 82716
rect 3116 82660 3172 82716
rect 3172 82660 3176 82716
rect 3112 82656 3176 82660
rect 3192 82716 3256 82720
rect 3192 82660 3196 82716
rect 3196 82660 3252 82716
rect 3252 82660 3256 82716
rect 3192 82656 3256 82660
rect 4552 82716 4616 82720
rect 4552 82660 4556 82716
rect 4556 82660 4612 82716
rect 4612 82660 4616 82716
rect 4552 82656 4616 82660
rect 4632 82716 4696 82720
rect 4632 82660 4636 82716
rect 4636 82660 4692 82716
rect 4692 82660 4696 82716
rect 4632 82656 4696 82660
rect 4712 82716 4776 82720
rect 4712 82660 4716 82716
rect 4716 82660 4772 82716
rect 4772 82660 4776 82716
rect 4712 82656 4776 82660
rect 4792 82716 4856 82720
rect 4792 82660 4796 82716
rect 4796 82660 4852 82716
rect 4852 82660 4856 82716
rect 4792 82656 4856 82660
rect 6152 82716 6216 82720
rect 6152 82660 6156 82716
rect 6156 82660 6212 82716
rect 6212 82660 6216 82716
rect 6152 82656 6216 82660
rect 6232 82716 6296 82720
rect 6232 82660 6236 82716
rect 6236 82660 6292 82716
rect 6292 82660 6296 82716
rect 6232 82656 6296 82660
rect 6312 82716 6376 82720
rect 6312 82660 6316 82716
rect 6316 82660 6372 82716
rect 6372 82660 6376 82716
rect 6312 82656 6376 82660
rect 6392 82716 6456 82720
rect 6392 82660 6396 82716
rect 6396 82660 6452 82716
rect 6452 82660 6456 82716
rect 6392 82656 6456 82660
rect 7752 82716 7816 82720
rect 7752 82660 7756 82716
rect 7756 82660 7812 82716
rect 7812 82660 7816 82716
rect 7752 82656 7816 82660
rect 7832 82716 7896 82720
rect 7832 82660 7836 82716
rect 7836 82660 7892 82716
rect 7892 82660 7896 82716
rect 7832 82656 7896 82660
rect 7912 82716 7976 82720
rect 7912 82660 7916 82716
rect 7916 82660 7972 82716
rect 7972 82660 7976 82716
rect 7912 82656 7976 82660
rect 7992 82716 8056 82720
rect 7992 82660 7996 82716
rect 7996 82660 8052 82716
rect 8052 82660 8056 82716
rect 7992 82656 8056 82660
rect 9352 82716 9416 82720
rect 9352 82660 9356 82716
rect 9356 82660 9412 82716
rect 9412 82660 9416 82716
rect 9352 82656 9416 82660
rect 9432 82716 9496 82720
rect 9432 82660 9436 82716
rect 9436 82660 9492 82716
rect 9492 82660 9496 82716
rect 9432 82656 9496 82660
rect 9512 82716 9576 82720
rect 9512 82660 9516 82716
rect 9516 82660 9572 82716
rect 9572 82660 9576 82716
rect 9512 82656 9576 82660
rect 9592 82716 9656 82720
rect 9592 82660 9596 82716
rect 9596 82660 9652 82716
rect 9652 82660 9656 82716
rect 9592 82656 9656 82660
rect 3612 82172 3676 82176
rect 3612 82116 3616 82172
rect 3616 82116 3672 82172
rect 3672 82116 3676 82172
rect 3612 82112 3676 82116
rect 3692 82172 3756 82176
rect 3692 82116 3696 82172
rect 3696 82116 3752 82172
rect 3752 82116 3756 82172
rect 3692 82112 3756 82116
rect 3772 82172 3836 82176
rect 3772 82116 3776 82172
rect 3776 82116 3832 82172
rect 3832 82116 3836 82172
rect 3772 82112 3836 82116
rect 3852 82172 3916 82176
rect 3852 82116 3856 82172
rect 3856 82116 3912 82172
rect 3912 82116 3916 82172
rect 3852 82112 3916 82116
rect 5212 82172 5276 82176
rect 5212 82116 5216 82172
rect 5216 82116 5272 82172
rect 5272 82116 5276 82172
rect 5212 82112 5276 82116
rect 5292 82172 5356 82176
rect 5292 82116 5296 82172
rect 5296 82116 5352 82172
rect 5352 82116 5356 82172
rect 5292 82112 5356 82116
rect 5372 82172 5436 82176
rect 5372 82116 5376 82172
rect 5376 82116 5432 82172
rect 5432 82116 5436 82172
rect 5372 82112 5436 82116
rect 5452 82172 5516 82176
rect 5452 82116 5456 82172
rect 5456 82116 5512 82172
rect 5512 82116 5516 82172
rect 5452 82112 5516 82116
rect 6812 82172 6876 82176
rect 6812 82116 6816 82172
rect 6816 82116 6872 82172
rect 6872 82116 6876 82172
rect 6812 82112 6876 82116
rect 6892 82172 6956 82176
rect 6892 82116 6896 82172
rect 6896 82116 6952 82172
rect 6952 82116 6956 82172
rect 6892 82112 6956 82116
rect 6972 82172 7036 82176
rect 6972 82116 6976 82172
rect 6976 82116 7032 82172
rect 7032 82116 7036 82172
rect 6972 82112 7036 82116
rect 7052 82172 7116 82176
rect 7052 82116 7056 82172
rect 7056 82116 7112 82172
rect 7112 82116 7116 82172
rect 7052 82112 7116 82116
rect 8412 82172 8476 82176
rect 8412 82116 8416 82172
rect 8416 82116 8472 82172
rect 8472 82116 8476 82172
rect 8412 82112 8476 82116
rect 8492 82172 8556 82176
rect 8492 82116 8496 82172
rect 8496 82116 8552 82172
rect 8552 82116 8556 82172
rect 8492 82112 8556 82116
rect 8572 82172 8636 82176
rect 8572 82116 8576 82172
rect 8576 82116 8632 82172
rect 8632 82116 8636 82172
rect 8572 82112 8636 82116
rect 8652 82172 8716 82176
rect 8652 82116 8656 82172
rect 8656 82116 8712 82172
rect 8712 82116 8716 82172
rect 8652 82112 8716 82116
rect 2952 81628 3016 81632
rect 2952 81572 2956 81628
rect 2956 81572 3012 81628
rect 3012 81572 3016 81628
rect 2952 81568 3016 81572
rect 3032 81628 3096 81632
rect 3032 81572 3036 81628
rect 3036 81572 3092 81628
rect 3092 81572 3096 81628
rect 3032 81568 3096 81572
rect 3112 81628 3176 81632
rect 3112 81572 3116 81628
rect 3116 81572 3172 81628
rect 3172 81572 3176 81628
rect 3112 81568 3176 81572
rect 3192 81628 3256 81632
rect 3192 81572 3196 81628
rect 3196 81572 3252 81628
rect 3252 81572 3256 81628
rect 3192 81568 3256 81572
rect 4552 81628 4616 81632
rect 4552 81572 4556 81628
rect 4556 81572 4612 81628
rect 4612 81572 4616 81628
rect 4552 81568 4616 81572
rect 4632 81628 4696 81632
rect 4632 81572 4636 81628
rect 4636 81572 4692 81628
rect 4692 81572 4696 81628
rect 4632 81568 4696 81572
rect 4712 81628 4776 81632
rect 4712 81572 4716 81628
rect 4716 81572 4772 81628
rect 4772 81572 4776 81628
rect 4712 81568 4776 81572
rect 4792 81628 4856 81632
rect 4792 81572 4796 81628
rect 4796 81572 4852 81628
rect 4852 81572 4856 81628
rect 4792 81568 4856 81572
rect 6152 81628 6216 81632
rect 6152 81572 6156 81628
rect 6156 81572 6212 81628
rect 6212 81572 6216 81628
rect 6152 81568 6216 81572
rect 6232 81628 6296 81632
rect 6232 81572 6236 81628
rect 6236 81572 6292 81628
rect 6292 81572 6296 81628
rect 6232 81568 6296 81572
rect 6312 81628 6376 81632
rect 6312 81572 6316 81628
rect 6316 81572 6372 81628
rect 6372 81572 6376 81628
rect 6312 81568 6376 81572
rect 6392 81628 6456 81632
rect 6392 81572 6396 81628
rect 6396 81572 6452 81628
rect 6452 81572 6456 81628
rect 6392 81568 6456 81572
rect 7752 81628 7816 81632
rect 7752 81572 7756 81628
rect 7756 81572 7812 81628
rect 7812 81572 7816 81628
rect 7752 81568 7816 81572
rect 7832 81628 7896 81632
rect 7832 81572 7836 81628
rect 7836 81572 7892 81628
rect 7892 81572 7896 81628
rect 7832 81568 7896 81572
rect 7912 81628 7976 81632
rect 7912 81572 7916 81628
rect 7916 81572 7972 81628
rect 7972 81572 7976 81628
rect 7912 81568 7976 81572
rect 7992 81628 8056 81632
rect 7992 81572 7996 81628
rect 7996 81572 8052 81628
rect 8052 81572 8056 81628
rect 7992 81568 8056 81572
rect 9352 81628 9416 81632
rect 9352 81572 9356 81628
rect 9356 81572 9412 81628
rect 9412 81572 9416 81628
rect 9352 81568 9416 81572
rect 9432 81628 9496 81632
rect 9432 81572 9436 81628
rect 9436 81572 9492 81628
rect 9492 81572 9496 81628
rect 9432 81568 9496 81572
rect 9512 81628 9576 81632
rect 9512 81572 9516 81628
rect 9516 81572 9572 81628
rect 9572 81572 9576 81628
rect 9512 81568 9576 81572
rect 9592 81628 9656 81632
rect 9592 81572 9596 81628
rect 9596 81572 9652 81628
rect 9652 81572 9656 81628
rect 9592 81568 9656 81572
rect 3612 81084 3676 81088
rect 3612 81028 3616 81084
rect 3616 81028 3672 81084
rect 3672 81028 3676 81084
rect 3612 81024 3676 81028
rect 3692 81084 3756 81088
rect 3692 81028 3696 81084
rect 3696 81028 3752 81084
rect 3752 81028 3756 81084
rect 3692 81024 3756 81028
rect 3772 81084 3836 81088
rect 3772 81028 3776 81084
rect 3776 81028 3832 81084
rect 3832 81028 3836 81084
rect 3772 81024 3836 81028
rect 3852 81084 3916 81088
rect 3852 81028 3856 81084
rect 3856 81028 3912 81084
rect 3912 81028 3916 81084
rect 3852 81024 3916 81028
rect 5212 81084 5276 81088
rect 5212 81028 5216 81084
rect 5216 81028 5272 81084
rect 5272 81028 5276 81084
rect 5212 81024 5276 81028
rect 5292 81084 5356 81088
rect 5292 81028 5296 81084
rect 5296 81028 5352 81084
rect 5352 81028 5356 81084
rect 5292 81024 5356 81028
rect 5372 81084 5436 81088
rect 5372 81028 5376 81084
rect 5376 81028 5432 81084
rect 5432 81028 5436 81084
rect 5372 81024 5436 81028
rect 5452 81084 5516 81088
rect 5452 81028 5456 81084
rect 5456 81028 5512 81084
rect 5512 81028 5516 81084
rect 5452 81024 5516 81028
rect 6812 81084 6876 81088
rect 6812 81028 6816 81084
rect 6816 81028 6872 81084
rect 6872 81028 6876 81084
rect 6812 81024 6876 81028
rect 6892 81084 6956 81088
rect 6892 81028 6896 81084
rect 6896 81028 6952 81084
rect 6952 81028 6956 81084
rect 6892 81024 6956 81028
rect 6972 81084 7036 81088
rect 6972 81028 6976 81084
rect 6976 81028 7032 81084
rect 7032 81028 7036 81084
rect 6972 81024 7036 81028
rect 7052 81084 7116 81088
rect 7052 81028 7056 81084
rect 7056 81028 7112 81084
rect 7112 81028 7116 81084
rect 7052 81024 7116 81028
rect 8412 81084 8476 81088
rect 8412 81028 8416 81084
rect 8416 81028 8472 81084
rect 8472 81028 8476 81084
rect 8412 81024 8476 81028
rect 8492 81084 8556 81088
rect 8492 81028 8496 81084
rect 8496 81028 8552 81084
rect 8552 81028 8556 81084
rect 8492 81024 8556 81028
rect 8572 81084 8636 81088
rect 8572 81028 8576 81084
rect 8576 81028 8632 81084
rect 8632 81028 8636 81084
rect 8572 81024 8636 81028
rect 8652 81084 8716 81088
rect 8652 81028 8656 81084
rect 8656 81028 8712 81084
rect 8712 81028 8716 81084
rect 8652 81024 8716 81028
rect 2952 80540 3016 80544
rect 2952 80484 2956 80540
rect 2956 80484 3012 80540
rect 3012 80484 3016 80540
rect 2952 80480 3016 80484
rect 3032 80540 3096 80544
rect 3032 80484 3036 80540
rect 3036 80484 3092 80540
rect 3092 80484 3096 80540
rect 3032 80480 3096 80484
rect 3112 80540 3176 80544
rect 3112 80484 3116 80540
rect 3116 80484 3172 80540
rect 3172 80484 3176 80540
rect 3112 80480 3176 80484
rect 3192 80540 3256 80544
rect 3192 80484 3196 80540
rect 3196 80484 3252 80540
rect 3252 80484 3256 80540
rect 3192 80480 3256 80484
rect 4552 80540 4616 80544
rect 4552 80484 4556 80540
rect 4556 80484 4612 80540
rect 4612 80484 4616 80540
rect 4552 80480 4616 80484
rect 4632 80540 4696 80544
rect 4632 80484 4636 80540
rect 4636 80484 4692 80540
rect 4692 80484 4696 80540
rect 4632 80480 4696 80484
rect 4712 80540 4776 80544
rect 4712 80484 4716 80540
rect 4716 80484 4772 80540
rect 4772 80484 4776 80540
rect 4712 80480 4776 80484
rect 4792 80540 4856 80544
rect 4792 80484 4796 80540
rect 4796 80484 4852 80540
rect 4852 80484 4856 80540
rect 4792 80480 4856 80484
rect 6152 80540 6216 80544
rect 6152 80484 6156 80540
rect 6156 80484 6212 80540
rect 6212 80484 6216 80540
rect 6152 80480 6216 80484
rect 6232 80540 6296 80544
rect 6232 80484 6236 80540
rect 6236 80484 6292 80540
rect 6292 80484 6296 80540
rect 6232 80480 6296 80484
rect 6312 80540 6376 80544
rect 6312 80484 6316 80540
rect 6316 80484 6372 80540
rect 6372 80484 6376 80540
rect 6312 80480 6376 80484
rect 6392 80540 6456 80544
rect 6392 80484 6396 80540
rect 6396 80484 6452 80540
rect 6452 80484 6456 80540
rect 6392 80480 6456 80484
rect 7752 80540 7816 80544
rect 7752 80484 7756 80540
rect 7756 80484 7812 80540
rect 7812 80484 7816 80540
rect 7752 80480 7816 80484
rect 7832 80540 7896 80544
rect 7832 80484 7836 80540
rect 7836 80484 7892 80540
rect 7892 80484 7896 80540
rect 7832 80480 7896 80484
rect 7912 80540 7976 80544
rect 7912 80484 7916 80540
rect 7916 80484 7972 80540
rect 7972 80484 7976 80540
rect 7912 80480 7976 80484
rect 7992 80540 8056 80544
rect 7992 80484 7996 80540
rect 7996 80484 8052 80540
rect 8052 80484 8056 80540
rect 7992 80480 8056 80484
rect 9352 80540 9416 80544
rect 9352 80484 9356 80540
rect 9356 80484 9412 80540
rect 9412 80484 9416 80540
rect 9352 80480 9416 80484
rect 9432 80540 9496 80544
rect 9432 80484 9436 80540
rect 9436 80484 9492 80540
rect 9492 80484 9496 80540
rect 9432 80480 9496 80484
rect 9512 80540 9576 80544
rect 9512 80484 9516 80540
rect 9516 80484 9572 80540
rect 9572 80484 9576 80540
rect 9512 80480 9576 80484
rect 9592 80540 9656 80544
rect 9592 80484 9596 80540
rect 9596 80484 9652 80540
rect 9652 80484 9656 80540
rect 9592 80480 9656 80484
rect 3612 79996 3676 80000
rect 3612 79940 3616 79996
rect 3616 79940 3672 79996
rect 3672 79940 3676 79996
rect 3612 79936 3676 79940
rect 3692 79996 3756 80000
rect 3692 79940 3696 79996
rect 3696 79940 3752 79996
rect 3752 79940 3756 79996
rect 3692 79936 3756 79940
rect 3772 79996 3836 80000
rect 3772 79940 3776 79996
rect 3776 79940 3832 79996
rect 3832 79940 3836 79996
rect 3772 79936 3836 79940
rect 3852 79996 3916 80000
rect 3852 79940 3856 79996
rect 3856 79940 3912 79996
rect 3912 79940 3916 79996
rect 3852 79936 3916 79940
rect 5212 79996 5276 80000
rect 5212 79940 5216 79996
rect 5216 79940 5272 79996
rect 5272 79940 5276 79996
rect 5212 79936 5276 79940
rect 5292 79996 5356 80000
rect 5292 79940 5296 79996
rect 5296 79940 5352 79996
rect 5352 79940 5356 79996
rect 5292 79936 5356 79940
rect 5372 79996 5436 80000
rect 5372 79940 5376 79996
rect 5376 79940 5432 79996
rect 5432 79940 5436 79996
rect 5372 79936 5436 79940
rect 5452 79996 5516 80000
rect 5452 79940 5456 79996
rect 5456 79940 5512 79996
rect 5512 79940 5516 79996
rect 5452 79936 5516 79940
rect 6812 79996 6876 80000
rect 6812 79940 6816 79996
rect 6816 79940 6872 79996
rect 6872 79940 6876 79996
rect 6812 79936 6876 79940
rect 6892 79996 6956 80000
rect 6892 79940 6896 79996
rect 6896 79940 6952 79996
rect 6952 79940 6956 79996
rect 6892 79936 6956 79940
rect 6972 79996 7036 80000
rect 6972 79940 6976 79996
rect 6976 79940 7032 79996
rect 7032 79940 7036 79996
rect 6972 79936 7036 79940
rect 7052 79996 7116 80000
rect 7052 79940 7056 79996
rect 7056 79940 7112 79996
rect 7112 79940 7116 79996
rect 7052 79936 7116 79940
rect 8412 79996 8476 80000
rect 8412 79940 8416 79996
rect 8416 79940 8472 79996
rect 8472 79940 8476 79996
rect 8412 79936 8476 79940
rect 8492 79996 8556 80000
rect 8492 79940 8496 79996
rect 8496 79940 8552 79996
rect 8552 79940 8556 79996
rect 8492 79936 8556 79940
rect 8572 79996 8636 80000
rect 8572 79940 8576 79996
rect 8576 79940 8632 79996
rect 8632 79940 8636 79996
rect 8572 79936 8636 79940
rect 8652 79996 8716 80000
rect 8652 79940 8656 79996
rect 8656 79940 8712 79996
rect 8712 79940 8716 79996
rect 8652 79936 8716 79940
rect 2952 79452 3016 79456
rect 2952 79396 2956 79452
rect 2956 79396 3012 79452
rect 3012 79396 3016 79452
rect 2952 79392 3016 79396
rect 3032 79452 3096 79456
rect 3032 79396 3036 79452
rect 3036 79396 3092 79452
rect 3092 79396 3096 79452
rect 3032 79392 3096 79396
rect 3112 79452 3176 79456
rect 3112 79396 3116 79452
rect 3116 79396 3172 79452
rect 3172 79396 3176 79452
rect 3112 79392 3176 79396
rect 3192 79452 3256 79456
rect 3192 79396 3196 79452
rect 3196 79396 3252 79452
rect 3252 79396 3256 79452
rect 3192 79392 3256 79396
rect 4552 79452 4616 79456
rect 4552 79396 4556 79452
rect 4556 79396 4612 79452
rect 4612 79396 4616 79452
rect 4552 79392 4616 79396
rect 4632 79452 4696 79456
rect 4632 79396 4636 79452
rect 4636 79396 4692 79452
rect 4692 79396 4696 79452
rect 4632 79392 4696 79396
rect 4712 79452 4776 79456
rect 4712 79396 4716 79452
rect 4716 79396 4772 79452
rect 4772 79396 4776 79452
rect 4712 79392 4776 79396
rect 4792 79452 4856 79456
rect 4792 79396 4796 79452
rect 4796 79396 4852 79452
rect 4852 79396 4856 79452
rect 4792 79392 4856 79396
rect 6152 79452 6216 79456
rect 6152 79396 6156 79452
rect 6156 79396 6212 79452
rect 6212 79396 6216 79452
rect 6152 79392 6216 79396
rect 6232 79452 6296 79456
rect 6232 79396 6236 79452
rect 6236 79396 6292 79452
rect 6292 79396 6296 79452
rect 6232 79392 6296 79396
rect 6312 79452 6376 79456
rect 6312 79396 6316 79452
rect 6316 79396 6372 79452
rect 6372 79396 6376 79452
rect 6312 79392 6376 79396
rect 6392 79452 6456 79456
rect 6392 79396 6396 79452
rect 6396 79396 6452 79452
rect 6452 79396 6456 79452
rect 6392 79392 6456 79396
rect 7752 79452 7816 79456
rect 7752 79396 7756 79452
rect 7756 79396 7812 79452
rect 7812 79396 7816 79452
rect 7752 79392 7816 79396
rect 7832 79452 7896 79456
rect 7832 79396 7836 79452
rect 7836 79396 7892 79452
rect 7892 79396 7896 79452
rect 7832 79392 7896 79396
rect 7912 79452 7976 79456
rect 7912 79396 7916 79452
rect 7916 79396 7972 79452
rect 7972 79396 7976 79452
rect 7912 79392 7976 79396
rect 7992 79452 8056 79456
rect 7992 79396 7996 79452
rect 7996 79396 8052 79452
rect 8052 79396 8056 79452
rect 7992 79392 8056 79396
rect 9352 79452 9416 79456
rect 9352 79396 9356 79452
rect 9356 79396 9412 79452
rect 9412 79396 9416 79452
rect 9352 79392 9416 79396
rect 9432 79452 9496 79456
rect 9432 79396 9436 79452
rect 9436 79396 9492 79452
rect 9492 79396 9496 79452
rect 9432 79392 9496 79396
rect 9512 79452 9576 79456
rect 9512 79396 9516 79452
rect 9516 79396 9572 79452
rect 9572 79396 9576 79452
rect 9512 79392 9576 79396
rect 9592 79452 9656 79456
rect 9592 79396 9596 79452
rect 9596 79396 9652 79452
rect 9652 79396 9656 79452
rect 9592 79392 9656 79396
rect 3612 78908 3676 78912
rect 3612 78852 3616 78908
rect 3616 78852 3672 78908
rect 3672 78852 3676 78908
rect 3612 78848 3676 78852
rect 3692 78908 3756 78912
rect 3692 78852 3696 78908
rect 3696 78852 3752 78908
rect 3752 78852 3756 78908
rect 3692 78848 3756 78852
rect 3772 78908 3836 78912
rect 3772 78852 3776 78908
rect 3776 78852 3832 78908
rect 3832 78852 3836 78908
rect 3772 78848 3836 78852
rect 3852 78908 3916 78912
rect 3852 78852 3856 78908
rect 3856 78852 3912 78908
rect 3912 78852 3916 78908
rect 3852 78848 3916 78852
rect 5212 78908 5276 78912
rect 5212 78852 5216 78908
rect 5216 78852 5272 78908
rect 5272 78852 5276 78908
rect 5212 78848 5276 78852
rect 5292 78908 5356 78912
rect 5292 78852 5296 78908
rect 5296 78852 5352 78908
rect 5352 78852 5356 78908
rect 5292 78848 5356 78852
rect 5372 78908 5436 78912
rect 5372 78852 5376 78908
rect 5376 78852 5432 78908
rect 5432 78852 5436 78908
rect 5372 78848 5436 78852
rect 5452 78908 5516 78912
rect 5452 78852 5456 78908
rect 5456 78852 5512 78908
rect 5512 78852 5516 78908
rect 5452 78848 5516 78852
rect 6812 78908 6876 78912
rect 6812 78852 6816 78908
rect 6816 78852 6872 78908
rect 6872 78852 6876 78908
rect 6812 78848 6876 78852
rect 6892 78908 6956 78912
rect 6892 78852 6896 78908
rect 6896 78852 6952 78908
rect 6952 78852 6956 78908
rect 6892 78848 6956 78852
rect 6972 78908 7036 78912
rect 6972 78852 6976 78908
rect 6976 78852 7032 78908
rect 7032 78852 7036 78908
rect 6972 78848 7036 78852
rect 7052 78908 7116 78912
rect 7052 78852 7056 78908
rect 7056 78852 7112 78908
rect 7112 78852 7116 78908
rect 7052 78848 7116 78852
rect 8412 78908 8476 78912
rect 8412 78852 8416 78908
rect 8416 78852 8472 78908
rect 8472 78852 8476 78908
rect 8412 78848 8476 78852
rect 8492 78908 8556 78912
rect 8492 78852 8496 78908
rect 8496 78852 8552 78908
rect 8552 78852 8556 78908
rect 8492 78848 8556 78852
rect 8572 78908 8636 78912
rect 8572 78852 8576 78908
rect 8576 78852 8632 78908
rect 8632 78852 8636 78908
rect 8572 78848 8636 78852
rect 8652 78908 8716 78912
rect 8652 78852 8656 78908
rect 8656 78852 8712 78908
rect 8712 78852 8716 78908
rect 8652 78848 8716 78852
rect 2952 78364 3016 78368
rect 2952 78308 2956 78364
rect 2956 78308 3012 78364
rect 3012 78308 3016 78364
rect 2952 78304 3016 78308
rect 3032 78364 3096 78368
rect 3032 78308 3036 78364
rect 3036 78308 3092 78364
rect 3092 78308 3096 78364
rect 3032 78304 3096 78308
rect 3112 78364 3176 78368
rect 3112 78308 3116 78364
rect 3116 78308 3172 78364
rect 3172 78308 3176 78364
rect 3112 78304 3176 78308
rect 3192 78364 3256 78368
rect 3192 78308 3196 78364
rect 3196 78308 3252 78364
rect 3252 78308 3256 78364
rect 3192 78304 3256 78308
rect 4552 78364 4616 78368
rect 4552 78308 4556 78364
rect 4556 78308 4612 78364
rect 4612 78308 4616 78364
rect 4552 78304 4616 78308
rect 4632 78364 4696 78368
rect 4632 78308 4636 78364
rect 4636 78308 4692 78364
rect 4692 78308 4696 78364
rect 4632 78304 4696 78308
rect 4712 78364 4776 78368
rect 4712 78308 4716 78364
rect 4716 78308 4772 78364
rect 4772 78308 4776 78364
rect 4712 78304 4776 78308
rect 4792 78364 4856 78368
rect 4792 78308 4796 78364
rect 4796 78308 4852 78364
rect 4852 78308 4856 78364
rect 4792 78304 4856 78308
rect 6152 78364 6216 78368
rect 6152 78308 6156 78364
rect 6156 78308 6212 78364
rect 6212 78308 6216 78364
rect 6152 78304 6216 78308
rect 6232 78364 6296 78368
rect 6232 78308 6236 78364
rect 6236 78308 6292 78364
rect 6292 78308 6296 78364
rect 6232 78304 6296 78308
rect 6312 78364 6376 78368
rect 6312 78308 6316 78364
rect 6316 78308 6372 78364
rect 6372 78308 6376 78364
rect 6312 78304 6376 78308
rect 6392 78364 6456 78368
rect 6392 78308 6396 78364
rect 6396 78308 6452 78364
rect 6452 78308 6456 78364
rect 6392 78304 6456 78308
rect 7752 78364 7816 78368
rect 7752 78308 7756 78364
rect 7756 78308 7812 78364
rect 7812 78308 7816 78364
rect 7752 78304 7816 78308
rect 7832 78364 7896 78368
rect 7832 78308 7836 78364
rect 7836 78308 7892 78364
rect 7892 78308 7896 78364
rect 7832 78304 7896 78308
rect 7912 78364 7976 78368
rect 7912 78308 7916 78364
rect 7916 78308 7972 78364
rect 7972 78308 7976 78364
rect 7912 78304 7976 78308
rect 7992 78364 8056 78368
rect 7992 78308 7996 78364
rect 7996 78308 8052 78364
rect 8052 78308 8056 78364
rect 7992 78304 8056 78308
rect 9352 78364 9416 78368
rect 9352 78308 9356 78364
rect 9356 78308 9412 78364
rect 9412 78308 9416 78364
rect 9352 78304 9416 78308
rect 9432 78364 9496 78368
rect 9432 78308 9436 78364
rect 9436 78308 9492 78364
rect 9492 78308 9496 78364
rect 9432 78304 9496 78308
rect 9512 78364 9576 78368
rect 9512 78308 9516 78364
rect 9516 78308 9572 78364
rect 9572 78308 9576 78364
rect 9512 78304 9576 78308
rect 9592 78364 9656 78368
rect 9592 78308 9596 78364
rect 9596 78308 9652 78364
rect 9652 78308 9656 78364
rect 9592 78304 9656 78308
rect 3612 77820 3676 77824
rect 3612 77764 3616 77820
rect 3616 77764 3672 77820
rect 3672 77764 3676 77820
rect 3612 77760 3676 77764
rect 3692 77820 3756 77824
rect 3692 77764 3696 77820
rect 3696 77764 3752 77820
rect 3752 77764 3756 77820
rect 3692 77760 3756 77764
rect 3772 77820 3836 77824
rect 3772 77764 3776 77820
rect 3776 77764 3832 77820
rect 3832 77764 3836 77820
rect 3772 77760 3836 77764
rect 3852 77820 3916 77824
rect 3852 77764 3856 77820
rect 3856 77764 3912 77820
rect 3912 77764 3916 77820
rect 3852 77760 3916 77764
rect 5212 77820 5276 77824
rect 5212 77764 5216 77820
rect 5216 77764 5272 77820
rect 5272 77764 5276 77820
rect 5212 77760 5276 77764
rect 5292 77820 5356 77824
rect 5292 77764 5296 77820
rect 5296 77764 5352 77820
rect 5352 77764 5356 77820
rect 5292 77760 5356 77764
rect 5372 77820 5436 77824
rect 5372 77764 5376 77820
rect 5376 77764 5432 77820
rect 5432 77764 5436 77820
rect 5372 77760 5436 77764
rect 5452 77820 5516 77824
rect 5452 77764 5456 77820
rect 5456 77764 5512 77820
rect 5512 77764 5516 77820
rect 5452 77760 5516 77764
rect 6812 77820 6876 77824
rect 6812 77764 6816 77820
rect 6816 77764 6872 77820
rect 6872 77764 6876 77820
rect 6812 77760 6876 77764
rect 6892 77820 6956 77824
rect 6892 77764 6896 77820
rect 6896 77764 6952 77820
rect 6952 77764 6956 77820
rect 6892 77760 6956 77764
rect 6972 77820 7036 77824
rect 6972 77764 6976 77820
rect 6976 77764 7032 77820
rect 7032 77764 7036 77820
rect 6972 77760 7036 77764
rect 7052 77820 7116 77824
rect 7052 77764 7056 77820
rect 7056 77764 7112 77820
rect 7112 77764 7116 77820
rect 7052 77760 7116 77764
rect 8412 77820 8476 77824
rect 8412 77764 8416 77820
rect 8416 77764 8472 77820
rect 8472 77764 8476 77820
rect 8412 77760 8476 77764
rect 8492 77820 8556 77824
rect 8492 77764 8496 77820
rect 8496 77764 8552 77820
rect 8552 77764 8556 77820
rect 8492 77760 8556 77764
rect 8572 77820 8636 77824
rect 8572 77764 8576 77820
rect 8576 77764 8632 77820
rect 8632 77764 8636 77820
rect 8572 77760 8636 77764
rect 8652 77820 8716 77824
rect 8652 77764 8656 77820
rect 8656 77764 8712 77820
rect 8712 77764 8716 77820
rect 8652 77760 8716 77764
rect 2952 77276 3016 77280
rect 2952 77220 2956 77276
rect 2956 77220 3012 77276
rect 3012 77220 3016 77276
rect 2952 77216 3016 77220
rect 3032 77276 3096 77280
rect 3032 77220 3036 77276
rect 3036 77220 3092 77276
rect 3092 77220 3096 77276
rect 3032 77216 3096 77220
rect 3112 77276 3176 77280
rect 3112 77220 3116 77276
rect 3116 77220 3172 77276
rect 3172 77220 3176 77276
rect 3112 77216 3176 77220
rect 3192 77276 3256 77280
rect 3192 77220 3196 77276
rect 3196 77220 3252 77276
rect 3252 77220 3256 77276
rect 3192 77216 3256 77220
rect 4552 77276 4616 77280
rect 4552 77220 4556 77276
rect 4556 77220 4612 77276
rect 4612 77220 4616 77276
rect 4552 77216 4616 77220
rect 4632 77276 4696 77280
rect 4632 77220 4636 77276
rect 4636 77220 4692 77276
rect 4692 77220 4696 77276
rect 4632 77216 4696 77220
rect 4712 77276 4776 77280
rect 4712 77220 4716 77276
rect 4716 77220 4772 77276
rect 4772 77220 4776 77276
rect 4712 77216 4776 77220
rect 4792 77276 4856 77280
rect 4792 77220 4796 77276
rect 4796 77220 4852 77276
rect 4852 77220 4856 77276
rect 4792 77216 4856 77220
rect 6152 77276 6216 77280
rect 6152 77220 6156 77276
rect 6156 77220 6212 77276
rect 6212 77220 6216 77276
rect 6152 77216 6216 77220
rect 6232 77276 6296 77280
rect 6232 77220 6236 77276
rect 6236 77220 6292 77276
rect 6292 77220 6296 77276
rect 6232 77216 6296 77220
rect 6312 77276 6376 77280
rect 6312 77220 6316 77276
rect 6316 77220 6372 77276
rect 6372 77220 6376 77276
rect 6312 77216 6376 77220
rect 6392 77276 6456 77280
rect 6392 77220 6396 77276
rect 6396 77220 6452 77276
rect 6452 77220 6456 77276
rect 6392 77216 6456 77220
rect 7752 77276 7816 77280
rect 7752 77220 7756 77276
rect 7756 77220 7812 77276
rect 7812 77220 7816 77276
rect 7752 77216 7816 77220
rect 7832 77276 7896 77280
rect 7832 77220 7836 77276
rect 7836 77220 7892 77276
rect 7892 77220 7896 77276
rect 7832 77216 7896 77220
rect 7912 77276 7976 77280
rect 7912 77220 7916 77276
rect 7916 77220 7972 77276
rect 7972 77220 7976 77276
rect 7912 77216 7976 77220
rect 7992 77276 8056 77280
rect 7992 77220 7996 77276
rect 7996 77220 8052 77276
rect 8052 77220 8056 77276
rect 7992 77216 8056 77220
rect 9352 77276 9416 77280
rect 9352 77220 9356 77276
rect 9356 77220 9412 77276
rect 9412 77220 9416 77276
rect 9352 77216 9416 77220
rect 9432 77276 9496 77280
rect 9432 77220 9436 77276
rect 9436 77220 9492 77276
rect 9492 77220 9496 77276
rect 9432 77216 9496 77220
rect 9512 77276 9576 77280
rect 9512 77220 9516 77276
rect 9516 77220 9572 77276
rect 9572 77220 9576 77276
rect 9512 77216 9576 77220
rect 9592 77276 9656 77280
rect 9592 77220 9596 77276
rect 9596 77220 9652 77276
rect 9652 77220 9656 77276
rect 9592 77216 9656 77220
rect 3612 76732 3676 76736
rect 3612 76676 3616 76732
rect 3616 76676 3672 76732
rect 3672 76676 3676 76732
rect 3612 76672 3676 76676
rect 3692 76732 3756 76736
rect 3692 76676 3696 76732
rect 3696 76676 3752 76732
rect 3752 76676 3756 76732
rect 3692 76672 3756 76676
rect 3772 76732 3836 76736
rect 3772 76676 3776 76732
rect 3776 76676 3832 76732
rect 3832 76676 3836 76732
rect 3772 76672 3836 76676
rect 3852 76732 3916 76736
rect 3852 76676 3856 76732
rect 3856 76676 3912 76732
rect 3912 76676 3916 76732
rect 3852 76672 3916 76676
rect 5212 76732 5276 76736
rect 5212 76676 5216 76732
rect 5216 76676 5272 76732
rect 5272 76676 5276 76732
rect 5212 76672 5276 76676
rect 5292 76732 5356 76736
rect 5292 76676 5296 76732
rect 5296 76676 5352 76732
rect 5352 76676 5356 76732
rect 5292 76672 5356 76676
rect 5372 76732 5436 76736
rect 5372 76676 5376 76732
rect 5376 76676 5432 76732
rect 5432 76676 5436 76732
rect 5372 76672 5436 76676
rect 5452 76732 5516 76736
rect 5452 76676 5456 76732
rect 5456 76676 5512 76732
rect 5512 76676 5516 76732
rect 5452 76672 5516 76676
rect 6812 76732 6876 76736
rect 6812 76676 6816 76732
rect 6816 76676 6872 76732
rect 6872 76676 6876 76732
rect 6812 76672 6876 76676
rect 6892 76732 6956 76736
rect 6892 76676 6896 76732
rect 6896 76676 6952 76732
rect 6952 76676 6956 76732
rect 6892 76672 6956 76676
rect 6972 76732 7036 76736
rect 6972 76676 6976 76732
rect 6976 76676 7032 76732
rect 7032 76676 7036 76732
rect 6972 76672 7036 76676
rect 7052 76732 7116 76736
rect 7052 76676 7056 76732
rect 7056 76676 7112 76732
rect 7112 76676 7116 76732
rect 7052 76672 7116 76676
rect 8412 76732 8476 76736
rect 8412 76676 8416 76732
rect 8416 76676 8472 76732
rect 8472 76676 8476 76732
rect 8412 76672 8476 76676
rect 8492 76732 8556 76736
rect 8492 76676 8496 76732
rect 8496 76676 8552 76732
rect 8552 76676 8556 76732
rect 8492 76672 8556 76676
rect 8572 76732 8636 76736
rect 8572 76676 8576 76732
rect 8576 76676 8632 76732
rect 8632 76676 8636 76732
rect 8572 76672 8636 76676
rect 8652 76732 8716 76736
rect 8652 76676 8656 76732
rect 8656 76676 8712 76732
rect 8712 76676 8716 76732
rect 8652 76672 8716 76676
rect 2952 76188 3016 76192
rect 2952 76132 2956 76188
rect 2956 76132 3012 76188
rect 3012 76132 3016 76188
rect 2952 76128 3016 76132
rect 3032 76188 3096 76192
rect 3032 76132 3036 76188
rect 3036 76132 3092 76188
rect 3092 76132 3096 76188
rect 3032 76128 3096 76132
rect 3112 76188 3176 76192
rect 3112 76132 3116 76188
rect 3116 76132 3172 76188
rect 3172 76132 3176 76188
rect 3112 76128 3176 76132
rect 3192 76188 3256 76192
rect 3192 76132 3196 76188
rect 3196 76132 3252 76188
rect 3252 76132 3256 76188
rect 3192 76128 3256 76132
rect 4552 76188 4616 76192
rect 4552 76132 4556 76188
rect 4556 76132 4612 76188
rect 4612 76132 4616 76188
rect 4552 76128 4616 76132
rect 4632 76188 4696 76192
rect 4632 76132 4636 76188
rect 4636 76132 4692 76188
rect 4692 76132 4696 76188
rect 4632 76128 4696 76132
rect 4712 76188 4776 76192
rect 4712 76132 4716 76188
rect 4716 76132 4772 76188
rect 4772 76132 4776 76188
rect 4712 76128 4776 76132
rect 4792 76188 4856 76192
rect 4792 76132 4796 76188
rect 4796 76132 4852 76188
rect 4852 76132 4856 76188
rect 4792 76128 4856 76132
rect 6152 76188 6216 76192
rect 6152 76132 6156 76188
rect 6156 76132 6212 76188
rect 6212 76132 6216 76188
rect 6152 76128 6216 76132
rect 6232 76188 6296 76192
rect 6232 76132 6236 76188
rect 6236 76132 6292 76188
rect 6292 76132 6296 76188
rect 6232 76128 6296 76132
rect 6312 76188 6376 76192
rect 6312 76132 6316 76188
rect 6316 76132 6372 76188
rect 6372 76132 6376 76188
rect 6312 76128 6376 76132
rect 6392 76188 6456 76192
rect 6392 76132 6396 76188
rect 6396 76132 6452 76188
rect 6452 76132 6456 76188
rect 6392 76128 6456 76132
rect 7752 76188 7816 76192
rect 7752 76132 7756 76188
rect 7756 76132 7812 76188
rect 7812 76132 7816 76188
rect 7752 76128 7816 76132
rect 7832 76188 7896 76192
rect 7832 76132 7836 76188
rect 7836 76132 7892 76188
rect 7892 76132 7896 76188
rect 7832 76128 7896 76132
rect 7912 76188 7976 76192
rect 7912 76132 7916 76188
rect 7916 76132 7972 76188
rect 7972 76132 7976 76188
rect 7912 76128 7976 76132
rect 7992 76188 8056 76192
rect 7992 76132 7996 76188
rect 7996 76132 8052 76188
rect 8052 76132 8056 76188
rect 7992 76128 8056 76132
rect 9352 76188 9416 76192
rect 9352 76132 9356 76188
rect 9356 76132 9412 76188
rect 9412 76132 9416 76188
rect 9352 76128 9416 76132
rect 9432 76188 9496 76192
rect 9432 76132 9436 76188
rect 9436 76132 9492 76188
rect 9492 76132 9496 76188
rect 9432 76128 9496 76132
rect 9512 76188 9576 76192
rect 9512 76132 9516 76188
rect 9516 76132 9572 76188
rect 9572 76132 9576 76188
rect 9512 76128 9576 76132
rect 9592 76188 9656 76192
rect 9592 76132 9596 76188
rect 9596 76132 9652 76188
rect 9652 76132 9656 76188
rect 9592 76128 9656 76132
rect 3612 75644 3676 75648
rect 3612 75588 3616 75644
rect 3616 75588 3672 75644
rect 3672 75588 3676 75644
rect 3612 75584 3676 75588
rect 3692 75644 3756 75648
rect 3692 75588 3696 75644
rect 3696 75588 3752 75644
rect 3752 75588 3756 75644
rect 3692 75584 3756 75588
rect 3772 75644 3836 75648
rect 3772 75588 3776 75644
rect 3776 75588 3832 75644
rect 3832 75588 3836 75644
rect 3772 75584 3836 75588
rect 3852 75644 3916 75648
rect 3852 75588 3856 75644
rect 3856 75588 3912 75644
rect 3912 75588 3916 75644
rect 3852 75584 3916 75588
rect 5212 75644 5276 75648
rect 5212 75588 5216 75644
rect 5216 75588 5272 75644
rect 5272 75588 5276 75644
rect 5212 75584 5276 75588
rect 5292 75644 5356 75648
rect 5292 75588 5296 75644
rect 5296 75588 5352 75644
rect 5352 75588 5356 75644
rect 5292 75584 5356 75588
rect 5372 75644 5436 75648
rect 5372 75588 5376 75644
rect 5376 75588 5432 75644
rect 5432 75588 5436 75644
rect 5372 75584 5436 75588
rect 5452 75644 5516 75648
rect 5452 75588 5456 75644
rect 5456 75588 5512 75644
rect 5512 75588 5516 75644
rect 5452 75584 5516 75588
rect 6812 75644 6876 75648
rect 6812 75588 6816 75644
rect 6816 75588 6872 75644
rect 6872 75588 6876 75644
rect 6812 75584 6876 75588
rect 6892 75644 6956 75648
rect 6892 75588 6896 75644
rect 6896 75588 6952 75644
rect 6952 75588 6956 75644
rect 6892 75584 6956 75588
rect 6972 75644 7036 75648
rect 6972 75588 6976 75644
rect 6976 75588 7032 75644
rect 7032 75588 7036 75644
rect 6972 75584 7036 75588
rect 7052 75644 7116 75648
rect 7052 75588 7056 75644
rect 7056 75588 7112 75644
rect 7112 75588 7116 75644
rect 7052 75584 7116 75588
rect 8412 75644 8476 75648
rect 8412 75588 8416 75644
rect 8416 75588 8472 75644
rect 8472 75588 8476 75644
rect 8412 75584 8476 75588
rect 8492 75644 8556 75648
rect 8492 75588 8496 75644
rect 8496 75588 8552 75644
rect 8552 75588 8556 75644
rect 8492 75584 8556 75588
rect 8572 75644 8636 75648
rect 8572 75588 8576 75644
rect 8576 75588 8632 75644
rect 8632 75588 8636 75644
rect 8572 75584 8636 75588
rect 8652 75644 8716 75648
rect 8652 75588 8656 75644
rect 8656 75588 8712 75644
rect 8712 75588 8716 75644
rect 8652 75584 8716 75588
rect 2952 75100 3016 75104
rect 2952 75044 2956 75100
rect 2956 75044 3012 75100
rect 3012 75044 3016 75100
rect 2952 75040 3016 75044
rect 3032 75100 3096 75104
rect 3032 75044 3036 75100
rect 3036 75044 3092 75100
rect 3092 75044 3096 75100
rect 3032 75040 3096 75044
rect 3112 75100 3176 75104
rect 3112 75044 3116 75100
rect 3116 75044 3172 75100
rect 3172 75044 3176 75100
rect 3112 75040 3176 75044
rect 3192 75100 3256 75104
rect 3192 75044 3196 75100
rect 3196 75044 3252 75100
rect 3252 75044 3256 75100
rect 3192 75040 3256 75044
rect 4552 75100 4616 75104
rect 4552 75044 4556 75100
rect 4556 75044 4612 75100
rect 4612 75044 4616 75100
rect 4552 75040 4616 75044
rect 4632 75100 4696 75104
rect 4632 75044 4636 75100
rect 4636 75044 4692 75100
rect 4692 75044 4696 75100
rect 4632 75040 4696 75044
rect 4712 75100 4776 75104
rect 4712 75044 4716 75100
rect 4716 75044 4772 75100
rect 4772 75044 4776 75100
rect 4712 75040 4776 75044
rect 4792 75100 4856 75104
rect 4792 75044 4796 75100
rect 4796 75044 4852 75100
rect 4852 75044 4856 75100
rect 4792 75040 4856 75044
rect 6152 75100 6216 75104
rect 6152 75044 6156 75100
rect 6156 75044 6212 75100
rect 6212 75044 6216 75100
rect 6152 75040 6216 75044
rect 6232 75100 6296 75104
rect 6232 75044 6236 75100
rect 6236 75044 6292 75100
rect 6292 75044 6296 75100
rect 6232 75040 6296 75044
rect 6312 75100 6376 75104
rect 6312 75044 6316 75100
rect 6316 75044 6372 75100
rect 6372 75044 6376 75100
rect 6312 75040 6376 75044
rect 6392 75100 6456 75104
rect 6392 75044 6396 75100
rect 6396 75044 6452 75100
rect 6452 75044 6456 75100
rect 6392 75040 6456 75044
rect 7752 75100 7816 75104
rect 7752 75044 7756 75100
rect 7756 75044 7812 75100
rect 7812 75044 7816 75100
rect 7752 75040 7816 75044
rect 7832 75100 7896 75104
rect 7832 75044 7836 75100
rect 7836 75044 7892 75100
rect 7892 75044 7896 75100
rect 7832 75040 7896 75044
rect 7912 75100 7976 75104
rect 7912 75044 7916 75100
rect 7916 75044 7972 75100
rect 7972 75044 7976 75100
rect 7912 75040 7976 75044
rect 7992 75100 8056 75104
rect 7992 75044 7996 75100
rect 7996 75044 8052 75100
rect 8052 75044 8056 75100
rect 7992 75040 8056 75044
rect 9352 75100 9416 75104
rect 9352 75044 9356 75100
rect 9356 75044 9412 75100
rect 9412 75044 9416 75100
rect 9352 75040 9416 75044
rect 9432 75100 9496 75104
rect 9432 75044 9436 75100
rect 9436 75044 9492 75100
rect 9492 75044 9496 75100
rect 9432 75040 9496 75044
rect 9512 75100 9576 75104
rect 9512 75044 9516 75100
rect 9516 75044 9572 75100
rect 9572 75044 9576 75100
rect 9512 75040 9576 75044
rect 9592 75100 9656 75104
rect 9592 75044 9596 75100
rect 9596 75044 9652 75100
rect 9652 75044 9656 75100
rect 9592 75040 9656 75044
rect 3612 74556 3676 74560
rect 3612 74500 3616 74556
rect 3616 74500 3672 74556
rect 3672 74500 3676 74556
rect 3612 74496 3676 74500
rect 3692 74556 3756 74560
rect 3692 74500 3696 74556
rect 3696 74500 3752 74556
rect 3752 74500 3756 74556
rect 3692 74496 3756 74500
rect 3772 74556 3836 74560
rect 3772 74500 3776 74556
rect 3776 74500 3832 74556
rect 3832 74500 3836 74556
rect 3772 74496 3836 74500
rect 3852 74556 3916 74560
rect 3852 74500 3856 74556
rect 3856 74500 3912 74556
rect 3912 74500 3916 74556
rect 3852 74496 3916 74500
rect 5212 74556 5276 74560
rect 5212 74500 5216 74556
rect 5216 74500 5272 74556
rect 5272 74500 5276 74556
rect 5212 74496 5276 74500
rect 5292 74556 5356 74560
rect 5292 74500 5296 74556
rect 5296 74500 5352 74556
rect 5352 74500 5356 74556
rect 5292 74496 5356 74500
rect 5372 74556 5436 74560
rect 5372 74500 5376 74556
rect 5376 74500 5432 74556
rect 5432 74500 5436 74556
rect 5372 74496 5436 74500
rect 5452 74556 5516 74560
rect 5452 74500 5456 74556
rect 5456 74500 5512 74556
rect 5512 74500 5516 74556
rect 5452 74496 5516 74500
rect 6812 74556 6876 74560
rect 6812 74500 6816 74556
rect 6816 74500 6872 74556
rect 6872 74500 6876 74556
rect 6812 74496 6876 74500
rect 6892 74556 6956 74560
rect 6892 74500 6896 74556
rect 6896 74500 6952 74556
rect 6952 74500 6956 74556
rect 6892 74496 6956 74500
rect 6972 74556 7036 74560
rect 6972 74500 6976 74556
rect 6976 74500 7032 74556
rect 7032 74500 7036 74556
rect 6972 74496 7036 74500
rect 7052 74556 7116 74560
rect 7052 74500 7056 74556
rect 7056 74500 7112 74556
rect 7112 74500 7116 74556
rect 7052 74496 7116 74500
rect 2952 74012 3016 74016
rect 2952 73956 2956 74012
rect 2956 73956 3012 74012
rect 3012 73956 3016 74012
rect 2952 73952 3016 73956
rect 3032 74012 3096 74016
rect 3032 73956 3036 74012
rect 3036 73956 3092 74012
rect 3092 73956 3096 74012
rect 3032 73952 3096 73956
rect 3112 74012 3176 74016
rect 3112 73956 3116 74012
rect 3116 73956 3172 74012
rect 3172 73956 3176 74012
rect 3112 73952 3176 73956
rect 3192 74012 3256 74016
rect 3192 73956 3196 74012
rect 3196 73956 3252 74012
rect 3252 73956 3256 74012
rect 3192 73952 3256 73956
rect 4552 74012 4616 74016
rect 4552 73956 4556 74012
rect 4556 73956 4612 74012
rect 4612 73956 4616 74012
rect 4552 73952 4616 73956
rect 4632 74012 4696 74016
rect 4632 73956 4636 74012
rect 4636 73956 4692 74012
rect 4692 73956 4696 74012
rect 4632 73952 4696 73956
rect 4712 74012 4776 74016
rect 4712 73956 4716 74012
rect 4716 73956 4772 74012
rect 4772 73956 4776 74012
rect 4712 73952 4776 73956
rect 4792 74012 4856 74016
rect 4792 73956 4796 74012
rect 4796 73956 4852 74012
rect 4852 73956 4856 74012
rect 4792 73952 4856 73956
rect 6152 74012 6216 74016
rect 6152 73956 6156 74012
rect 6156 73956 6212 74012
rect 6212 73956 6216 74012
rect 6152 73952 6216 73956
rect 6232 74012 6296 74016
rect 6232 73956 6236 74012
rect 6236 73956 6292 74012
rect 6292 73956 6296 74012
rect 6232 73952 6296 73956
rect 6312 74012 6376 74016
rect 6312 73956 6316 74012
rect 6316 73956 6372 74012
rect 6372 73956 6376 74012
rect 6312 73952 6376 73956
rect 6392 74012 6456 74016
rect 6392 73956 6396 74012
rect 6396 73956 6452 74012
rect 6452 73956 6456 74012
rect 6392 73952 6456 73956
rect 8412 74556 8476 74560
rect 8412 74500 8416 74556
rect 8416 74500 8472 74556
rect 8472 74500 8476 74556
rect 8412 74496 8476 74500
rect 8492 74556 8556 74560
rect 8492 74500 8496 74556
rect 8496 74500 8552 74556
rect 8552 74500 8556 74556
rect 8492 74496 8556 74500
rect 8572 74556 8636 74560
rect 8572 74500 8576 74556
rect 8576 74500 8632 74556
rect 8632 74500 8636 74556
rect 8572 74496 8636 74500
rect 8652 74556 8716 74560
rect 8652 74500 8656 74556
rect 8656 74500 8712 74556
rect 8712 74500 8716 74556
rect 8652 74496 8716 74500
rect 10916 74292 10980 74356
rect 7752 74012 7816 74016
rect 7752 73956 7756 74012
rect 7756 73956 7812 74012
rect 7812 73956 7816 74012
rect 7752 73952 7816 73956
rect 7832 74012 7896 74016
rect 7832 73956 7836 74012
rect 7836 73956 7892 74012
rect 7892 73956 7896 74012
rect 7832 73952 7896 73956
rect 7912 74012 7976 74016
rect 7912 73956 7916 74012
rect 7916 73956 7972 74012
rect 7972 73956 7976 74012
rect 7912 73952 7976 73956
rect 7992 74012 8056 74016
rect 7992 73956 7996 74012
rect 7996 73956 8052 74012
rect 8052 73956 8056 74012
rect 7992 73952 8056 73956
rect 9352 74012 9416 74016
rect 9352 73956 9356 74012
rect 9356 73956 9412 74012
rect 9412 73956 9416 74012
rect 9352 73952 9416 73956
rect 9432 74012 9496 74016
rect 9432 73956 9436 74012
rect 9436 73956 9492 74012
rect 9492 73956 9496 74012
rect 9432 73952 9496 73956
rect 9512 74012 9576 74016
rect 9512 73956 9516 74012
rect 9516 73956 9572 74012
rect 9572 73956 9576 74012
rect 9512 73952 9576 73956
rect 9592 74012 9656 74016
rect 9592 73956 9596 74012
rect 9596 73956 9652 74012
rect 9652 73956 9656 74012
rect 9592 73952 9656 73956
rect 3612 73468 3676 73472
rect 3612 73412 3616 73468
rect 3616 73412 3672 73468
rect 3672 73412 3676 73468
rect 3612 73408 3676 73412
rect 3692 73468 3756 73472
rect 3692 73412 3696 73468
rect 3696 73412 3752 73468
rect 3752 73412 3756 73468
rect 3692 73408 3756 73412
rect 3772 73468 3836 73472
rect 3772 73412 3776 73468
rect 3776 73412 3832 73468
rect 3832 73412 3836 73468
rect 3772 73408 3836 73412
rect 3852 73468 3916 73472
rect 3852 73412 3856 73468
rect 3856 73412 3912 73468
rect 3912 73412 3916 73468
rect 3852 73408 3916 73412
rect 5212 73468 5276 73472
rect 5212 73412 5216 73468
rect 5216 73412 5272 73468
rect 5272 73412 5276 73468
rect 5212 73408 5276 73412
rect 5292 73468 5356 73472
rect 5292 73412 5296 73468
rect 5296 73412 5352 73468
rect 5352 73412 5356 73468
rect 5292 73408 5356 73412
rect 5372 73468 5436 73472
rect 5372 73412 5376 73468
rect 5376 73412 5432 73468
rect 5432 73412 5436 73468
rect 5372 73408 5436 73412
rect 5452 73468 5516 73472
rect 5452 73412 5456 73468
rect 5456 73412 5512 73468
rect 5512 73412 5516 73468
rect 5452 73408 5516 73412
rect 6812 73468 6876 73472
rect 6812 73412 6816 73468
rect 6816 73412 6872 73468
rect 6872 73412 6876 73468
rect 6812 73408 6876 73412
rect 6892 73468 6956 73472
rect 6892 73412 6896 73468
rect 6896 73412 6952 73468
rect 6952 73412 6956 73468
rect 6892 73408 6956 73412
rect 6972 73468 7036 73472
rect 6972 73412 6976 73468
rect 6976 73412 7032 73468
rect 7032 73412 7036 73468
rect 6972 73408 7036 73412
rect 7052 73468 7116 73472
rect 7052 73412 7056 73468
rect 7056 73412 7112 73468
rect 7112 73412 7116 73468
rect 7052 73408 7116 73412
rect 8412 73468 8476 73472
rect 8412 73412 8416 73468
rect 8416 73412 8472 73468
rect 8472 73412 8476 73468
rect 8412 73408 8476 73412
rect 8492 73468 8556 73472
rect 8492 73412 8496 73468
rect 8496 73412 8552 73468
rect 8552 73412 8556 73468
rect 8492 73408 8556 73412
rect 8572 73468 8636 73472
rect 8572 73412 8576 73468
rect 8576 73412 8632 73468
rect 8632 73412 8636 73468
rect 8572 73408 8636 73412
rect 8652 73468 8716 73472
rect 8652 73412 8656 73468
rect 8656 73412 8712 73468
rect 8712 73412 8716 73468
rect 8652 73408 8716 73412
rect 2952 72924 3016 72928
rect 2952 72868 2956 72924
rect 2956 72868 3012 72924
rect 3012 72868 3016 72924
rect 2952 72864 3016 72868
rect 3032 72924 3096 72928
rect 3032 72868 3036 72924
rect 3036 72868 3092 72924
rect 3092 72868 3096 72924
rect 3032 72864 3096 72868
rect 3112 72924 3176 72928
rect 3112 72868 3116 72924
rect 3116 72868 3172 72924
rect 3172 72868 3176 72924
rect 3112 72864 3176 72868
rect 3192 72924 3256 72928
rect 3192 72868 3196 72924
rect 3196 72868 3252 72924
rect 3252 72868 3256 72924
rect 3192 72864 3256 72868
rect 4552 72924 4616 72928
rect 4552 72868 4556 72924
rect 4556 72868 4612 72924
rect 4612 72868 4616 72924
rect 4552 72864 4616 72868
rect 4632 72924 4696 72928
rect 4632 72868 4636 72924
rect 4636 72868 4692 72924
rect 4692 72868 4696 72924
rect 4632 72864 4696 72868
rect 4712 72924 4776 72928
rect 4712 72868 4716 72924
rect 4716 72868 4772 72924
rect 4772 72868 4776 72924
rect 4712 72864 4776 72868
rect 4792 72924 4856 72928
rect 4792 72868 4796 72924
rect 4796 72868 4852 72924
rect 4852 72868 4856 72924
rect 4792 72864 4856 72868
rect 6152 72924 6216 72928
rect 6152 72868 6156 72924
rect 6156 72868 6212 72924
rect 6212 72868 6216 72924
rect 6152 72864 6216 72868
rect 6232 72924 6296 72928
rect 6232 72868 6236 72924
rect 6236 72868 6292 72924
rect 6292 72868 6296 72924
rect 6232 72864 6296 72868
rect 6312 72924 6376 72928
rect 6312 72868 6316 72924
rect 6316 72868 6372 72924
rect 6372 72868 6376 72924
rect 6312 72864 6376 72868
rect 6392 72924 6456 72928
rect 6392 72868 6396 72924
rect 6396 72868 6452 72924
rect 6452 72868 6456 72924
rect 6392 72864 6456 72868
rect 7752 72924 7816 72928
rect 7752 72868 7756 72924
rect 7756 72868 7812 72924
rect 7812 72868 7816 72924
rect 7752 72864 7816 72868
rect 7832 72924 7896 72928
rect 7832 72868 7836 72924
rect 7836 72868 7892 72924
rect 7892 72868 7896 72924
rect 7832 72864 7896 72868
rect 7912 72924 7976 72928
rect 7912 72868 7916 72924
rect 7916 72868 7972 72924
rect 7972 72868 7976 72924
rect 7912 72864 7976 72868
rect 7992 72924 8056 72928
rect 7992 72868 7996 72924
rect 7996 72868 8052 72924
rect 8052 72868 8056 72924
rect 7992 72864 8056 72868
rect 9352 72924 9416 72928
rect 9352 72868 9356 72924
rect 9356 72868 9412 72924
rect 9412 72868 9416 72924
rect 9352 72864 9416 72868
rect 9432 72924 9496 72928
rect 9432 72868 9436 72924
rect 9436 72868 9492 72924
rect 9492 72868 9496 72924
rect 9432 72864 9496 72868
rect 9512 72924 9576 72928
rect 9512 72868 9516 72924
rect 9516 72868 9572 72924
rect 9572 72868 9576 72924
rect 9512 72864 9576 72868
rect 9592 72924 9656 72928
rect 9592 72868 9596 72924
rect 9596 72868 9652 72924
rect 9652 72868 9656 72924
rect 9592 72864 9656 72868
rect 3612 72380 3676 72384
rect 3612 72324 3616 72380
rect 3616 72324 3672 72380
rect 3672 72324 3676 72380
rect 3612 72320 3676 72324
rect 3692 72380 3756 72384
rect 3692 72324 3696 72380
rect 3696 72324 3752 72380
rect 3752 72324 3756 72380
rect 3692 72320 3756 72324
rect 3772 72380 3836 72384
rect 3772 72324 3776 72380
rect 3776 72324 3832 72380
rect 3832 72324 3836 72380
rect 3772 72320 3836 72324
rect 3852 72380 3916 72384
rect 3852 72324 3856 72380
rect 3856 72324 3912 72380
rect 3912 72324 3916 72380
rect 3852 72320 3916 72324
rect 5212 72380 5276 72384
rect 5212 72324 5216 72380
rect 5216 72324 5272 72380
rect 5272 72324 5276 72380
rect 5212 72320 5276 72324
rect 5292 72380 5356 72384
rect 5292 72324 5296 72380
rect 5296 72324 5352 72380
rect 5352 72324 5356 72380
rect 5292 72320 5356 72324
rect 5372 72380 5436 72384
rect 5372 72324 5376 72380
rect 5376 72324 5432 72380
rect 5432 72324 5436 72380
rect 5372 72320 5436 72324
rect 5452 72380 5516 72384
rect 5452 72324 5456 72380
rect 5456 72324 5512 72380
rect 5512 72324 5516 72380
rect 5452 72320 5516 72324
rect 6812 72380 6876 72384
rect 6812 72324 6816 72380
rect 6816 72324 6872 72380
rect 6872 72324 6876 72380
rect 6812 72320 6876 72324
rect 6892 72380 6956 72384
rect 6892 72324 6896 72380
rect 6896 72324 6952 72380
rect 6952 72324 6956 72380
rect 6892 72320 6956 72324
rect 6972 72380 7036 72384
rect 6972 72324 6976 72380
rect 6976 72324 7032 72380
rect 7032 72324 7036 72380
rect 6972 72320 7036 72324
rect 7052 72380 7116 72384
rect 7052 72324 7056 72380
rect 7056 72324 7112 72380
rect 7112 72324 7116 72380
rect 7052 72320 7116 72324
rect 8412 72380 8476 72384
rect 8412 72324 8416 72380
rect 8416 72324 8472 72380
rect 8472 72324 8476 72380
rect 8412 72320 8476 72324
rect 8492 72380 8556 72384
rect 8492 72324 8496 72380
rect 8496 72324 8552 72380
rect 8552 72324 8556 72380
rect 8492 72320 8556 72324
rect 8572 72380 8636 72384
rect 8572 72324 8576 72380
rect 8576 72324 8632 72380
rect 8632 72324 8636 72380
rect 8572 72320 8636 72324
rect 8652 72380 8716 72384
rect 8652 72324 8656 72380
rect 8656 72324 8712 72380
rect 8712 72324 8716 72380
rect 8652 72320 8716 72324
rect 796 71844 860 71908
rect 2952 71836 3016 71840
rect 2952 71780 2956 71836
rect 2956 71780 3012 71836
rect 3012 71780 3016 71836
rect 2952 71776 3016 71780
rect 3032 71836 3096 71840
rect 3032 71780 3036 71836
rect 3036 71780 3092 71836
rect 3092 71780 3096 71836
rect 3032 71776 3096 71780
rect 3112 71836 3176 71840
rect 3112 71780 3116 71836
rect 3116 71780 3172 71836
rect 3172 71780 3176 71836
rect 3112 71776 3176 71780
rect 3192 71836 3256 71840
rect 3192 71780 3196 71836
rect 3196 71780 3252 71836
rect 3252 71780 3256 71836
rect 3192 71776 3256 71780
rect 4552 71836 4616 71840
rect 4552 71780 4556 71836
rect 4556 71780 4612 71836
rect 4612 71780 4616 71836
rect 4552 71776 4616 71780
rect 4632 71836 4696 71840
rect 4632 71780 4636 71836
rect 4636 71780 4692 71836
rect 4692 71780 4696 71836
rect 4632 71776 4696 71780
rect 4712 71836 4776 71840
rect 4712 71780 4716 71836
rect 4716 71780 4772 71836
rect 4772 71780 4776 71836
rect 4712 71776 4776 71780
rect 4792 71836 4856 71840
rect 4792 71780 4796 71836
rect 4796 71780 4852 71836
rect 4852 71780 4856 71836
rect 4792 71776 4856 71780
rect 6152 71836 6216 71840
rect 6152 71780 6156 71836
rect 6156 71780 6212 71836
rect 6212 71780 6216 71836
rect 6152 71776 6216 71780
rect 6232 71836 6296 71840
rect 6232 71780 6236 71836
rect 6236 71780 6292 71836
rect 6292 71780 6296 71836
rect 6232 71776 6296 71780
rect 6312 71836 6376 71840
rect 6312 71780 6316 71836
rect 6316 71780 6372 71836
rect 6372 71780 6376 71836
rect 6312 71776 6376 71780
rect 6392 71836 6456 71840
rect 6392 71780 6396 71836
rect 6396 71780 6452 71836
rect 6452 71780 6456 71836
rect 6392 71776 6456 71780
rect 7752 71836 7816 71840
rect 7752 71780 7756 71836
rect 7756 71780 7812 71836
rect 7812 71780 7816 71836
rect 7752 71776 7816 71780
rect 7832 71836 7896 71840
rect 7832 71780 7836 71836
rect 7836 71780 7892 71836
rect 7892 71780 7896 71836
rect 7832 71776 7896 71780
rect 7912 71836 7976 71840
rect 7912 71780 7916 71836
rect 7916 71780 7972 71836
rect 7972 71780 7976 71836
rect 7912 71776 7976 71780
rect 7992 71836 8056 71840
rect 7992 71780 7996 71836
rect 7996 71780 8052 71836
rect 8052 71780 8056 71836
rect 7992 71776 8056 71780
rect 9352 71836 9416 71840
rect 9352 71780 9356 71836
rect 9356 71780 9412 71836
rect 9412 71780 9416 71836
rect 9352 71776 9416 71780
rect 9432 71836 9496 71840
rect 9432 71780 9436 71836
rect 9436 71780 9492 71836
rect 9492 71780 9496 71836
rect 9432 71776 9496 71780
rect 9512 71836 9576 71840
rect 9512 71780 9516 71836
rect 9516 71780 9572 71836
rect 9572 71780 9576 71836
rect 9512 71776 9576 71780
rect 9592 71836 9656 71840
rect 9592 71780 9596 71836
rect 9596 71780 9652 71836
rect 9652 71780 9656 71836
rect 9592 71776 9656 71780
rect 3612 71292 3676 71296
rect 3612 71236 3616 71292
rect 3616 71236 3672 71292
rect 3672 71236 3676 71292
rect 3612 71232 3676 71236
rect 3692 71292 3756 71296
rect 3692 71236 3696 71292
rect 3696 71236 3752 71292
rect 3752 71236 3756 71292
rect 3692 71232 3756 71236
rect 3772 71292 3836 71296
rect 3772 71236 3776 71292
rect 3776 71236 3832 71292
rect 3832 71236 3836 71292
rect 3772 71232 3836 71236
rect 3852 71292 3916 71296
rect 3852 71236 3856 71292
rect 3856 71236 3912 71292
rect 3912 71236 3916 71292
rect 3852 71232 3916 71236
rect 5212 71292 5276 71296
rect 5212 71236 5216 71292
rect 5216 71236 5272 71292
rect 5272 71236 5276 71292
rect 5212 71232 5276 71236
rect 5292 71292 5356 71296
rect 5292 71236 5296 71292
rect 5296 71236 5352 71292
rect 5352 71236 5356 71292
rect 5292 71232 5356 71236
rect 5372 71292 5436 71296
rect 5372 71236 5376 71292
rect 5376 71236 5432 71292
rect 5432 71236 5436 71292
rect 5372 71232 5436 71236
rect 5452 71292 5516 71296
rect 5452 71236 5456 71292
rect 5456 71236 5512 71292
rect 5512 71236 5516 71292
rect 5452 71232 5516 71236
rect 6812 71292 6876 71296
rect 6812 71236 6816 71292
rect 6816 71236 6872 71292
rect 6872 71236 6876 71292
rect 6812 71232 6876 71236
rect 6892 71292 6956 71296
rect 6892 71236 6896 71292
rect 6896 71236 6952 71292
rect 6952 71236 6956 71292
rect 6892 71232 6956 71236
rect 6972 71292 7036 71296
rect 6972 71236 6976 71292
rect 6976 71236 7032 71292
rect 7032 71236 7036 71292
rect 6972 71232 7036 71236
rect 7052 71292 7116 71296
rect 7052 71236 7056 71292
rect 7056 71236 7112 71292
rect 7112 71236 7116 71292
rect 7052 71232 7116 71236
rect 8412 71292 8476 71296
rect 8412 71236 8416 71292
rect 8416 71236 8472 71292
rect 8472 71236 8476 71292
rect 8412 71232 8476 71236
rect 8492 71292 8556 71296
rect 8492 71236 8496 71292
rect 8496 71236 8552 71292
rect 8552 71236 8556 71292
rect 8492 71232 8556 71236
rect 8572 71292 8636 71296
rect 8572 71236 8576 71292
rect 8576 71236 8632 71292
rect 8632 71236 8636 71292
rect 8572 71232 8636 71236
rect 8652 71292 8716 71296
rect 8652 71236 8656 71292
rect 8656 71236 8712 71292
rect 8712 71236 8716 71292
rect 8652 71232 8716 71236
rect 2952 70748 3016 70752
rect 2952 70692 2956 70748
rect 2956 70692 3012 70748
rect 3012 70692 3016 70748
rect 2952 70688 3016 70692
rect 3032 70748 3096 70752
rect 3032 70692 3036 70748
rect 3036 70692 3092 70748
rect 3092 70692 3096 70748
rect 3032 70688 3096 70692
rect 3112 70748 3176 70752
rect 3112 70692 3116 70748
rect 3116 70692 3172 70748
rect 3172 70692 3176 70748
rect 3112 70688 3176 70692
rect 3192 70748 3256 70752
rect 3192 70692 3196 70748
rect 3196 70692 3252 70748
rect 3252 70692 3256 70748
rect 3192 70688 3256 70692
rect 4552 70748 4616 70752
rect 4552 70692 4556 70748
rect 4556 70692 4612 70748
rect 4612 70692 4616 70748
rect 4552 70688 4616 70692
rect 4632 70748 4696 70752
rect 4632 70692 4636 70748
rect 4636 70692 4692 70748
rect 4692 70692 4696 70748
rect 4632 70688 4696 70692
rect 4712 70748 4776 70752
rect 4712 70692 4716 70748
rect 4716 70692 4772 70748
rect 4772 70692 4776 70748
rect 4712 70688 4776 70692
rect 4792 70748 4856 70752
rect 4792 70692 4796 70748
rect 4796 70692 4852 70748
rect 4852 70692 4856 70748
rect 4792 70688 4856 70692
rect 6152 70748 6216 70752
rect 6152 70692 6156 70748
rect 6156 70692 6212 70748
rect 6212 70692 6216 70748
rect 6152 70688 6216 70692
rect 6232 70748 6296 70752
rect 6232 70692 6236 70748
rect 6236 70692 6292 70748
rect 6292 70692 6296 70748
rect 6232 70688 6296 70692
rect 6312 70748 6376 70752
rect 6312 70692 6316 70748
rect 6316 70692 6372 70748
rect 6372 70692 6376 70748
rect 6312 70688 6376 70692
rect 6392 70748 6456 70752
rect 6392 70692 6396 70748
rect 6396 70692 6452 70748
rect 6452 70692 6456 70748
rect 6392 70688 6456 70692
rect 7752 70748 7816 70752
rect 7752 70692 7756 70748
rect 7756 70692 7812 70748
rect 7812 70692 7816 70748
rect 7752 70688 7816 70692
rect 7832 70748 7896 70752
rect 7832 70692 7836 70748
rect 7836 70692 7892 70748
rect 7892 70692 7896 70748
rect 7832 70688 7896 70692
rect 7912 70748 7976 70752
rect 7912 70692 7916 70748
rect 7916 70692 7972 70748
rect 7972 70692 7976 70748
rect 7912 70688 7976 70692
rect 7992 70748 8056 70752
rect 7992 70692 7996 70748
rect 7996 70692 8052 70748
rect 8052 70692 8056 70748
rect 7992 70688 8056 70692
rect 3612 70204 3676 70208
rect 3612 70148 3616 70204
rect 3616 70148 3672 70204
rect 3672 70148 3676 70204
rect 3612 70144 3676 70148
rect 3692 70204 3756 70208
rect 3692 70148 3696 70204
rect 3696 70148 3752 70204
rect 3752 70148 3756 70204
rect 3692 70144 3756 70148
rect 3772 70204 3836 70208
rect 3772 70148 3776 70204
rect 3776 70148 3832 70204
rect 3832 70148 3836 70204
rect 3772 70144 3836 70148
rect 3852 70204 3916 70208
rect 3852 70148 3856 70204
rect 3856 70148 3912 70204
rect 3912 70148 3916 70204
rect 3852 70144 3916 70148
rect 5212 70204 5276 70208
rect 5212 70148 5216 70204
rect 5216 70148 5272 70204
rect 5272 70148 5276 70204
rect 5212 70144 5276 70148
rect 5292 70204 5356 70208
rect 5292 70148 5296 70204
rect 5296 70148 5352 70204
rect 5352 70148 5356 70204
rect 5292 70144 5356 70148
rect 5372 70204 5436 70208
rect 5372 70148 5376 70204
rect 5376 70148 5432 70204
rect 5432 70148 5436 70204
rect 5372 70144 5436 70148
rect 5452 70204 5516 70208
rect 5452 70148 5456 70204
rect 5456 70148 5512 70204
rect 5512 70148 5516 70204
rect 5452 70144 5516 70148
rect 6812 70204 6876 70208
rect 6812 70148 6816 70204
rect 6816 70148 6872 70204
rect 6872 70148 6876 70204
rect 6812 70144 6876 70148
rect 6892 70204 6956 70208
rect 6892 70148 6896 70204
rect 6896 70148 6952 70204
rect 6952 70148 6956 70204
rect 6892 70144 6956 70148
rect 6972 70204 7036 70208
rect 6972 70148 6976 70204
rect 6976 70148 7032 70204
rect 7032 70148 7036 70204
rect 6972 70144 7036 70148
rect 7052 70204 7116 70208
rect 7052 70148 7056 70204
rect 7056 70148 7112 70204
rect 7112 70148 7116 70204
rect 7052 70144 7116 70148
rect 8412 70204 8476 70208
rect 8412 70148 8416 70204
rect 8416 70148 8472 70204
rect 8472 70148 8476 70204
rect 8412 70144 8476 70148
rect 8492 70204 8556 70208
rect 8492 70148 8496 70204
rect 8496 70148 8552 70204
rect 8552 70148 8556 70204
rect 8492 70144 8556 70148
rect 8572 70204 8636 70208
rect 8572 70148 8576 70204
rect 8576 70148 8632 70204
rect 8632 70148 8636 70204
rect 8572 70144 8636 70148
rect 8652 70204 8716 70208
rect 8652 70148 8656 70204
rect 8656 70148 8712 70204
rect 8712 70148 8716 70204
rect 8652 70144 8716 70148
rect 9352 70748 9416 70752
rect 9352 70692 9356 70748
rect 9356 70692 9412 70748
rect 9412 70692 9416 70748
rect 9352 70688 9416 70692
rect 9432 70748 9496 70752
rect 9432 70692 9436 70748
rect 9436 70692 9492 70748
rect 9492 70692 9496 70748
rect 9432 70688 9496 70692
rect 9512 70748 9576 70752
rect 9512 70692 9516 70748
rect 9516 70692 9572 70748
rect 9572 70692 9576 70748
rect 9512 70688 9576 70692
rect 9592 70748 9656 70752
rect 9592 70692 9596 70748
rect 9596 70692 9652 70748
rect 9652 70692 9656 70748
rect 9592 70688 9656 70692
rect 10548 69804 10612 69868
rect 2952 69660 3016 69664
rect 2952 69604 2956 69660
rect 2956 69604 3012 69660
rect 3012 69604 3016 69660
rect 2952 69600 3016 69604
rect 3032 69660 3096 69664
rect 3032 69604 3036 69660
rect 3036 69604 3092 69660
rect 3092 69604 3096 69660
rect 3032 69600 3096 69604
rect 3112 69660 3176 69664
rect 3112 69604 3116 69660
rect 3116 69604 3172 69660
rect 3172 69604 3176 69660
rect 3112 69600 3176 69604
rect 3192 69660 3256 69664
rect 3192 69604 3196 69660
rect 3196 69604 3252 69660
rect 3252 69604 3256 69660
rect 3192 69600 3256 69604
rect 4552 69660 4616 69664
rect 4552 69604 4556 69660
rect 4556 69604 4612 69660
rect 4612 69604 4616 69660
rect 4552 69600 4616 69604
rect 4632 69660 4696 69664
rect 4632 69604 4636 69660
rect 4636 69604 4692 69660
rect 4692 69604 4696 69660
rect 4632 69600 4696 69604
rect 4712 69660 4776 69664
rect 4712 69604 4716 69660
rect 4716 69604 4772 69660
rect 4772 69604 4776 69660
rect 4712 69600 4776 69604
rect 4792 69660 4856 69664
rect 4792 69604 4796 69660
rect 4796 69604 4852 69660
rect 4852 69604 4856 69660
rect 4792 69600 4856 69604
rect 6152 69660 6216 69664
rect 6152 69604 6156 69660
rect 6156 69604 6212 69660
rect 6212 69604 6216 69660
rect 6152 69600 6216 69604
rect 6232 69660 6296 69664
rect 6232 69604 6236 69660
rect 6236 69604 6292 69660
rect 6292 69604 6296 69660
rect 6232 69600 6296 69604
rect 6312 69660 6376 69664
rect 6312 69604 6316 69660
rect 6316 69604 6372 69660
rect 6372 69604 6376 69660
rect 6312 69600 6376 69604
rect 6392 69660 6456 69664
rect 6392 69604 6396 69660
rect 6396 69604 6452 69660
rect 6452 69604 6456 69660
rect 6392 69600 6456 69604
rect 7752 69660 7816 69664
rect 7752 69604 7756 69660
rect 7756 69604 7812 69660
rect 7812 69604 7816 69660
rect 7752 69600 7816 69604
rect 7832 69660 7896 69664
rect 7832 69604 7836 69660
rect 7836 69604 7892 69660
rect 7892 69604 7896 69660
rect 7832 69600 7896 69604
rect 7912 69660 7976 69664
rect 7912 69604 7916 69660
rect 7916 69604 7972 69660
rect 7972 69604 7976 69660
rect 7912 69600 7976 69604
rect 7992 69660 8056 69664
rect 7992 69604 7996 69660
rect 7996 69604 8052 69660
rect 8052 69604 8056 69660
rect 7992 69600 8056 69604
rect 9352 69660 9416 69664
rect 9352 69604 9356 69660
rect 9356 69604 9412 69660
rect 9412 69604 9416 69660
rect 9352 69600 9416 69604
rect 9432 69660 9496 69664
rect 9432 69604 9436 69660
rect 9436 69604 9492 69660
rect 9492 69604 9496 69660
rect 9432 69600 9496 69604
rect 9512 69660 9576 69664
rect 9512 69604 9516 69660
rect 9516 69604 9572 69660
rect 9572 69604 9576 69660
rect 9512 69600 9576 69604
rect 9592 69660 9656 69664
rect 9592 69604 9596 69660
rect 9596 69604 9652 69660
rect 9652 69604 9656 69660
rect 9592 69600 9656 69604
rect 11100 69396 11164 69460
rect 3612 69116 3676 69120
rect 3612 69060 3616 69116
rect 3616 69060 3672 69116
rect 3672 69060 3676 69116
rect 3612 69056 3676 69060
rect 3692 69116 3756 69120
rect 3692 69060 3696 69116
rect 3696 69060 3752 69116
rect 3752 69060 3756 69116
rect 3692 69056 3756 69060
rect 3772 69116 3836 69120
rect 3772 69060 3776 69116
rect 3776 69060 3832 69116
rect 3832 69060 3836 69116
rect 3772 69056 3836 69060
rect 3852 69116 3916 69120
rect 3852 69060 3856 69116
rect 3856 69060 3912 69116
rect 3912 69060 3916 69116
rect 3852 69056 3916 69060
rect 5212 69116 5276 69120
rect 5212 69060 5216 69116
rect 5216 69060 5272 69116
rect 5272 69060 5276 69116
rect 5212 69056 5276 69060
rect 5292 69116 5356 69120
rect 5292 69060 5296 69116
rect 5296 69060 5352 69116
rect 5352 69060 5356 69116
rect 5292 69056 5356 69060
rect 5372 69116 5436 69120
rect 5372 69060 5376 69116
rect 5376 69060 5432 69116
rect 5432 69060 5436 69116
rect 5372 69056 5436 69060
rect 5452 69116 5516 69120
rect 5452 69060 5456 69116
rect 5456 69060 5512 69116
rect 5512 69060 5516 69116
rect 5452 69056 5516 69060
rect 6812 69116 6876 69120
rect 6812 69060 6816 69116
rect 6816 69060 6872 69116
rect 6872 69060 6876 69116
rect 6812 69056 6876 69060
rect 6892 69116 6956 69120
rect 6892 69060 6896 69116
rect 6896 69060 6952 69116
rect 6952 69060 6956 69116
rect 6892 69056 6956 69060
rect 6972 69116 7036 69120
rect 6972 69060 6976 69116
rect 6976 69060 7032 69116
rect 7032 69060 7036 69116
rect 6972 69056 7036 69060
rect 7052 69116 7116 69120
rect 7052 69060 7056 69116
rect 7056 69060 7112 69116
rect 7112 69060 7116 69116
rect 7052 69056 7116 69060
rect 8412 69116 8476 69120
rect 8412 69060 8416 69116
rect 8416 69060 8472 69116
rect 8472 69060 8476 69116
rect 8412 69056 8476 69060
rect 8492 69116 8556 69120
rect 8492 69060 8496 69116
rect 8496 69060 8552 69116
rect 8552 69060 8556 69116
rect 8492 69056 8556 69060
rect 8572 69116 8636 69120
rect 8572 69060 8576 69116
rect 8576 69060 8632 69116
rect 8632 69060 8636 69116
rect 8572 69056 8636 69060
rect 8652 69116 8716 69120
rect 8652 69060 8656 69116
rect 8656 69060 8712 69116
rect 8712 69060 8716 69116
rect 8652 69056 8716 69060
rect 11468 68852 11532 68916
rect 2952 68572 3016 68576
rect 2952 68516 2956 68572
rect 2956 68516 3012 68572
rect 3012 68516 3016 68572
rect 2952 68512 3016 68516
rect 3032 68572 3096 68576
rect 3032 68516 3036 68572
rect 3036 68516 3092 68572
rect 3092 68516 3096 68572
rect 3032 68512 3096 68516
rect 3112 68572 3176 68576
rect 3112 68516 3116 68572
rect 3116 68516 3172 68572
rect 3172 68516 3176 68572
rect 3112 68512 3176 68516
rect 3192 68572 3256 68576
rect 3192 68516 3196 68572
rect 3196 68516 3252 68572
rect 3252 68516 3256 68572
rect 3192 68512 3256 68516
rect 4552 68572 4616 68576
rect 4552 68516 4556 68572
rect 4556 68516 4612 68572
rect 4612 68516 4616 68572
rect 4552 68512 4616 68516
rect 4632 68572 4696 68576
rect 4632 68516 4636 68572
rect 4636 68516 4692 68572
rect 4692 68516 4696 68572
rect 4632 68512 4696 68516
rect 4712 68572 4776 68576
rect 4712 68516 4716 68572
rect 4716 68516 4772 68572
rect 4772 68516 4776 68572
rect 4712 68512 4776 68516
rect 4792 68572 4856 68576
rect 4792 68516 4796 68572
rect 4796 68516 4852 68572
rect 4852 68516 4856 68572
rect 4792 68512 4856 68516
rect 6152 68572 6216 68576
rect 6152 68516 6156 68572
rect 6156 68516 6212 68572
rect 6212 68516 6216 68572
rect 6152 68512 6216 68516
rect 6232 68572 6296 68576
rect 6232 68516 6236 68572
rect 6236 68516 6292 68572
rect 6292 68516 6296 68572
rect 6232 68512 6296 68516
rect 6312 68572 6376 68576
rect 6312 68516 6316 68572
rect 6316 68516 6372 68572
rect 6372 68516 6376 68572
rect 6312 68512 6376 68516
rect 6392 68572 6456 68576
rect 6392 68516 6396 68572
rect 6396 68516 6452 68572
rect 6452 68516 6456 68572
rect 6392 68512 6456 68516
rect 7752 68572 7816 68576
rect 7752 68516 7756 68572
rect 7756 68516 7812 68572
rect 7812 68516 7816 68572
rect 7752 68512 7816 68516
rect 7832 68572 7896 68576
rect 7832 68516 7836 68572
rect 7836 68516 7892 68572
rect 7892 68516 7896 68572
rect 7832 68512 7896 68516
rect 7912 68572 7976 68576
rect 7912 68516 7916 68572
rect 7916 68516 7972 68572
rect 7972 68516 7976 68572
rect 7912 68512 7976 68516
rect 7992 68572 8056 68576
rect 7992 68516 7996 68572
rect 7996 68516 8052 68572
rect 8052 68516 8056 68572
rect 7992 68512 8056 68516
rect 9352 68572 9416 68576
rect 9352 68516 9356 68572
rect 9356 68516 9412 68572
rect 9412 68516 9416 68572
rect 9352 68512 9416 68516
rect 9432 68572 9496 68576
rect 9432 68516 9436 68572
rect 9436 68516 9492 68572
rect 9492 68516 9496 68572
rect 9432 68512 9496 68516
rect 9512 68572 9576 68576
rect 9512 68516 9516 68572
rect 9516 68516 9572 68572
rect 9572 68516 9576 68572
rect 9512 68512 9576 68516
rect 9592 68572 9656 68576
rect 9592 68516 9596 68572
rect 9596 68516 9652 68572
rect 9652 68516 9656 68572
rect 9592 68512 9656 68516
rect 3612 68028 3676 68032
rect 3612 67972 3616 68028
rect 3616 67972 3672 68028
rect 3672 67972 3676 68028
rect 3612 67968 3676 67972
rect 3692 68028 3756 68032
rect 3692 67972 3696 68028
rect 3696 67972 3752 68028
rect 3752 67972 3756 68028
rect 3692 67968 3756 67972
rect 3772 68028 3836 68032
rect 3772 67972 3776 68028
rect 3776 67972 3832 68028
rect 3832 67972 3836 68028
rect 3772 67968 3836 67972
rect 3852 68028 3916 68032
rect 3852 67972 3856 68028
rect 3856 67972 3912 68028
rect 3912 67972 3916 68028
rect 3852 67968 3916 67972
rect 5212 68028 5276 68032
rect 5212 67972 5216 68028
rect 5216 67972 5272 68028
rect 5272 67972 5276 68028
rect 5212 67968 5276 67972
rect 5292 68028 5356 68032
rect 5292 67972 5296 68028
rect 5296 67972 5352 68028
rect 5352 67972 5356 68028
rect 5292 67968 5356 67972
rect 5372 68028 5436 68032
rect 5372 67972 5376 68028
rect 5376 67972 5432 68028
rect 5432 67972 5436 68028
rect 5372 67968 5436 67972
rect 5452 68028 5516 68032
rect 5452 67972 5456 68028
rect 5456 67972 5512 68028
rect 5512 67972 5516 68028
rect 5452 67968 5516 67972
rect 6812 68028 6876 68032
rect 6812 67972 6816 68028
rect 6816 67972 6872 68028
rect 6872 67972 6876 68028
rect 6812 67968 6876 67972
rect 6892 68028 6956 68032
rect 6892 67972 6896 68028
rect 6896 67972 6952 68028
rect 6952 67972 6956 68028
rect 6892 67968 6956 67972
rect 6972 68028 7036 68032
rect 6972 67972 6976 68028
rect 6976 67972 7032 68028
rect 7032 67972 7036 68028
rect 6972 67968 7036 67972
rect 7052 68028 7116 68032
rect 7052 67972 7056 68028
rect 7056 67972 7112 68028
rect 7112 67972 7116 68028
rect 7052 67968 7116 67972
rect 8412 68028 8476 68032
rect 8412 67972 8416 68028
rect 8416 67972 8472 68028
rect 8472 67972 8476 68028
rect 8412 67968 8476 67972
rect 8492 68028 8556 68032
rect 8492 67972 8496 68028
rect 8496 67972 8552 68028
rect 8552 67972 8556 68028
rect 8492 67968 8556 67972
rect 8572 68028 8636 68032
rect 8572 67972 8576 68028
rect 8576 67972 8632 68028
rect 8632 67972 8636 68028
rect 8572 67968 8636 67972
rect 8652 68028 8716 68032
rect 8652 67972 8656 68028
rect 8656 67972 8712 68028
rect 8712 67972 8716 68028
rect 8652 67968 8716 67972
rect 2952 67484 3016 67488
rect 2952 67428 2956 67484
rect 2956 67428 3012 67484
rect 3012 67428 3016 67484
rect 2952 67424 3016 67428
rect 3032 67484 3096 67488
rect 3032 67428 3036 67484
rect 3036 67428 3092 67484
rect 3092 67428 3096 67484
rect 3032 67424 3096 67428
rect 3112 67484 3176 67488
rect 3112 67428 3116 67484
rect 3116 67428 3172 67484
rect 3172 67428 3176 67484
rect 3112 67424 3176 67428
rect 3192 67484 3256 67488
rect 3192 67428 3196 67484
rect 3196 67428 3252 67484
rect 3252 67428 3256 67484
rect 3192 67424 3256 67428
rect 4552 67484 4616 67488
rect 4552 67428 4556 67484
rect 4556 67428 4612 67484
rect 4612 67428 4616 67484
rect 4552 67424 4616 67428
rect 4632 67484 4696 67488
rect 4632 67428 4636 67484
rect 4636 67428 4692 67484
rect 4692 67428 4696 67484
rect 4632 67424 4696 67428
rect 4712 67484 4776 67488
rect 4712 67428 4716 67484
rect 4716 67428 4772 67484
rect 4772 67428 4776 67484
rect 4712 67424 4776 67428
rect 4792 67484 4856 67488
rect 4792 67428 4796 67484
rect 4796 67428 4852 67484
rect 4852 67428 4856 67484
rect 4792 67424 4856 67428
rect 6152 67484 6216 67488
rect 6152 67428 6156 67484
rect 6156 67428 6212 67484
rect 6212 67428 6216 67484
rect 6152 67424 6216 67428
rect 6232 67484 6296 67488
rect 6232 67428 6236 67484
rect 6236 67428 6292 67484
rect 6292 67428 6296 67484
rect 6232 67424 6296 67428
rect 6312 67484 6376 67488
rect 6312 67428 6316 67484
rect 6316 67428 6372 67484
rect 6372 67428 6376 67484
rect 6312 67424 6376 67428
rect 6392 67484 6456 67488
rect 6392 67428 6396 67484
rect 6396 67428 6452 67484
rect 6452 67428 6456 67484
rect 6392 67424 6456 67428
rect 7752 67484 7816 67488
rect 7752 67428 7756 67484
rect 7756 67428 7812 67484
rect 7812 67428 7816 67484
rect 7752 67424 7816 67428
rect 7832 67484 7896 67488
rect 7832 67428 7836 67484
rect 7836 67428 7892 67484
rect 7892 67428 7896 67484
rect 7832 67424 7896 67428
rect 7912 67484 7976 67488
rect 7912 67428 7916 67484
rect 7916 67428 7972 67484
rect 7972 67428 7976 67484
rect 7912 67424 7976 67428
rect 7992 67484 8056 67488
rect 7992 67428 7996 67484
rect 7996 67428 8052 67484
rect 8052 67428 8056 67484
rect 7992 67424 8056 67428
rect 9352 67484 9416 67488
rect 9352 67428 9356 67484
rect 9356 67428 9412 67484
rect 9412 67428 9416 67484
rect 9352 67424 9416 67428
rect 9432 67484 9496 67488
rect 9432 67428 9436 67484
rect 9436 67428 9492 67484
rect 9492 67428 9496 67484
rect 9432 67424 9496 67428
rect 9512 67484 9576 67488
rect 9512 67428 9516 67484
rect 9516 67428 9572 67484
rect 9572 67428 9576 67484
rect 9512 67424 9576 67428
rect 9592 67484 9656 67488
rect 9592 67428 9596 67484
rect 9596 67428 9652 67484
rect 9652 67428 9656 67484
rect 9592 67424 9656 67428
rect 3612 66940 3676 66944
rect 3612 66884 3616 66940
rect 3616 66884 3672 66940
rect 3672 66884 3676 66940
rect 3612 66880 3676 66884
rect 3692 66940 3756 66944
rect 3692 66884 3696 66940
rect 3696 66884 3752 66940
rect 3752 66884 3756 66940
rect 3692 66880 3756 66884
rect 3772 66940 3836 66944
rect 3772 66884 3776 66940
rect 3776 66884 3832 66940
rect 3832 66884 3836 66940
rect 3772 66880 3836 66884
rect 3852 66940 3916 66944
rect 3852 66884 3856 66940
rect 3856 66884 3912 66940
rect 3912 66884 3916 66940
rect 3852 66880 3916 66884
rect 5212 66940 5276 66944
rect 5212 66884 5216 66940
rect 5216 66884 5272 66940
rect 5272 66884 5276 66940
rect 5212 66880 5276 66884
rect 5292 66940 5356 66944
rect 5292 66884 5296 66940
rect 5296 66884 5352 66940
rect 5352 66884 5356 66940
rect 5292 66880 5356 66884
rect 5372 66940 5436 66944
rect 5372 66884 5376 66940
rect 5376 66884 5432 66940
rect 5432 66884 5436 66940
rect 5372 66880 5436 66884
rect 5452 66940 5516 66944
rect 5452 66884 5456 66940
rect 5456 66884 5512 66940
rect 5512 66884 5516 66940
rect 5452 66880 5516 66884
rect 6812 66940 6876 66944
rect 6812 66884 6816 66940
rect 6816 66884 6872 66940
rect 6872 66884 6876 66940
rect 6812 66880 6876 66884
rect 6892 66940 6956 66944
rect 6892 66884 6896 66940
rect 6896 66884 6952 66940
rect 6952 66884 6956 66940
rect 6892 66880 6956 66884
rect 6972 66940 7036 66944
rect 6972 66884 6976 66940
rect 6976 66884 7032 66940
rect 7032 66884 7036 66940
rect 6972 66880 7036 66884
rect 7052 66940 7116 66944
rect 7052 66884 7056 66940
rect 7056 66884 7112 66940
rect 7112 66884 7116 66940
rect 7052 66880 7116 66884
rect 8412 66940 8476 66944
rect 8412 66884 8416 66940
rect 8416 66884 8472 66940
rect 8472 66884 8476 66940
rect 8412 66880 8476 66884
rect 8492 66940 8556 66944
rect 8492 66884 8496 66940
rect 8496 66884 8552 66940
rect 8552 66884 8556 66940
rect 8492 66880 8556 66884
rect 8572 66940 8636 66944
rect 8572 66884 8576 66940
rect 8576 66884 8632 66940
rect 8632 66884 8636 66940
rect 8572 66880 8636 66884
rect 8652 66940 8716 66944
rect 8652 66884 8656 66940
rect 8656 66884 8712 66940
rect 8712 66884 8716 66940
rect 8652 66880 8716 66884
rect 2952 66396 3016 66400
rect 2952 66340 2956 66396
rect 2956 66340 3012 66396
rect 3012 66340 3016 66396
rect 2952 66336 3016 66340
rect 3032 66396 3096 66400
rect 3032 66340 3036 66396
rect 3036 66340 3092 66396
rect 3092 66340 3096 66396
rect 3032 66336 3096 66340
rect 3112 66396 3176 66400
rect 3112 66340 3116 66396
rect 3116 66340 3172 66396
rect 3172 66340 3176 66396
rect 3112 66336 3176 66340
rect 3192 66396 3256 66400
rect 3192 66340 3196 66396
rect 3196 66340 3252 66396
rect 3252 66340 3256 66396
rect 3192 66336 3256 66340
rect 4552 66396 4616 66400
rect 4552 66340 4556 66396
rect 4556 66340 4612 66396
rect 4612 66340 4616 66396
rect 4552 66336 4616 66340
rect 4632 66396 4696 66400
rect 4632 66340 4636 66396
rect 4636 66340 4692 66396
rect 4692 66340 4696 66396
rect 4632 66336 4696 66340
rect 4712 66396 4776 66400
rect 4712 66340 4716 66396
rect 4716 66340 4772 66396
rect 4772 66340 4776 66396
rect 4712 66336 4776 66340
rect 4792 66396 4856 66400
rect 4792 66340 4796 66396
rect 4796 66340 4852 66396
rect 4852 66340 4856 66396
rect 4792 66336 4856 66340
rect 3612 65852 3676 65856
rect 3612 65796 3616 65852
rect 3616 65796 3672 65852
rect 3672 65796 3676 65852
rect 3612 65792 3676 65796
rect 3692 65852 3756 65856
rect 3692 65796 3696 65852
rect 3696 65796 3752 65852
rect 3752 65796 3756 65852
rect 3692 65792 3756 65796
rect 3772 65852 3836 65856
rect 3772 65796 3776 65852
rect 3776 65796 3832 65852
rect 3832 65796 3836 65852
rect 3772 65792 3836 65796
rect 3852 65852 3916 65856
rect 3852 65796 3856 65852
rect 3856 65796 3912 65852
rect 3912 65796 3916 65852
rect 3852 65792 3916 65796
rect 11836 66540 11900 66604
rect 6152 66396 6216 66400
rect 6152 66340 6156 66396
rect 6156 66340 6212 66396
rect 6212 66340 6216 66396
rect 6152 66336 6216 66340
rect 6232 66396 6296 66400
rect 6232 66340 6236 66396
rect 6236 66340 6292 66396
rect 6292 66340 6296 66396
rect 6232 66336 6296 66340
rect 6312 66396 6376 66400
rect 6312 66340 6316 66396
rect 6316 66340 6372 66396
rect 6372 66340 6376 66396
rect 6312 66336 6376 66340
rect 6392 66396 6456 66400
rect 6392 66340 6396 66396
rect 6396 66340 6452 66396
rect 6452 66340 6456 66396
rect 6392 66336 6456 66340
rect 7752 66396 7816 66400
rect 7752 66340 7756 66396
rect 7756 66340 7812 66396
rect 7812 66340 7816 66396
rect 7752 66336 7816 66340
rect 7832 66396 7896 66400
rect 7832 66340 7836 66396
rect 7836 66340 7892 66396
rect 7892 66340 7896 66396
rect 7832 66336 7896 66340
rect 7912 66396 7976 66400
rect 7912 66340 7916 66396
rect 7916 66340 7972 66396
rect 7972 66340 7976 66396
rect 7912 66336 7976 66340
rect 7992 66396 8056 66400
rect 7992 66340 7996 66396
rect 7996 66340 8052 66396
rect 8052 66340 8056 66396
rect 7992 66336 8056 66340
rect 9352 66396 9416 66400
rect 9352 66340 9356 66396
rect 9356 66340 9412 66396
rect 9412 66340 9416 66396
rect 9352 66336 9416 66340
rect 9432 66396 9496 66400
rect 9432 66340 9436 66396
rect 9436 66340 9492 66396
rect 9492 66340 9496 66396
rect 9432 66336 9496 66340
rect 9512 66396 9576 66400
rect 9512 66340 9516 66396
rect 9516 66340 9572 66396
rect 9572 66340 9576 66396
rect 9512 66336 9576 66340
rect 9592 66396 9656 66400
rect 9592 66340 9596 66396
rect 9596 66340 9652 66396
rect 9652 66340 9656 66396
rect 9592 66336 9656 66340
rect 5212 65852 5276 65856
rect 5212 65796 5216 65852
rect 5216 65796 5272 65852
rect 5272 65796 5276 65852
rect 5212 65792 5276 65796
rect 5292 65852 5356 65856
rect 5292 65796 5296 65852
rect 5296 65796 5352 65852
rect 5352 65796 5356 65852
rect 5292 65792 5356 65796
rect 5372 65852 5436 65856
rect 5372 65796 5376 65852
rect 5376 65796 5432 65852
rect 5432 65796 5436 65852
rect 5372 65792 5436 65796
rect 5452 65852 5516 65856
rect 5452 65796 5456 65852
rect 5456 65796 5512 65852
rect 5512 65796 5516 65852
rect 5452 65792 5516 65796
rect 6812 65852 6876 65856
rect 6812 65796 6816 65852
rect 6816 65796 6872 65852
rect 6872 65796 6876 65852
rect 6812 65792 6876 65796
rect 6892 65852 6956 65856
rect 6892 65796 6896 65852
rect 6896 65796 6952 65852
rect 6952 65796 6956 65852
rect 6892 65792 6956 65796
rect 6972 65852 7036 65856
rect 6972 65796 6976 65852
rect 6976 65796 7032 65852
rect 7032 65796 7036 65852
rect 6972 65792 7036 65796
rect 7052 65852 7116 65856
rect 7052 65796 7056 65852
rect 7056 65796 7112 65852
rect 7112 65796 7116 65852
rect 7052 65792 7116 65796
rect 8412 65852 8476 65856
rect 8412 65796 8416 65852
rect 8416 65796 8472 65852
rect 8472 65796 8476 65852
rect 8412 65792 8476 65796
rect 8492 65852 8556 65856
rect 8492 65796 8496 65852
rect 8496 65796 8552 65852
rect 8552 65796 8556 65852
rect 8492 65792 8556 65796
rect 8572 65852 8636 65856
rect 8572 65796 8576 65852
rect 8576 65796 8632 65852
rect 8632 65796 8636 65852
rect 8572 65792 8636 65796
rect 8652 65852 8716 65856
rect 8652 65796 8656 65852
rect 8656 65796 8712 65852
rect 8712 65796 8716 65852
rect 8652 65792 8716 65796
rect 2952 65308 3016 65312
rect 2952 65252 2956 65308
rect 2956 65252 3012 65308
rect 3012 65252 3016 65308
rect 2952 65248 3016 65252
rect 3032 65308 3096 65312
rect 3032 65252 3036 65308
rect 3036 65252 3092 65308
rect 3092 65252 3096 65308
rect 3032 65248 3096 65252
rect 3112 65308 3176 65312
rect 3112 65252 3116 65308
rect 3116 65252 3172 65308
rect 3172 65252 3176 65308
rect 3112 65248 3176 65252
rect 3192 65308 3256 65312
rect 3192 65252 3196 65308
rect 3196 65252 3252 65308
rect 3252 65252 3256 65308
rect 3192 65248 3256 65252
rect 4552 65308 4616 65312
rect 4552 65252 4556 65308
rect 4556 65252 4612 65308
rect 4612 65252 4616 65308
rect 4552 65248 4616 65252
rect 4632 65308 4696 65312
rect 4632 65252 4636 65308
rect 4636 65252 4692 65308
rect 4692 65252 4696 65308
rect 4632 65248 4696 65252
rect 4712 65308 4776 65312
rect 4712 65252 4716 65308
rect 4716 65252 4772 65308
rect 4772 65252 4776 65308
rect 4712 65248 4776 65252
rect 4792 65308 4856 65312
rect 4792 65252 4796 65308
rect 4796 65252 4852 65308
rect 4852 65252 4856 65308
rect 4792 65248 4856 65252
rect 6152 65308 6216 65312
rect 6152 65252 6156 65308
rect 6156 65252 6212 65308
rect 6212 65252 6216 65308
rect 6152 65248 6216 65252
rect 6232 65308 6296 65312
rect 6232 65252 6236 65308
rect 6236 65252 6292 65308
rect 6292 65252 6296 65308
rect 6232 65248 6296 65252
rect 6312 65308 6376 65312
rect 6312 65252 6316 65308
rect 6316 65252 6372 65308
rect 6372 65252 6376 65308
rect 6312 65248 6376 65252
rect 6392 65308 6456 65312
rect 6392 65252 6396 65308
rect 6396 65252 6452 65308
rect 6452 65252 6456 65308
rect 6392 65248 6456 65252
rect 7752 65308 7816 65312
rect 7752 65252 7756 65308
rect 7756 65252 7812 65308
rect 7812 65252 7816 65308
rect 7752 65248 7816 65252
rect 7832 65308 7896 65312
rect 7832 65252 7836 65308
rect 7836 65252 7892 65308
rect 7892 65252 7896 65308
rect 7832 65248 7896 65252
rect 7912 65308 7976 65312
rect 7912 65252 7916 65308
rect 7916 65252 7972 65308
rect 7972 65252 7976 65308
rect 7912 65248 7976 65252
rect 7992 65308 8056 65312
rect 7992 65252 7996 65308
rect 7996 65252 8052 65308
rect 8052 65252 8056 65308
rect 7992 65248 8056 65252
rect 9352 65308 9416 65312
rect 9352 65252 9356 65308
rect 9356 65252 9412 65308
rect 9412 65252 9416 65308
rect 9352 65248 9416 65252
rect 9432 65308 9496 65312
rect 9432 65252 9436 65308
rect 9436 65252 9492 65308
rect 9492 65252 9496 65308
rect 9432 65248 9496 65252
rect 9512 65308 9576 65312
rect 9512 65252 9516 65308
rect 9516 65252 9572 65308
rect 9572 65252 9576 65308
rect 9512 65248 9576 65252
rect 9592 65308 9656 65312
rect 9592 65252 9596 65308
rect 9596 65252 9652 65308
rect 9652 65252 9656 65308
rect 9592 65248 9656 65252
rect 3612 64764 3676 64768
rect 3612 64708 3616 64764
rect 3616 64708 3672 64764
rect 3672 64708 3676 64764
rect 3612 64704 3676 64708
rect 3692 64764 3756 64768
rect 3692 64708 3696 64764
rect 3696 64708 3752 64764
rect 3752 64708 3756 64764
rect 3692 64704 3756 64708
rect 3772 64764 3836 64768
rect 3772 64708 3776 64764
rect 3776 64708 3832 64764
rect 3832 64708 3836 64764
rect 3772 64704 3836 64708
rect 3852 64764 3916 64768
rect 3852 64708 3856 64764
rect 3856 64708 3912 64764
rect 3912 64708 3916 64764
rect 3852 64704 3916 64708
rect 5212 64764 5276 64768
rect 5212 64708 5216 64764
rect 5216 64708 5272 64764
rect 5272 64708 5276 64764
rect 5212 64704 5276 64708
rect 5292 64764 5356 64768
rect 5292 64708 5296 64764
rect 5296 64708 5352 64764
rect 5352 64708 5356 64764
rect 5292 64704 5356 64708
rect 5372 64764 5436 64768
rect 5372 64708 5376 64764
rect 5376 64708 5432 64764
rect 5432 64708 5436 64764
rect 5372 64704 5436 64708
rect 5452 64764 5516 64768
rect 5452 64708 5456 64764
rect 5456 64708 5512 64764
rect 5512 64708 5516 64764
rect 5452 64704 5516 64708
rect 6812 64764 6876 64768
rect 6812 64708 6816 64764
rect 6816 64708 6872 64764
rect 6872 64708 6876 64764
rect 6812 64704 6876 64708
rect 6892 64764 6956 64768
rect 6892 64708 6896 64764
rect 6896 64708 6952 64764
rect 6952 64708 6956 64764
rect 6892 64704 6956 64708
rect 6972 64764 7036 64768
rect 6972 64708 6976 64764
rect 6976 64708 7032 64764
rect 7032 64708 7036 64764
rect 6972 64704 7036 64708
rect 7052 64764 7116 64768
rect 7052 64708 7056 64764
rect 7056 64708 7112 64764
rect 7112 64708 7116 64764
rect 7052 64704 7116 64708
rect 8412 64764 8476 64768
rect 8412 64708 8416 64764
rect 8416 64708 8472 64764
rect 8472 64708 8476 64764
rect 8412 64704 8476 64708
rect 8492 64764 8556 64768
rect 8492 64708 8496 64764
rect 8496 64708 8552 64764
rect 8552 64708 8556 64764
rect 8492 64704 8556 64708
rect 8572 64764 8636 64768
rect 8572 64708 8576 64764
rect 8576 64708 8632 64764
rect 8632 64708 8636 64764
rect 8572 64704 8636 64708
rect 8652 64764 8716 64768
rect 8652 64708 8656 64764
rect 8656 64708 8712 64764
rect 8712 64708 8716 64764
rect 8652 64704 8716 64708
rect 2952 64220 3016 64224
rect 2952 64164 2956 64220
rect 2956 64164 3012 64220
rect 3012 64164 3016 64220
rect 2952 64160 3016 64164
rect 3032 64220 3096 64224
rect 3032 64164 3036 64220
rect 3036 64164 3092 64220
rect 3092 64164 3096 64220
rect 3032 64160 3096 64164
rect 3112 64220 3176 64224
rect 3112 64164 3116 64220
rect 3116 64164 3172 64220
rect 3172 64164 3176 64220
rect 3112 64160 3176 64164
rect 3192 64220 3256 64224
rect 3192 64164 3196 64220
rect 3196 64164 3252 64220
rect 3252 64164 3256 64220
rect 3192 64160 3256 64164
rect 4552 64220 4616 64224
rect 4552 64164 4556 64220
rect 4556 64164 4612 64220
rect 4612 64164 4616 64220
rect 4552 64160 4616 64164
rect 4632 64220 4696 64224
rect 4632 64164 4636 64220
rect 4636 64164 4692 64220
rect 4692 64164 4696 64220
rect 4632 64160 4696 64164
rect 4712 64220 4776 64224
rect 4712 64164 4716 64220
rect 4716 64164 4772 64220
rect 4772 64164 4776 64220
rect 4712 64160 4776 64164
rect 4792 64220 4856 64224
rect 4792 64164 4796 64220
rect 4796 64164 4852 64220
rect 4852 64164 4856 64220
rect 4792 64160 4856 64164
rect 6152 64220 6216 64224
rect 6152 64164 6156 64220
rect 6156 64164 6212 64220
rect 6212 64164 6216 64220
rect 6152 64160 6216 64164
rect 6232 64220 6296 64224
rect 6232 64164 6236 64220
rect 6236 64164 6292 64220
rect 6292 64164 6296 64220
rect 6232 64160 6296 64164
rect 6312 64220 6376 64224
rect 6312 64164 6316 64220
rect 6316 64164 6372 64220
rect 6372 64164 6376 64220
rect 6312 64160 6376 64164
rect 6392 64220 6456 64224
rect 6392 64164 6396 64220
rect 6396 64164 6452 64220
rect 6452 64164 6456 64220
rect 6392 64160 6456 64164
rect 7752 64220 7816 64224
rect 7752 64164 7756 64220
rect 7756 64164 7812 64220
rect 7812 64164 7816 64220
rect 7752 64160 7816 64164
rect 7832 64220 7896 64224
rect 7832 64164 7836 64220
rect 7836 64164 7892 64220
rect 7892 64164 7896 64220
rect 7832 64160 7896 64164
rect 7912 64220 7976 64224
rect 7912 64164 7916 64220
rect 7916 64164 7972 64220
rect 7972 64164 7976 64220
rect 7912 64160 7976 64164
rect 7992 64220 8056 64224
rect 7992 64164 7996 64220
rect 7996 64164 8052 64220
rect 8052 64164 8056 64220
rect 7992 64160 8056 64164
rect 9352 64220 9416 64224
rect 9352 64164 9356 64220
rect 9356 64164 9412 64220
rect 9412 64164 9416 64220
rect 9352 64160 9416 64164
rect 9432 64220 9496 64224
rect 9432 64164 9436 64220
rect 9436 64164 9492 64220
rect 9492 64164 9496 64220
rect 9432 64160 9496 64164
rect 9512 64220 9576 64224
rect 9512 64164 9516 64220
rect 9516 64164 9572 64220
rect 9572 64164 9576 64220
rect 9512 64160 9576 64164
rect 9592 64220 9656 64224
rect 9592 64164 9596 64220
rect 9596 64164 9652 64220
rect 9652 64164 9656 64220
rect 9592 64160 9656 64164
rect 3612 63676 3676 63680
rect 3612 63620 3616 63676
rect 3616 63620 3672 63676
rect 3672 63620 3676 63676
rect 3612 63616 3676 63620
rect 3692 63676 3756 63680
rect 3692 63620 3696 63676
rect 3696 63620 3752 63676
rect 3752 63620 3756 63676
rect 3692 63616 3756 63620
rect 3772 63676 3836 63680
rect 3772 63620 3776 63676
rect 3776 63620 3832 63676
rect 3832 63620 3836 63676
rect 3772 63616 3836 63620
rect 3852 63676 3916 63680
rect 3852 63620 3856 63676
rect 3856 63620 3912 63676
rect 3912 63620 3916 63676
rect 3852 63616 3916 63620
rect 5212 63676 5276 63680
rect 5212 63620 5216 63676
rect 5216 63620 5272 63676
rect 5272 63620 5276 63676
rect 5212 63616 5276 63620
rect 5292 63676 5356 63680
rect 5292 63620 5296 63676
rect 5296 63620 5352 63676
rect 5352 63620 5356 63676
rect 5292 63616 5356 63620
rect 5372 63676 5436 63680
rect 5372 63620 5376 63676
rect 5376 63620 5432 63676
rect 5432 63620 5436 63676
rect 5372 63616 5436 63620
rect 5452 63676 5516 63680
rect 5452 63620 5456 63676
rect 5456 63620 5512 63676
rect 5512 63620 5516 63676
rect 5452 63616 5516 63620
rect 6812 63676 6876 63680
rect 6812 63620 6816 63676
rect 6816 63620 6872 63676
rect 6872 63620 6876 63676
rect 6812 63616 6876 63620
rect 6892 63676 6956 63680
rect 6892 63620 6896 63676
rect 6896 63620 6952 63676
rect 6952 63620 6956 63676
rect 6892 63616 6956 63620
rect 6972 63676 7036 63680
rect 6972 63620 6976 63676
rect 6976 63620 7032 63676
rect 7032 63620 7036 63676
rect 6972 63616 7036 63620
rect 7052 63676 7116 63680
rect 7052 63620 7056 63676
rect 7056 63620 7112 63676
rect 7112 63620 7116 63676
rect 7052 63616 7116 63620
rect 8412 63676 8476 63680
rect 8412 63620 8416 63676
rect 8416 63620 8472 63676
rect 8472 63620 8476 63676
rect 8412 63616 8476 63620
rect 8492 63676 8556 63680
rect 8492 63620 8496 63676
rect 8496 63620 8552 63676
rect 8552 63620 8556 63676
rect 8492 63616 8556 63620
rect 8572 63676 8636 63680
rect 8572 63620 8576 63676
rect 8576 63620 8632 63676
rect 8632 63620 8636 63676
rect 8572 63616 8636 63620
rect 8652 63676 8716 63680
rect 8652 63620 8656 63676
rect 8656 63620 8712 63676
rect 8712 63620 8716 63676
rect 8652 63616 8716 63620
rect 2952 63132 3016 63136
rect 2952 63076 2956 63132
rect 2956 63076 3012 63132
rect 3012 63076 3016 63132
rect 2952 63072 3016 63076
rect 3032 63132 3096 63136
rect 3032 63076 3036 63132
rect 3036 63076 3092 63132
rect 3092 63076 3096 63132
rect 3032 63072 3096 63076
rect 3112 63132 3176 63136
rect 3112 63076 3116 63132
rect 3116 63076 3172 63132
rect 3172 63076 3176 63132
rect 3112 63072 3176 63076
rect 3192 63132 3256 63136
rect 3192 63076 3196 63132
rect 3196 63076 3252 63132
rect 3252 63076 3256 63132
rect 3192 63072 3256 63076
rect 4552 63132 4616 63136
rect 4552 63076 4556 63132
rect 4556 63076 4612 63132
rect 4612 63076 4616 63132
rect 4552 63072 4616 63076
rect 4632 63132 4696 63136
rect 4632 63076 4636 63132
rect 4636 63076 4692 63132
rect 4692 63076 4696 63132
rect 4632 63072 4696 63076
rect 4712 63132 4776 63136
rect 4712 63076 4716 63132
rect 4716 63076 4772 63132
rect 4772 63076 4776 63132
rect 4712 63072 4776 63076
rect 4792 63132 4856 63136
rect 4792 63076 4796 63132
rect 4796 63076 4852 63132
rect 4852 63076 4856 63132
rect 4792 63072 4856 63076
rect 6152 63132 6216 63136
rect 6152 63076 6156 63132
rect 6156 63076 6212 63132
rect 6212 63076 6216 63132
rect 6152 63072 6216 63076
rect 6232 63132 6296 63136
rect 6232 63076 6236 63132
rect 6236 63076 6292 63132
rect 6292 63076 6296 63132
rect 6232 63072 6296 63076
rect 6312 63132 6376 63136
rect 6312 63076 6316 63132
rect 6316 63076 6372 63132
rect 6372 63076 6376 63132
rect 6312 63072 6376 63076
rect 6392 63132 6456 63136
rect 6392 63076 6396 63132
rect 6396 63076 6452 63132
rect 6452 63076 6456 63132
rect 6392 63072 6456 63076
rect 7752 63132 7816 63136
rect 7752 63076 7756 63132
rect 7756 63076 7812 63132
rect 7812 63076 7816 63132
rect 7752 63072 7816 63076
rect 7832 63132 7896 63136
rect 7832 63076 7836 63132
rect 7836 63076 7892 63132
rect 7892 63076 7896 63132
rect 7832 63072 7896 63076
rect 7912 63132 7976 63136
rect 7912 63076 7916 63132
rect 7916 63076 7972 63132
rect 7972 63076 7976 63132
rect 7912 63072 7976 63076
rect 7992 63132 8056 63136
rect 7992 63076 7996 63132
rect 7996 63076 8052 63132
rect 8052 63076 8056 63132
rect 7992 63072 8056 63076
rect 9352 63132 9416 63136
rect 9352 63076 9356 63132
rect 9356 63076 9412 63132
rect 9412 63076 9416 63132
rect 9352 63072 9416 63076
rect 9432 63132 9496 63136
rect 9432 63076 9436 63132
rect 9436 63076 9492 63132
rect 9492 63076 9496 63132
rect 9432 63072 9496 63076
rect 9512 63132 9576 63136
rect 9512 63076 9516 63132
rect 9516 63076 9572 63132
rect 9572 63076 9576 63132
rect 9512 63072 9576 63076
rect 9592 63132 9656 63136
rect 9592 63076 9596 63132
rect 9596 63076 9652 63132
rect 9652 63076 9656 63132
rect 9592 63072 9656 63076
rect 3612 62588 3676 62592
rect 3612 62532 3616 62588
rect 3616 62532 3672 62588
rect 3672 62532 3676 62588
rect 3612 62528 3676 62532
rect 3692 62588 3756 62592
rect 3692 62532 3696 62588
rect 3696 62532 3752 62588
rect 3752 62532 3756 62588
rect 3692 62528 3756 62532
rect 3772 62588 3836 62592
rect 3772 62532 3776 62588
rect 3776 62532 3832 62588
rect 3832 62532 3836 62588
rect 3772 62528 3836 62532
rect 3852 62588 3916 62592
rect 3852 62532 3856 62588
rect 3856 62532 3912 62588
rect 3912 62532 3916 62588
rect 3852 62528 3916 62532
rect 5212 62588 5276 62592
rect 5212 62532 5216 62588
rect 5216 62532 5272 62588
rect 5272 62532 5276 62588
rect 5212 62528 5276 62532
rect 5292 62588 5356 62592
rect 5292 62532 5296 62588
rect 5296 62532 5352 62588
rect 5352 62532 5356 62588
rect 5292 62528 5356 62532
rect 5372 62588 5436 62592
rect 5372 62532 5376 62588
rect 5376 62532 5432 62588
rect 5432 62532 5436 62588
rect 5372 62528 5436 62532
rect 5452 62588 5516 62592
rect 5452 62532 5456 62588
rect 5456 62532 5512 62588
rect 5512 62532 5516 62588
rect 5452 62528 5516 62532
rect 6812 62588 6876 62592
rect 6812 62532 6816 62588
rect 6816 62532 6872 62588
rect 6872 62532 6876 62588
rect 6812 62528 6876 62532
rect 6892 62588 6956 62592
rect 6892 62532 6896 62588
rect 6896 62532 6952 62588
rect 6952 62532 6956 62588
rect 6892 62528 6956 62532
rect 6972 62588 7036 62592
rect 6972 62532 6976 62588
rect 6976 62532 7032 62588
rect 7032 62532 7036 62588
rect 6972 62528 7036 62532
rect 7052 62588 7116 62592
rect 7052 62532 7056 62588
rect 7056 62532 7112 62588
rect 7112 62532 7116 62588
rect 7052 62528 7116 62532
rect 8412 62588 8476 62592
rect 8412 62532 8416 62588
rect 8416 62532 8472 62588
rect 8472 62532 8476 62588
rect 8412 62528 8476 62532
rect 8492 62588 8556 62592
rect 8492 62532 8496 62588
rect 8496 62532 8552 62588
rect 8552 62532 8556 62588
rect 8492 62528 8556 62532
rect 8572 62588 8636 62592
rect 8572 62532 8576 62588
rect 8576 62532 8632 62588
rect 8632 62532 8636 62588
rect 8572 62528 8636 62532
rect 8652 62588 8716 62592
rect 8652 62532 8656 62588
rect 8656 62532 8712 62588
rect 8712 62532 8716 62588
rect 8652 62528 8716 62532
rect 2952 62044 3016 62048
rect 2952 61988 2956 62044
rect 2956 61988 3012 62044
rect 3012 61988 3016 62044
rect 2952 61984 3016 61988
rect 3032 62044 3096 62048
rect 3032 61988 3036 62044
rect 3036 61988 3092 62044
rect 3092 61988 3096 62044
rect 3032 61984 3096 61988
rect 3112 62044 3176 62048
rect 3112 61988 3116 62044
rect 3116 61988 3172 62044
rect 3172 61988 3176 62044
rect 3112 61984 3176 61988
rect 3192 62044 3256 62048
rect 3192 61988 3196 62044
rect 3196 61988 3252 62044
rect 3252 61988 3256 62044
rect 3192 61984 3256 61988
rect 4552 62044 4616 62048
rect 4552 61988 4556 62044
rect 4556 61988 4612 62044
rect 4612 61988 4616 62044
rect 4552 61984 4616 61988
rect 4632 62044 4696 62048
rect 4632 61988 4636 62044
rect 4636 61988 4692 62044
rect 4692 61988 4696 62044
rect 4632 61984 4696 61988
rect 4712 62044 4776 62048
rect 4712 61988 4716 62044
rect 4716 61988 4772 62044
rect 4772 61988 4776 62044
rect 4712 61984 4776 61988
rect 4792 62044 4856 62048
rect 4792 61988 4796 62044
rect 4796 61988 4852 62044
rect 4852 61988 4856 62044
rect 4792 61984 4856 61988
rect 6152 62044 6216 62048
rect 6152 61988 6156 62044
rect 6156 61988 6212 62044
rect 6212 61988 6216 62044
rect 6152 61984 6216 61988
rect 6232 62044 6296 62048
rect 6232 61988 6236 62044
rect 6236 61988 6292 62044
rect 6292 61988 6296 62044
rect 6232 61984 6296 61988
rect 6312 62044 6376 62048
rect 6312 61988 6316 62044
rect 6316 61988 6372 62044
rect 6372 61988 6376 62044
rect 6312 61984 6376 61988
rect 6392 62044 6456 62048
rect 6392 61988 6396 62044
rect 6396 61988 6452 62044
rect 6452 61988 6456 62044
rect 6392 61984 6456 61988
rect 7752 62044 7816 62048
rect 7752 61988 7756 62044
rect 7756 61988 7812 62044
rect 7812 61988 7816 62044
rect 7752 61984 7816 61988
rect 7832 62044 7896 62048
rect 7832 61988 7836 62044
rect 7836 61988 7892 62044
rect 7892 61988 7896 62044
rect 7832 61984 7896 61988
rect 7912 62044 7976 62048
rect 7912 61988 7916 62044
rect 7916 61988 7972 62044
rect 7972 61988 7976 62044
rect 7912 61984 7976 61988
rect 7992 62044 8056 62048
rect 7992 61988 7996 62044
rect 7996 61988 8052 62044
rect 8052 61988 8056 62044
rect 7992 61984 8056 61988
rect 9352 62044 9416 62048
rect 9352 61988 9356 62044
rect 9356 61988 9412 62044
rect 9412 61988 9416 62044
rect 9352 61984 9416 61988
rect 9432 62044 9496 62048
rect 9432 61988 9436 62044
rect 9436 61988 9492 62044
rect 9492 61988 9496 62044
rect 9432 61984 9496 61988
rect 9512 62044 9576 62048
rect 9512 61988 9516 62044
rect 9516 61988 9572 62044
rect 9572 61988 9576 62044
rect 9512 61984 9576 61988
rect 9592 62044 9656 62048
rect 9592 61988 9596 62044
rect 9596 61988 9652 62044
rect 9652 61988 9656 62044
rect 9592 61984 9656 61988
rect 3612 61500 3676 61504
rect 3612 61444 3616 61500
rect 3616 61444 3672 61500
rect 3672 61444 3676 61500
rect 3612 61440 3676 61444
rect 3692 61500 3756 61504
rect 3692 61444 3696 61500
rect 3696 61444 3752 61500
rect 3752 61444 3756 61500
rect 3692 61440 3756 61444
rect 3772 61500 3836 61504
rect 3772 61444 3776 61500
rect 3776 61444 3832 61500
rect 3832 61444 3836 61500
rect 3772 61440 3836 61444
rect 3852 61500 3916 61504
rect 3852 61444 3856 61500
rect 3856 61444 3912 61500
rect 3912 61444 3916 61500
rect 3852 61440 3916 61444
rect 5212 61500 5276 61504
rect 5212 61444 5216 61500
rect 5216 61444 5272 61500
rect 5272 61444 5276 61500
rect 5212 61440 5276 61444
rect 5292 61500 5356 61504
rect 5292 61444 5296 61500
rect 5296 61444 5352 61500
rect 5352 61444 5356 61500
rect 5292 61440 5356 61444
rect 5372 61500 5436 61504
rect 5372 61444 5376 61500
rect 5376 61444 5432 61500
rect 5432 61444 5436 61500
rect 5372 61440 5436 61444
rect 5452 61500 5516 61504
rect 5452 61444 5456 61500
rect 5456 61444 5512 61500
rect 5512 61444 5516 61500
rect 5452 61440 5516 61444
rect 6812 61500 6876 61504
rect 6812 61444 6816 61500
rect 6816 61444 6872 61500
rect 6872 61444 6876 61500
rect 6812 61440 6876 61444
rect 6892 61500 6956 61504
rect 6892 61444 6896 61500
rect 6896 61444 6952 61500
rect 6952 61444 6956 61500
rect 6892 61440 6956 61444
rect 6972 61500 7036 61504
rect 6972 61444 6976 61500
rect 6976 61444 7032 61500
rect 7032 61444 7036 61500
rect 6972 61440 7036 61444
rect 7052 61500 7116 61504
rect 7052 61444 7056 61500
rect 7056 61444 7112 61500
rect 7112 61444 7116 61500
rect 7052 61440 7116 61444
rect 8412 61500 8476 61504
rect 8412 61444 8416 61500
rect 8416 61444 8472 61500
rect 8472 61444 8476 61500
rect 8412 61440 8476 61444
rect 8492 61500 8556 61504
rect 8492 61444 8496 61500
rect 8496 61444 8552 61500
rect 8552 61444 8556 61500
rect 8492 61440 8556 61444
rect 8572 61500 8636 61504
rect 8572 61444 8576 61500
rect 8576 61444 8632 61500
rect 8632 61444 8636 61500
rect 8572 61440 8636 61444
rect 8652 61500 8716 61504
rect 8652 61444 8656 61500
rect 8656 61444 8712 61500
rect 8712 61444 8716 61500
rect 8652 61440 8716 61444
rect 2952 60956 3016 60960
rect 2952 60900 2956 60956
rect 2956 60900 3012 60956
rect 3012 60900 3016 60956
rect 2952 60896 3016 60900
rect 3032 60956 3096 60960
rect 3032 60900 3036 60956
rect 3036 60900 3092 60956
rect 3092 60900 3096 60956
rect 3032 60896 3096 60900
rect 3112 60956 3176 60960
rect 3112 60900 3116 60956
rect 3116 60900 3172 60956
rect 3172 60900 3176 60956
rect 3112 60896 3176 60900
rect 3192 60956 3256 60960
rect 3192 60900 3196 60956
rect 3196 60900 3252 60956
rect 3252 60900 3256 60956
rect 3192 60896 3256 60900
rect 4552 60956 4616 60960
rect 4552 60900 4556 60956
rect 4556 60900 4612 60956
rect 4612 60900 4616 60956
rect 4552 60896 4616 60900
rect 4632 60956 4696 60960
rect 4632 60900 4636 60956
rect 4636 60900 4692 60956
rect 4692 60900 4696 60956
rect 4632 60896 4696 60900
rect 4712 60956 4776 60960
rect 4712 60900 4716 60956
rect 4716 60900 4772 60956
rect 4772 60900 4776 60956
rect 4712 60896 4776 60900
rect 4792 60956 4856 60960
rect 4792 60900 4796 60956
rect 4796 60900 4852 60956
rect 4852 60900 4856 60956
rect 4792 60896 4856 60900
rect 6152 60956 6216 60960
rect 6152 60900 6156 60956
rect 6156 60900 6212 60956
rect 6212 60900 6216 60956
rect 6152 60896 6216 60900
rect 6232 60956 6296 60960
rect 6232 60900 6236 60956
rect 6236 60900 6292 60956
rect 6292 60900 6296 60956
rect 6232 60896 6296 60900
rect 6312 60956 6376 60960
rect 6312 60900 6316 60956
rect 6316 60900 6372 60956
rect 6372 60900 6376 60956
rect 6312 60896 6376 60900
rect 6392 60956 6456 60960
rect 6392 60900 6396 60956
rect 6396 60900 6452 60956
rect 6452 60900 6456 60956
rect 6392 60896 6456 60900
rect 7752 60956 7816 60960
rect 7752 60900 7756 60956
rect 7756 60900 7812 60956
rect 7812 60900 7816 60956
rect 7752 60896 7816 60900
rect 7832 60956 7896 60960
rect 7832 60900 7836 60956
rect 7836 60900 7892 60956
rect 7892 60900 7896 60956
rect 7832 60896 7896 60900
rect 7912 60956 7976 60960
rect 7912 60900 7916 60956
rect 7916 60900 7972 60956
rect 7972 60900 7976 60956
rect 7912 60896 7976 60900
rect 7992 60956 8056 60960
rect 7992 60900 7996 60956
rect 7996 60900 8052 60956
rect 8052 60900 8056 60956
rect 7992 60896 8056 60900
rect 9352 60956 9416 60960
rect 9352 60900 9356 60956
rect 9356 60900 9412 60956
rect 9412 60900 9416 60956
rect 9352 60896 9416 60900
rect 9432 60956 9496 60960
rect 9432 60900 9436 60956
rect 9436 60900 9492 60956
rect 9492 60900 9496 60956
rect 9432 60896 9496 60900
rect 9512 60956 9576 60960
rect 9512 60900 9516 60956
rect 9516 60900 9572 60956
rect 9572 60900 9576 60956
rect 9512 60896 9576 60900
rect 9592 60956 9656 60960
rect 9592 60900 9596 60956
rect 9596 60900 9652 60956
rect 9652 60900 9656 60956
rect 9592 60896 9656 60900
rect 3612 60412 3676 60416
rect 3612 60356 3616 60412
rect 3616 60356 3672 60412
rect 3672 60356 3676 60412
rect 3612 60352 3676 60356
rect 3692 60412 3756 60416
rect 3692 60356 3696 60412
rect 3696 60356 3752 60412
rect 3752 60356 3756 60412
rect 3692 60352 3756 60356
rect 3772 60412 3836 60416
rect 3772 60356 3776 60412
rect 3776 60356 3832 60412
rect 3832 60356 3836 60412
rect 3772 60352 3836 60356
rect 3852 60412 3916 60416
rect 3852 60356 3856 60412
rect 3856 60356 3912 60412
rect 3912 60356 3916 60412
rect 3852 60352 3916 60356
rect 5212 60412 5276 60416
rect 5212 60356 5216 60412
rect 5216 60356 5272 60412
rect 5272 60356 5276 60412
rect 5212 60352 5276 60356
rect 5292 60412 5356 60416
rect 5292 60356 5296 60412
rect 5296 60356 5352 60412
rect 5352 60356 5356 60412
rect 5292 60352 5356 60356
rect 5372 60412 5436 60416
rect 5372 60356 5376 60412
rect 5376 60356 5432 60412
rect 5432 60356 5436 60412
rect 5372 60352 5436 60356
rect 5452 60412 5516 60416
rect 5452 60356 5456 60412
rect 5456 60356 5512 60412
rect 5512 60356 5516 60412
rect 5452 60352 5516 60356
rect 6812 60412 6876 60416
rect 6812 60356 6816 60412
rect 6816 60356 6872 60412
rect 6872 60356 6876 60412
rect 6812 60352 6876 60356
rect 6892 60412 6956 60416
rect 6892 60356 6896 60412
rect 6896 60356 6952 60412
rect 6952 60356 6956 60412
rect 6892 60352 6956 60356
rect 6972 60412 7036 60416
rect 6972 60356 6976 60412
rect 6976 60356 7032 60412
rect 7032 60356 7036 60412
rect 6972 60352 7036 60356
rect 7052 60412 7116 60416
rect 7052 60356 7056 60412
rect 7056 60356 7112 60412
rect 7112 60356 7116 60412
rect 7052 60352 7116 60356
rect 8412 60412 8476 60416
rect 8412 60356 8416 60412
rect 8416 60356 8472 60412
rect 8472 60356 8476 60412
rect 8412 60352 8476 60356
rect 8492 60412 8556 60416
rect 8492 60356 8496 60412
rect 8496 60356 8552 60412
rect 8552 60356 8556 60412
rect 8492 60352 8556 60356
rect 8572 60412 8636 60416
rect 8572 60356 8576 60412
rect 8576 60356 8632 60412
rect 8632 60356 8636 60412
rect 8572 60352 8636 60356
rect 8652 60412 8716 60416
rect 8652 60356 8656 60412
rect 8656 60356 8712 60412
rect 8712 60356 8716 60412
rect 8652 60352 8716 60356
rect 2952 59868 3016 59872
rect 2952 59812 2956 59868
rect 2956 59812 3012 59868
rect 3012 59812 3016 59868
rect 2952 59808 3016 59812
rect 3032 59868 3096 59872
rect 3032 59812 3036 59868
rect 3036 59812 3092 59868
rect 3092 59812 3096 59868
rect 3032 59808 3096 59812
rect 3112 59868 3176 59872
rect 3112 59812 3116 59868
rect 3116 59812 3172 59868
rect 3172 59812 3176 59868
rect 3112 59808 3176 59812
rect 3192 59868 3256 59872
rect 3192 59812 3196 59868
rect 3196 59812 3252 59868
rect 3252 59812 3256 59868
rect 3192 59808 3256 59812
rect 4552 59868 4616 59872
rect 4552 59812 4556 59868
rect 4556 59812 4612 59868
rect 4612 59812 4616 59868
rect 4552 59808 4616 59812
rect 4632 59868 4696 59872
rect 4632 59812 4636 59868
rect 4636 59812 4692 59868
rect 4692 59812 4696 59868
rect 4632 59808 4696 59812
rect 4712 59868 4776 59872
rect 4712 59812 4716 59868
rect 4716 59812 4772 59868
rect 4772 59812 4776 59868
rect 4712 59808 4776 59812
rect 4792 59868 4856 59872
rect 4792 59812 4796 59868
rect 4796 59812 4852 59868
rect 4852 59812 4856 59868
rect 4792 59808 4856 59812
rect 6152 59868 6216 59872
rect 6152 59812 6156 59868
rect 6156 59812 6212 59868
rect 6212 59812 6216 59868
rect 6152 59808 6216 59812
rect 6232 59868 6296 59872
rect 6232 59812 6236 59868
rect 6236 59812 6292 59868
rect 6292 59812 6296 59868
rect 6232 59808 6296 59812
rect 6312 59868 6376 59872
rect 6312 59812 6316 59868
rect 6316 59812 6372 59868
rect 6372 59812 6376 59868
rect 6312 59808 6376 59812
rect 6392 59868 6456 59872
rect 6392 59812 6396 59868
rect 6396 59812 6452 59868
rect 6452 59812 6456 59868
rect 6392 59808 6456 59812
rect 7752 59868 7816 59872
rect 7752 59812 7756 59868
rect 7756 59812 7812 59868
rect 7812 59812 7816 59868
rect 7752 59808 7816 59812
rect 7832 59868 7896 59872
rect 7832 59812 7836 59868
rect 7836 59812 7892 59868
rect 7892 59812 7896 59868
rect 7832 59808 7896 59812
rect 7912 59868 7976 59872
rect 7912 59812 7916 59868
rect 7916 59812 7972 59868
rect 7972 59812 7976 59868
rect 7912 59808 7976 59812
rect 7992 59868 8056 59872
rect 7992 59812 7996 59868
rect 7996 59812 8052 59868
rect 8052 59812 8056 59868
rect 7992 59808 8056 59812
rect 9352 59868 9416 59872
rect 9352 59812 9356 59868
rect 9356 59812 9412 59868
rect 9412 59812 9416 59868
rect 9352 59808 9416 59812
rect 9432 59868 9496 59872
rect 9432 59812 9436 59868
rect 9436 59812 9492 59868
rect 9492 59812 9496 59868
rect 9432 59808 9496 59812
rect 9512 59868 9576 59872
rect 9512 59812 9516 59868
rect 9516 59812 9572 59868
rect 9572 59812 9576 59868
rect 9512 59808 9576 59812
rect 9592 59868 9656 59872
rect 9592 59812 9596 59868
rect 9596 59812 9652 59868
rect 9652 59812 9656 59868
rect 9592 59808 9656 59812
rect 3612 59324 3676 59328
rect 3612 59268 3616 59324
rect 3616 59268 3672 59324
rect 3672 59268 3676 59324
rect 3612 59264 3676 59268
rect 3692 59324 3756 59328
rect 3692 59268 3696 59324
rect 3696 59268 3752 59324
rect 3752 59268 3756 59324
rect 3692 59264 3756 59268
rect 3772 59324 3836 59328
rect 3772 59268 3776 59324
rect 3776 59268 3832 59324
rect 3832 59268 3836 59324
rect 3772 59264 3836 59268
rect 3852 59324 3916 59328
rect 3852 59268 3856 59324
rect 3856 59268 3912 59324
rect 3912 59268 3916 59324
rect 3852 59264 3916 59268
rect 5212 59324 5276 59328
rect 5212 59268 5216 59324
rect 5216 59268 5272 59324
rect 5272 59268 5276 59324
rect 5212 59264 5276 59268
rect 5292 59324 5356 59328
rect 5292 59268 5296 59324
rect 5296 59268 5352 59324
rect 5352 59268 5356 59324
rect 5292 59264 5356 59268
rect 5372 59324 5436 59328
rect 5372 59268 5376 59324
rect 5376 59268 5432 59324
rect 5432 59268 5436 59324
rect 5372 59264 5436 59268
rect 5452 59324 5516 59328
rect 5452 59268 5456 59324
rect 5456 59268 5512 59324
rect 5512 59268 5516 59324
rect 5452 59264 5516 59268
rect 6812 59324 6876 59328
rect 6812 59268 6816 59324
rect 6816 59268 6872 59324
rect 6872 59268 6876 59324
rect 6812 59264 6876 59268
rect 6892 59324 6956 59328
rect 6892 59268 6896 59324
rect 6896 59268 6952 59324
rect 6952 59268 6956 59324
rect 6892 59264 6956 59268
rect 6972 59324 7036 59328
rect 6972 59268 6976 59324
rect 6976 59268 7032 59324
rect 7032 59268 7036 59324
rect 6972 59264 7036 59268
rect 7052 59324 7116 59328
rect 7052 59268 7056 59324
rect 7056 59268 7112 59324
rect 7112 59268 7116 59324
rect 7052 59264 7116 59268
rect 8412 59324 8476 59328
rect 8412 59268 8416 59324
rect 8416 59268 8472 59324
rect 8472 59268 8476 59324
rect 8412 59264 8476 59268
rect 8492 59324 8556 59328
rect 8492 59268 8496 59324
rect 8496 59268 8552 59324
rect 8552 59268 8556 59324
rect 8492 59264 8556 59268
rect 8572 59324 8636 59328
rect 8572 59268 8576 59324
rect 8576 59268 8632 59324
rect 8632 59268 8636 59324
rect 8572 59264 8636 59268
rect 8652 59324 8716 59328
rect 8652 59268 8656 59324
rect 8656 59268 8712 59324
rect 8712 59268 8716 59324
rect 8652 59264 8716 59268
rect 2952 58780 3016 58784
rect 2952 58724 2956 58780
rect 2956 58724 3012 58780
rect 3012 58724 3016 58780
rect 2952 58720 3016 58724
rect 3032 58780 3096 58784
rect 3032 58724 3036 58780
rect 3036 58724 3092 58780
rect 3092 58724 3096 58780
rect 3032 58720 3096 58724
rect 3112 58780 3176 58784
rect 3112 58724 3116 58780
rect 3116 58724 3172 58780
rect 3172 58724 3176 58780
rect 3112 58720 3176 58724
rect 3192 58780 3256 58784
rect 3192 58724 3196 58780
rect 3196 58724 3252 58780
rect 3252 58724 3256 58780
rect 3192 58720 3256 58724
rect 4552 58780 4616 58784
rect 4552 58724 4556 58780
rect 4556 58724 4612 58780
rect 4612 58724 4616 58780
rect 4552 58720 4616 58724
rect 4632 58780 4696 58784
rect 4632 58724 4636 58780
rect 4636 58724 4692 58780
rect 4692 58724 4696 58780
rect 4632 58720 4696 58724
rect 4712 58780 4776 58784
rect 4712 58724 4716 58780
rect 4716 58724 4772 58780
rect 4772 58724 4776 58780
rect 4712 58720 4776 58724
rect 4792 58780 4856 58784
rect 4792 58724 4796 58780
rect 4796 58724 4852 58780
rect 4852 58724 4856 58780
rect 4792 58720 4856 58724
rect 6152 58780 6216 58784
rect 6152 58724 6156 58780
rect 6156 58724 6212 58780
rect 6212 58724 6216 58780
rect 6152 58720 6216 58724
rect 6232 58780 6296 58784
rect 6232 58724 6236 58780
rect 6236 58724 6292 58780
rect 6292 58724 6296 58780
rect 6232 58720 6296 58724
rect 6312 58780 6376 58784
rect 6312 58724 6316 58780
rect 6316 58724 6372 58780
rect 6372 58724 6376 58780
rect 6312 58720 6376 58724
rect 6392 58780 6456 58784
rect 6392 58724 6396 58780
rect 6396 58724 6452 58780
rect 6452 58724 6456 58780
rect 6392 58720 6456 58724
rect 7752 58780 7816 58784
rect 7752 58724 7756 58780
rect 7756 58724 7812 58780
rect 7812 58724 7816 58780
rect 7752 58720 7816 58724
rect 7832 58780 7896 58784
rect 7832 58724 7836 58780
rect 7836 58724 7892 58780
rect 7892 58724 7896 58780
rect 7832 58720 7896 58724
rect 7912 58780 7976 58784
rect 7912 58724 7916 58780
rect 7916 58724 7972 58780
rect 7972 58724 7976 58780
rect 7912 58720 7976 58724
rect 7992 58780 8056 58784
rect 7992 58724 7996 58780
rect 7996 58724 8052 58780
rect 8052 58724 8056 58780
rect 7992 58720 8056 58724
rect 9352 58780 9416 58784
rect 9352 58724 9356 58780
rect 9356 58724 9412 58780
rect 9412 58724 9416 58780
rect 9352 58720 9416 58724
rect 9432 58780 9496 58784
rect 9432 58724 9436 58780
rect 9436 58724 9492 58780
rect 9492 58724 9496 58780
rect 9432 58720 9496 58724
rect 9512 58780 9576 58784
rect 9512 58724 9516 58780
rect 9516 58724 9572 58780
rect 9572 58724 9576 58780
rect 9512 58720 9576 58724
rect 9592 58780 9656 58784
rect 9592 58724 9596 58780
rect 9596 58724 9652 58780
rect 9652 58724 9656 58780
rect 9592 58720 9656 58724
rect 3612 58236 3676 58240
rect 3612 58180 3616 58236
rect 3616 58180 3672 58236
rect 3672 58180 3676 58236
rect 3612 58176 3676 58180
rect 3692 58236 3756 58240
rect 3692 58180 3696 58236
rect 3696 58180 3752 58236
rect 3752 58180 3756 58236
rect 3692 58176 3756 58180
rect 3772 58236 3836 58240
rect 3772 58180 3776 58236
rect 3776 58180 3832 58236
rect 3832 58180 3836 58236
rect 3772 58176 3836 58180
rect 3852 58236 3916 58240
rect 3852 58180 3856 58236
rect 3856 58180 3912 58236
rect 3912 58180 3916 58236
rect 3852 58176 3916 58180
rect 5212 58236 5276 58240
rect 5212 58180 5216 58236
rect 5216 58180 5272 58236
rect 5272 58180 5276 58236
rect 5212 58176 5276 58180
rect 5292 58236 5356 58240
rect 5292 58180 5296 58236
rect 5296 58180 5352 58236
rect 5352 58180 5356 58236
rect 5292 58176 5356 58180
rect 5372 58236 5436 58240
rect 5372 58180 5376 58236
rect 5376 58180 5432 58236
rect 5432 58180 5436 58236
rect 5372 58176 5436 58180
rect 5452 58236 5516 58240
rect 5452 58180 5456 58236
rect 5456 58180 5512 58236
rect 5512 58180 5516 58236
rect 5452 58176 5516 58180
rect 6812 58236 6876 58240
rect 6812 58180 6816 58236
rect 6816 58180 6872 58236
rect 6872 58180 6876 58236
rect 6812 58176 6876 58180
rect 6892 58236 6956 58240
rect 6892 58180 6896 58236
rect 6896 58180 6952 58236
rect 6952 58180 6956 58236
rect 6892 58176 6956 58180
rect 6972 58236 7036 58240
rect 6972 58180 6976 58236
rect 6976 58180 7032 58236
rect 7032 58180 7036 58236
rect 6972 58176 7036 58180
rect 7052 58236 7116 58240
rect 7052 58180 7056 58236
rect 7056 58180 7112 58236
rect 7112 58180 7116 58236
rect 7052 58176 7116 58180
rect 8412 58236 8476 58240
rect 8412 58180 8416 58236
rect 8416 58180 8472 58236
rect 8472 58180 8476 58236
rect 8412 58176 8476 58180
rect 8492 58236 8556 58240
rect 8492 58180 8496 58236
rect 8496 58180 8552 58236
rect 8552 58180 8556 58236
rect 8492 58176 8556 58180
rect 8572 58236 8636 58240
rect 8572 58180 8576 58236
rect 8576 58180 8632 58236
rect 8632 58180 8636 58236
rect 8572 58176 8636 58180
rect 8652 58236 8716 58240
rect 8652 58180 8656 58236
rect 8656 58180 8712 58236
rect 8712 58180 8716 58236
rect 8652 58176 8716 58180
rect 2952 57692 3016 57696
rect 2952 57636 2956 57692
rect 2956 57636 3012 57692
rect 3012 57636 3016 57692
rect 2952 57632 3016 57636
rect 3032 57692 3096 57696
rect 3032 57636 3036 57692
rect 3036 57636 3092 57692
rect 3092 57636 3096 57692
rect 3032 57632 3096 57636
rect 3112 57692 3176 57696
rect 3112 57636 3116 57692
rect 3116 57636 3172 57692
rect 3172 57636 3176 57692
rect 3112 57632 3176 57636
rect 3192 57692 3256 57696
rect 3192 57636 3196 57692
rect 3196 57636 3252 57692
rect 3252 57636 3256 57692
rect 3192 57632 3256 57636
rect 4552 57692 4616 57696
rect 4552 57636 4556 57692
rect 4556 57636 4612 57692
rect 4612 57636 4616 57692
rect 4552 57632 4616 57636
rect 4632 57692 4696 57696
rect 4632 57636 4636 57692
rect 4636 57636 4692 57692
rect 4692 57636 4696 57692
rect 4632 57632 4696 57636
rect 4712 57692 4776 57696
rect 4712 57636 4716 57692
rect 4716 57636 4772 57692
rect 4772 57636 4776 57692
rect 4712 57632 4776 57636
rect 4792 57692 4856 57696
rect 4792 57636 4796 57692
rect 4796 57636 4852 57692
rect 4852 57636 4856 57692
rect 4792 57632 4856 57636
rect 6152 57692 6216 57696
rect 6152 57636 6156 57692
rect 6156 57636 6212 57692
rect 6212 57636 6216 57692
rect 6152 57632 6216 57636
rect 6232 57692 6296 57696
rect 6232 57636 6236 57692
rect 6236 57636 6292 57692
rect 6292 57636 6296 57692
rect 6232 57632 6296 57636
rect 6312 57692 6376 57696
rect 6312 57636 6316 57692
rect 6316 57636 6372 57692
rect 6372 57636 6376 57692
rect 6312 57632 6376 57636
rect 6392 57692 6456 57696
rect 6392 57636 6396 57692
rect 6396 57636 6452 57692
rect 6452 57636 6456 57692
rect 6392 57632 6456 57636
rect 7752 57692 7816 57696
rect 7752 57636 7756 57692
rect 7756 57636 7812 57692
rect 7812 57636 7816 57692
rect 7752 57632 7816 57636
rect 7832 57692 7896 57696
rect 7832 57636 7836 57692
rect 7836 57636 7892 57692
rect 7892 57636 7896 57692
rect 7832 57632 7896 57636
rect 7912 57692 7976 57696
rect 7912 57636 7916 57692
rect 7916 57636 7972 57692
rect 7972 57636 7976 57692
rect 7912 57632 7976 57636
rect 7992 57692 8056 57696
rect 7992 57636 7996 57692
rect 7996 57636 8052 57692
rect 8052 57636 8056 57692
rect 7992 57632 8056 57636
rect 9352 57692 9416 57696
rect 9352 57636 9356 57692
rect 9356 57636 9412 57692
rect 9412 57636 9416 57692
rect 9352 57632 9416 57636
rect 9432 57692 9496 57696
rect 9432 57636 9436 57692
rect 9436 57636 9492 57692
rect 9492 57636 9496 57692
rect 9432 57632 9496 57636
rect 9512 57692 9576 57696
rect 9512 57636 9516 57692
rect 9516 57636 9572 57692
rect 9572 57636 9576 57692
rect 9512 57632 9576 57636
rect 9592 57692 9656 57696
rect 9592 57636 9596 57692
rect 9596 57636 9652 57692
rect 9652 57636 9656 57692
rect 9592 57632 9656 57636
rect 3612 57148 3676 57152
rect 3612 57092 3616 57148
rect 3616 57092 3672 57148
rect 3672 57092 3676 57148
rect 3612 57088 3676 57092
rect 3692 57148 3756 57152
rect 3692 57092 3696 57148
rect 3696 57092 3752 57148
rect 3752 57092 3756 57148
rect 3692 57088 3756 57092
rect 3772 57148 3836 57152
rect 3772 57092 3776 57148
rect 3776 57092 3832 57148
rect 3832 57092 3836 57148
rect 3772 57088 3836 57092
rect 3852 57148 3916 57152
rect 3852 57092 3856 57148
rect 3856 57092 3912 57148
rect 3912 57092 3916 57148
rect 3852 57088 3916 57092
rect 5212 57148 5276 57152
rect 5212 57092 5216 57148
rect 5216 57092 5272 57148
rect 5272 57092 5276 57148
rect 5212 57088 5276 57092
rect 5292 57148 5356 57152
rect 5292 57092 5296 57148
rect 5296 57092 5352 57148
rect 5352 57092 5356 57148
rect 5292 57088 5356 57092
rect 5372 57148 5436 57152
rect 5372 57092 5376 57148
rect 5376 57092 5432 57148
rect 5432 57092 5436 57148
rect 5372 57088 5436 57092
rect 5452 57148 5516 57152
rect 5452 57092 5456 57148
rect 5456 57092 5512 57148
rect 5512 57092 5516 57148
rect 5452 57088 5516 57092
rect 6812 57148 6876 57152
rect 6812 57092 6816 57148
rect 6816 57092 6872 57148
rect 6872 57092 6876 57148
rect 6812 57088 6876 57092
rect 6892 57148 6956 57152
rect 6892 57092 6896 57148
rect 6896 57092 6952 57148
rect 6952 57092 6956 57148
rect 6892 57088 6956 57092
rect 6972 57148 7036 57152
rect 6972 57092 6976 57148
rect 6976 57092 7032 57148
rect 7032 57092 7036 57148
rect 6972 57088 7036 57092
rect 7052 57148 7116 57152
rect 7052 57092 7056 57148
rect 7056 57092 7112 57148
rect 7112 57092 7116 57148
rect 7052 57088 7116 57092
rect 8412 57148 8476 57152
rect 8412 57092 8416 57148
rect 8416 57092 8472 57148
rect 8472 57092 8476 57148
rect 8412 57088 8476 57092
rect 8492 57148 8556 57152
rect 8492 57092 8496 57148
rect 8496 57092 8552 57148
rect 8552 57092 8556 57148
rect 8492 57088 8556 57092
rect 8572 57148 8636 57152
rect 8572 57092 8576 57148
rect 8576 57092 8632 57148
rect 8632 57092 8636 57148
rect 8572 57088 8636 57092
rect 8652 57148 8716 57152
rect 8652 57092 8656 57148
rect 8656 57092 8712 57148
rect 8712 57092 8716 57148
rect 8652 57088 8716 57092
rect 2952 56604 3016 56608
rect 2952 56548 2956 56604
rect 2956 56548 3012 56604
rect 3012 56548 3016 56604
rect 2952 56544 3016 56548
rect 3032 56604 3096 56608
rect 3032 56548 3036 56604
rect 3036 56548 3092 56604
rect 3092 56548 3096 56604
rect 3032 56544 3096 56548
rect 3112 56604 3176 56608
rect 3112 56548 3116 56604
rect 3116 56548 3172 56604
rect 3172 56548 3176 56604
rect 3112 56544 3176 56548
rect 3192 56604 3256 56608
rect 3192 56548 3196 56604
rect 3196 56548 3252 56604
rect 3252 56548 3256 56604
rect 3192 56544 3256 56548
rect 4552 56604 4616 56608
rect 4552 56548 4556 56604
rect 4556 56548 4612 56604
rect 4612 56548 4616 56604
rect 4552 56544 4616 56548
rect 4632 56604 4696 56608
rect 4632 56548 4636 56604
rect 4636 56548 4692 56604
rect 4692 56548 4696 56604
rect 4632 56544 4696 56548
rect 4712 56604 4776 56608
rect 4712 56548 4716 56604
rect 4716 56548 4772 56604
rect 4772 56548 4776 56604
rect 4712 56544 4776 56548
rect 4792 56604 4856 56608
rect 4792 56548 4796 56604
rect 4796 56548 4852 56604
rect 4852 56548 4856 56604
rect 4792 56544 4856 56548
rect 6152 56604 6216 56608
rect 6152 56548 6156 56604
rect 6156 56548 6212 56604
rect 6212 56548 6216 56604
rect 6152 56544 6216 56548
rect 6232 56604 6296 56608
rect 6232 56548 6236 56604
rect 6236 56548 6292 56604
rect 6292 56548 6296 56604
rect 6232 56544 6296 56548
rect 6312 56604 6376 56608
rect 6312 56548 6316 56604
rect 6316 56548 6372 56604
rect 6372 56548 6376 56604
rect 6312 56544 6376 56548
rect 6392 56604 6456 56608
rect 6392 56548 6396 56604
rect 6396 56548 6452 56604
rect 6452 56548 6456 56604
rect 6392 56544 6456 56548
rect 7752 56604 7816 56608
rect 7752 56548 7756 56604
rect 7756 56548 7812 56604
rect 7812 56548 7816 56604
rect 7752 56544 7816 56548
rect 7832 56604 7896 56608
rect 7832 56548 7836 56604
rect 7836 56548 7892 56604
rect 7892 56548 7896 56604
rect 7832 56544 7896 56548
rect 7912 56604 7976 56608
rect 7912 56548 7916 56604
rect 7916 56548 7972 56604
rect 7972 56548 7976 56604
rect 7912 56544 7976 56548
rect 7992 56604 8056 56608
rect 7992 56548 7996 56604
rect 7996 56548 8052 56604
rect 8052 56548 8056 56604
rect 7992 56544 8056 56548
rect 9352 56604 9416 56608
rect 9352 56548 9356 56604
rect 9356 56548 9412 56604
rect 9412 56548 9416 56604
rect 9352 56544 9416 56548
rect 9432 56604 9496 56608
rect 9432 56548 9436 56604
rect 9436 56548 9492 56604
rect 9492 56548 9496 56604
rect 9432 56544 9496 56548
rect 9512 56604 9576 56608
rect 9512 56548 9516 56604
rect 9516 56548 9572 56604
rect 9572 56548 9576 56604
rect 9512 56544 9576 56548
rect 9592 56604 9656 56608
rect 9592 56548 9596 56604
rect 9596 56548 9652 56604
rect 9652 56548 9656 56604
rect 9592 56544 9656 56548
rect 3612 56060 3676 56064
rect 3612 56004 3616 56060
rect 3616 56004 3672 56060
rect 3672 56004 3676 56060
rect 3612 56000 3676 56004
rect 3692 56060 3756 56064
rect 3692 56004 3696 56060
rect 3696 56004 3752 56060
rect 3752 56004 3756 56060
rect 3692 56000 3756 56004
rect 3772 56060 3836 56064
rect 3772 56004 3776 56060
rect 3776 56004 3832 56060
rect 3832 56004 3836 56060
rect 3772 56000 3836 56004
rect 3852 56060 3916 56064
rect 3852 56004 3856 56060
rect 3856 56004 3912 56060
rect 3912 56004 3916 56060
rect 3852 56000 3916 56004
rect 5212 56060 5276 56064
rect 5212 56004 5216 56060
rect 5216 56004 5272 56060
rect 5272 56004 5276 56060
rect 5212 56000 5276 56004
rect 5292 56060 5356 56064
rect 5292 56004 5296 56060
rect 5296 56004 5352 56060
rect 5352 56004 5356 56060
rect 5292 56000 5356 56004
rect 5372 56060 5436 56064
rect 5372 56004 5376 56060
rect 5376 56004 5432 56060
rect 5432 56004 5436 56060
rect 5372 56000 5436 56004
rect 5452 56060 5516 56064
rect 5452 56004 5456 56060
rect 5456 56004 5512 56060
rect 5512 56004 5516 56060
rect 5452 56000 5516 56004
rect 6812 56060 6876 56064
rect 6812 56004 6816 56060
rect 6816 56004 6872 56060
rect 6872 56004 6876 56060
rect 6812 56000 6876 56004
rect 6892 56060 6956 56064
rect 6892 56004 6896 56060
rect 6896 56004 6952 56060
rect 6952 56004 6956 56060
rect 6892 56000 6956 56004
rect 6972 56060 7036 56064
rect 6972 56004 6976 56060
rect 6976 56004 7032 56060
rect 7032 56004 7036 56060
rect 6972 56000 7036 56004
rect 7052 56060 7116 56064
rect 7052 56004 7056 56060
rect 7056 56004 7112 56060
rect 7112 56004 7116 56060
rect 7052 56000 7116 56004
rect 8412 56060 8476 56064
rect 8412 56004 8416 56060
rect 8416 56004 8472 56060
rect 8472 56004 8476 56060
rect 8412 56000 8476 56004
rect 8492 56060 8556 56064
rect 8492 56004 8496 56060
rect 8496 56004 8552 56060
rect 8552 56004 8556 56060
rect 8492 56000 8556 56004
rect 8572 56060 8636 56064
rect 8572 56004 8576 56060
rect 8576 56004 8632 56060
rect 8632 56004 8636 56060
rect 8572 56000 8636 56004
rect 8652 56060 8716 56064
rect 8652 56004 8656 56060
rect 8656 56004 8712 56060
rect 8712 56004 8716 56060
rect 8652 56000 8716 56004
rect 2952 55516 3016 55520
rect 2952 55460 2956 55516
rect 2956 55460 3012 55516
rect 3012 55460 3016 55516
rect 2952 55456 3016 55460
rect 3032 55516 3096 55520
rect 3032 55460 3036 55516
rect 3036 55460 3092 55516
rect 3092 55460 3096 55516
rect 3032 55456 3096 55460
rect 3112 55516 3176 55520
rect 3112 55460 3116 55516
rect 3116 55460 3172 55516
rect 3172 55460 3176 55516
rect 3112 55456 3176 55460
rect 3192 55516 3256 55520
rect 3192 55460 3196 55516
rect 3196 55460 3252 55516
rect 3252 55460 3256 55516
rect 3192 55456 3256 55460
rect 4552 55516 4616 55520
rect 4552 55460 4556 55516
rect 4556 55460 4612 55516
rect 4612 55460 4616 55516
rect 4552 55456 4616 55460
rect 4632 55516 4696 55520
rect 4632 55460 4636 55516
rect 4636 55460 4692 55516
rect 4692 55460 4696 55516
rect 4632 55456 4696 55460
rect 4712 55516 4776 55520
rect 4712 55460 4716 55516
rect 4716 55460 4772 55516
rect 4772 55460 4776 55516
rect 4712 55456 4776 55460
rect 4792 55516 4856 55520
rect 4792 55460 4796 55516
rect 4796 55460 4852 55516
rect 4852 55460 4856 55516
rect 4792 55456 4856 55460
rect 6152 55516 6216 55520
rect 6152 55460 6156 55516
rect 6156 55460 6212 55516
rect 6212 55460 6216 55516
rect 6152 55456 6216 55460
rect 6232 55516 6296 55520
rect 6232 55460 6236 55516
rect 6236 55460 6292 55516
rect 6292 55460 6296 55516
rect 6232 55456 6296 55460
rect 6312 55516 6376 55520
rect 6312 55460 6316 55516
rect 6316 55460 6372 55516
rect 6372 55460 6376 55516
rect 6312 55456 6376 55460
rect 6392 55516 6456 55520
rect 6392 55460 6396 55516
rect 6396 55460 6452 55516
rect 6452 55460 6456 55516
rect 6392 55456 6456 55460
rect 7752 55516 7816 55520
rect 7752 55460 7756 55516
rect 7756 55460 7812 55516
rect 7812 55460 7816 55516
rect 7752 55456 7816 55460
rect 7832 55516 7896 55520
rect 7832 55460 7836 55516
rect 7836 55460 7892 55516
rect 7892 55460 7896 55516
rect 7832 55456 7896 55460
rect 7912 55516 7976 55520
rect 7912 55460 7916 55516
rect 7916 55460 7972 55516
rect 7972 55460 7976 55516
rect 7912 55456 7976 55460
rect 7992 55516 8056 55520
rect 7992 55460 7996 55516
rect 7996 55460 8052 55516
rect 8052 55460 8056 55516
rect 7992 55456 8056 55460
rect 9352 55516 9416 55520
rect 9352 55460 9356 55516
rect 9356 55460 9412 55516
rect 9412 55460 9416 55516
rect 9352 55456 9416 55460
rect 9432 55516 9496 55520
rect 9432 55460 9436 55516
rect 9436 55460 9492 55516
rect 9492 55460 9496 55516
rect 9432 55456 9496 55460
rect 9512 55516 9576 55520
rect 9512 55460 9516 55516
rect 9516 55460 9572 55516
rect 9572 55460 9576 55516
rect 9512 55456 9576 55460
rect 9592 55516 9656 55520
rect 9592 55460 9596 55516
rect 9596 55460 9652 55516
rect 9652 55460 9656 55516
rect 9592 55456 9656 55460
rect 3612 54972 3676 54976
rect 3612 54916 3616 54972
rect 3616 54916 3672 54972
rect 3672 54916 3676 54972
rect 3612 54912 3676 54916
rect 3692 54972 3756 54976
rect 3692 54916 3696 54972
rect 3696 54916 3752 54972
rect 3752 54916 3756 54972
rect 3692 54912 3756 54916
rect 3772 54972 3836 54976
rect 3772 54916 3776 54972
rect 3776 54916 3832 54972
rect 3832 54916 3836 54972
rect 3772 54912 3836 54916
rect 3852 54972 3916 54976
rect 3852 54916 3856 54972
rect 3856 54916 3912 54972
rect 3912 54916 3916 54972
rect 3852 54912 3916 54916
rect 5212 54972 5276 54976
rect 5212 54916 5216 54972
rect 5216 54916 5272 54972
rect 5272 54916 5276 54972
rect 5212 54912 5276 54916
rect 5292 54972 5356 54976
rect 5292 54916 5296 54972
rect 5296 54916 5352 54972
rect 5352 54916 5356 54972
rect 5292 54912 5356 54916
rect 5372 54972 5436 54976
rect 5372 54916 5376 54972
rect 5376 54916 5432 54972
rect 5432 54916 5436 54972
rect 5372 54912 5436 54916
rect 5452 54972 5516 54976
rect 5452 54916 5456 54972
rect 5456 54916 5512 54972
rect 5512 54916 5516 54972
rect 5452 54912 5516 54916
rect 6812 54972 6876 54976
rect 6812 54916 6816 54972
rect 6816 54916 6872 54972
rect 6872 54916 6876 54972
rect 6812 54912 6876 54916
rect 6892 54972 6956 54976
rect 6892 54916 6896 54972
rect 6896 54916 6952 54972
rect 6952 54916 6956 54972
rect 6892 54912 6956 54916
rect 6972 54972 7036 54976
rect 6972 54916 6976 54972
rect 6976 54916 7032 54972
rect 7032 54916 7036 54972
rect 6972 54912 7036 54916
rect 7052 54972 7116 54976
rect 7052 54916 7056 54972
rect 7056 54916 7112 54972
rect 7112 54916 7116 54972
rect 7052 54912 7116 54916
rect 8412 54972 8476 54976
rect 8412 54916 8416 54972
rect 8416 54916 8472 54972
rect 8472 54916 8476 54972
rect 8412 54912 8476 54916
rect 8492 54972 8556 54976
rect 8492 54916 8496 54972
rect 8496 54916 8552 54972
rect 8552 54916 8556 54972
rect 8492 54912 8556 54916
rect 8572 54972 8636 54976
rect 8572 54916 8576 54972
rect 8576 54916 8632 54972
rect 8632 54916 8636 54972
rect 8572 54912 8636 54916
rect 8652 54972 8716 54976
rect 8652 54916 8656 54972
rect 8656 54916 8712 54972
rect 8712 54916 8716 54972
rect 8652 54912 8716 54916
rect 2952 54428 3016 54432
rect 2952 54372 2956 54428
rect 2956 54372 3012 54428
rect 3012 54372 3016 54428
rect 2952 54368 3016 54372
rect 3032 54428 3096 54432
rect 3032 54372 3036 54428
rect 3036 54372 3092 54428
rect 3092 54372 3096 54428
rect 3032 54368 3096 54372
rect 3112 54428 3176 54432
rect 3112 54372 3116 54428
rect 3116 54372 3172 54428
rect 3172 54372 3176 54428
rect 3112 54368 3176 54372
rect 3192 54428 3256 54432
rect 3192 54372 3196 54428
rect 3196 54372 3252 54428
rect 3252 54372 3256 54428
rect 3192 54368 3256 54372
rect 4552 54428 4616 54432
rect 4552 54372 4556 54428
rect 4556 54372 4612 54428
rect 4612 54372 4616 54428
rect 4552 54368 4616 54372
rect 4632 54428 4696 54432
rect 4632 54372 4636 54428
rect 4636 54372 4692 54428
rect 4692 54372 4696 54428
rect 4632 54368 4696 54372
rect 4712 54428 4776 54432
rect 4712 54372 4716 54428
rect 4716 54372 4772 54428
rect 4772 54372 4776 54428
rect 4712 54368 4776 54372
rect 4792 54428 4856 54432
rect 4792 54372 4796 54428
rect 4796 54372 4852 54428
rect 4852 54372 4856 54428
rect 4792 54368 4856 54372
rect 6152 54428 6216 54432
rect 6152 54372 6156 54428
rect 6156 54372 6212 54428
rect 6212 54372 6216 54428
rect 6152 54368 6216 54372
rect 6232 54428 6296 54432
rect 6232 54372 6236 54428
rect 6236 54372 6292 54428
rect 6292 54372 6296 54428
rect 6232 54368 6296 54372
rect 6312 54428 6376 54432
rect 6312 54372 6316 54428
rect 6316 54372 6372 54428
rect 6372 54372 6376 54428
rect 6312 54368 6376 54372
rect 6392 54428 6456 54432
rect 6392 54372 6396 54428
rect 6396 54372 6452 54428
rect 6452 54372 6456 54428
rect 6392 54368 6456 54372
rect 7752 54428 7816 54432
rect 7752 54372 7756 54428
rect 7756 54372 7812 54428
rect 7812 54372 7816 54428
rect 7752 54368 7816 54372
rect 7832 54428 7896 54432
rect 7832 54372 7836 54428
rect 7836 54372 7892 54428
rect 7892 54372 7896 54428
rect 7832 54368 7896 54372
rect 7912 54428 7976 54432
rect 7912 54372 7916 54428
rect 7916 54372 7972 54428
rect 7972 54372 7976 54428
rect 7912 54368 7976 54372
rect 7992 54428 8056 54432
rect 7992 54372 7996 54428
rect 7996 54372 8052 54428
rect 8052 54372 8056 54428
rect 7992 54368 8056 54372
rect 9352 54428 9416 54432
rect 9352 54372 9356 54428
rect 9356 54372 9412 54428
rect 9412 54372 9416 54428
rect 9352 54368 9416 54372
rect 9432 54428 9496 54432
rect 9432 54372 9436 54428
rect 9436 54372 9492 54428
rect 9492 54372 9496 54428
rect 9432 54368 9496 54372
rect 9512 54428 9576 54432
rect 9512 54372 9516 54428
rect 9516 54372 9572 54428
rect 9572 54372 9576 54428
rect 9512 54368 9576 54372
rect 9592 54428 9656 54432
rect 9592 54372 9596 54428
rect 9596 54372 9652 54428
rect 9652 54372 9656 54428
rect 9592 54368 9656 54372
rect 3612 53884 3676 53888
rect 3612 53828 3616 53884
rect 3616 53828 3672 53884
rect 3672 53828 3676 53884
rect 3612 53824 3676 53828
rect 3692 53884 3756 53888
rect 3692 53828 3696 53884
rect 3696 53828 3752 53884
rect 3752 53828 3756 53884
rect 3692 53824 3756 53828
rect 3772 53884 3836 53888
rect 3772 53828 3776 53884
rect 3776 53828 3832 53884
rect 3832 53828 3836 53884
rect 3772 53824 3836 53828
rect 3852 53884 3916 53888
rect 3852 53828 3856 53884
rect 3856 53828 3912 53884
rect 3912 53828 3916 53884
rect 3852 53824 3916 53828
rect 5212 53884 5276 53888
rect 5212 53828 5216 53884
rect 5216 53828 5272 53884
rect 5272 53828 5276 53884
rect 5212 53824 5276 53828
rect 5292 53884 5356 53888
rect 5292 53828 5296 53884
rect 5296 53828 5352 53884
rect 5352 53828 5356 53884
rect 5292 53824 5356 53828
rect 5372 53884 5436 53888
rect 5372 53828 5376 53884
rect 5376 53828 5432 53884
rect 5432 53828 5436 53884
rect 5372 53824 5436 53828
rect 5452 53884 5516 53888
rect 5452 53828 5456 53884
rect 5456 53828 5512 53884
rect 5512 53828 5516 53884
rect 5452 53824 5516 53828
rect 6812 53884 6876 53888
rect 6812 53828 6816 53884
rect 6816 53828 6872 53884
rect 6872 53828 6876 53884
rect 6812 53824 6876 53828
rect 6892 53884 6956 53888
rect 6892 53828 6896 53884
rect 6896 53828 6952 53884
rect 6952 53828 6956 53884
rect 6892 53824 6956 53828
rect 6972 53884 7036 53888
rect 6972 53828 6976 53884
rect 6976 53828 7032 53884
rect 7032 53828 7036 53884
rect 6972 53824 7036 53828
rect 7052 53884 7116 53888
rect 7052 53828 7056 53884
rect 7056 53828 7112 53884
rect 7112 53828 7116 53884
rect 7052 53824 7116 53828
rect 8412 53884 8476 53888
rect 8412 53828 8416 53884
rect 8416 53828 8472 53884
rect 8472 53828 8476 53884
rect 8412 53824 8476 53828
rect 8492 53884 8556 53888
rect 8492 53828 8496 53884
rect 8496 53828 8552 53884
rect 8552 53828 8556 53884
rect 8492 53824 8556 53828
rect 8572 53884 8636 53888
rect 8572 53828 8576 53884
rect 8576 53828 8632 53884
rect 8632 53828 8636 53884
rect 8572 53824 8636 53828
rect 8652 53884 8716 53888
rect 8652 53828 8656 53884
rect 8656 53828 8712 53884
rect 8712 53828 8716 53884
rect 8652 53824 8716 53828
rect 2952 53340 3016 53344
rect 2952 53284 2956 53340
rect 2956 53284 3012 53340
rect 3012 53284 3016 53340
rect 2952 53280 3016 53284
rect 3032 53340 3096 53344
rect 3032 53284 3036 53340
rect 3036 53284 3092 53340
rect 3092 53284 3096 53340
rect 3032 53280 3096 53284
rect 3112 53340 3176 53344
rect 3112 53284 3116 53340
rect 3116 53284 3172 53340
rect 3172 53284 3176 53340
rect 3112 53280 3176 53284
rect 3192 53340 3256 53344
rect 3192 53284 3196 53340
rect 3196 53284 3252 53340
rect 3252 53284 3256 53340
rect 3192 53280 3256 53284
rect 4552 53340 4616 53344
rect 4552 53284 4556 53340
rect 4556 53284 4612 53340
rect 4612 53284 4616 53340
rect 4552 53280 4616 53284
rect 4632 53340 4696 53344
rect 4632 53284 4636 53340
rect 4636 53284 4692 53340
rect 4692 53284 4696 53340
rect 4632 53280 4696 53284
rect 4712 53340 4776 53344
rect 4712 53284 4716 53340
rect 4716 53284 4772 53340
rect 4772 53284 4776 53340
rect 4712 53280 4776 53284
rect 4792 53340 4856 53344
rect 4792 53284 4796 53340
rect 4796 53284 4852 53340
rect 4852 53284 4856 53340
rect 4792 53280 4856 53284
rect 6152 53340 6216 53344
rect 6152 53284 6156 53340
rect 6156 53284 6212 53340
rect 6212 53284 6216 53340
rect 6152 53280 6216 53284
rect 6232 53340 6296 53344
rect 6232 53284 6236 53340
rect 6236 53284 6292 53340
rect 6292 53284 6296 53340
rect 6232 53280 6296 53284
rect 6312 53340 6376 53344
rect 6312 53284 6316 53340
rect 6316 53284 6372 53340
rect 6372 53284 6376 53340
rect 6312 53280 6376 53284
rect 6392 53340 6456 53344
rect 6392 53284 6396 53340
rect 6396 53284 6452 53340
rect 6452 53284 6456 53340
rect 6392 53280 6456 53284
rect 7752 53340 7816 53344
rect 7752 53284 7756 53340
rect 7756 53284 7812 53340
rect 7812 53284 7816 53340
rect 7752 53280 7816 53284
rect 7832 53340 7896 53344
rect 7832 53284 7836 53340
rect 7836 53284 7892 53340
rect 7892 53284 7896 53340
rect 7832 53280 7896 53284
rect 7912 53340 7976 53344
rect 7912 53284 7916 53340
rect 7916 53284 7972 53340
rect 7972 53284 7976 53340
rect 7912 53280 7976 53284
rect 7992 53340 8056 53344
rect 7992 53284 7996 53340
rect 7996 53284 8052 53340
rect 8052 53284 8056 53340
rect 7992 53280 8056 53284
rect 9352 53340 9416 53344
rect 9352 53284 9356 53340
rect 9356 53284 9412 53340
rect 9412 53284 9416 53340
rect 9352 53280 9416 53284
rect 9432 53340 9496 53344
rect 9432 53284 9436 53340
rect 9436 53284 9492 53340
rect 9492 53284 9496 53340
rect 9432 53280 9496 53284
rect 9512 53340 9576 53344
rect 9512 53284 9516 53340
rect 9516 53284 9572 53340
rect 9572 53284 9576 53340
rect 9512 53280 9576 53284
rect 9592 53340 9656 53344
rect 9592 53284 9596 53340
rect 9596 53284 9652 53340
rect 9652 53284 9656 53340
rect 9592 53280 9656 53284
rect 3612 52796 3676 52800
rect 3612 52740 3616 52796
rect 3616 52740 3672 52796
rect 3672 52740 3676 52796
rect 3612 52736 3676 52740
rect 3692 52796 3756 52800
rect 3692 52740 3696 52796
rect 3696 52740 3752 52796
rect 3752 52740 3756 52796
rect 3692 52736 3756 52740
rect 3772 52796 3836 52800
rect 3772 52740 3776 52796
rect 3776 52740 3832 52796
rect 3832 52740 3836 52796
rect 3772 52736 3836 52740
rect 3852 52796 3916 52800
rect 3852 52740 3856 52796
rect 3856 52740 3912 52796
rect 3912 52740 3916 52796
rect 3852 52736 3916 52740
rect 5212 52796 5276 52800
rect 5212 52740 5216 52796
rect 5216 52740 5272 52796
rect 5272 52740 5276 52796
rect 5212 52736 5276 52740
rect 5292 52796 5356 52800
rect 5292 52740 5296 52796
rect 5296 52740 5352 52796
rect 5352 52740 5356 52796
rect 5292 52736 5356 52740
rect 5372 52796 5436 52800
rect 5372 52740 5376 52796
rect 5376 52740 5432 52796
rect 5432 52740 5436 52796
rect 5372 52736 5436 52740
rect 5452 52796 5516 52800
rect 5452 52740 5456 52796
rect 5456 52740 5512 52796
rect 5512 52740 5516 52796
rect 5452 52736 5516 52740
rect 6812 52796 6876 52800
rect 6812 52740 6816 52796
rect 6816 52740 6872 52796
rect 6872 52740 6876 52796
rect 6812 52736 6876 52740
rect 6892 52796 6956 52800
rect 6892 52740 6896 52796
rect 6896 52740 6952 52796
rect 6952 52740 6956 52796
rect 6892 52736 6956 52740
rect 6972 52796 7036 52800
rect 6972 52740 6976 52796
rect 6976 52740 7032 52796
rect 7032 52740 7036 52796
rect 6972 52736 7036 52740
rect 7052 52796 7116 52800
rect 7052 52740 7056 52796
rect 7056 52740 7112 52796
rect 7112 52740 7116 52796
rect 7052 52736 7116 52740
rect 8412 52796 8476 52800
rect 8412 52740 8416 52796
rect 8416 52740 8472 52796
rect 8472 52740 8476 52796
rect 8412 52736 8476 52740
rect 8492 52796 8556 52800
rect 8492 52740 8496 52796
rect 8496 52740 8552 52796
rect 8552 52740 8556 52796
rect 8492 52736 8556 52740
rect 8572 52796 8636 52800
rect 8572 52740 8576 52796
rect 8576 52740 8632 52796
rect 8632 52740 8636 52796
rect 8572 52736 8636 52740
rect 8652 52796 8716 52800
rect 8652 52740 8656 52796
rect 8656 52740 8712 52796
rect 8712 52740 8716 52796
rect 8652 52736 8716 52740
rect 2952 52252 3016 52256
rect 2952 52196 2956 52252
rect 2956 52196 3012 52252
rect 3012 52196 3016 52252
rect 2952 52192 3016 52196
rect 3032 52252 3096 52256
rect 3032 52196 3036 52252
rect 3036 52196 3092 52252
rect 3092 52196 3096 52252
rect 3032 52192 3096 52196
rect 3112 52252 3176 52256
rect 3112 52196 3116 52252
rect 3116 52196 3172 52252
rect 3172 52196 3176 52252
rect 3112 52192 3176 52196
rect 3192 52252 3256 52256
rect 3192 52196 3196 52252
rect 3196 52196 3252 52252
rect 3252 52196 3256 52252
rect 3192 52192 3256 52196
rect 4552 52252 4616 52256
rect 4552 52196 4556 52252
rect 4556 52196 4612 52252
rect 4612 52196 4616 52252
rect 4552 52192 4616 52196
rect 4632 52252 4696 52256
rect 4632 52196 4636 52252
rect 4636 52196 4692 52252
rect 4692 52196 4696 52252
rect 4632 52192 4696 52196
rect 4712 52252 4776 52256
rect 4712 52196 4716 52252
rect 4716 52196 4772 52252
rect 4772 52196 4776 52252
rect 4712 52192 4776 52196
rect 4792 52252 4856 52256
rect 4792 52196 4796 52252
rect 4796 52196 4852 52252
rect 4852 52196 4856 52252
rect 4792 52192 4856 52196
rect 6152 52252 6216 52256
rect 6152 52196 6156 52252
rect 6156 52196 6212 52252
rect 6212 52196 6216 52252
rect 6152 52192 6216 52196
rect 6232 52252 6296 52256
rect 6232 52196 6236 52252
rect 6236 52196 6292 52252
rect 6292 52196 6296 52252
rect 6232 52192 6296 52196
rect 6312 52252 6376 52256
rect 6312 52196 6316 52252
rect 6316 52196 6372 52252
rect 6372 52196 6376 52252
rect 6312 52192 6376 52196
rect 6392 52252 6456 52256
rect 6392 52196 6396 52252
rect 6396 52196 6452 52252
rect 6452 52196 6456 52252
rect 6392 52192 6456 52196
rect 7752 52252 7816 52256
rect 7752 52196 7756 52252
rect 7756 52196 7812 52252
rect 7812 52196 7816 52252
rect 7752 52192 7816 52196
rect 7832 52252 7896 52256
rect 7832 52196 7836 52252
rect 7836 52196 7892 52252
rect 7892 52196 7896 52252
rect 7832 52192 7896 52196
rect 7912 52252 7976 52256
rect 7912 52196 7916 52252
rect 7916 52196 7972 52252
rect 7972 52196 7976 52252
rect 7912 52192 7976 52196
rect 7992 52252 8056 52256
rect 7992 52196 7996 52252
rect 7996 52196 8052 52252
rect 8052 52196 8056 52252
rect 7992 52192 8056 52196
rect 9352 52252 9416 52256
rect 9352 52196 9356 52252
rect 9356 52196 9412 52252
rect 9412 52196 9416 52252
rect 9352 52192 9416 52196
rect 9432 52252 9496 52256
rect 9432 52196 9436 52252
rect 9436 52196 9492 52252
rect 9492 52196 9496 52252
rect 9432 52192 9496 52196
rect 9512 52252 9576 52256
rect 9512 52196 9516 52252
rect 9516 52196 9572 52252
rect 9572 52196 9576 52252
rect 9512 52192 9576 52196
rect 9592 52252 9656 52256
rect 9592 52196 9596 52252
rect 9596 52196 9652 52252
rect 9652 52196 9656 52252
rect 9592 52192 9656 52196
rect 3612 51708 3676 51712
rect 3612 51652 3616 51708
rect 3616 51652 3672 51708
rect 3672 51652 3676 51708
rect 3612 51648 3676 51652
rect 3692 51708 3756 51712
rect 3692 51652 3696 51708
rect 3696 51652 3752 51708
rect 3752 51652 3756 51708
rect 3692 51648 3756 51652
rect 3772 51708 3836 51712
rect 3772 51652 3776 51708
rect 3776 51652 3832 51708
rect 3832 51652 3836 51708
rect 3772 51648 3836 51652
rect 3852 51708 3916 51712
rect 3852 51652 3856 51708
rect 3856 51652 3912 51708
rect 3912 51652 3916 51708
rect 3852 51648 3916 51652
rect 5212 51708 5276 51712
rect 5212 51652 5216 51708
rect 5216 51652 5272 51708
rect 5272 51652 5276 51708
rect 5212 51648 5276 51652
rect 5292 51708 5356 51712
rect 5292 51652 5296 51708
rect 5296 51652 5352 51708
rect 5352 51652 5356 51708
rect 5292 51648 5356 51652
rect 5372 51708 5436 51712
rect 5372 51652 5376 51708
rect 5376 51652 5432 51708
rect 5432 51652 5436 51708
rect 5372 51648 5436 51652
rect 5452 51708 5516 51712
rect 5452 51652 5456 51708
rect 5456 51652 5512 51708
rect 5512 51652 5516 51708
rect 5452 51648 5516 51652
rect 6812 51708 6876 51712
rect 6812 51652 6816 51708
rect 6816 51652 6872 51708
rect 6872 51652 6876 51708
rect 6812 51648 6876 51652
rect 6892 51708 6956 51712
rect 6892 51652 6896 51708
rect 6896 51652 6952 51708
rect 6952 51652 6956 51708
rect 6892 51648 6956 51652
rect 6972 51708 7036 51712
rect 6972 51652 6976 51708
rect 6976 51652 7032 51708
rect 7032 51652 7036 51708
rect 6972 51648 7036 51652
rect 7052 51708 7116 51712
rect 7052 51652 7056 51708
rect 7056 51652 7112 51708
rect 7112 51652 7116 51708
rect 7052 51648 7116 51652
rect 8412 51708 8476 51712
rect 8412 51652 8416 51708
rect 8416 51652 8472 51708
rect 8472 51652 8476 51708
rect 8412 51648 8476 51652
rect 8492 51708 8556 51712
rect 8492 51652 8496 51708
rect 8496 51652 8552 51708
rect 8552 51652 8556 51708
rect 8492 51648 8556 51652
rect 8572 51708 8636 51712
rect 8572 51652 8576 51708
rect 8576 51652 8632 51708
rect 8632 51652 8636 51708
rect 8572 51648 8636 51652
rect 8652 51708 8716 51712
rect 8652 51652 8656 51708
rect 8656 51652 8712 51708
rect 8712 51652 8716 51708
rect 8652 51648 8716 51652
rect 2952 51164 3016 51168
rect 2952 51108 2956 51164
rect 2956 51108 3012 51164
rect 3012 51108 3016 51164
rect 2952 51104 3016 51108
rect 3032 51164 3096 51168
rect 3032 51108 3036 51164
rect 3036 51108 3092 51164
rect 3092 51108 3096 51164
rect 3032 51104 3096 51108
rect 3112 51164 3176 51168
rect 3112 51108 3116 51164
rect 3116 51108 3172 51164
rect 3172 51108 3176 51164
rect 3112 51104 3176 51108
rect 3192 51164 3256 51168
rect 3192 51108 3196 51164
rect 3196 51108 3252 51164
rect 3252 51108 3256 51164
rect 3192 51104 3256 51108
rect 4552 51164 4616 51168
rect 4552 51108 4556 51164
rect 4556 51108 4612 51164
rect 4612 51108 4616 51164
rect 4552 51104 4616 51108
rect 4632 51164 4696 51168
rect 4632 51108 4636 51164
rect 4636 51108 4692 51164
rect 4692 51108 4696 51164
rect 4632 51104 4696 51108
rect 4712 51164 4776 51168
rect 4712 51108 4716 51164
rect 4716 51108 4772 51164
rect 4772 51108 4776 51164
rect 4712 51104 4776 51108
rect 4792 51164 4856 51168
rect 4792 51108 4796 51164
rect 4796 51108 4852 51164
rect 4852 51108 4856 51164
rect 4792 51104 4856 51108
rect 6152 51164 6216 51168
rect 6152 51108 6156 51164
rect 6156 51108 6212 51164
rect 6212 51108 6216 51164
rect 6152 51104 6216 51108
rect 6232 51164 6296 51168
rect 6232 51108 6236 51164
rect 6236 51108 6292 51164
rect 6292 51108 6296 51164
rect 6232 51104 6296 51108
rect 6312 51164 6376 51168
rect 6312 51108 6316 51164
rect 6316 51108 6372 51164
rect 6372 51108 6376 51164
rect 6312 51104 6376 51108
rect 6392 51164 6456 51168
rect 6392 51108 6396 51164
rect 6396 51108 6452 51164
rect 6452 51108 6456 51164
rect 6392 51104 6456 51108
rect 7752 51164 7816 51168
rect 7752 51108 7756 51164
rect 7756 51108 7812 51164
rect 7812 51108 7816 51164
rect 7752 51104 7816 51108
rect 7832 51164 7896 51168
rect 7832 51108 7836 51164
rect 7836 51108 7892 51164
rect 7892 51108 7896 51164
rect 7832 51104 7896 51108
rect 7912 51164 7976 51168
rect 7912 51108 7916 51164
rect 7916 51108 7972 51164
rect 7972 51108 7976 51164
rect 7912 51104 7976 51108
rect 7992 51164 8056 51168
rect 7992 51108 7996 51164
rect 7996 51108 8052 51164
rect 8052 51108 8056 51164
rect 7992 51104 8056 51108
rect 9352 51164 9416 51168
rect 9352 51108 9356 51164
rect 9356 51108 9412 51164
rect 9412 51108 9416 51164
rect 9352 51104 9416 51108
rect 9432 51164 9496 51168
rect 9432 51108 9436 51164
rect 9436 51108 9492 51164
rect 9492 51108 9496 51164
rect 9432 51104 9496 51108
rect 9512 51164 9576 51168
rect 9512 51108 9516 51164
rect 9516 51108 9572 51164
rect 9572 51108 9576 51164
rect 9512 51104 9576 51108
rect 9592 51164 9656 51168
rect 9592 51108 9596 51164
rect 9596 51108 9652 51164
rect 9652 51108 9656 51164
rect 9592 51104 9656 51108
rect 3612 50620 3676 50624
rect 3612 50564 3616 50620
rect 3616 50564 3672 50620
rect 3672 50564 3676 50620
rect 3612 50560 3676 50564
rect 3692 50620 3756 50624
rect 3692 50564 3696 50620
rect 3696 50564 3752 50620
rect 3752 50564 3756 50620
rect 3692 50560 3756 50564
rect 3772 50620 3836 50624
rect 3772 50564 3776 50620
rect 3776 50564 3832 50620
rect 3832 50564 3836 50620
rect 3772 50560 3836 50564
rect 3852 50620 3916 50624
rect 3852 50564 3856 50620
rect 3856 50564 3912 50620
rect 3912 50564 3916 50620
rect 3852 50560 3916 50564
rect 5212 50620 5276 50624
rect 5212 50564 5216 50620
rect 5216 50564 5272 50620
rect 5272 50564 5276 50620
rect 5212 50560 5276 50564
rect 5292 50620 5356 50624
rect 5292 50564 5296 50620
rect 5296 50564 5352 50620
rect 5352 50564 5356 50620
rect 5292 50560 5356 50564
rect 5372 50620 5436 50624
rect 5372 50564 5376 50620
rect 5376 50564 5432 50620
rect 5432 50564 5436 50620
rect 5372 50560 5436 50564
rect 5452 50620 5516 50624
rect 5452 50564 5456 50620
rect 5456 50564 5512 50620
rect 5512 50564 5516 50620
rect 5452 50560 5516 50564
rect 6812 50620 6876 50624
rect 6812 50564 6816 50620
rect 6816 50564 6872 50620
rect 6872 50564 6876 50620
rect 6812 50560 6876 50564
rect 6892 50620 6956 50624
rect 6892 50564 6896 50620
rect 6896 50564 6952 50620
rect 6952 50564 6956 50620
rect 6892 50560 6956 50564
rect 6972 50620 7036 50624
rect 6972 50564 6976 50620
rect 6976 50564 7032 50620
rect 7032 50564 7036 50620
rect 6972 50560 7036 50564
rect 7052 50620 7116 50624
rect 7052 50564 7056 50620
rect 7056 50564 7112 50620
rect 7112 50564 7116 50620
rect 7052 50560 7116 50564
rect 8412 50620 8476 50624
rect 8412 50564 8416 50620
rect 8416 50564 8472 50620
rect 8472 50564 8476 50620
rect 8412 50560 8476 50564
rect 8492 50620 8556 50624
rect 8492 50564 8496 50620
rect 8496 50564 8552 50620
rect 8552 50564 8556 50620
rect 8492 50560 8556 50564
rect 8572 50620 8636 50624
rect 8572 50564 8576 50620
rect 8576 50564 8632 50620
rect 8632 50564 8636 50620
rect 8572 50560 8636 50564
rect 8652 50620 8716 50624
rect 8652 50564 8656 50620
rect 8656 50564 8712 50620
rect 8712 50564 8716 50620
rect 8652 50560 8716 50564
rect 2952 50076 3016 50080
rect 2952 50020 2956 50076
rect 2956 50020 3012 50076
rect 3012 50020 3016 50076
rect 2952 50016 3016 50020
rect 3032 50076 3096 50080
rect 3032 50020 3036 50076
rect 3036 50020 3092 50076
rect 3092 50020 3096 50076
rect 3032 50016 3096 50020
rect 3112 50076 3176 50080
rect 3112 50020 3116 50076
rect 3116 50020 3172 50076
rect 3172 50020 3176 50076
rect 3112 50016 3176 50020
rect 3192 50076 3256 50080
rect 3192 50020 3196 50076
rect 3196 50020 3252 50076
rect 3252 50020 3256 50076
rect 3192 50016 3256 50020
rect 4552 50076 4616 50080
rect 4552 50020 4556 50076
rect 4556 50020 4612 50076
rect 4612 50020 4616 50076
rect 4552 50016 4616 50020
rect 4632 50076 4696 50080
rect 4632 50020 4636 50076
rect 4636 50020 4692 50076
rect 4692 50020 4696 50076
rect 4632 50016 4696 50020
rect 4712 50076 4776 50080
rect 4712 50020 4716 50076
rect 4716 50020 4772 50076
rect 4772 50020 4776 50076
rect 4712 50016 4776 50020
rect 4792 50076 4856 50080
rect 4792 50020 4796 50076
rect 4796 50020 4852 50076
rect 4852 50020 4856 50076
rect 4792 50016 4856 50020
rect 6152 50076 6216 50080
rect 6152 50020 6156 50076
rect 6156 50020 6212 50076
rect 6212 50020 6216 50076
rect 6152 50016 6216 50020
rect 6232 50076 6296 50080
rect 6232 50020 6236 50076
rect 6236 50020 6292 50076
rect 6292 50020 6296 50076
rect 6232 50016 6296 50020
rect 6312 50076 6376 50080
rect 6312 50020 6316 50076
rect 6316 50020 6372 50076
rect 6372 50020 6376 50076
rect 6312 50016 6376 50020
rect 6392 50076 6456 50080
rect 6392 50020 6396 50076
rect 6396 50020 6452 50076
rect 6452 50020 6456 50076
rect 6392 50016 6456 50020
rect 7752 50076 7816 50080
rect 7752 50020 7756 50076
rect 7756 50020 7812 50076
rect 7812 50020 7816 50076
rect 7752 50016 7816 50020
rect 7832 50076 7896 50080
rect 7832 50020 7836 50076
rect 7836 50020 7892 50076
rect 7892 50020 7896 50076
rect 7832 50016 7896 50020
rect 7912 50076 7976 50080
rect 7912 50020 7916 50076
rect 7916 50020 7972 50076
rect 7972 50020 7976 50076
rect 7912 50016 7976 50020
rect 7992 50076 8056 50080
rect 7992 50020 7996 50076
rect 7996 50020 8052 50076
rect 8052 50020 8056 50076
rect 7992 50016 8056 50020
rect 3612 49532 3676 49536
rect 3612 49476 3616 49532
rect 3616 49476 3672 49532
rect 3672 49476 3676 49532
rect 3612 49472 3676 49476
rect 3692 49532 3756 49536
rect 3692 49476 3696 49532
rect 3696 49476 3752 49532
rect 3752 49476 3756 49532
rect 3692 49472 3756 49476
rect 3772 49532 3836 49536
rect 3772 49476 3776 49532
rect 3776 49476 3832 49532
rect 3832 49476 3836 49532
rect 3772 49472 3836 49476
rect 3852 49532 3916 49536
rect 3852 49476 3856 49532
rect 3856 49476 3912 49532
rect 3912 49476 3916 49532
rect 3852 49472 3916 49476
rect 5212 49532 5276 49536
rect 5212 49476 5216 49532
rect 5216 49476 5272 49532
rect 5272 49476 5276 49532
rect 5212 49472 5276 49476
rect 5292 49532 5356 49536
rect 5292 49476 5296 49532
rect 5296 49476 5352 49532
rect 5352 49476 5356 49532
rect 5292 49472 5356 49476
rect 5372 49532 5436 49536
rect 5372 49476 5376 49532
rect 5376 49476 5432 49532
rect 5432 49476 5436 49532
rect 5372 49472 5436 49476
rect 5452 49532 5516 49536
rect 5452 49476 5456 49532
rect 5456 49476 5512 49532
rect 5512 49476 5516 49532
rect 5452 49472 5516 49476
rect 6812 49532 6876 49536
rect 6812 49476 6816 49532
rect 6816 49476 6872 49532
rect 6872 49476 6876 49532
rect 6812 49472 6876 49476
rect 6892 49532 6956 49536
rect 6892 49476 6896 49532
rect 6896 49476 6952 49532
rect 6952 49476 6956 49532
rect 6892 49472 6956 49476
rect 6972 49532 7036 49536
rect 6972 49476 6976 49532
rect 6976 49476 7032 49532
rect 7032 49476 7036 49532
rect 6972 49472 7036 49476
rect 7052 49532 7116 49536
rect 7052 49476 7056 49532
rect 7056 49476 7112 49532
rect 7112 49476 7116 49532
rect 7052 49472 7116 49476
rect 8412 49532 8476 49536
rect 8412 49476 8416 49532
rect 8416 49476 8472 49532
rect 8472 49476 8476 49532
rect 8412 49472 8476 49476
rect 8492 49532 8556 49536
rect 8492 49476 8496 49532
rect 8496 49476 8552 49532
rect 8552 49476 8556 49532
rect 8492 49472 8556 49476
rect 8572 49532 8636 49536
rect 8572 49476 8576 49532
rect 8576 49476 8632 49532
rect 8632 49476 8636 49532
rect 8572 49472 8636 49476
rect 8652 49532 8716 49536
rect 8652 49476 8656 49532
rect 8656 49476 8712 49532
rect 8712 49476 8716 49532
rect 8652 49472 8716 49476
rect 2952 48988 3016 48992
rect 2952 48932 2956 48988
rect 2956 48932 3012 48988
rect 3012 48932 3016 48988
rect 2952 48928 3016 48932
rect 3032 48988 3096 48992
rect 3032 48932 3036 48988
rect 3036 48932 3092 48988
rect 3092 48932 3096 48988
rect 3032 48928 3096 48932
rect 3112 48988 3176 48992
rect 3112 48932 3116 48988
rect 3116 48932 3172 48988
rect 3172 48932 3176 48988
rect 3112 48928 3176 48932
rect 3192 48988 3256 48992
rect 3192 48932 3196 48988
rect 3196 48932 3252 48988
rect 3252 48932 3256 48988
rect 3192 48928 3256 48932
rect 4552 48988 4616 48992
rect 4552 48932 4556 48988
rect 4556 48932 4612 48988
rect 4612 48932 4616 48988
rect 4552 48928 4616 48932
rect 4632 48988 4696 48992
rect 4632 48932 4636 48988
rect 4636 48932 4692 48988
rect 4692 48932 4696 48988
rect 4632 48928 4696 48932
rect 4712 48988 4776 48992
rect 4712 48932 4716 48988
rect 4716 48932 4772 48988
rect 4772 48932 4776 48988
rect 4712 48928 4776 48932
rect 4792 48988 4856 48992
rect 4792 48932 4796 48988
rect 4796 48932 4852 48988
rect 4852 48932 4856 48988
rect 4792 48928 4856 48932
rect 6152 48988 6216 48992
rect 6152 48932 6156 48988
rect 6156 48932 6212 48988
rect 6212 48932 6216 48988
rect 6152 48928 6216 48932
rect 6232 48988 6296 48992
rect 6232 48932 6236 48988
rect 6236 48932 6292 48988
rect 6292 48932 6296 48988
rect 6232 48928 6296 48932
rect 6312 48988 6376 48992
rect 6312 48932 6316 48988
rect 6316 48932 6372 48988
rect 6372 48932 6376 48988
rect 6312 48928 6376 48932
rect 6392 48988 6456 48992
rect 6392 48932 6396 48988
rect 6396 48932 6452 48988
rect 6452 48932 6456 48988
rect 6392 48928 6456 48932
rect 7752 48988 7816 48992
rect 7752 48932 7756 48988
rect 7756 48932 7812 48988
rect 7812 48932 7816 48988
rect 7752 48928 7816 48932
rect 7832 48988 7896 48992
rect 7832 48932 7836 48988
rect 7836 48932 7892 48988
rect 7892 48932 7896 48988
rect 7832 48928 7896 48932
rect 7912 48988 7976 48992
rect 7912 48932 7916 48988
rect 7916 48932 7972 48988
rect 7972 48932 7976 48988
rect 7912 48928 7976 48932
rect 7992 48988 8056 48992
rect 7992 48932 7996 48988
rect 7996 48932 8052 48988
rect 8052 48932 8056 48988
rect 7992 48928 8056 48932
rect 9352 50076 9416 50080
rect 9352 50020 9356 50076
rect 9356 50020 9412 50076
rect 9412 50020 9416 50076
rect 9352 50016 9416 50020
rect 9432 50076 9496 50080
rect 9432 50020 9436 50076
rect 9436 50020 9492 50076
rect 9492 50020 9496 50076
rect 9432 50016 9496 50020
rect 9512 50076 9576 50080
rect 9512 50020 9516 50076
rect 9516 50020 9572 50076
rect 9572 50020 9576 50076
rect 9512 50016 9576 50020
rect 9592 50076 9656 50080
rect 9592 50020 9596 50076
rect 9596 50020 9652 50076
rect 9652 50020 9656 50076
rect 9592 50016 9656 50020
rect 9352 48988 9416 48992
rect 9352 48932 9356 48988
rect 9356 48932 9412 48988
rect 9412 48932 9416 48988
rect 9352 48928 9416 48932
rect 9432 48988 9496 48992
rect 9432 48932 9436 48988
rect 9436 48932 9492 48988
rect 9492 48932 9496 48988
rect 9432 48928 9496 48932
rect 9512 48988 9576 48992
rect 9512 48932 9516 48988
rect 9516 48932 9572 48988
rect 9572 48932 9576 48988
rect 9512 48928 9576 48932
rect 9592 48988 9656 48992
rect 9592 48932 9596 48988
rect 9596 48932 9652 48988
rect 9652 48932 9656 48988
rect 9592 48928 9656 48932
rect 3612 48444 3676 48448
rect 3612 48388 3616 48444
rect 3616 48388 3672 48444
rect 3672 48388 3676 48444
rect 3612 48384 3676 48388
rect 3692 48444 3756 48448
rect 3692 48388 3696 48444
rect 3696 48388 3752 48444
rect 3752 48388 3756 48444
rect 3692 48384 3756 48388
rect 3772 48444 3836 48448
rect 3772 48388 3776 48444
rect 3776 48388 3832 48444
rect 3832 48388 3836 48444
rect 3772 48384 3836 48388
rect 3852 48444 3916 48448
rect 3852 48388 3856 48444
rect 3856 48388 3912 48444
rect 3912 48388 3916 48444
rect 3852 48384 3916 48388
rect 5212 48444 5276 48448
rect 5212 48388 5216 48444
rect 5216 48388 5272 48444
rect 5272 48388 5276 48444
rect 5212 48384 5276 48388
rect 5292 48444 5356 48448
rect 5292 48388 5296 48444
rect 5296 48388 5352 48444
rect 5352 48388 5356 48444
rect 5292 48384 5356 48388
rect 5372 48444 5436 48448
rect 5372 48388 5376 48444
rect 5376 48388 5432 48444
rect 5432 48388 5436 48444
rect 5372 48384 5436 48388
rect 5452 48444 5516 48448
rect 5452 48388 5456 48444
rect 5456 48388 5512 48444
rect 5512 48388 5516 48444
rect 5452 48384 5516 48388
rect 6812 48444 6876 48448
rect 6812 48388 6816 48444
rect 6816 48388 6872 48444
rect 6872 48388 6876 48444
rect 6812 48384 6876 48388
rect 6892 48444 6956 48448
rect 6892 48388 6896 48444
rect 6896 48388 6952 48444
rect 6952 48388 6956 48444
rect 6892 48384 6956 48388
rect 6972 48444 7036 48448
rect 6972 48388 6976 48444
rect 6976 48388 7032 48444
rect 7032 48388 7036 48444
rect 6972 48384 7036 48388
rect 7052 48444 7116 48448
rect 7052 48388 7056 48444
rect 7056 48388 7112 48444
rect 7112 48388 7116 48444
rect 7052 48384 7116 48388
rect 8412 48444 8476 48448
rect 8412 48388 8416 48444
rect 8416 48388 8472 48444
rect 8472 48388 8476 48444
rect 8412 48384 8476 48388
rect 8492 48444 8556 48448
rect 8492 48388 8496 48444
rect 8496 48388 8552 48444
rect 8552 48388 8556 48444
rect 8492 48384 8556 48388
rect 8572 48444 8636 48448
rect 8572 48388 8576 48444
rect 8576 48388 8632 48444
rect 8632 48388 8636 48444
rect 8572 48384 8636 48388
rect 8652 48444 8716 48448
rect 8652 48388 8656 48444
rect 8656 48388 8712 48444
rect 8712 48388 8716 48444
rect 8652 48384 8716 48388
rect 2952 47900 3016 47904
rect 2952 47844 2956 47900
rect 2956 47844 3012 47900
rect 3012 47844 3016 47900
rect 2952 47840 3016 47844
rect 3032 47900 3096 47904
rect 3032 47844 3036 47900
rect 3036 47844 3092 47900
rect 3092 47844 3096 47900
rect 3032 47840 3096 47844
rect 3112 47900 3176 47904
rect 3112 47844 3116 47900
rect 3116 47844 3172 47900
rect 3172 47844 3176 47900
rect 3112 47840 3176 47844
rect 3192 47900 3256 47904
rect 3192 47844 3196 47900
rect 3196 47844 3252 47900
rect 3252 47844 3256 47900
rect 3192 47840 3256 47844
rect 4552 47900 4616 47904
rect 4552 47844 4556 47900
rect 4556 47844 4612 47900
rect 4612 47844 4616 47900
rect 4552 47840 4616 47844
rect 4632 47900 4696 47904
rect 4632 47844 4636 47900
rect 4636 47844 4692 47900
rect 4692 47844 4696 47900
rect 4632 47840 4696 47844
rect 4712 47900 4776 47904
rect 4712 47844 4716 47900
rect 4716 47844 4772 47900
rect 4772 47844 4776 47900
rect 4712 47840 4776 47844
rect 4792 47900 4856 47904
rect 4792 47844 4796 47900
rect 4796 47844 4852 47900
rect 4852 47844 4856 47900
rect 4792 47840 4856 47844
rect 6152 47900 6216 47904
rect 6152 47844 6156 47900
rect 6156 47844 6212 47900
rect 6212 47844 6216 47900
rect 6152 47840 6216 47844
rect 6232 47900 6296 47904
rect 6232 47844 6236 47900
rect 6236 47844 6292 47900
rect 6292 47844 6296 47900
rect 6232 47840 6296 47844
rect 6312 47900 6376 47904
rect 6312 47844 6316 47900
rect 6316 47844 6372 47900
rect 6372 47844 6376 47900
rect 6312 47840 6376 47844
rect 6392 47900 6456 47904
rect 6392 47844 6396 47900
rect 6396 47844 6452 47900
rect 6452 47844 6456 47900
rect 6392 47840 6456 47844
rect 7752 47900 7816 47904
rect 7752 47844 7756 47900
rect 7756 47844 7812 47900
rect 7812 47844 7816 47900
rect 7752 47840 7816 47844
rect 7832 47900 7896 47904
rect 7832 47844 7836 47900
rect 7836 47844 7892 47900
rect 7892 47844 7896 47900
rect 7832 47840 7896 47844
rect 7912 47900 7976 47904
rect 7912 47844 7916 47900
rect 7916 47844 7972 47900
rect 7972 47844 7976 47900
rect 7912 47840 7976 47844
rect 7992 47900 8056 47904
rect 7992 47844 7996 47900
rect 7996 47844 8052 47900
rect 8052 47844 8056 47900
rect 7992 47840 8056 47844
rect 3612 47356 3676 47360
rect 3612 47300 3616 47356
rect 3616 47300 3672 47356
rect 3672 47300 3676 47356
rect 3612 47296 3676 47300
rect 3692 47356 3756 47360
rect 3692 47300 3696 47356
rect 3696 47300 3752 47356
rect 3752 47300 3756 47356
rect 3692 47296 3756 47300
rect 3772 47356 3836 47360
rect 3772 47300 3776 47356
rect 3776 47300 3832 47356
rect 3832 47300 3836 47356
rect 3772 47296 3836 47300
rect 3852 47356 3916 47360
rect 3852 47300 3856 47356
rect 3856 47300 3912 47356
rect 3912 47300 3916 47356
rect 3852 47296 3916 47300
rect 5212 47356 5276 47360
rect 5212 47300 5216 47356
rect 5216 47300 5272 47356
rect 5272 47300 5276 47356
rect 5212 47296 5276 47300
rect 5292 47356 5356 47360
rect 5292 47300 5296 47356
rect 5296 47300 5352 47356
rect 5352 47300 5356 47356
rect 5292 47296 5356 47300
rect 5372 47356 5436 47360
rect 5372 47300 5376 47356
rect 5376 47300 5432 47356
rect 5432 47300 5436 47356
rect 5372 47296 5436 47300
rect 5452 47356 5516 47360
rect 5452 47300 5456 47356
rect 5456 47300 5512 47356
rect 5512 47300 5516 47356
rect 5452 47296 5516 47300
rect 6812 47356 6876 47360
rect 6812 47300 6816 47356
rect 6816 47300 6872 47356
rect 6872 47300 6876 47356
rect 6812 47296 6876 47300
rect 6892 47356 6956 47360
rect 6892 47300 6896 47356
rect 6896 47300 6952 47356
rect 6952 47300 6956 47356
rect 6892 47296 6956 47300
rect 6972 47356 7036 47360
rect 6972 47300 6976 47356
rect 6976 47300 7032 47356
rect 7032 47300 7036 47356
rect 6972 47296 7036 47300
rect 7052 47356 7116 47360
rect 7052 47300 7056 47356
rect 7056 47300 7112 47356
rect 7112 47300 7116 47356
rect 7052 47296 7116 47300
rect 8412 47356 8476 47360
rect 8412 47300 8416 47356
rect 8416 47300 8472 47356
rect 8472 47300 8476 47356
rect 8412 47296 8476 47300
rect 8492 47356 8556 47360
rect 8492 47300 8496 47356
rect 8496 47300 8552 47356
rect 8552 47300 8556 47356
rect 8492 47296 8556 47300
rect 8572 47356 8636 47360
rect 8572 47300 8576 47356
rect 8576 47300 8632 47356
rect 8632 47300 8636 47356
rect 8572 47296 8636 47300
rect 8652 47356 8716 47360
rect 8652 47300 8656 47356
rect 8656 47300 8712 47356
rect 8712 47300 8716 47356
rect 8652 47296 8716 47300
rect 2952 46812 3016 46816
rect 2952 46756 2956 46812
rect 2956 46756 3012 46812
rect 3012 46756 3016 46812
rect 2952 46752 3016 46756
rect 3032 46812 3096 46816
rect 3032 46756 3036 46812
rect 3036 46756 3092 46812
rect 3092 46756 3096 46812
rect 3032 46752 3096 46756
rect 3112 46812 3176 46816
rect 3112 46756 3116 46812
rect 3116 46756 3172 46812
rect 3172 46756 3176 46812
rect 3112 46752 3176 46756
rect 3192 46812 3256 46816
rect 3192 46756 3196 46812
rect 3196 46756 3252 46812
rect 3252 46756 3256 46812
rect 3192 46752 3256 46756
rect 4552 46812 4616 46816
rect 4552 46756 4556 46812
rect 4556 46756 4612 46812
rect 4612 46756 4616 46812
rect 4552 46752 4616 46756
rect 4632 46812 4696 46816
rect 4632 46756 4636 46812
rect 4636 46756 4692 46812
rect 4692 46756 4696 46812
rect 4632 46752 4696 46756
rect 4712 46812 4776 46816
rect 4712 46756 4716 46812
rect 4716 46756 4772 46812
rect 4772 46756 4776 46812
rect 4712 46752 4776 46756
rect 4792 46812 4856 46816
rect 4792 46756 4796 46812
rect 4796 46756 4852 46812
rect 4852 46756 4856 46812
rect 4792 46752 4856 46756
rect 6152 46812 6216 46816
rect 6152 46756 6156 46812
rect 6156 46756 6212 46812
rect 6212 46756 6216 46812
rect 6152 46752 6216 46756
rect 6232 46812 6296 46816
rect 6232 46756 6236 46812
rect 6236 46756 6292 46812
rect 6292 46756 6296 46812
rect 6232 46752 6296 46756
rect 6312 46812 6376 46816
rect 6312 46756 6316 46812
rect 6316 46756 6372 46812
rect 6372 46756 6376 46812
rect 6312 46752 6376 46756
rect 6392 46812 6456 46816
rect 6392 46756 6396 46812
rect 6396 46756 6452 46812
rect 6452 46756 6456 46812
rect 6392 46752 6456 46756
rect 7752 46812 7816 46816
rect 7752 46756 7756 46812
rect 7756 46756 7812 46812
rect 7812 46756 7816 46812
rect 7752 46752 7816 46756
rect 7832 46812 7896 46816
rect 7832 46756 7836 46812
rect 7836 46756 7892 46812
rect 7892 46756 7896 46812
rect 7832 46752 7896 46756
rect 7912 46812 7976 46816
rect 7912 46756 7916 46812
rect 7916 46756 7972 46812
rect 7972 46756 7976 46812
rect 7912 46752 7976 46756
rect 7992 46812 8056 46816
rect 7992 46756 7996 46812
rect 7996 46756 8052 46812
rect 8052 46756 8056 46812
rect 7992 46752 8056 46756
rect 9352 47900 9416 47904
rect 9352 47844 9356 47900
rect 9356 47844 9412 47900
rect 9412 47844 9416 47900
rect 9352 47840 9416 47844
rect 9432 47900 9496 47904
rect 9432 47844 9436 47900
rect 9436 47844 9492 47900
rect 9492 47844 9496 47900
rect 9432 47840 9496 47844
rect 9512 47900 9576 47904
rect 9512 47844 9516 47900
rect 9516 47844 9572 47900
rect 9572 47844 9576 47900
rect 9512 47840 9576 47844
rect 9592 47900 9656 47904
rect 9592 47844 9596 47900
rect 9596 47844 9652 47900
rect 9652 47844 9656 47900
rect 9592 47840 9656 47844
rect 9352 46812 9416 46816
rect 9352 46756 9356 46812
rect 9356 46756 9412 46812
rect 9412 46756 9416 46812
rect 9352 46752 9416 46756
rect 9432 46812 9496 46816
rect 9432 46756 9436 46812
rect 9436 46756 9492 46812
rect 9492 46756 9496 46812
rect 9432 46752 9496 46756
rect 9512 46812 9576 46816
rect 9512 46756 9516 46812
rect 9516 46756 9572 46812
rect 9572 46756 9576 46812
rect 9512 46752 9576 46756
rect 9592 46812 9656 46816
rect 9592 46756 9596 46812
rect 9596 46756 9652 46812
rect 9652 46756 9656 46812
rect 9592 46752 9656 46756
rect 3612 46268 3676 46272
rect 3612 46212 3616 46268
rect 3616 46212 3672 46268
rect 3672 46212 3676 46268
rect 3612 46208 3676 46212
rect 3692 46268 3756 46272
rect 3692 46212 3696 46268
rect 3696 46212 3752 46268
rect 3752 46212 3756 46268
rect 3692 46208 3756 46212
rect 3772 46268 3836 46272
rect 3772 46212 3776 46268
rect 3776 46212 3832 46268
rect 3832 46212 3836 46268
rect 3772 46208 3836 46212
rect 3852 46268 3916 46272
rect 3852 46212 3856 46268
rect 3856 46212 3912 46268
rect 3912 46212 3916 46268
rect 3852 46208 3916 46212
rect 5212 46268 5276 46272
rect 5212 46212 5216 46268
rect 5216 46212 5272 46268
rect 5272 46212 5276 46268
rect 5212 46208 5276 46212
rect 5292 46268 5356 46272
rect 5292 46212 5296 46268
rect 5296 46212 5352 46268
rect 5352 46212 5356 46268
rect 5292 46208 5356 46212
rect 5372 46268 5436 46272
rect 5372 46212 5376 46268
rect 5376 46212 5432 46268
rect 5432 46212 5436 46268
rect 5372 46208 5436 46212
rect 5452 46268 5516 46272
rect 5452 46212 5456 46268
rect 5456 46212 5512 46268
rect 5512 46212 5516 46268
rect 5452 46208 5516 46212
rect 6812 46268 6876 46272
rect 6812 46212 6816 46268
rect 6816 46212 6872 46268
rect 6872 46212 6876 46268
rect 6812 46208 6876 46212
rect 6892 46268 6956 46272
rect 6892 46212 6896 46268
rect 6896 46212 6952 46268
rect 6952 46212 6956 46268
rect 6892 46208 6956 46212
rect 6972 46268 7036 46272
rect 6972 46212 6976 46268
rect 6976 46212 7032 46268
rect 7032 46212 7036 46268
rect 6972 46208 7036 46212
rect 7052 46268 7116 46272
rect 7052 46212 7056 46268
rect 7056 46212 7112 46268
rect 7112 46212 7116 46268
rect 7052 46208 7116 46212
rect 2952 45724 3016 45728
rect 2952 45668 2956 45724
rect 2956 45668 3012 45724
rect 3012 45668 3016 45724
rect 2952 45664 3016 45668
rect 3032 45724 3096 45728
rect 3032 45668 3036 45724
rect 3036 45668 3092 45724
rect 3092 45668 3096 45724
rect 3032 45664 3096 45668
rect 3112 45724 3176 45728
rect 3112 45668 3116 45724
rect 3116 45668 3172 45724
rect 3172 45668 3176 45724
rect 3112 45664 3176 45668
rect 3192 45724 3256 45728
rect 3192 45668 3196 45724
rect 3196 45668 3252 45724
rect 3252 45668 3256 45724
rect 3192 45664 3256 45668
rect 4552 45724 4616 45728
rect 4552 45668 4556 45724
rect 4556 45668 4612 45724
rect 4612 45668 4616 45724
rect 4552 45664 4616 45668
rect 4632 45724 4696 45728
rect 4632 45668 4636 45724
rect 4636 45668 4692 45724
rect 4692 45668 4696 45724
rect 4632 45664 4696 45668
rect 4712 45724 4776 45728
rect 4712 45668 4716 45724
rect 4716 45668 4772 45724
rect 4772 45668 4776 45724
rect 4712 45664 4776 45668
rect 4792 45724 4856 45728
rect 4792 45668 4796 45724
rect 4796 45668 4852 45724
rect 4852 45668 4856 45724
rect 4792 45664 4856 45668
rect 6152 45724 6216 45728
rect 6152 45668 6156 45724
rect 6156 45668 6212 45724
rect 6212 45668 6216 45724
rect 6152 45664 6216 45668
rect 6232 45724 6296 45728
rect 6232 45668 6236 45724
rect 6236 45668 6292 45724
rect 6292 45668 6296 45724
rect 6232 45664 6296 45668
rect 6312 45724 6376 45728
rect 6312 45668 6316 45724
rect 6316 45668 6372 45724
rect 6372 45668 6376 45724
rect 6312 45664 6376 45668
rect 6392 45724 6456 45728
rect 6392 45668 6396 45724
rect 6396 45668 6452 45724
rect 6452 45668 6456 45724
rect 6392 45664 6456 45668
rect 7752 45724 7816 45728
rect 7752 45668 7756 45724
rect 7756 45668 7812 45724
rect 7812 45668 7816 45724
rect 7752 45664 7816 45668
rect 7832 45724 7896 45728
rect 7832 45668 7836 45724
rect 7836 45668 7892 45724
rect 7892 45668 7896 45724
rect 7832 45664 7896 45668
rect 7912 45724 7976 45728
rect 7912 45668 7916 45724
rect 7916 45668 7972 45724
rect 7972 45668 7976 45724
rect 7912 45664 7976 45668
rect 7992 45724 8056 45728
rect 7992 45668 7996 45724
rect 7996 45668 8052 45724
rect 8052 45668 8056 45724
rect 7992 45664 8056 45668
rect 8412 46268 8476 46272
rect 8412 46212 8416 46268
rect 8416 46212 8472 46268
rect 8472 46212 8476 46268
rect 8412 46208 8476 46212
rect 8492 46268 8556 46272
rect 8492 46212 8496 46268
rect 8496 46212 8552 46268
rect 8552 46212 8556 46268
rect 8492 46208 8556 46212
rect 8572 46268 8636 46272
rect 8572 46212 8576 46268
rect 8576 46212 8632 46268
rect 8632 46212 8636 46268
rect 8572 46208 8636 46212
rect 8652 46268 8716 46272
rect 8652 46212 8656 46268
rect 8656 46212 8712 46268
rect 8712 46212 8716 46268
rect 8652 46208 8716 46212
rect 9352 45724 9416 45728
rect 9352 45668 9356 45724
rect 9356 45668 9412 45724
rect 9412 45668 9416 45724
rect 9352 45664 9416 45668
rect 9432 45724 9496 45728
rect 9432 45668 9436 45724
rect 9436 45668 9492 45724
rect 9492 45668 9496 45724
rect 9432 45664 9496 45668
rect 9512 45724 9576 45728
rect 9512 45668 9516 45724
rect 9516 45668 9572 45724
rect 9572 45668 9576 45724
rect 9512 45664 9576 45668
rect 9592 45724 9656 45728
rect 9592 45668 9596 45724
rect 9596 45668 9652 45724
rect 9652 45668 9656 45724
rect 9592 45664 9656 45668
rect 3612 45180 3676 45184
rect 3612 45124 3616 45180
rect 3616 45124 3672 45180
rect 3672 45124 3676 45180
rect 3612 45120 3676 45124
rect 3692 45180 3756 45184
rect 3692 45124 3696 45180
rect 3696 45124 3752 45180
rect 3752 45124 3756 45180
rect 3692 45120 3756 45124
rect 3772 45180 3836 45184
rect 3772 45124 3776 45180
rect 3776 45124 3832 45180
rect 3832 45124 3836 45180
rect 3772 45120 3836 45124
rect 3852 45180 3916 45184
rect 3852 45124 3856 45180
rect 3856 45124 3912 45180
rect 3912 45124 3916 45180
rect 3852 45120 3916 45124
rect 5212 45180 5276 45184
rect 5212 45124 5216 45180
rect 5216 45124 5272 45180
rect 5272 45124 5276 45180
rect 5212 45120 5276 45124
rect 5292 45180 5356 45184
rect 5292 45124 5296 45180
rect 5296 45124 5352 45180
rect 5352 45124 5356 45180
rect 5292 45120 5356 45124
rect 5372 45180 5436 45184
rect 5372 45124 5376 45180
rect 5376 45124 5432 45180
rect 5432 45124 5436 45180
rect 5372 45120 5436 45124
rect 5452 45180 5516 45184
rect 5452 45124 5456 45180
rect 5456 45124 5512 45180
rect 5512 45124 5516 45180
rect 5452 45120 5516 45124
rect 6812 45180 6876 45184
rect 6812 45124 6816 45180
rect 6816 45124 6872 45180
rect 6872 45124 6876 45180
rect 6812 45120 6876 45124
rect 6892 45180 6956 45184
rect 6892 45124 6896 45180
rect 6896 45124 6952 45180
rect 6952 45124 6956 45180
rect 6892 45120 6956 45124
rect 6972 45180 7036 45184
rect 6972 45124 6976 45180
rect 6976 45124 7032 45180
rect 7032 45124 7036 45180
rect 6972 45120 7036 45124
rect 7052 45180 7116 45184
rect 7052 45124 7056 45180
rect 7056 45124 7112 45180
rect 7112 45124 7116 45180
rect 7052 45120 7116 45124
rect 8412 45180 8476 45184
rect 8412 45124 8416 45180
rect 8416 45124 8472 45180
rect 8472 45124 8476 45180
rect 8412 45120 8476 45124
rect 8492 45180 8556 45184
rect 8492 45124 8496 45180
rect 8496 45124 8552 45180
rect 8552 45124 8556 45180
rect 8492 45120 8556 45124
rect 8572 45180 8636 45184
rect 8572 45124 8576 45180
rect 8576 45124 8632 45180
rect 8632 45124 8636 45180
rect 8572 45120 8636 45124
rect 8652 45180 8716 45184
rect 8652 45124 8656 45180
rect 8656 45124 8712 45180
rect 8712 45124 8716 45180
rect 8652 45120 8716 45124
rect 2952 44636 3016 44640
rect 2952 44580 2956 44636
rect 2956 44580 3012 44636
rect 3012 44580 3016 44636
rect 2952 44576 3016 44580
rect 3032 44636 3096 44640
rect 3032 44580 3036 44636
rect 3036 44580 3092 44636
rect 3092 44580 3096 44636
rect 3032 44576 3096 44580
rect 3112 44636 3176 44640
rect 3112 44580 3116 44636
rect 3116 44580 3172 44636
rect 3172 44580 3176 44636
rect 3112 44576 3176 44580
rect 3192 44636 3256 44640
rect 3192 44580 3196 44636
rect 3196 44580 3252 44636
rect 3252 44580 3256 44636
rect 3192 44576 3256 44580
rect 4552 44636 4616 44640
rect 4552 44580 4556 44636
rect 4556 44580 4612 44636
rect 4612 44580 4616 44636
rect 4552 44576 4616 44580
rect 4632 44636 4696 44640
rect 4632 44580 4636 44636
rect 4636 44580 4692 44636
rect 4692 44580 4696 44636
rect 4632 44576 4696 44580
rect 4712 44636 4776 44640
rect 4712 44580 4716 44636
rect 4716 44580 4772 44636
rect 4772 44580 4776 44636
rect 4712 44576 4776 44580
rect 4792 44636 4856 44640
rect 4792 44580 4796 44636
rect 4796 44580 4852 44636
rect 4852 44580 4856 44636
rect 4792 44576 4856 44580
rect 6152 44636 6216 44640
rect 6152 44580 6156 44636
rect 6156 44580 6212 44636
rect 6212 44580 6216 44636
rect 6152 44576 6216 44580
rect 6232 44636 6296 44640
rect 6232 44580 6236 44636
rect 6236 44580 6292 44636
rect 6292 44580 6296 44636
rect 6232 44576 6296 44580
rect 6312 44636 6376 44640
rect 6312 44580 6316 44636
rect 6316 44580 6372 44636
rect 6372 44580 6376 44636
rect 6312 44576 6376 44580
rect 6392 44636 6456 44640
rect 6392 44580 6396 44636
rect 6396 44580 6452 44636
rect 6452 44580 6456 44636
rect 6392 44576 6456 44580
rect 7752 44636 7816 44640
rect 7752 44580 7756 44636
rect 7756 44580 7812 44636
rect 7812 44580 7816 44636
rect 7752 44576 7816 44580
rect 7832 44636 7896 44640
rect 7832 44580 7836 44636
rect 7836 44580 7892 44636
rect 7892 44580 7896 44636
rect 7832 44576 7896 44580
rect 7912 44636 7976 44640
rect 7912 44580 7916 44636
rect 7916 44580 7972 44636
rect 7972 44580 7976 44636
rect 7912 44576 7976 44580
rect 7992 44636 8056 44640
rect 7992 44580 7996 44636
rect 7996 44580 8052 44636
rect 8052 44580 8056 44636
rect 7992 44576 8056 44580
rect 9352 44636 9416 44640
rect 9352 44580 9356 44636
rect 9356 44580 9412 44636
rect 9412 44580 9416 44636
rect 9352 44576 9416 44580
rect 9432 44636 9496 44640
rect 9432 44580 9436 44636
rect 9436 44580 9492 44636
rect 9492 44580 9496 44636
rect 9432 44576 9496 44580
rect 9512 44636 9576 44640
rect 9512 44580 9516 44636
rect 9516 44580 9572 44636
rect 9572 44580 9576 44636
rect 9512 44576 9576 44580
rect 9592 44636 9656 44640
rect 9592 44580 9596 44636
rect 9596 44580 9652 44636
rect 9652 44580 9656 44636
rect 9592 44576 9656 44580
rect 3612 44092 3676 44096
rect 3612 44036 3616 44092
rect 3616 44036 3672 44092
rect 3672 44036 3676 44092
rect 3612 44032 3676 44036
rect 3692 44092 3756 44096
rect 3692 44036 3696 44092
rect 3696 44036 3752 44092
rect 3752 44036 3756 44092
rect 3692 44032 3756 44036
rect 3772 44092 3836 44096
rect 3772 44036 3776 44092
rect 3776 44036 3832 44092
rect 3832 44036 3836 44092
rect 3772 44032 3836 44036
rect 3852 44092 3916 44096
rect 3852 44036 3856 44092
rect 3856 44036 3912 44092
rect 3912 44036 3916 44092
rect 3852 44032 3916 44036
rect 5212 44092 5276 44096
rect 5212 44036 5216 44092
rect 5216 44036 5272 44092
rect 5272 44036 5276 44092
rect 5212 44032 5276 44036
rect 5292 44092 5356 44096
rect 5292 44036 5296 44092
rect 5296 44036 5352 44092
rect 5352 44036 5356 44092
rect 5292 44032 5356 44036
rect 5372 44092 5436 44096
rect 5372 44036 5376 44092
rect 5376 44036 5432 44092
rect 5432 44036 5436 44092
rect 5372 44032 5436 44036
rect 5452 44092 5516 44096
rect 5452 44036 5456 44092
rect 5456 44036 5512 44092
rect 5512 44036 5516 44092
rect 5452 44032 5516 44036
rect 6812 44092 6876 44096
rect 6812 44036 6816 44092
rect 6816 44036 6872 44092
rect 6872 44036 6876 44092
rect 6812 44032 6876 44036
rect 6892 44092 6956 44096
rect 6892 44036 6896 44092
rect 6896 44036 6952 44092
rect 6952 44036 6956 44092
rect 6892 44032 6956 44036
rect 6972 44092 7036 44096
rect 6972 44036 6976 44092
rect 6976 44036 7032 44092
rect 7032 44036 7036 44092
rect 6972 44032 7036 44036
rect 7052 44092 7116 44096
rect 7052 44036 7056 44092
rect 7056 44036 7112 44092
rect 7112 44036 7116 44092
rect 7052 44032 7116 44036
rect 8412 44092 8476 44096
rect 8412 44036 8416 44092
rect 8416 44036 8472 44092
rect 8472 44036 8476 44092
rect 8412 44032 8476 44036
rect 8492 44092 8556 44096
rect 8492 44036 8496 44092
rect 8496 44036 8552 44092
rect 8552 44036 8556 44092
rect 8492 44032 8556 44036
rect 8572 44092 8636 44096
rect 8572 44036 8576 44092
rect 8576 44036 8632 44092
rect 8632 44036 8636 44092
rect 8572 44032 8636 44036
rect 8652 44092 8716 44096
rect 8652 44036 8656 44092
rect 8656 44036 8712 44092
rect 8712 44036 8716 44092
rect 8652 44032 8716 44036
rect 2952 43548 3016 43552
rect 2952 43492 2956 43548
rect 2956 43492 3012 43548
rect 3012 43492 3016 43548
rect 2952 43488 3016 43492
rect 3032 43548 3096 43552
rect 3032 43492 3036 43548
rect 3036 43492 3092 43548
rect 3092 43492 3096 43548
rect 3032 43488 3096 43492
rect 3112 43548 3176 43552
rect 3112 43492 3116 43548
rect 3116 43492 3172 43548
rect 3172 43492 3176 43548
rect 3112 43488 3176 43492
rect 3192 43548 3256 43552
rect 3192 43492 3196 43548
rect 3196 43492 3252 43548
rect 3252 43492 3256 43548
rect 3192 43488 3256 43492
rect 4552 43548 4616 43552
rect 4552 43492 4556 43548
rect 4556 43492 4612 43548
rect 4612 43492 4616 43548
rect 4552 43488 4616 43492
rect 4632 43548 4696 43552
rect 4632 43492 4636 43548
rect 4636 43492 4692 43548
rect 4692 43492 4696 43548
rect 4632 43488 4696 43492
rect 4712 43548 4776 43552
rect 4712 43492 4716 43548
rect 4716 43492 4772 43548
rect 4772 43492 4776 43548
rect 4712 43488 4776 43492
rect 4792 43548 4856 43552
rect 4792 43492 4796 43548
rect 4796 43492 4852 43548
rect 4852 43492 4856 43548
rect 4792 43488 4856 43492
rect 6152 43548 6216 43552
rect 6152 43492 6156 43548
rect 6156 43492 6212 43548
rect 6212 43492 6216 43548
rect 6152 43488 6216 43492
rect 6232 43548 6296 43552
rect 6232 43492 6236 43548
rect 6236 43492 6292 43548
rect 6292 43492 6296 43548
rect 6232 43488 6296 43492
rect 6312 43548 6376 43552
rect 6312 43492 6316 43548
rect 6316 43492 6372 43548
rect 6372 43492 6376 43548
rect 6312 43488 6376 43492
rect 6392 43548 6456 43552
rect 6392 43492 6396 43548
rect 6396 43492 6452 43548
rect 6452 43492 6456 43548
rect 6392 43488 6456 43492
rect 7752 43548 7816 43552
rect 7752 43492 7756 43548
rect 7756 43492 7812 43548
rect 7812 43492 7816 43548
rect 7752 43488 7816 43492
rect 7832 43548 7896 43552
rect 7832 43492 7836 43548
rect 7836 43492 7892 43548
rect 7892 43492 7896 43548
rect 7832 43488 7896 43492
rect 7912 43548 7976 43552
rect 7912 43492 7916 43548
rect 7916 43492 7972 43548
rect 7972 43492 7976 43548
rect 7912 43488 7976 43492
rect 7992 43548 8056 43552
rect 7992 43492 7996 43548
rect 7996 43492 8052 43548
rect 8052 43492 8056 43548
rect 7992 43488 8056 43492
rect 9352 43548 9416 43552
rect 9352 43492 9356 43548
rect 9356 43492 9412 43548
rect 9412 43492 9416 43548
rect 9352 43488 9416 43492
rect 9432 43548 9496 43552
rect 9432 43492 9436 43548
rect 9436 43492 9492 43548
rect 9492 43492 9496 43548
rect 9432 43488 9496 43492
rect 9512 43548 9576 43552
rect 9512 43492 9516 43548
rect 9516 43492 9572 43548
rect 9572 43492 9576 43548
rect 9512 43488 9576 43492
rect 9592 43548 9656 43552
rect 9592 43492 9596 43548
rect 9596 43492 9652 43548
rect 9652 43492 9656 43548
rect 9592 43488 9656 43492
rect 3612 43004 3676 43008
rect 3612 42948 3616 43004
rect 3616 42948 3672 43004
rect 3672 42948 3676 43004
rect 3612 42944 3676 42948
rect 3692 43004 3756 43008
rect 3692 42948 3696 43004
rect 3696 42948 3752 43004
rect 3752 42948 3756 43004
rect 3692 42944 3756 42948
rect 3772 43004 3836 43008
rect 3772 42948 3776 43004
rect 3776 42948 3832 43004
rect 3832 42948 3836 43004
rect 3772 42944 3836 42948
rect 3852 43004 3916 43008
rect 3852 42948 3856 43004
rect 3856 42948 3912 43004
rect 3912 42948 3916 43004
rect 3852 42944 3916 42948
rect 5212 43004 5276 43008
rect 5212 42948 5216 43004
rect 5216 42948 5272 43004
rect 5272 42948 5276 43004
rect 5212 42944 5276 42948
rect 5292 43004 5356 43008
rect 5292 42948 5296 43004
rect 5296 42948 5352 43004
rect 5352 42948 5356 43004
rect 5292 42944 5356 42948
rect 5372 43004 5436 43008
rect 5372 42948 5376 43004
rect 5376 42948 5432 43004
rect 5432 42948 5436 43004
rect 5372 42944 5436 42948
rect 5452 43004 5516 43008
rect 5452 42948 5456 43004
rect 5456 42948 5512 43004
rect 5512 42948 5516 43004
rect 5452 42944 5516 42948
rect 6812 43004 6876 43008
rect 6812 42948 6816 43004
rect 6816 42948 6872 43004
rect 6872 42948 6876 43004
rect 6812 42944 6876 42948
rect 6892 43004 6956 43008
rect 6892 42948 6896 43004
rect 6896 42948 6952 43004
rect 6952 42948 6956 43004
rect 6892 42944 6956 42948
rect 6972 43004 7036 43008
rect 6972 42948 6976 43004
rect 6976 42948 7032 43004
rect 7032 42948 7036 43004
rect 6972 42944 7036 42948
rect 7052 43004 7116 43008
rect 7052 42948 7056 43004
rect 7056 42948 7112 43004
rect 7112 42948 7116 43004
rect 7052 42944 7116 42948
rect 8412 43004 8476 43008
rect 8412 42948 8416 43004
rect 8416 42948 8472 43004
rect 8472 42948 8476 43004
rect 8412 42944 8476 42948
rect 8492 43004 8556 43008
rect 8492 42948 8496 43004
rect 8496 42948 8552 43004
rect 8552 42948 8556 43004
rect 8492 42944 8556 42948
rect 8572 43004 8636 43008
rect 8572 42948 8576 43004
rect 8576 42948 8632 43004
rect 8632 42948 8636 43004
rect 8572 42944 8636 42948
rect 8652 43004 8716 43008
rect 8652 42948 8656 43004
rect 8656 42948 8712 43004
rect 8712 42948 8716 43004
rect 8652 42944 8716 42948
rect 2952 42460 3016 42464
rect 2952 42404 2956 42460
rect 2956 42404 3012 42460
rect 3012 42404 3016 42460
rect 2952 42400 3016 42404
rect 3032 42460 3096 42464
rect 3032 42404 3036 42460
rect 3036 42404 3092 42460
rect 3092 42404 3096 42460
rect 3032 42400 3096 42404
rect 3112 42460 3176 42464
rect 3112 42404 3116 42460
rect 3116 42404 3172 42460
rect 3172 42404 3176 42460
rect 3112 42400 3176 42404
rect 3192 42460 3256 42464
rect 3192 42404 3196 42460
rect 3196 42404 3252 42460
rect 3252 42404 3256 42460
rect 3192 42400 3256 42404
rect 4552 42460 4616 42464
rect 4552 42404 4556 42460
rect 4556 42404 4612 42460
rect 4612 42404 4616 42460
rect 4552 42400 4616 42404
rect 4632 42460 4696 42464
rect 4632 42404 4636 42460
rect 4636 42404 4692 42460
rect 4692 42404 4696 42460
rect 4632 42400 4696 42404
rect 4712 42460 4776 42464
rect 4712 42404 4716 42460
rect 4716 42404 4772 42460
rect 4772 42404 4776 42460
rect 4712 42400 4776 42404
rect 4792 42460 4856 42464
rect 4792 42404 4796 42460
rect 4796 42404 4852 42460
rect 4852 42404 4856 42460
rect 4792 42400 4856 42404
rect 6152 42460 6216 42464
rect 6152 42404 6156 42460
rect 6156 42404 6212 42460
rect 6212 42404 6216 42460
rect 6152 42400 6216 42404
rect 6232 42460 6296 42464
rect 6232 42404 6236 42460
rect 6236 42404 6292 42460
rect 6292 42404 6296 42460
rect 6232 42400 6296 42404
rect 6312 42460 6376 42464
rect 6312 42404 6316 42460
rect 6316 42404 6372 42460
rect 6372 42404 6376 42460
rect 6312 42400 6376 42404
rect 6392 42460 6456 42464
rect 6392 42404 6396 42460
rect 6396 42404 6452 42460
rect 6452 42404 6456 42460
rect 6392 42400 6456 42404
rect 7752 42460 7816 42464
rect 7752 42404 7756 42460
rect 7756 42404 7812 42460
rect 7812 42404 7816 42460
rect 7752 42400 7816 42404
rect 7832 42460 7896 42464
rect 7832 42404 7836 42460
rect 7836 42404 7892 42460
rect 7892 42404 7896 42460
rect 7832 42400 7896 42404
rect 7912 42460 7976 42464
rect 7912 42404 7916 42460
rect 7916 42404 7972 42460
rect 7972 42404 7976 42460
rect 7912 42400 7976 42404
rect 7992 42460 8056 42464
rect 7992 42404 7996 42460
rect 7996 42404 8052 42460
rect 8052 42404 8056 42460
rect 7992 42400 8056 42404
rect 9352 42460 9416 42464
rect 9352 42404 9356 42460
rect 9356 42404 9412 42460
rect 9412 42404 9416 42460
rect 9352 42400 9416 42404
rect 9432 42460 9496 42464
rect 9432 42404 9436 42460
rect 9436 42404 9492 42460
rect 9492 42404 9496 42460
rect 9432 42400 9496 42404
rect 9512 42460 9576 42464
rect 9512 42404 9516 42460
rect 9516 42404 9572 42460
rect 9572 42404 9576 42460
rect 9512 42400 9576 42404
rect 9592 42460 9656 42464
rect 9592 42404 9596 42460
rect 9596 42404 9652 42460
rect 9652 42404 9656 42460
rect 9592 42400 9656 42404
rect 3612 41916 3676 41920
rect 3612 41860 3616 41916
rect 3616 41860 3672 41916
rect 3672 41860 3676 41916
rect 3612 41856 3676 41860
rect 3692 41916 3756 41920
rect 3692 41860 3696 41916
rect 3696 41860 3752 41916
rect 3752 41860 3756 41916
rect 3692 41856 3756 41860
rect 3772 41916 3836 41920
rect 3772 41860 3776 41916
rect 3776 41860 3832 41916
rect 3832 41860 3836 41916
rect 3772 41856 3836 41860
rect 3852 41916 3916 41920
rect 3852 41860 3856 41916
rect 3856 41860 3912 41916
rect 3912 41860 3916 41916
rect 3852 41856 3916 41860
rect 5212 41916 5276 41920
rect 5212 41860 5216 41916
rect 5216 41860 5272 41916
rect 5272 41860 5276 41916
rect 5212 41856 5276 41860
rect 5292 41916 5356 41920
rect 5292 41860 5296 41916
rect 5296 41860 5352 41916
rect 5352 41860 5356 41916
rect 5292 41856 5356 41860
rect 5372 41916 5436 41920
rect 5372 41860 5376 41916
rect 5376 41860 5432 41916
rect 5432 41860 5436 41916
rect 5372 41856 5436 41860
rect 5452 41916 5516 41920
rect 5452 41860 5456 41916
rect 5456 41860 5512 41916
rect 5512 41860 5516 41916
rect 5452 41856 5516 41860
rect 6812 41916 6876 41920
rect 6812 41860 6816 41916
rect 6816 41860 6872 41916
rect 6872 41860 6876 41916
rect 6812 41856 6876 41860
rect 6892 41916 6956 41920
rect 6892 41860 6896 41916
rect 6896 41860 6952 41916
rect 6952 41860 6956 41916
rect 6892 41856 6956 41860
rect 6972 41916 7036 41920
rect 6972 41860 6976 41916
rect 6976 41860 7032 41916
rect 7032 41860 7036 41916
rect 6972 41856 7036 41860
rect 7052 41916 7116 41920
rect 7052 41860 7056 41916
rect 7056 41860 7112 41916
rect 7112 41860 7116 41916
rect 7052 41856 7116 41860
rect 8412 41916 8476 41920
rect 8412 41860 8416 41916
rect 8416 41860 8472 41916
rect 8472 41860 8476 41916
rect 8412 41856 8476 41860
rect 8492 41916 8556 41920
rect 8492 41860 8496 41916
rect 8496 41860 8552 41916
rect 8552 41860 8556 41916
rect 8492 41856 8556 41860
rect 8572 41916 8636 41920
rect 8572 41860 8576 41916
rect 8576 41860 8632 41916
rect 8632 41860 8636 41916
rect 8572 41856 8636 41860
rect 8652 41916 8716 41920
rect 8652 41860 8656 41916
rect 8656 41860 8712 41916
rect 8712 41860 8716 41916
rect 8652 41856 8716 41860
rect 2952 41372 3016 41376
rect 2952 41316 2956 41372
rect 2956 41316 3012 41372
rect 3012 41316 3016 41372
rect 2952 41312 3016 41316
rect 3032 41372 3096 41376
rect 3032 41316 3036 41372
rect 3036 41316 3092 41372
rect 3092 41316 3096 41372
rect 3032 41312 3096 41316
rect 3112 41372 3176 41376
rect 3112 41316 3116 41372
rect 3116 41316 3172 41372
rect 3172 41316 3176 41372
rect 3112 41312 3176 41316
rect 3192 41372 3256 41376
rect 3192 41316 3196 41372
rect 3196 41316 3252 41372
rect 3252 41316 3256 41372
rect 3192 41312 3256 41316
rect 4552 41372 4616 41376
rect 4552 41316 4556 41372
rect 4556 41316 4612 41372
rect 4612 41316 4616 41372
rect 4552 41312 4616 41316
rect 4632 41372 4696 41376
rect 4632 41316 4636 41372
rect 4636 41316 4692 41372
rect 4692 41316 4696 41372
rect 4632 41312 4696 41316
rect 4712 41372 4776 41376
rect 4712 41316 4716 41372
rect 4716 41316 4772 41372
rect 4772 41316 4776 41372
rect 4712 41312 4776 41316
rect 4792 41372 4856 41376
rect 4792 41316 4796 41372
rect 4796 41316 4852 41372
rect 4852 41316 4856 41372
rect 4792 41312 4856 41316
rect 6152 41372 6216 41376
rect 6152 41316 6156 41372
rect 6156 41316 6212 41372
rect 6212 41316 6216 41372
rect 6152 41312 6216 41316
rect 6232 41372 6296 41376
rect 6232 41316 6236 41372
rect 6236 41316 6292 41372
rect 6292 41316 6296 41372
rect 6232 41312 6296 41316
rect 6312 41372 6376 41376
rect 6312 41316 6316 41372
rect 6316 41316 6372 41372
rect 6372 41316 6376 41372
rect 6312 41312 6376 41316
rect 6392 41372 6456 41376
rect 6392 41316 6396 41372
rect 6396 41316 6452 41372
rect 6452 41316 6456 41372
rect 6392 41312 6456 41316
rect 7752 41372 7816 41376
rect 7752 41316 7756 41372
rect 7756 41316 7812 41372
rect 7812 41316 7816 41372
rect 7752 41312 7816 41316
rect 7832 41372 7896 41376
rect 7832 41316 7836 41372
rect 7836 41316 7892 41372
rect 7892 41316 7896 41372
rect 7832 41312 7896 41316
rect 7912 41372 7976 41376
rect 7912 41316 7916 41372
rect 7916 41316 7972 41372
rect 7972 41316 7976 41372
rect 7912 41312 7976 41316
rect 7992 41372 8056 41376
rect 7992 41316 7996 41372
rect 7996 41316 8052 41372
rect 8052 41316 8056 41372
rect 7992 41312 8056 41316
rect 9352 41372 9416 41376
rect 9352 41316 9356 41372
rect 9356 41316 9412 41372
rect 9412 41316 9416 41372
rect 9352 41312 9416 41316
rect 9432 41372 9496 41376
rect 9432 41316 9436 41372
rect 9436 41316 9492 41372
rect 9492 41316 9496 41372
rect 9432 41312 9496 41316
rect 9512 41372 9576 41376
rect 9512 41316 9516 41372
rect 9516 41316 9572 41372
rect 9572 41316 9576 41372
rect 9512 41312 9576 41316
rect 9592 41372 9656 41376
rect 9592 41316 9596 41372
rect 9596 41316 9652 41372
rect 9652 41316 9656 41372
rect 9592 41312 9656 41316
rect 3612 40828 3676 40832
rect 3612 40772 3616 40828
rect 3616 40772 3672 40828
rect 3672 40772 3676 40828
rect 3612 40768 3676 40772
rect 3692 40828 3756 40832
rect 3692 40772 3696 40828
rect 3696 40772 3752 40828
rect 3752 40772 3756 40828
rect 3692 40768 3756 40772
rect 3772 40828 3836 40832
rect 3772 40772 3776 40828
rect 3776 40772 3832 40828
rect 3832 40772 3836 40828
rect 3772 40768 3836 40772
rect 3852 40828 3916 40832
rect 3852 40772 3856 40828
rect 3856 40772 3912 40828
rect 3912 40772 3916 40828
rect 3852 40768 3916 40772
rect 5212 40828 5276 40832
rect 5212 40772 5216 40828
rect 5216 40772 5272 40828
rect 5272 40772 5276 40828
rect 5212 40768 5276 40772
rect 5292 40828 5356 40832
rect 5292 40772 5296 40828
rect 5296 40772 5352 40828
rect 5352 40772 5356 40828
rect 5292 40768 5356 40772
rect 5372 40828 5436 40832
rect 5372 40772 5376 40828
rect 5376 40772 5432 40828
rect 5432 40772 5436 40828
rect 5372 40768 5436 40772
rect 5452 40828 5516 40832
rect 5452 40772 5456 40828
rect 5456 40772 5512 40828
rect 5512 40772 5516 40828
rect 5452 40768 5516 40772
rect 6812 40828 6876 40832
rect 6812 40772 6816 40828
rect 6816 40772 6872 40828
rect 6872 40772 6876 40828
rect 6812 40768 6876 40772
rect 6892 40828 6956 40832
rect 6892 40772 6896 40828
rect 6896 40772 6952 40828
rect 6952 40772 6956 40828
rect 6892 40768 6956 40772
rect 6972 40828 7036 40832
rect 6972 40772 6976 40828
rect 6976 40772 7032 40828
rect 7032 40772 7036 40828
rect 6972 40768 7036 40772
rect 7052 40828 7116 40832
rect 7052 40772 7056 40828
rect 7056 40772 7112 40828
rect 7112 40772 7116 40828
rect 7052 40768 7116 40772
rect 8412 40828 8476 40832
rect 8412 40772 8416 40828
rect 8416 40772 8472 40828
rect 8472 40772 8476 40828
rect 8412 40768 8476 40772
rect 8492 40828 8556 40832
rect 8492 40772 8496 40828
rect 8496 40772 8552 40828
rect 8552 40772 8556 40828
rect 8492 40768 8556 40772
rect 8572 40828 8636 40832
rect 8572 40772 8576 40828
rect 8576 40772 8632 40828
rect 8632 40772 8636 40828
rect 8572 40768 8636 40772
rect 8652 40828 8716 40832
rect 8652 40772 8656 40828
rect 8656 40772 8712 40828
rect 8712 40772 8716 40828
rect 8652 40768 8716 40772
rect 2952 40284 3016 40288
rect 2952 40228 2956 40284
rect 2956 40228 3012 40284
rect 3012 40228 3016 40284
rect 2952 40224 3016 40228
rect 3032 40284 3096 40288
rect 3032 40228 3036 40284
rect 3036 40228 3092 40284
rect 3092 40228 3096 40284
rect 3032 40224 3096 40228
rect 3112 40284 3176 40288
rect 3112 40228 3116 40284
rect 3116 40228 3172 40284
rect 3172 40228 3176 40284
rect 3112 40224 3176 40228
rect 3192 40284 3256 40288
rect 3192 40228 3196 40284
rect 3196 40228 3252 40284
rect 3252 40228 3256 40284
rect 3192 40224 3256 40228
rect 4552 40284 4616 40288
rect 4552 40228 4556 40284
rect 4556 40228 4612 40284
rect 4612 40228 4616 40284
rect 4552 40224 4616 40228
rect 4632 40284 4696 40288
rect 4632 40228 4636 40284
rect 4636 40228 4692 40284
rect 4692 40228 4696 40284
rect 4632 40224 4696 40228
rect 4712 40284 4776 40288
rect 4712 40228 4716 40284
rect 4716 40228 4772 40284
rect 4772 40228 4776 40284
rect 4712 40224 4776 40228
rect 4792 40284 4856 40288
rect 4792 40228 4796 40284
rect 4796 40228 4852 40284
rect 4852 40228 4856 40284
rect 4792 40224 4856 40228
rect 6152 40284 6216 40288
rect 6152 40228 6156 40284
rect 6156 40228 6212 40284
rect 6212 40228 6216 40284
rect 6152 40224 6216 40228
rect 6232 40284 6296 40288
rect 6232 40228 6236 40284
rect 6236 40228 6292 40284
rect 6292 40228 6296 40284
rect 6232 40224 6296 40228
rect 6312 40284 6376 40288
rect 6312 40228 6316 40284
rect 6316 40228 6372 40284
rect 6372 40228 6376 40284
rect 6312 40224 6376 40228
rect 6392 40284 6456 40288
rect 6392 40228 6396 40284
rect 6396 40228 6452 40284
rect 6452 40228 6456 40284
rect 6392 40224 6456 40228
rect 7752 40284 7816 40288
rect 7752 40228 7756 40284
rect 7756 40228 7812 40284
rect 7812 40228 7816 40284
rect 7752 40224 7816 40228
rect 7832 40284 7896 40288
rect 7832 40228 7836 40284
rect 7836 40228 7892 40284
rect 7892 40228 7896 40284
rect 7832 40224 7896 40228
rect 7912 40284 7976 40288
rect 7912 40228 7916 40284
rect 7916 40228 7972 40284
rect 7972 40228 7976 40284
rect 7912 40224 7976 40228
rect 7992 40284 8056 40288
rect 7992 40228 7996 40284
rect 7996 40228 8052 40284
rect 8052 40228 8056 40284
rect 7992 40224 8056 40228
rect 9352 40284 9416 40288
rect 9352 40228 9356 40284
rect 9356 40228 9412 40284
rect 9412 40228 9416 40284
rect 9352 40224 9416 40228
rect 9432 40284 9496 40288
rect 9432 40228 9436 40284
rect 9436 40228 9492 40284
rect 9492 40228 9496 40284
rect 9432 40224 9496 40228
rect 9512 40284 9576 40288
rect 9512 40228 9516 40284
rect 9516 40228 9572 40284
rect 9572 40228 9576 40284
rect 9512 40224 9576 40228
rect 9592 40284 9656 40288
rect 9592 40228 9596 40284
rect 9596 40228 9652 40284
rect 9652 40228 9656 40284
rect 9592 40224 9656 40228
rect 11100 39884 11164 39948
rect 3612 39740 3676 39744
rect 3612 39684 3616 39740
rect 3616 39684 3672 39740
rect 3672 39684 3676 39740
rect 3612 39680 3676 39684
rect 3692 39740 3756 39744
rect 3692 39684 3696 39740
rect 3696 39684 3752 39740
rect 3752 39684 3756 39740
rect 3692 39680 3756 39684
rect 3772 39740 3836 39744
rect 3772 39684 3776 39740
rect 3776 39684 3832 39740
rect 3832 39684 3836 39740
rect 3772 39680 3836 39684
rect 3852 39740 3916 39744
rect 3852 39684 3856 39740
rect 3856 39684 3912 39740
rect 3912 39684 3916 39740
rect 3852 39680 3916 39684
rect 5212 39740 5276 39744
rect 5212 39684 5216 39740
rect 5216 39684 5272 39740
rect 5272 39684 5276 39740
rect 5212 39680 5276 39684
rect 5292 39740 5356 39744
rect 5292 39684 5296 39740
rect 5296 39684 5352 39740
rect 5352 39684 5356 39740
rect 5292 39680 5356 39684
rect 5372 39740 5436 39744
rect 5372 39684 5376 39740
rect 5376 39684 5432 39740
rect 5432 39684 5436 39740
rect 5372 39680 5436 39684
rect 5452 39740 5516 39744
rect 5452 39684 5456 39740
rect 5456 39684 5512 39740
rect 5512 39684 5516 39740
rect 5452 39680 5516 39684
rect 6812 39740 6876 39744
rect 6812 39684 6816 39740
rect 6816 39684 6872 39740
rect 6872 39684 6876 39740
rect 6812 39680 6876 39684
rect 6892 39740 6956 39744
rect 6892 39684 6896 39740
rect 6896 39684 6952 39740
rect 6952 39684 6956 39740
rect 6892 39680 6956 39684
rect 6972 39740 7036 39744
rect 6972 39684 6976 39740
rect 6976 39684 7032 39740
rect 7032 39684 7036 39740
rect 6972 39680 7036 39684
rect 7052 39740 7116 39744
rect 7052 39684 7056 39740
rect 7056 39684 7112 39740
rect 7112 39684 7116 39740
rect 7052 39680 7116 39684
rect 8412 39740 8476 39744
rect 8412 39684 8416 39740
rect 8416 39684 8472 39740
rect 8472 39684 8476 39740
rect 8412 39680 8476 39684
rect 8492 39740 8556 39744
rect 8492 39684 8496 39740
rect 8496 39684 8552 39740
rect 8552 39684 8556 39740
rect 8492 39680 8556 39684
rect 8572 39740 8636 39744
rect 8572 39684 8576 39740
rect 8576 39684 8632 39740
rect 8632 39684 8636 39740
rect 8572 39680 8636 39684
rect 8652 39740 8716 39744
rect 8652 39684 8656 39740
rect 8656 39684 8712 39740
rect 8712 39684 8716 39740
rect 8652 39680 8716 39684
rect 2952 39196 3016 39200
rect 2952 39140 2956 39196
rect 2956 39140 3012 39196
rect 3012 39140 3016 39196
rect 2952 39136 3016 39140
rect 3032 39196 3096 39200
rect 3032 39140 3036 39196
rect 3036 39140 3092 39196
rect 3092 39140 3096 39196
rect 3032 39136 3096 39140
rect 3112 39196 3176 39200
rect 3112 39140 3116 39196
rect 3116 39140 3172 39196
rect 3172 39140 3176 39196
rect 3112 39136 3176 39140
rect 3192 39196 3256 39200
rect 3192 39140 3196 39196
rect 3196 39140 3252 39196
rect 3252 39140 3256 39196
rect 3192 39136 3256 39140
rect 4552 39196 4616 39200
rect 4552 39140 4556 39196
rect 4556 39140 4612 39196
rect 4612 39140 4616 39196
rect 4552 39136 4616 39140
rect 4632 39196 4696 39200
rect 4632 39140 4636 39196
rect 4636 39140 4692 39196
rect 4692 39140 4696 39196
rect 4632 39136 4696 39140
rect 4712 39196 4776 39200
rect 4712 39140 4716 39196
rect 4716 39140 4772 39196
rect 4772 39140 4776 39196
rect 4712 39136 4776 39140
rect 4792 39196 4856 39200
rect 4792 39140 4796 39196
rect 4796 39140 4852 39196
rect 4852 39140 4856 39196
rect 4792 39136 4856 39140
rect 6152 39196 6216 39200
rect 6152 39140 6156 39196
rect 6156 39140 6212 39196
rect 6212 39140 6216 39196
rect 6152 39136 6216 39140
rect 6232 39196 6296 39200
rect 6232 39140 6236 39196
rect 6236 39140 6292 39196
rect 6292 39140 6296 39196
rect 6232 39136 6296 39140
rect 6312 39196 6376 39200
rect 6312 39140 6316 39196
rect 6316 39140 6372 39196
rect 6372 39140 6376 39196
rect 6312 39136 6376 39140
rect 6392 39196 6456 39200
rect 6392 39140 6396 39196
rect 6396 39140 6452 39196
rect 6452 39140 6456 39196
rect 6392 39136 6456 39140
rect 7752 39196 7816 39200
rect 7752 39140 7756 39196
rect 7756 39140 7812 39196
rect 7812 39140 7816 39196
rect 7752 39136 7816 39140
rect 7832 39196 7896 39200
rect 7832 39140 7836 39196
rect 7836 39140 7892 39196
rect 7892 39140 7896 39196
rect 7832 39136 7896 39140
rect 7912 39196 7976 39200
rect 7912 39140 7916 39196
rect 7916 39140 7972 39196
rect 7972 39140 7976 39196
rect 7912 39136 7976 39140
rect 7992 39196 8056 39200
rect 7992 39140 7996 39196
rect 7996 39140 8052 39196
rect 8052 39140 8056 39196
rect 7992 39136 8056 39140
rect 9352 39196 9416 39200
rect 9352 39140 9356 39196
rect 9356 39140 9412 39196
rect 9412 39140 9416 39196
rect 9352 39136 9416 39140
rect 9432 39196 9496 39200
rect 9432 39140 9436 39196
rect 9436 39140 9492 39196
rect 9492 39140 9496 39196
rect 9432 39136 9496 39140
rect 9512 39196 9576 39200
rect 9512 39140 9516 39196
rect 9516 39140 9572 39196
rect 9572 39140 9576 39196
rect 9512 39136 9576 39140
rect 9592 39196 9656 39200
rect 9592 39140 9596 39196
rect 9596 39140 9652 39196
rect 9652 39140 9656 39196
rect 9592 39136 9656 39140
rect 3612 38652 3676 38656
rect 3612 38596 3616 38652
rect 3616 38596 3672 38652
rect 3672 38596 3676 38652
rect 3612 38592 3676 38596
rect 3692 38652 3756 38656
rect 3692 38596 3696 38652
rect 3696 38596 3752 38652
rect 3752 38596 3756 38652
rect 3692 38592 3756 38596
rect 3772 38652 3836 38656
rect 3772 38596 3776 38652
rect 3776 38596 3832 38652
rect 3832 38596 3836 38652
rect 3772 38592 3836 38596
rect 3852 38652 3916 38656
rect 3852 38596 3856 38652
rect 3856 38596 3912 38652
rect 3912 38596 3916 38652
rect 3852 38592 3916 38596
rect 5212 38652 5276 38656
rect 5212 38596 5216 38652
rect 5216 38596 5272 38652
rect 5272 38596 5276 38652
rect 5212 38592 5276 38596
rect 5292 38652 5356 38656
rect 5292 38596 5296 38652
rect 5296 38596 5352 38652
rect 5352 38596 5356 38652
rect 5292 38592 5356 38596
rect 5372 38652 5436 38656
rect 5372 38596 5376 38652
rect 5376 38596 5432 38652
rect 5432 38596 5436 38652
rect 5372 38592 5436 38596
rect 5452 38652 5516 38656
rect 5452 38596 5456 38652
rect 5456 38596 5512 38652
rect 5512 38596 5516 38652
rect 5452 38592 5516 38596
rect 6812 38652 6876 38656
rect 6812 38596 6816 38652
rect 6816 38596 6872 38652
rect 6872 38596 6876 38652
rect 6812 38592 6876 38596
rect 6892 38652 6956 38656
rect 6892 38596 6896 38652
rect 6896 38596 6952 38652
rect 6952 38596 6956 38652
rect 6892 38592 6956 38596
rect 6972 38652 7036 38656
rect 6972 38596 6976 38652
rect 6976 38596 7032 38652
rect 7032 38596 7036 38652
rect 6972 38592 7036 38596
rect 7052 38652 7116 38656
rect 7052 38596 7056 38652
rect 7056 38596 7112 38652
rect 7112 38596 7116 38652
rect 7052 38592 7116 38596
rect 8412 38652 8476 38656
rect 8412 38596 8416 38652
rect 8416 38596 8472 38652
rect 8472 38596 8476 38652
rect 8412 38592 8476 38596
rect 8492 38652 8556 38656
rect 8492 38596 8496 38652
rect 8496 38596 8552 38652
rect 8552 38596 8556 38652
rect 8492 38592 8556 38596
rect 8572 38652 8636 38656
rect 8572 38596 8576 38652
rect 8576 38596 8632 38652
rect 8632 38596 8636 38652
rect 8572 38592 8636 38596
rect 8652 38652 8716 38656
rect 8652 38596 8656 38652
rect 8656 38596 8712 38652
rect 8712 38596 8716 38652
rect 8652 38592 8716 38596
rect 10548 38388 10612 38452
rect 2952 38108 3016 38112
rect 2952 38052 2956 38108
rect 2956 38052 3012 38108
rect 3012 38052 3016 38108
rect 2952 38048 3016 38052
rect 3032 38108 3096 38112
rect 3032 38052 3036 38108
rect 3036 38052 3092 38108
rect 3092 38052 3096 38108
rect 3032 38048 3096 38052
rect 3112 38108 3176 38112
rect 3112 38052 3116 38108
rect 3116 38052 3172 38108
rect 3172 38052 3176 38108
rect 3112 38048 3176 38052
rect 3192 38108 3256 38112
rect 3192 38052 3196 38108
rect 3196 38052 3252 38108
rect 3252 38052 3256 38108
rect 3192 38048 3256 38052
rect 4552 38108 4616 38112
rect 4552 38052 4556 38108
rect 4556 38052 4612 38108
rect 4612 38052 4616 38108
rect 4552 38048 4616 38052
rect 4632 38108 4696 38112
rect 4632 38052 4636 38108
rect 4636 38052 4692 38108
rect 4692 38052 4696 38108
rect 4632 38048 4696 38052
rect 4712 38108 4776 38112
rect 4712 38052 4716 38108
rect 4716 38052 4772 38108
rect 4772 38052 4776 38108
rect 4712 38048 4776 38052
rect 4792 38108 4856 38112
rect 4792 38052 4796 38108
rect 4796 38052 4852 38108
rect 4852 38052 4856 38108
rect 4792 38048 4856 38052
rect 6152 38108 6216 38112
rect 6152 38052 6156 38108
rect 6156 38052 6212 38108
rect 6212 38052 6216 38108
rect 6152 38048 6216 38052
rect 6232 38108 6296 38112
rect 6232 38052 6236 38108
rect 6236 38052 6292 38108
rect 6292 38052 6296 38108
rect 6232 38048 6296 38052
rect 6312 38108 6376 38112
rect 6312 38052 6316 38108
rect 6316 38052 6372 38108
rect 6372 38052 6376 38108
rect 6312 38048 6376 38052
rect 6392 38108 6456 38112
rect 6392 38052 6396 38108
rect 6396 38052 6452 38108
rect 6452 38052 6456 38108
rect 6392 38048 6456 38052
rect 7752 38108 7816 38112
rect 7752 38052 7756 38108
rect 7756 38052 7812 38108
rect 7812 38052 7816 38108
rect 7752 38048 7816 38052
rect 7832 38108 7896 38112
rect 7832 38052 7836 38108
rect 7836 38052 7892 38108
rect 7892 38052 7896 38108
rect 7832 38048 7896 38052
rect 7912 38108 7976 38112
rect 7912 38052 7916 38108
rect 7916 38052 7972 38108
rect 7972 38052 7976 38108
rect 7912 38048 7976 38052
rect 7992 38108 8056 38112
rect 7992 38052 7996 38108
rect 7996 38052 8052 38108
rect 8052 38052 8056 38108
rect 7992 38048 8056 38052
rect 9352 38108 9416 38112
rect 9352 38052 9356 38108
rect 9356 38052 9412 38108
rect 9412 38052 9416 38108
rect 9352 38048 9416 38052
rect 9432 38108 9496 38112
rect 9432 38052 9436 38108
rect 9436 38052 9492 38108
rect 9492 38052 9496 38108
rect 9432 38048 9496 38052
rect 9512 38108 9576 38112
rect 9512 38052 9516 38108
rect 9516 38052 9572 38108
rect 9572 38052 9576 38108
rect 9512 38048 9576 38052
rect 9592 38108 9656 38112
rect 9592 38052 9596 38108
rect 9596 38052 9652 38108
rect 9652 38052 9656 38108
rect 9592 38048 9656 38052
rect 3612 37564 3676 37568
rect 3612 37508 3616 37564
rect 3616 37508 3672 37564
rect 3672 37508 3676 37564
rect 3612 37504 3676 37508
rect 3692 37564 3756 37568
rect 3692 37508 3696 37564
rect 3696 37508 3752 37564
rect 3752 37508 3756 37564
rect 3692 37504 3756 37508
rect 3772 37564 3836 37568
rect 3772 37508 3776 37564
rect 3776 37508 3832 37564
rect 3832 37508 3836 37564
rect 3772 37504 3836 37508
rect 3852 37564 3916 37568
rect 3852 37508 3856 37564
rect 3856 37508 3912 37564
rect 3912 37508 3916 37564
rect 3852 37504 3916 37508
rect 5212 37564 5276 37568
rect 5212 37508 5216 37564
rect 5216 37508 5272 37564
rect 5272 37508 5276 37564
rect 5212 37504 5276 37508
rect 5292 37564 5356 37568
rect 5292 37508 5296 37564
rect 5296 37508 5352 37564
rect 5352 37508 5356 37564
rect 5292 37504 5356 37508
rect 5372 37564 5436 37568
rect 5372 37508 5376 37564
rect 5376 37508 5432 37564
rect 5432 37508 5436 37564
rect 5372 37504 5436 37508
rect 5452 37564 5516 37568
rect 5452 37508 5456 37564
rect 5456 37508 5512 37564
rect 5512 37508 5516 37564
rect 5452 37504 5516 37508
rect 6812 37564 6876 37568
rect 6812 37508 6816 37564
rect 6816 37508 6872 37564
rect 6872 37508 6876 37564
rect 6812 37504 6876 37508
rect 6892 37564 6956 37568
rect 6892 37508 6896 37564
rect 6896 37508 6952 37564
rect 6952 37508 6956 37564
rect 6892 37504 6956 37508
rect 6972 37564 7036 37568
rect 6972 37508 6976 37564
rect 6976 37508 7032 37564
rect 7032 37508 7036 37564
rect 6972 37504 7036 37508
rect 7052 37564 7116 37568
rect 7052 37508 7056 37564
rect 7056 37508 7112 37564
rect 7112 37508 7116 37564
rect 7052 37504 7116 37508
rect 8412 37564 8476 37568
rect 8412 37508 8416 37564
rect 8416 37508 8472 37564
rect 8472 37508 8476 37564
rect 8412 37504 8476 37508
rect 8492 37564 8556 37568
rect 8492 37508 8496 37564
rect 8496 37508 8552 37564
rect 8552 37508 8556 37564
rect 8492 37504 8556 37508
rect 8572 37564 8636 37568
rect 8572 37508 8576 37564
rect 8576 37508 8632 37564
rect 8632 37508 8636 37564
rect 8572 37504 8636 37508
rect 8652 37564 8716 37568
rect 8652 37508 8656 37564
rect 8656 37508 8712 37564
rect 8712 37508 8716 37564
rect 8652 37504 8716 37508
rect 796 37300 860 37364
rect 10732 37300 10796 37364
rect 2952 37020 3016 37024
rect 2952 36964 2956 37020
rect 2956 36964 3012 37020
rect 3012 36964 3016 37020
rect 2952 36960 3016 36964
rect 3032 37020 3096 37024
rect 3032 36964 3036 37020
rect 3036 36964 3092 37020
rect 3092 36964 3096 37020
rect 3032 36960 3096 36964
rect 3112 37020 3176 37024
rect 3112 36964 3116 37020
rect 3116 36964 3172 37020
rect 3172 36964 3176 37020
rect 3112 36960 3176 36964
rect 3192 37020 3256 37024
rect 3192 36964 3196 37020
rect 3196 36964 3252 37020
rect 3252 36964 3256 37020
rect 3192 36960 3256 36964
rect 4552 37020 4616 37024
rect 4552 36964 4556 37020
rect 4556 36964 4612 37020
rect 4612 36964 4616 37020
rect 4552 36960 4616 36964
rect 4632 37020 4696 37024
rect 4632 36964 4636 37020
rect 4636 36964 4692 37020
rect 4692 36964 4696 37020
rect 4632 36960 4696 36964
rect 4712 37020 4776 37024
rect 4712 36964 4716 37020
rect 4716 36964 4772 37020
rect 4772 36964 4776 37020
rect 4712 36960 4776 36964
rect 4792 37020 4856 37024
rect 4792 36964 4796 37020
rect 4796 36964 4852 37020
rect 4852 36964 4856 37020
rect 4792 36960 4856 36964
rect 6152 37020 6216 37024
rect 6152 36964 6156 37020
rect 6156 36964 6212 37020
rect 6212 36964 6216 37020
rect 6152 36960 6216 36964
rect 6232 37020 6296 37024
rect 6232 36964 6236 37020
rect 6236 36964 6292 37020
rect 6292 36964 6296 37020
rect 6232 36960 6296 36964
rect 6312 37020 6376 37024
rect 6312 36964 6316 37020
rect 6316 36964 6372 37020
rect 6372 36964 6376 37020
rect 6312 36960 6376 36964
rect 6392 37020 6456 37024
rect 6392 36964 6396 37020
rect 6396 36964 6452 37020
rect 6452 36964 6456 37020
rect 6392 36960 6456 36964
rect 7752 37020 7816 37024
rect 7752 36964 7756 37020
rect 7756 36964 7812 37020
rect 7812 36964 7816 37020
rect 7752 36960 7816 36964
rect 7832 37020 7896 37024
rect 7832 36964 7836 37020
rect 7836 36964 7892 37020
rect 7892 36964 7896 37020
rect 7832 36960 7896 36964
rect 7912 37020 7976 37024
rect 7912 36964 7916 37020
rect 7916 36964 7972 37020
rect 7972 36964 7976 37020
rect 7912 36960 7976 36964
rect 7992 37020 8056 37024
rect 7992 36964 7996 37020
rect 7996 36964 8052 37020
rect 8052 36964 8056 37020
rect 7992 36960 8056 36964
rect 9352 37020 9416 37024
rect 9352 36964 9356 37020
rect 9356 36964 9412 37020
rect 9412 36964 9416 37020
rect 9352 36960 9416 36964
rect 9432 37020 9496 37024
rect 9432 36964 9436 37020
rect 9436 36964 9492 37020
rect 9492 36964 9496 37020
rect 9432 36960 9496 36964
rect 9512 37020 9576 37024
rect 9512 36964 9516 37020
rect 9516 36964 9572 37020
rect 9572 36964 9576 37020
rect 9512 36960 9576 36964
rect 9592 37020 9656 37024
rect 9592 36964 9596 37020
rect 9596 36964 9652 37020
rect 9652 36964 9656 37020
rect 9592 36960 9656 36964
rect 3612 36476 3676 36480
rect 3612 36420 3616 36476
rect 3616 36420 3672 36476
rect 3672 36420 3676 36476
rect 3612 36416 3676 36420
rect 3692 36476 3756 36480
rect 3692 36420 3696 36476
rect 3696 36420 3752 36476
rect 3752 36420 3756 36476
rect 3692 36416 3756 36420
rect 3772 36476 3836 36480
rect 3772 36420 3776 36476
rect 3776 36420 3832 36476
rect 3832 36420 3836 36476
rect 3772 36416 3836 36420
rect 3852 36476 3916 36480
rect 3852 36420 3856 36476
rect 3856 36420 3912 36476
rect 3912 36420 3916 36476
rect 3852 36416 3916 36420
rect 5212 36476 5276 36480
rect 5212 36420 5216 36476
rect 5216 36420 5272 36476
rect 5272 36420 5276 36476
rect 5212 36416 5276 36420
rect 5292 36476 5356 36480
rect 5292 36420 5296 36476
rect 5296 36420 5352 36476
rect 5352 36420 5356 36476
rect 5292 36416 5356 36420
rect 5372 36476 5436 36480
rect 5372 36420 5376 36476
rect 5376 36420 5432 36476
rect 5432 36420 5436 36476
rect 5372 36416 5436 36420
rect 5452 36476 5516 36480
rect 5452 36420 5456 36476
rect 5456 36420 5512 36476
rect 5512 36420 5516 36476
rect 5452 36416 5516 36420
rect 6812 36476 6876 36480
rect 6812 36420 6816 36476
rect 6816 36420 6872 36476
rect 6872 36420 6876 36476
rect 6812 36416 6876 36420
rect 6892 36476 6956 36480
rect 6892 36420 6896 36476
rect 6896 36420 6952 36476
rect 6952 36420 6956 36476
rect 6892 36416 6956 36420
rect 6972 36476 7036 36480
rect 6972 36420 6976 36476
rect 6976 36420 7032 36476
rect 7032 36420 7036 36476
rect 6972 36416 7036 36420
rect 7052 36476 7116 36480
rect 7052 36420 7056 36476
rect 7056 36420 7112 36476
rect 7112 36420 7116 36476
rect 7052 36416 7116 36420
rect 8412 36476 8476 36480
rect 8412 36420 8416 36476
rect 8416 36420 8472 36476
rect 8472 36420 8476 36476
rect 8412 36416 8476 36420
rect 8492 36476 8556 36480
rect 8492 36420 8496 36476
rect 8496 36420 8552 36476
rect 8552 36420 8556 36476
rect 8492 36416 8556 36420
rect 8572 36476 8636 36480
rect 8572 36420 8576 36476
rect 8576 36420 8632 36476
rect 8632 36420 8636 36476
rect 8572 36416 8636 36420
rect 8652 36476 8716 36480
rect 8652 36420 8656 36476
rect 8656 36420 8712 36476
rect 8712 36420 8716 36476
rect 8652 36416 8716 36420
rect 11652 36348 11716 36412
rect 2952 35932 3016 35936
rect 2952 35876 2956 35932
rect 2956 35876 3012 35932
rect 3012 35876 3016 35932
rect 2952 35872 3016 35876
rect 3032 35932 3096 35936
rect 3032 35876 3036 35932
rect 3036 35876 3092 35932
rect 3092 35876 3096 35932
rect 3032 35872 3096 35876
rect 3112 35932 3176 35936
rect 3112 35876 3116 35932
rect 3116 35876 3172 35932
rect 3172 35876 3176 35932
rect 3112 35872 3176 35876
rect 3192 35932 3256 35936
rect 3192 35876 3196 35932
rect 3196 35876 3252 35932
rect 3252 35876 3256 35932
rect 3192 35872 3256 35876
rect 4552 35932 4616 35936
rect 4552 35876 4556 35932
rect 4556 35876 4612 35932
rect 4612 35876 4616 35932
rect 4552 35872 4616 35876
rect 4632 35932 4696 35936
rect 4632 35876 4636 35932
rect 4636 35876 4692 35932
rect 4692 35876 4696 35932
rect 4632 35872 4696 35876
rect 4712 35932 4776 35936
rect 4712 35876 4716 35932
rect 4716 35876 4772 35932
rect 4772 35876 4776 35932
rect 4712 35872 4776 35876
rect 4792 35932 4856 35936
rect 4792 35876 4796 35932
rect 4796 35876 4852 35932
rect 4852 35876 4856 35932
rect 4792 35872 4856 35876
rect 6152 35932 6216 35936
rect 6152 35876 6156 35932
rect 6156 35876 6212 35932
rect 6212 35876 6216 35932
rect 6152 35872 6216 35876
rect 6232 35932 6296 35936
rect 6232 35876 6236 35932
rect 6236 35876 6292 35932
rect 6292 35876 6296 35932
rect 6232 35872 6296 35876
rect 6312 35932 6376 35936
rect 6312 35876 6316 35932
rect 6316 35876 6372 35932
rect 6372 35876 6376 35932
rect 6312 35872 6376 35876
rect 6392 35932 6456 35936
rect 6392 35876 6396 35932
rect 6396 35876 6452 35932
rect 6452 35876 6456 35932
rect 6392 35872 6456 35876
rect 7752 35932 7816 35936
rect 7752 35876 7756 35932
rect 7756 35876 7812 35932
rect 7812 35876 7816 35932
rect 7752 35872 7816 35876
rect 7832 35932 7896 35936
rect 7832 35876 7836 35932
rect 7836 35876 7892 35932
rect 7892 35876 7896 35932
rect 7832 35872 7896 35876
rect 7912 35932 7976 35936
rect 7912 35876 7916 35932
rect 7916 35876 7972 35932
rect 7972 35876 7976 35932
rect 7912 35872 7976 35876
rect 7992 35932 8056 35936
rect 7992 35876 7996 35932
rect 7996 35876 8052 35932
rect 8052 35876 8056 35932
rect 7992 35872 8056 35876
rect 9352 35932 9416 35936
rect 9352 35876 9356 35932
rect 9356 35876 9412 35932
rect 9412 35876 9416 35932
rect 9352 35872 9416 35876
rect 9432 35932 9496 35936
rect 9432 35876 9436 35932
rect 9436 35876 9492 35932
rect 9492 35876 9496 35932
rect 9432 35872 9496 35876
rect 9512 35932 9576 35936
rect 9512 35876 9516 35932
rect 9516 35876 9572 35932
rect 9572 35876 9576 35932
rect 9512 35872 9576 35876
rect 9592 35932 9656 35936
rect 9592 35876 9596 35932
rect 9596 35876 9652 35932
rect 9652 35876 9656 35932
rect 9592 35872 9656 35876
rect 3612 35388 3676 35392
rect 3612 35332 3616 35388
rect 3616 35332 3672 35388
rect 3672 35332 3676 35388
rect 3612 35328 3676 35332
rect 3692 35388 3756 35392
rect 3692 35332 3696 35388
rect 3696 35332 3752 35388
rect 3752 35332 3756 35388
rect 3692 35328 3756 35332
rect 3772 35388 3836 35392
rect 3772 35332 3776 35388
rect 3776 35332 3832 35388
rect 3832 35332 3836 35388
rect 3772 35328 3836 35332
rect 3852 35388 3916 35392
rect 3852 35332 3856 35388
rect 3856 35332 3912 35388
rect 3912 35332 3916 35388
rect 3852 35328 3916 35332
rect 5212 35388 5276 35392
rect 5212 35332 5216 35388
rect 5216 35332 5272 35388
rect 5272 35332 5276 35388
rect 5212 35328 5276 35332
rect 5292 35388 5356 35392
rect 5292 35332 5296 35388
rect 5296 35332 5352 35388
rect 5352 35332 5356 35388
rect 5292 35328 5356 35332
rect 5372 35388 5436 35392
rect 5372 35332 5376 35388
rect 5376 35332 5432 35388
rect 5432 35332 5436 35388
rect 5372 35328 5436 35332
rect 5452 35388 5516 35392
rect 5452 35332 5456 35388
rect 5456 35332 5512 35388
rect 5512 35332 5516 35388
rect 5452 35328 5516 35332
rect 6812 35388 6876 35392
rect 6812 35332 6816 35388
rect 6816 35332 6872 35388
rect 6872 35332 6876 35388
rect 6812 35328 6876 35332
rect 6892 35388 6956 35392
rect 6892 35332 6896 35388
rect 6896 35332 6952 35388
rect 6952 35332 6956 35388
rect 6892 35328 6956 35332
rect 6972 35388 7036 35392
rect 6972 35332 6976 35388
rect 6976 35332 7032 35388
rect 7032 35332 7036 35388
rect 6972 35328 7036 35332
rect 7052 35388 7116 35392
rect 7052 35332 7056 35388
rect 7056 35332 7112 35388
rect 7112 35332 7116 35388
rect 7052 35328 7116 35332
rect 8412 35388 8476 35392
rect 8412 35332 8416 35388
rect 8416 35332 8472 35388
rect 8472 35332 8476 35388
rect 8412 35328 8476 35332
rect 8492 35388 8556 35392
rect 8492 35332 8496 35388
rect 8496 35332 8552 35388
rect 8552 35332 8556 35388
rect 8492 35328 8556 35332
rect 8572 35388 8636 35392
rect 8572 35332 8576 35388
rect 8576 35332 8632 35388
rect 8632 35332 8636 35388
rect 8572 35328 8636 35332
rect 8652 35388 8716 35392
rect 8652 35332 8656 35388
rect 8656 35332 8712 35388
rect 8712 35332 8716 35388
rect 8652 35328 8716 35332
rect 2952 34844 3016 34848
rect 2952 34788 2956 34844
rect 2956 34788 3012 34844
rect 3012 34788 3016 34844
rect 2952 34784 3016 34788
rect 3032 34844 3096 34848
rect 3032 34788 3036 34844
rect 3036 34788 3092 34844
rect 3092 34788 3096 34844
rect 3032 34784 3096 34788
rect 3112 34844 3176 34848
rect 3112 34788 3116 34844
rect 3116 34788 3172 34844
rect 3172 34788 3176 34844
rect 3112 34784 3176 34788
rect 3192 34844 3256 34848
rect 3192 34788 3196 34844
rect 3196 34788 3252 34844
rect 3252 34788 3256 34844
rect 3192 34784 3256 34788
rect 4552 34844 4616 34848
rect 4552 34788 4556 34844
rect 4556 34788 4612 34844
rect 4612 34788 4616 34844
rect 4552 34784 4616 34788
rect 4632 34844 4696 34848
rect 4632 34788 4636 34844
rect 4636 34788 4692 34844
rect 4692 34788 4696 34844
rect 4632 34784 4696 34788
rect 4712 34844 4776 34848
rect 4712 34788 4716 34844
rect 4716 34788 4772 34844
rect 4772 34788 4776 34844
rect 4712 34784 4776 34788
rect 4792 34844 4856 34848
rect 4792 34788 4796 34844
rect 4796 34788 4852 34844
rect 4852 34788 4856 34844
rect 4792 34784 4856 34788
rect 6152 34844 6216 34848
rect 6152 34788 6156 34844
rect 6156 34788 6212 34844
rect 6212 34788 6216 34844
rect 6152 34784 6216 34788
rect 6232 34844 6296 34848
rect 6232 34788 6236 34844
rect 6236 34788 6292 34844
rect 6292 34788 6296 34844
rect 6232 34784 6296 34788
rect 6312 34844 6376 34848
rect 6312 34788 6316 34844
rect 6316 34788 6372 34844
rect 6372 34788 6376 34844
rect 6312 34784 6376 34788
rect 6392 34844 6456 34848
rect 6392 34788 6396 34844
rect 6396 34788 6452 34844
rect 6452 34788 6456 34844
rect 6392 34784 6456 34788
rect 7752 34844 7816 34848
rect 7752 34788 7756 34844
rect 7756 34788 7812 34844
rect 7812 34788 7816 34844
rect 7752 34784 7816 34788
rect 7832 34844 7896 34848
rect 7832 34788 7836 34844
rect 7836 34788 7892 34844
rect 7892 34788 7896 34844
rect 7832 34784 7896 34788
rect 7912 34844 7976 34848
rect 7912 34788 7916 34844
rect 7916 34788 7972 34844
rect 7972 34788 7976 34844
rect 7912 34784 7976 34788
rect 7992 34844 8056 34848
rect 7992 34788 7996 34844
rect 7996 34788 8052 34844
rect 8052 34788 8056 34844
rect 7992 34784 8056 34788
rect 9352 34844 9416 34848
rect 9352 34788 9356 34844
rect 9356 34788 9412 34844
rect 9412 34788 9416 34844
rect 9352 34784 9416 34788
rect 9432 34844 9496 34848
rect 9432 34788 9436 34844
rect 9436 34788 9492 34844
rect 9492 34788 9496 34844
rect 9432 34784 9496 34788
rect 9512 34844 9576 34848
rect 9512 34788 9516 34844
rect 9516 34788 9572 34844
rect 9572 34788 9576 34844
rect 9512 34784 9576 34788
rect 9592 34844 9656 34848
rect 9592 34788 9596 34844
rect 9596 34788 9652 34844
rect 9652 34788 9656 34844
rect 9592 34784 9656 34788
rect 3612 34300 3676 34304
rect 3612 34244 3616 34300
rect 3616 34244 3672 34300
rect 3672 34244 3676 34300
rect 3612 34240 3676 34244
rect 3692 34300 3756 34304
rect 3692 34244 3696 34300
rect 3696 34244 3752 34300
rect 3752 34244 3756 34300
rect 3692 34240 3756 34244
rect 3772 34300 3836 34304
rect 3772 34244 3776 34300
rect 3776 34244 3832 34300
rect 3832 34244 3836 34300
rect 3772 34240 3836 34244
rect 3852 34300 3916 34304
rect 3852 34244 3856 34300
rect 3856 34244 3912 34300
rect 3912 34244 3916 34300
rect 3852 34240 3916 34244
rect 5212 34300 5276 34304
rect 5212 34244 5216 34300
rect 5216 34244 5272 34300
rect 5272 34244 5276 34300
rect 5212 34240 5276 34244
rect 5292 34300 5356 34304
rect 5292 34244 5296 34300
rect 5296 34244 5352 34300
rect 5352 34244 5356 34300
rect 5292 34240 5356 34244
rect 5372 34300 5436 34304
rect 5372 34244 5376 34300
rect 5376 34244 5432 34300
rect 5432 34244 5436 34300
rect 5372 34240 5436 34244
rect 5452 34300 5516 34304
rect 5452 34244 5456 34300
rect 5456 34244 5512 34300
rect 5512 34244 5516 34300
rect 5452 34240 5516 34244
rect 6812 34300 6876 34304
rect 6812 34244 6816 34300
rect 6816 34244 6872 34300
rect 6872 34244 6876 34300
rect 6812 34240 6876 34244
rect 6892 34300 6956 34304
rect 6892 34244 6896 34300
rect 6896 34244 6952 34300
rect 6952 34244 6956 34300
rect 6892 34240 6956 34244
rect 6972 34300 7036 34304
rect 6972 34244 6976 34300
rect 6976 34244 7032 34300
rect 7032 34244 7036 34300
rect 6972 34240 7036 34244
rect 7052 34300 7116 34304
rect 7052 34244 7056 34300
rect 7056 34244 7112 34300
rect 7112 34244 7116 34300
rect 7052 34240 7116 34244
rect 8412 34300 8476 34304
rect 8412 34244 8416 34300
rect 8416 34244 8472 34300
rect 8472 34244 8476 34300
rect 8412 34240 8476 34244
rect 8492 34300 8556 34304
rect 8492 34244 8496 34300
rect 8496 34244 8552 34300
rect 8552 34244 8556 34300
rect 8492 34240 8556 34244
rect 8572 34300 8636 34304
rect 8572 34244 8576 34300
rect 8576 34244 8632 34300
rect 8632 34244 8636 34300
rect 8572 34240 8636 34244
rect 8652 34300 8716 34304
rect 8652 34244 8656 34300
rect 8656 34244 8712 34300
rect 8712 34244 8716 34300
rect 8652 34240 8716 34244
rect 11836 34062 11900 34126
rect 2952 33756 3016 33760
rect 2952 33700 2956 33756
rect 2956 33700 3012 33756
rect 3012 33700 3016 33756
rect 2952 33696 3016 33700
rect 3032 33756 3096 33760
rect 3032 33700 3036 33756
rect 3036 33700 3092 33756
rect 3092 33700 3096 33756
rect 3032 33696 3096 33700
rect 3112 33756 3176 33760
rect 3112 33700 3116 33756
rect 3116 33700 3172 33756
rect 3172 33700 3176 33756
rect 3112 33696 3176 33700
rect 3192 33756 3256 33760
rect 3192 33700 3196 33756
rect 3196 33700 3252 33756
rect 3252 33700 3256 33756
rect 3192 33696 3256 33700
rect 4552 33756 4616 33760
rect 4552 33700 4556 33756
rect 4556 33700 4612 33756
rect 4612 33700 4616 33756
rect 4552 33696 4616 33700
rect 4632 33756 4696 33760
rect 4632 33700 4636 33756
rect 4636 33700 4692 33756
rect 4692 33700 4696 33756
rect 4632 33696 4696 33700
rect 4712 33756 4776 33760
rect 4712 33700 4716 33756
rect 4716 33700 4772 33756
rect 4772 33700 4776 33756
rect 4712 33696 4776 33700
rect 4792 33756 4856 33760
rect 4792 33700 4796 33756
rect 4796 33700 4852 33756
rect 4852 33700 4856 33756
rect 4792 33696 4856 33700
rect 6152 33756 6216 33760
rect 6152 33700 6156 33756
rect 6156 33700 6212 33756
rect 6212 33700 6216 33756
rect 6152 33696 6216 33700
rect 6232 33756 6296 33760
rect 6232 33700 6236 33756
rect 6236 33700 6292 33756
rect 6292 33700 6296 33756
rect 6232 33696 6296 33700
rect 6312 33756 6376 33760
rect 6312 33700 6316 33756
rect 6316 33700 6372 33756
rect 6372 33700 6376 33756
rect 6312 33696 6376 33700
rect 6392 33756 6456 33760
rect 6392 33700 6396 33756
rect 6396 33700 6452 33756
rect 6452 33700 6456 33756
rect 6392 33696 6456 33700
rect 7752 33756 7816 33760
rect 7752 33700 7756 33756
rect 7756 33700 7812 33756
rect 7812 33700 7816 33756
rect 7752 33696 7816 33700
rect 7832 33756 7896 33760
rect 7832 33700 7836 33756
rect 7836 33700 7892 33756
rect 7892 33700 7896 33756
rect 7832 33696 7896 33700
rect 7912 33756 7976 33760
rect 7912 33700 7916 33756
rect 7916 33700 7972 33756
rect 7972 33700 7976 33756
rect 7912 33696 7976 33700
rect 7992 33756 8056 33760
rect 7992 33700 7996 33756
rect 7996 33700 8052 33756
rect 8052 33700 8056 33756
rect 7992 33696 8056 33700
rect 9352 33756 9416 33760
rect 9352 33700 9356 33756
rect 9356 33700 9412 33756
rect 9412 33700 9416 33756
rect 9352 33696 9416 33700
rect 9432 33756 9496 33760
rect 9432 33700 9436 33756
rect 9436 33700 9492 33756
rect 9492 33700 9496 33756
rect 9432 33696 9496 33700
rect 9512 33756 9576 33760
rect 9512 33700 9516 33756
rect 9516 33700 9572 33756
rect 9572 33700 9576 33756
rect 9512 33696 9576 33700
rect 9592 33756 9656 33760
rect 9592 33700 9596 33756
rect 9596 33700 9652 33756
rect 9652 33700 9656 33756
rect 9592 33696 9656 33700
rect 3612 33212 3676 33216
rect 3612 33156 3616 33212
rect 3616 33156 3672 33212
rect 3672 33156 3676 33212
rect 3612 33152 3676 33156
rect 3692 33212 3756 33216
rect 3692 33156 3696 33212
rect 3696 33156 3752 33212
rect 3752 33156 3756 33212
rect 3692 33152 3756 33156
rect 3772 33212 3836 33216
rect 3772 33156 3776 33212
rect 3776 33156 3832 33212
rect 3832 33156 3836 33212
rect 3772 33152 3836 33156
rect 3852 33212 3916 33216
rect 3852 33156 3856 33212
rect 3856 33156 3912 33212
rect 3912 33156 3916 33212
rect 3852 33152 3916 33156
rect 5212 33212 5276 33216
rect 5212 33156 5216 33212
rect 5216 33156 5272 33212
rect 5272 33156 5276 33212
rect 5212 33152 5276 33156
rect 5292 33212 5356 33216
rect 5292 33156 5296 33212
rect 5296 33156 5352 33212
rect 5352 33156 5356 33212
rect 5292 33152 5356 33156
rect 5372 33212 5436 33216
rect 5372 33156 5376 33212
rect 5376 33156 5432 33212
rect 5432 33156 5436 33212
rect 5372 33152 5436 33156
rect 5452 33212 5516 33216
rect 5452 33156 5456 33212
rect 5456 33156 5512 33212
rect 5512 33156 5516 33212
rect 5452 33152 5516 33156
rect 6812 33212 6876 33216
rect 6812 33156 6816 33212
rect 6816 33156 6872 33212
rect 6872 33156 6876 33212
rect 6812 33152 6876 33156
rect 6892 33212 6956 33216
rect 6892 33156 6896 33212
rect 6896 33156 6952 33212
rect 6952 33156 6956 33212
rect 6892 33152 6956 33156
rect 6972 33212 7036 33216
rect 6972 33156 6976 33212
rect 6976 33156 7032 33212
rect 7032 33156 7036 33212
rect 6972 33152 7036 33156
rect 7052 33212 7116 33216
rect 7052 33156 7056 33212
rect 7056 33156 7112 33212
rect 7112 33156 7116 33212
rect 7052 33152 7116 33156
rect 8412 33212 8476 33216
rect 8412 33156 8416 33212
rect 8416 33156 8472 33212
rect 8472 33156 8476 33212
rect 8412 33152 8476 33156
rect 8492 33212 8556 33216
rect 8492 33156 8496 33212
rect 8496 33156 8552 33212
rect 8552 33156 8556 33212
rect 8492 33152 8556 33156
rect 8572 33212 8636 33216
rect 8572 33156 8576 33212
rect 8576 33156 8632 33212
rect 8632 33156 8636 33212
rect 8572 33152 8636 33156
rect 8652 33212 8716 33216
rect 8652 33156 8656 33212
rect 8656 33156 8712 33212
rect 8712 33156 8716 33212
rect 8652 33152 8716 33156
rect 2952 32668 3016 32672
rect 2952 32612 2956 32668
rect 2956 32612 3012 32668
rect 3012 32612 3016 32668
rect 2952 32608 3016 32612
rect 3032 32668 3096 32672
rect 3032 32612 3036 32668
rect 3036 32612 3092 32668
rect 3092 32612 3096 32668
rect 3032 32608 3096 32612
rect 3112 32668 3176 32672
rect 3112 32612 3116 32668
rect 3116 32612 3172 32668
rect 3172 32612 3176 32668
rect 3112 32608 3176 32612
rect 3192 32668 3256 32672
rect 3192 32612 3196 32668
rect 3196 32612 3252 32668
rect 3252 32612 3256 32668
rect 3192 32608 3256 32612
rect 4552 32668 4616 32672
rect 4552 32612 4556 32668
rect 4556 32612 4612 32668
rect 4612 32612 4616 32668
rect 4552 32608 4616 32612
rect 4632 32668 4696 32672
rect 4632 32612 4636 32668
rect 4636 32612 4692 32668
rect 4692 32612 4696 32668
rect 4632 32608 4696 32612
rect 4712 32668 4776 32672
rect 4712 32612 4716 32668
rect 4716 32612 4772 32668
rect 4772 32612 4776 32668
rect 4712 32608 4776 32612
rect 4792 32668 4856 32672
rect 4792 32612 4796 32668
rect 4796 32612 4852 32668
rect 4852 32612 4856 32668
rect 4792 32608 4856 32612
rect 6152 32668 6216 32672
rect 6152 32612 6156 32668
rect 6156 32612 6212 32668
rect 6212 32612 6216 32668
rect 6152 32608 6216 32612
rect 6232 32668 6296 32672
rect 6232 32612 6236 32668
rect 6236 32612 6292 32668
rect 6292 32612 6296 32668
rect 6232 32608 6296 32612
rect 6312 32668 6376 32672
rect 6312 32612 6316 32668
rect 6316 32612 6372 32668
rect 6372 32612 6376 32668
rect 6312 32608 6376 32612
rect 6392 32668 6456 32672
rect 6392 32612 6396 32668
rect 6396 32612 6452 32668
rect 6452 32612 6456 32668
rect 6392 32608 6456 32612
rect 7752 32668 7816 32672
rect 7752 32612 7756 32668
rect 7756 32612 7812 32668
rect 7812 32612 7816 32668
rect 7752 32608 7816 32612
rect 7832 32668 7896 32672
rect 7832 32612 7836 32668
rect 7836 32612 7892 32668
rect 7892 32612 7896 32668
rect 7832 32608 7896 32612
rect 7912 32668 7976 32672
rect 7912 32612 7916 32668
rect 7916 32612 7972 32668
rect 7972 32612 7976 32668
rect 7912 32608 7976 32612
rect 7992 32668 8056 32672
rect 7992 32612 7996 32668
rect 7996 32612 8052 32668
rect 8052 32612 8056 32668
rect 7992 32608 8056 32612
rect 9352 32668 9416 32672
rect 9352 32612 9356 32668
rect 9356 32612 9412 32668
rect 9412 32612 9416 32668
rect 9352 32608 9416 32612
rect 9432 32668 9496 32672
rect 9432 32612 9436 32668
rect 9436 32612 9492 32668
rect 9492 32612 9496 32668
rect 9432 32608 9496 32612
rect 9512 32668 9576 32672
rect 9512 32612 9516 32668
rect 9516 32612 9572 32668
rect 9572 32612 9576 32668
rect 9512 32608 9576 32612
rect 9592 32668 9656 32672
rect 9592 32612 9596 32668
rect 9596 32612 9652 32668
rect 9652 32612 9656 32668
rect 9592 32608 9656 32612
rect 3612 32124 3676 32128
rect 3612 32068 3616 32124
rect 3616 32068 3672 32124
rect 3672 32068 3676 32124
rect 3612 32064 3676 32068
rect 3692 32124 3756 32128
rect 3692 32068 3696 32124
rect 3696 32068 3752 32124
rect 3752 32068 3756 32124
rect 3692 32064 3756 32068
rect 3772 32124 3836 32128
rect 3772 32068 3776 32124
rect 3776 32068 3832 32124
rect 3832 32068 3836 32124
rect 3772 32064 3836 32068
rect 3852 32124 3916 32128
rect 3852 32068 3856 32124
rect 3856 32068 3912 32124
rect 3912 32068 3916 32124
rect 3852 32064 3916 32068
rect 5212 32124 5276 32128
rect 5212 32068 5216 32124
rect 5216 32068 5272 32124
rect 5272 32068 5276 32124
rect 5212 32064 5276 32068
rect 5292 32124 5356 32128
rect 5292 32068 5296 32124
rect 5296 32068 5352 32124
rect 5352 32068 5356 32124
rect 5292 32064 5356 32068
rect 5372 32124 5436 32128
rect 5372 32068 5376 32124
rect 5376 32068 5432 32124
rect 5432 32068 5436 32124
rect 5372 32064 5436 32068
rect 5452 32124 5516 32128
rect 5452 32068 5456 32124
rect 5456 32068 5512 32124
rect 5512 32068 5516 32124
rect 5452 32064 5516 32068
rect 6812 32124 6876 32128
rect 6812 32068 6816 32124
rect 6816 32068 6872 32124
rect 6872 32068 6876 32124
rect 6812 32064 6876 32068
rect 6892 32124 6956 32128
rect 6892 32068 6896 32124
rect 6896 32068 6952 32124
rect 6952 32068 6956 32124
rect 6892 32064 6956 32068
rect 6972 32124 7036 32128
rect 6972 32068 6976 32124
rect 6976 32068 7032 32124
rect 7032 32068 7036 32124
rect 6972 32064 7036 32068
rect 7052 32124 7116 32128
rect 7052 32068 7056 32124
rect 7056 32068 7112 32124
rect 7112 32068 7116 32124
rect 7052 32064 7116 32068
rect 8412 32124 8476 32128
rect 8412 32068 8416 32124
rect 8416 32068 8472 32124
rect 8472 32068 8476 32124
rect 8412 32064 8476 32068
rect 8492 32124 8556 32128
rect 8492 32068 8496 32124
rect 8496 32068 8552 32124
rect 8552 32068 8556 32124
rect 8492 32064 8556 32068
rect 8572 32124 8636 32128
rect 8572 32068 8576 32124
rect 8576 32068 8632 32124
rect 8632 32068 8636 32124
rect 8572 32064 8636 32068
rect 8652 32124 8716 32128
rect 8652 32068 8656 32124
rect 8656 32068 8712 32124
rect 8712 32068 8716 32124
rect 8652 32064 8716 32068
rect 2952 31580 3016 31584
rect 2952 31524 2956 31580
rect 2956 31524 3012 31580
rect 3012 31524 3016 31580
rect 2952 31520 3016 31524
rect 3032 31580 3096 31584
rect 3032 31524 3036 31580
rect 3036 31524 3092 31580
rect 3092 31524 3096 31580
rect 3032 31520 3096 31524
rect 3112 31580 3176 31584
rect 3112 31524 3116 31580
rect 3116 31524 3172 31580
rect 3172 31524 3176 31580
rect 3112 31520 3176 31524
rect 3192 31580 3256 31584
rect 3192 31524 3196 31580
rect 3196 31524 3252 31580
rect 3252 31524 3256 31580
rect 3192 31520 3256 31524
rect 4552 31580 4616 31584
rect 4552 31524 4556 31580
rect 4556 31524 4612 31580
rect 4612 31524 4616 31580
rect 4552 31520 4616 31524
rect 4632 31580 4696 31584
rect 4632 31524 4636 31580
rect 4636 31524 4692 31580
rect 4692 31524 4696 31580
rect 4632 31520 4696 31524
rect 4712 31580 4776 31584
rect 4712 31524 4716 31580
rect 4716 31524 4772 31580
rect 4772 31524 4776 31580
rect 4712 31520 4776 31524
rect 4792 31580 4856 31584
rect 4792 31524 4796 31580
rect 4796 31524 4852 31580
rect 4852 31524 4856 31580
rect 4792 31520 4856 31524
rect 6152 31580 6216 31584
rect 6152 31524 6156 31580
rect 6156 31524 6212 31580
rect 6212 31524 6216 31580
rect 6152 31520 6216 31524
rect 6232 31580 6296 31584
rect 6232 31524 6236 31580
rect 6236 31524 6292 31580
rect 6292 31524 6296 31580
rect 6232 31520 6296 31524
rect 6312 31580 6376 31584
rect 6312 31524 6316 31580
rect 6316 31524 6372 31580
rect 6372 31524 6376 31580
rect 6312 31520 6376 31524
rect 6392 31580 6456 31584
rect 6392 31524 6396 31580
rect 6396 31524 6452 31580
rect 6452 31524 6456 31580
rect 6392 31520 6456 31524
rect 7752 31580 7816 31584
rect 7752 31524 7756 31580
rect 7756 31524 7812 31580
rect 7812 31524 7816 31580
rect 7752 31520 7816 31524
rect 7832 31580 7896 31584
rect 7832 31524 7836 31580
rect 7836 31524 7892 31580
rect 7892 31524 7896 31580
rect 7832 31520 7896 31524
rect 7912 31580 7976 31584
rect 7912 31524 7916 31580
rect 7916 31524 7972 31580
rect 7972 31524 7976 31580
rect 7912 31520 7976 31524
rect 7992 31580 8056 31584
rect 7992 31524 7996 31580
rect 7996 31524 8052 31580
rect 8052 31524 8056 31580
rect 7992 31520 8056 31524
rect 9352 31580 9416 31584
rect 9352 31524 9356 31580
rect 9356 31524 9412 31580
rect 9412 31524 9416 31580
rect 9352 31520 9416 31524
rect 9432 31580 9496 31584
rect 9432 31524 9436 31580
rect 9436 31524 9492 31580
rect 9492 31524 9496 31580
rect 9432 31520 9496 31524
rect 9512 31580 9576 31584
rect 9512 31524 9516 31580
rect 9516 31524 9572 31580
rect 9572 31524 9576 31580
rect 9512 31520 9576 31524
rect 9592 31580 9656 31584
rect 9592 31524 9596 31580
rect 9596 31524 9652 31580
rect 9652 31524 9656 31580
rect 9592 31520 9656 31524
rect 3612 31036 3676 31040
rect 3612 30980 3616 31036
rect 3616 30980 3672 31036
rect 3672 30980 3676 31036
rect 3612 30976 3676 30980
rect 3692 31036 3756 31040
rect 3692 30980 3696 31036
rect 3696 30980 3752 31036
rect 3752 30980 3756 31036
rect 3692 30976 3756 30980
rect 3772 31036 3836 31040
rect 3772 30980 3776 31036
rect 3776 30980 3832 31036
rect 3832 30980 3836 31036
rect 3772 30976 3836 30980
rect 3852 31036 3916 31040
rect 3852 30980 3856 31036
rect 3856 30980 3912 31036
rect 3912 30980 3916 31036
rect 3852 30976 3916 30980
rect 5212 31036 5276 31040
rect 5212 30980 5216 31036
rect 5216 30980 5272 31036
rect 5272 30980 5276 31036
rect 5212 30976 5276 30980
rect 5292 31036 5356 31040
rect 5292 30980 5296 31036
rect 5296 30980 5352 31036
rect 5352 30980 5356 31036
rect 5292 30976 5356 30980
rect 5372 31036 5436 31040
rect 5372 30980 5376 31036
rect 5376 30980 5432 31036
rect 5432 30980 5436 31036
rect 5372 30976 5436 30980
rect 5452 31036 5516 31040
rect 5452 30980 5456 31036
rect 5456 30980 5512 31036
rect 5512 30980 5516 31036
rect 5452 30976 5516 30980
rect 6812 31036 6876 31040
rect 6812 30980 6816 31036
rect 6816 30980 6872 31036
rect 6872 30980 6876 31036
rect 6812 30976 6876 30980
rect 6892 31036 6956 31040
rect 6892 30980 6896 31036
rect 6896 30980 6952 31036
rect 6952 30980 6956 31036
rect 6892 30976 6956 30980
rect 6972 31036 7036 31040
rect 6972 30980 6976 31036
rect 6976 30980 7032 31036
rect 7032 30980 7036 31036
rect 6972 30976 7036 30980
rect 7052 31036 7116 31040
rect 7052 30980 7056 31036
rect 7056 30980 7112 31036
rect 7112 30980 7116 31036
rect 7052 30976 7116 30980
rect 8412 31036 8476 31040
rect 8412 30980 8416 31036
rect 8416 30980 8472 31036
rect 8472 30980 8476 31036
rect 8412 30976 8476 30980
rect 8492 31036 8556 31040
rect 8492 30980 8496 31036
rect 8496 30980 8552 31036
rect 8552 30980 8556 31036
rect 8492 30976 8556 30980
rect 8572 31036 8636 31040
rect 8572 30980 8576 31036
rect 8576 30980 8632 31036
rect 8632 30980 8636 31036
rect 8572 30976 8636 30980
rect 8652 31036 8716 31040
rect 8652 30980 8656 31036
rect 8656 30980 8712 31036
rect 8712 30980 8716 31036
rect 8652 30976 8716 30980
rect 2952 30492 3016 30496
rect 2952 30436 2956 30492
rect 2956 30436 3012 30492
rect 3012 30436 3016 30492
rect 2952 30432 3016 30436
rect 3032 30492 3096 30496
rect 3032 30436 3036 30492
rect 3036 30436 3092 30492
rect 3092 30436 3096 30492
rect 3032 30432 3096 30436
rect 3112 30492 3176 30496
rect 3112 30436 3116 30492
rect 3116 30436 3172 30492
rect 3172 30436 3176 30492
rect 3112 30432 3176 30436
rect 3192 30492 3256 30496
rect 3192 30436 3196 30492
rect 3196 30436 3252 30492
rect 3252 30436 3256 30492
rect 3192 30432 3256 30436
rect 4552 30492 4616 30496
rect 4552 30436 4556 30492
rect 4556 30436 4612 30492
rect 4612 30436 4616 30492
rect 4552 30432 4616 30436
rect 4632 30492 4696 30496
rect 4632 30436 4636 30492
rect 4636 30436 4692 30492
rect 4692 30436 4696 30492
rect 4632 30432 4696 30436
rect 4712 30492 4776 30496
rect 4712 30436 4716 30492
rect 4716 30436 4772 30492
rect 4772 30436 4776 30492
rect 4712 30432 4776 30436
rect 4792 30492 4856 30496
rect 4792 30436 4796 30492
rect 4796 30436 4852 30492
rect 4852 30436 4856 30492
rect 4792 30432 4856 30436
rect 3612 29948 3676 29952
rect 3612 29892 3616 29948
rect 3616 29892 3672 29948
rect 3672 29892 3676 29948
rect 3612 29888 3676 29892
rect 3692 29948 3756 29952
rect 3692 29892 3696 29948
rect 3696 29892 3752 29948
rect 3752 29892 3756 29948
rect 3692 29888 3756 29892
rect 3772 29948 3836 29952
rect 3772 29892 3776 29948
rect 3776 29892 3832 29948
rect 3832 29892 3836 29948
rect 3772 29888 3836 29892
rect 3852 29948 3916 29952
rect 3852 29892 3856 29948
rect 3856 29892 3912 29948
rect 3912 29892 3916 29948
rect 3852 29888 3916 29892
rect 5212 29948 5276 29952
rect 5212 29892 5216 29948
rect 5216 29892 5272 29948
rect 5272 29892 5276 29948
rect 5212 29888 5276 29892
rect 5292 29948 5356 29952
rect 5292 29892 5296 29948
rect 5296 29892 5352 29948
rect 5352 29892 5356 29948
rect 5292 29888 5356 29892
rect 5372 29948 5436 29952
rect 5372 29892 5376 29948
rect 5376 29892 5432 29948
rect 5432 29892 5436 29948
rect 5372 29888 5436 29892
rect 5452 29948 5516 29952
rect 5452 29892 5456 29948
rect 5456 29892 5512 29948
rect 5512 29892 5516 29948
rect 5452 29888 5516 29892
rect 2952 29404 3016 29408
rect 2952 29348 2956 29404
rect 2956 29348 3012 29404
rect 3012 29348 3016 29404
rect 2952 29344 3016 29348
rect 3032 29404 3096 29408
rect 3032 29348 3036 29404
rect 3036 29348 3092 29404
rect 3092 29348 3096 29404
rect 3032 29344 3096 29348
rect 3112 29404 3176 29408
rect 3112 29348 3116 29404
rect 3116 29348 3172 29404
rect 3172 29348 3176 29404
rect 3112 29344 3176 29348
rect 3192 29404 3256 29408
rect 3192 29348 3196 29404
rect 3196 29348 3252 29404
rect 3252 29348 3256 29404
rect 3192 29344 3256 29348
rect 4552 29404 4616 29408
rect 4552 29348 4556 29404
rect 4556 29348 4612 29404
rect 4612 29348 4616 29404
rect 4552 29344 4616 29348
rect 4632 29404 4696 29408
rect 4632 29348 4636 29404
rect 4636 29348 4692 29404
rect 4692 29348 4696 29404
rect 4632 29344 4696 29348
rect 4712 29404 4776 29408
rect 4712 29348 4716 29404
rect 4716 29348 4772 29404
rect 4772 29348 4776 29404
rect 4712 29344 4776 29348
rect 4792 29404 4856 29408
rect 4792 29348 4796 29404
rect 4796 29348 4852 29404
rect 4852 29348 4856 29404
rect 4792 29344 4856 29348
rect 6152 30492 6216 30496
rect 6152 30436 6156 30492
rect 6156 30436 6212 30492
rect 6212 30436 6216 30492
rect 6152 30432 6216 30436
rect 6232 30492 6296 30496
rect 6232 30436 6236 30492
rect 6236 30436 6292 30492
rect 6292 30436 6296 30492
rect 6232 30432 6296 30436
rect 6312 30492 6376 30496
rect 6312 30436 6316 30492
rect 6316 30436 6372 30492
rect 6372 30436 6376 30492
rect 6312 30432 6376 30436
rect 6392 30492 6456 30496
rect 6392 30436 6396 30492
rect 6396 30436 6452 30492
rect 6452 30436 6456 30492
rect 6392 30432 6456 30436
rect 7752 30492 7816 30496
rect 7752 30436 7756 30492
rect 7756 30436 7812 30492
rect 7812 30436 7816 30492
rect 7752 30432 7816 30436
rect 7832 30492 7896 30496
rect 7832 30436 7836 30492
rect 7836 30436 7892 30492
rect 7892 30436 7896 30492
rect 7832 30432 7896 30436
rect 7912 30492 7976 30496
rect 7912 30436 7916 30492
rect 7916 30436 7972 30492
rect 7972 30436 7976 30492
rect 7912 30432 7976 30436
rect 7992 30492 8056 30496
rect 7992 30436 7996 30492
rect 7996 30436 8052 30492
rect 8052 30436 8056 30492
rect 7992 30432 8056 30436
rect 9352 30492 9416 30496
rect 9352 30436 9356 30492
rect 9356 30436 9412 30492
rect 9412 30436 9416 30492
rect 9352 30432 9416 30436
rect 9432 30492 9496 30496
rect 9432 30436 9436 30492
rect 9436 30436 9492 30492
rect 9492 30436 9496 30492
rect 9432 30432 9496 30436
rect 9512 30492 9576 30496
rect 9512 30436 9516 30492
rect 9516 30436 9572 30492
rect 9572 30436 9576 30492
rect 9512 30432 9576 30436
rect 9592 30492 9656 30496
rect 9592 30436 9596 30492
rect 9596 30436 9652 30492
rect 9652 30436 9656 30492
rect 9592 30432 9656 30436
rect 6812 29948 6876 29952
rect 6812 29892 6816 29948
rect 6816 29892 6872 29948
rect 6872 29892 6876 29948
rect 6812 29888 6876 29892
rect 6892 29948 6956 29952
rect 6892 29892 6896 29948
rect 6896 29892 6952 29948
rect 6952 29892 6956 29948
rect 6892 29888 6956 29892
rect 6972 29948 7036 29952
rect 6972 29892 6976 29948
rect 6976 29892 7032 29948
rect 7032 29892 7036 29948
rect 6972 29888 7036 29892
rect 7052 29948 7116 29952
rect 7052 29892 7056 29948
rect 7056 29892 7112 29948
rect 7112 29892 7116 29948
rect 7052 29888 7116 29892
rect 8412 29948 8476 29952
rect 8412 29892 8416 29948
rect 8416 29892 8472 29948
rect 8472 29892 8476 29948
rect 8412 29888 8476 29892
rect 8492 29948 8556 29952
rect 8492 29892 8496 29948
rect 8496 29892 8552 29948
rect 8552 29892 8556 29948
rect 8492 29888 8556 29892
rect 8572 29948 8636 29952
rect 8572 29892 8576 29948
rect 8576 29892 8632 29948
rect 8632 29892 8636 29948
rect 8572 29888 8636 29892
rect 8652 29948 8716 29952
rect 8652 29892 8656 29948
rect 8656 29892 8712 29948
rect 8712 29892 8716 29948
rect 8652 29888 8716 29892
rect 6152 29404 6216 29408
rect 6152 29348 6156 29404
rect 6156 29348 6212 29404
rect 6212 29348 6216 29404
rect 6152 29344 6216 29348
rect 6232 29404 6296 29408
rect 6232 29348 6236 29404
rect 6236 29348 6292 29404
rect 6292 29348 6296 29404
rect 6232 29344 6296 29348
rect 6312 29404 6376 29408
rect 6312 29348 6316 29404
rect 6316 29348 6372 29404
rect 6372 29348 6376 29404
rect 6312 29344 6376 29348
rect 6392 29404 6456 29408
rect 6392 29348 6396 29404
rect 6396 29348 6452 29404
rect 6452 29348 6456 29404
rect 6392 29344 6456 29348
rect 7752 29404 7816 29408
rect 7752 29348 7756 29404
rect 7756 29348 7812 29404
rect 7812 29348 7816 29404
rect 7752 29344 7816 29348
rect 7832 29404 7896 29408
rect 7832 29348 7836 29404
rect 7836 29348 7892 29404
rect 7892 29348 7896 29404
rect 7832 29344 7896 29348
rect 7912 29404 7976 29408
rect 7912 29348 7916 29404
rect 7916 29348 7972 29404
rect 7972 29348 7976 29404
rect 7912 29344 7976 29348
rect 7992 29404 8056 29408
rect 7992 29348 7996 29404
rect 7996 29348 8052 29404
rect 8052 29348 8056 29404
rect 7992 29344 8056 29348
rect 9352 29404 9416 29408
rect 9352 29348 9356 29404
rect 9356 29348 9412 29404
rect 9412 29348 9416 29404
rect 9352 29344 9416 29348
rect 9432 29404 9496 29408
rect 9432 29348 9436 29404
rect 9436 29348 9492 29404
rect 9492 29348 9496 29404
rect 9432 29344 9496 29348
rect 9512 29404 9576 29408
rect 9512 29348 9516 29404
rect 9516 29348 9572 29404
rect 9572 29348 9576 29404
rect 9512 29344 9576 29348
rect 9592 29404 9656 29408
rect 9592 29348 9596 29404
rect 9596 29348 9652 29404
rect 9652 29348 9656 29404
rect 9592 29344 9656 29348
rect 3612 28860 3676 28864
rect 3612 28804 3616 28860
rect 3616 28804 3672 28860
rect 3672 28804 3676 28860
rect 3612 28800 3676 28804
rect 3692 28860 3756 28864
rect 3692 28804 3696 28860
rect 3696 28804 3752 28860
rect 3752 28804 3756 28860
rect 3692 28800 3756 28804
rect 3772 28860 3836 28864
rect 3772 28804 3776 28860
rect 3776 28804 3832 28860
rect 3832 28804 3836 28860
rect 3772 28800 3836 28804
rect 3852 28860 3916 28864
rect 3852 28804 3856 28860
rect 3856 28804 3912 28860
rect 3912 28804 3916 28860
rect 3852 28800 3916 28804
rect 5212 28860 5276 28864
rect 5212 28804 5216 28860
rect 5216 28804 5272 28860
rect 5272 28804 5276 28860
rect 5212 28800 5276 28804
rect 5292 28860 5356 28864
rect 5292 28804 5296 28860
rect 5296 28804 5352 28860
rect 5352 28804 5356 28860
rect 5292 28800 5356 28804
rect 5372 28860 5436 28864
rect 5372 28804 5376 28860
rect 5376 28804 5432 28860
rect 5432 28804 5436 28860
rect 5372 28800 5436 28804
rect 5452 28860 5516 28864
rect 5452 28804 5456 28860
rect 5456 28804 5512 28860
rect 5512 28804 5516 28860
rect 5452 28800 5516 28804
rect 6812 28860 6876 28864
rect 6812 28804 6816 28860
rect 6816 28804 6872 28860
rect 6872 28804 6876 28860
rect 6812 28800 6876 28804
rect 6892 28860 6956 28864
rect 6892 28804 6896 28860
rect 6896 28804 6952 28860
rect 6952 28804 6956 28860
rect 6892 28800 6956 28804
rect 6972 28860 7036 28864
rect 6972 28804 6976 28860
rect 6976 28804 7032 28860
rect 7032 28804 7036 28860
rect 6972 28800 7036 28804
rect 7052 28860 7116 28864
rect 7052 28804 7056 28860
rect 7056 28804 7112 28860
rect 7112 28804 7116 28860
rect 7052 28800 7116 28804
rect 8412 28860 8476 28864
rect 8412 28804 8416 28860
rect 8416 28804 8472 28860
rect 8472 28804 8476 28860
rect 8412 28800 8476 28804
rect 8492 28860 8556 28864
rect 8492 28804 8496 28860
rect 8496 28804 8552 28860
rect 8552 28804 8556 28860
rect 8492 28800 8556 28804
rect 8572 28860 8636 28864
rect 8572 28804 8576 28860
rect 8576 28804 8632 28860
rect 8632 28804 8636 28860
rect 8572 28800 8636 28804
rect 8652 28860 8716 28864
rect 8652 28804 8656 28860
rect 8656 28804 8712 28860
rect 8712 28804 8716 28860
rect 8652 28800 8716 28804
rect 2952 28316 3016 28320
rect 2952 28260 2956 28316
rect 2956 28260 3012 28316
rect 3012 28260 3016 28316
rect 2952 28256 3016 28260
rect 3032 28316 3096 28320
rect 3032 28260 3036 28316
rect 3036 28260 3092 28316
rect 3092 28260 3096 28316
rect 3032 28256 3096 28260
rect 3112 28316 3176 28320
rect 3112 28260 3116 28316
rect 3116 28260 3172 28316
rect 3172 28260 3176 28316
rect 3112 28256 3176 28260
rect 3192 28316 3256 28320
rect 3192 28260 3196 28316
rect 3196 28260 3252 28316
rect 3252 28260 3256 28316
rect 3192 28256 3256 28260
rect 4552 28316 4616 28320
rect 4552 28260 4556 28316
rect 4556 28260 4612 28316
rect 4612 28260 4616 28316
rect 4552 28256 4616 28260
rect 4632 28316 4696 28320
rect 4632 28260 4636 28316
rect 4636 28260 4692 28316
rect 4692 28260 4696 28316
rect 4632 28256 4696 28260
rect 4712 28316 4776 28320
rect 4712 28260 4716 28316
rect 4716 28260 4772 28316
rect 4772 28260 4776 28316
rect 4712 28256 4776 28260
rect 4792 28316 4856 28320
rect 4792 28260 4796 28316
rect 4796 28260 4852 28316
rect 4852 28260 4856 28316
rect 4792 28256 4856 28260
rect 6152 28316 6216 28320
rect 6152 28260 6156 28316
rect 6156 28260 6212 28316
rect 6212 28260 6216 28316
rect 6152 28256 6216 28260
rect 6232 28316 6296 28320
rect 6232 28260 6236 28316
rect 6236 28260 6292 28316
rect 6292 28260 6296 28316
rect 6232 28256 6296 28260
rect 6312 28316 6376 28320
rect 6312 28260 6316 28316
rect 6316 28260 6372 28316
rect 6372 28260 6376 28316
rect 6312 28256 6376 28260
rect 6392 28316 6456 28320
rect 6392 28260 6396 28316
rect 6396 28260 6452 28316
rect 6452 28260 6456 28316
rect 6392 28256 6456 28260
rect 7752 28316 7816 28320
rect 7752 28260 7756 28316
rect 7756 28260 7812 28316
rect 7812 28260 7816 28316
rect 7752 28256 7816 28260
rect 7832 28316 7896 28320
rect 7832 28260 7836 28316
rect 7836 28260 7892 28316
rect 7892 28260 7896 28316
rect 7832 28256 7896 28260
rect 7912 28316 7976 28320
rect 7912 28260 7916 28316
rect 7916 28260 7972 28316
rect 7972 28260 7976 28316
rect 7912 28256 7976 28260
rect 7992 28316 8056 28320
rect 7992 28260 7996 28316
rect 7996 28260 8052 28316
rect 8052 28260 8056 28316
rect 7992 28256 8056 28260
rect 9352 28316 9416 28320
rect 9352 28260 9356 28316
rect 9356 28260 9412 28316
rect 9412 28260 9416 28316
rect 9352 28256 9416 28260
rect 9432 28316 9496 28320
rect 9432 28260 9436 28316
rect 9436 28260 9492 28316
rect 9492 28260 9496 28316
rect 9432 28256 9496 28260
rect 9512 28316 9576 28320
rect 9512 28260 9516 28316
rect 9516 28260 9572 28316
rect 9572 28260 9576 28316
rect 9512 28256 9576 28260
rect 9592 28316 9656 28320
rect 9592 28260 9596 28316
rect 9596 28260 9652 28316
rect 9652 28260 9656 28316
rect 9592 28256 9656 28260
rect 3612 27772 3676 27776
rect 3612 27716 3616 27772
rect 3616 27716 3672 27772
rect 3672 27716 3676 27772
rect 3612 27712 3676 27716
rect 3692 27772 3756 27776
rect 3692 27716 3696 27772
rect 3696 27716 3752 27772
rect 3752 27716 3756 27772
rect 3692 27712 3756 27716
rect 3772 27772 3836 27776
rect 3772 27716 3776 27772
rect 3776 27716 3832 27772
rect 3832 27716 3836 27772
rect 3772 27712 3836 27716
rect 3852 27772 3916 27776
rect 3852 27716 3856 27772
rect 3856 27716 3912 27772
rect 3912 27716 3916 27772
rect 3852 27712 3916 27716
rect 5212 27772 5276 27776
rect 5212 27716 5216 27772
rect 5216 27716 5272 27772
rect 5272 27716 5276 27772
rect 5212 27712 5276 27716
rect 5292 27772 5356 27776
rect 5292 27716 5296 27772
rect 5296 27716 5352 27772
rect 5352 27716 5356 27772
rect 5292 27712 5356 27716
rect 5372 27772 5436 27776
rect 5372 27716 5376 27772
rect 5376 27716 5432 27772
rect 5432 27716 5436 27772
rect 5372 27712 5436 27716
rect 5452 27772 5516 27776
rect 5452 27716 5456 27772
rect 5456 27716 5512 27772
rect 5512 27716 5516 27772
rect 5452 27712 5516 27716
rect 6812 27772 6876 27776
rect 6812 27716 6816 27772
rect 6816 27716 6872 27772
rect 6872 27716 6876 27772
rect 6812 27712 6876 27716
rect 6892 27772 6956 27776
rect 6892 27716 6896 27772
rect 6896 27716 6952 27772
rect 6952 27716 6956 27772
rect 6892 27712 6956 27716
rect 6972 27772 7036 27776
rect 6972 27716 6976 27772
rect 6976 27716 7032 27772
rect 7032 27716 7036 27772
rect 6972 27712 7036 27716
rect 7052 27772 7116 27776
rect 7052 27716 7056 27772
rect 7056 27716 7112 27772
rect 7112 27716 7116 27772
rect 7052 27712 7116 27716
rect 8412 27772 8476 27776
rect 8412 27716 8416 27772
rect 8416 27716 8472 27772
rect 8472 27716 8476 27772
rect 8412 27712 8476 27716
rect 8492 27772 8556 27776
rect 8492 27716 8496 27772
rect 8496 27716 8552 27772
rect 8552 27716 8556 27772
rect 8492 27712 8556 27716
rect 8572 27772 8636 27776
rect 8572 27716 8576 27772
rect 8576 27716 8632 27772
rect 8632 27716 8636 27772
rect 8572 27712 8636 27716
rect 8652 27772 8716 27776
rect 8652 27716 8656 27772
rect 8656 27716 8712 27772
rect 8712 27716 8716 27772
rect 8652 27712 8716 27716
rect 2952 27228 3016 27232
rect 2952 27172 2956 27228
rect 2956 27172 3012 27228
rect 3012 27172 3016 27228
rect 2952 27168 3016 27172
rect 3032 27228 3096 27232
rect 3032 27172 3036 27228
rect 3036 27172 3092 27228
rect 3092 27172 3096 27228
rect 3032 27168 3096 27172
rect 3112 27228 3176 27232
rect 3112 27172 3116 27228
rect 3116 27172 3172 27228
rect 3172 27172 3176 27228
rect 3112 27168 3176 27172
rect 3192 27228 3256 27232
rect 3192 27172 3196 27228
rect 3196 27172 3252 27228
rect 3252 27172 3256 27228
rect 3192 27168 3256 27172
rect 4552 27228 4616 27232
rect 4552 27172 4556 27228
rect 4556 27172 4612 27228
rect 4612 27172 4616 27228
rect 4552 27168 4616 27172
rect 4632 27228 4696 27232
rect 4632 27172 4636 27228
rect 4636 27172 4692 27228
rect 4692 27172 4696 27228
rect 4632 27168 4696 27172
rect 4712 27228 4776 27232
rect 4712 27172 4716 27228
rect 4716 27172 4772 27228
rect 4772 27172 4776 27228
rect 4712 27168 4776 27172
rect 4792 27228 4856 27232
rect 4792 27172 4796 27228
rect 4796 27172 4852 27228
rect 4852 27172 4856 27228
rect 4792 27168 4856 27172
rect 6152 27228 6216 27232
rect 6152 27172 6156 27228
rect 6156 27172 6212 27228
rect 6212 27172 6216 27228
rect 6152 27168 6216 27172
rect 6232 27228 6296 27232
rect 6232 27172 6236 27228
rect 6236 27172 6292 27228
rect 6292 27172 6296 27228
rect 6232 27168 6296 27172
rect 6312 27228 6376 27232
rect 6312 27172 6316 27228
rect 6316 27172 6372 27228
rect 6372 27172 6376 27228
rect 6312 27168 6376 27172
rect 6392 27228 6456 27232
rect 6392 27172 6396 27228
rect 6396 27172 6452 27228
rect 6452 27172 6456 27228
rect 6392 27168 6456 27172
rect 7752 27228 7816 27232
rect 7752 27172 7756 27228
rect 7756 27172 7812 27228
rect 7812 27172 7816 27228
rect 7752 27168 7816 27172
rect 7832 27228 7896 27232
rect 7832 27172 7836 27228
rect 7836 27172 7892 27228
rect 7892 27172 7896 27228
rect 7832 27168 7896 27172
rect 7912 27228 7976 27232
rect 7912 27172 7916 27228
rect 7916 27172 7972 27228
rect 7972 27172 7976 27228
rect 7912 27168 7976 27172
rect 7992 27228 8056 27232
rect 7992 27172 7996 27228
rect 7996 27172 8052 27228
rect 8052 27172 8056 27228
rect 7992 27168 8056 27172
rect 9352 27228 9416 27232
rect 9352 27172 9356 27228
rect 9356 27172 9412 27228
rect 9412 27172 9416 27228
rect 9352 27168 9416 27172
rect 9432 27228 9496 27232
rect 9432 27172 9436 27228
rect 9436 27172 9492 27228
rect 9492 27172 9496 27228
rect 9432 27168 9496 27172
rect 9512 27228 9576 27232
rect 9512 27172 9516 27228
rect 9516 27172 9572 27228
rect 9572 27172 9576 27228
rect 9512 27168 9576 27172
rect 9592 27228 9656 27232
rect 9592 27172 9596 27228
rect 9596 27172 9652 27228
rect 9652 27172 9656 27228
rect 9592 27168 9656 27172
rect 3612 26684 3676 26688
rect 3612 26628 3616 26684
rect 3616 26628 3672 26684
rect 3672 26628 3676 26684
rect 3612 26624 3676 26628
rect 3692 26684 3756 26688
rect 3692 26628 3696 26684
rect 3696 26628 3752 26684
rect 3752 26628 3756 26684
rect 3692 26624 3756 26628
rect 3772 26684 3836 26688
rect 3772 26628 3776 26684
rect 3776 26628 3832 26684
rect 3832 26628 3836 26684
rect 3772 26624 3836 26628
rect 3852 26684 3916 26688
rect 3852 26628 3856 26684
rect 3856 26628 3912 26684
rect 3912 26628 3916 26684
rect 3852 26624 3916 26628
rect 5212 26684 5276 26688
rect 5212 26628 5216 26684
rect 5216 26628 5272 26684
rect 5272 26628 5276 26684
rect 5212 26624 5276 26628
rect 5292 26684 5356 26688
rect 5292 26628 5296 26684
rect 5296 26628 5352 26684
rect 5352 26628 5356 26684
rect 5292 26624 5356 26628
rect 5372 26684 5436 26688
rect 5372 26628 5376 26684
rect 5376 26628 5432 26684
rect 5432 26628 5436 26684
rect 5372 26624 5436 26628
rect 5452 26684 5516 26688
rect 5452 26628 5456 26684
rect 5456 26628 5512 26684
rect 5512 26628 5516 26684
rect 5452 26624 5516 26628
rect 6812 26684 6876 26688
rect 6812 26628 6816 26684
rect 6816 26628 6872 26684
rect 6872 26628 6876 26684
rect 6812 26624 6876 26628
rect 6892 26684 6956 26688
rect 6892 26628 6896 26684
rect 6896 26628 6952 26684
rect 6952 26628 6956 26684
rect 6892 26624 6956 26628
rect 6972 26684 7036 26688
rect 6972 26628 6976 26684
rect 6976 26628 7032 26684
rect 7032 26628 7036 26684
rect 6972 26624 7036 26628
rect 7052 26684 7116 26688
rect 7052 26628 7056 26684
rect 7056 26628 7112 26684
rect 7112 26628 7116 26684
rect 7052 26624 7116 26628
rect 8412 26684 8476 26688
rect 8412 26628 8416 26684
rect 8416 26628 8472 26684
rect 8472 26628 8476 26684
rect 8412 26624 8476 26628
rect 8492 26684 8556 26688
rect 8492 26628 8496 26684
rect 8496 26628 8552 26684
rect 8552 26628 8556 26684
rect 8492 26624 8556 26628
rect 8572 26684 8636 26688
rect 8572 26628 8576 26684
rect 8576 26628 8632 26684
rect 8632 26628 8636 26684
rect 8572 26624 8636 26628
rect 8652 26684 8716 26688
rect 8652 26628 8656 26684
rect 8656 26628 8712 26684
rect 8712 26628 8716 26684
rect 8652 26624 8716 26628
rect 2952 26140 3016 26144
rect 2952 26084 2956 26140
rect 2956 26084 3012 26140
rect 3012 26084 3016 26140
rect 2952 26080 3016 26084
rect 3032 26140 3096 26144
rect 3032 26084 3036 26140
rect 3036 26084 3092 26140
rect 3092 26084 3096 26140
rect 3032 26080 3096 26084
rect 3112 26140 3176 26144
rect 3112 26084 3116 26140
rect 3116 26084 3172 26140
rect 3172 26084 3176 26140
rect 3112 26080 3176 26084
rect 3192 26140 3256 26144
rect 3192 26084 3196 26140
rect 3196 26084 3252 26140
rect 3252 26084 3256 26140
rect 3192 26080 3256 26084
rect 4552 26140 4616 26144
rect 4552 26084 4556 26140
rect 4556 26084 4612 26140
rect 4612 26084 4616 26140
rect 4552 26080 4616 26084
rect 4632 26140 4696 26144
rect 4632 26084 4636 26140
rect 4636 26084 4692 26140
rect 4692 26084 4696 26140
rect 4632 26080 4696 26084
rect 4712 26140 4776 26144
rect 4712 26084 4716 26140
rect 4716 26084 4772 26140
rect 4772 26084 4776 26140
rect 4712 26080 4776 26084
rect 4792 26140 4856 26144
rect 4792 26084 4796 26140
rect 4796 26084 4852 26140
rect 4852 26084 4856 26140
rect 4792 26080 4856 26084
rect 6152 26140 6216 26144
rect 6152 26084 6156 26140
rect 6156 26084 6212 26140
rect 6212 26084 6216 26140
rect 6152 26080 6216 26084
rect 6232 26140 6296 26144
rect 6232 26084 6236 26140
rect 6236 26084 6292 26140
rect 6292 26084 6296 26140
rect 6232 26080 6296 26084
rect 6312 26140 6376 26144
rect 6312 26084 6316 26140
rect 6316 26084 6372 26140
rect 6372 26084 6376 26140
rect 6312 26080 6376 26084
rect 6392 26140 6456 26144
rect 6392 26084 6396 26140
rect 6396 26084 6452 26140
rect 6452 26084 6456 26140
rect 6392 26080 6456 26084
rect 7752 26140 7816 26144
rect 7752 26084 7756 26140
rect 7756 26084 7812 26140
rect 7812 26084 7816 26140
rect 7752 26080 7816 26084
rect 7832 26140 7896 26144
rect 7832 26084 7836 26140
rect 7836 26084 7892 26140
rect 7892 26084 7896 26140
rect 7832 26080 7896 26084
rect 7912 26140 7976 26144
rect 7912 26084 7916 26140
rect 7916 26084 7972 26140
rect 7972 26084 7976 26140
rect 7912 26080 7976 26084
rect 7992 26140 8056 26144
rect 7992 26084 7996 26140
rect 7996 26084 8052 26140
rect 8052 26084 8056 26140
rect 7992 26080 8056 26084
rect 9352 26140 9416 26144
rect 9352 26084 9356 26140
rect 9356 26084 9412 26140
rect 9412 26084 9416 26140
rect 9352 26080 9416 26084
rect 9432 26140 9496 26144
rect 9432 26084 9436 26140
rect 9436 26084 9492 26140
rect 9492 26084 9496 26140
rect 9432 26080 9496 26084
rect 9512 26140 9576 26144
rect 9512 26084 9516 26140
rect 9516 26084 9572 26140
rect 9572 26084 9576 26140
rect 9512 26080 9576 26084
rect 9592 26140 9656 26144
rect 9592 26084 9596 26140
rect 9596 26084 9652 26140
rect 9652 26084 9656 26140
rect 9592 26080 9656 26084
rect 11836 25740 11900 25804
rect 3612 25596 3676 25600
rect 3612 25540 3616 25596
rect 3616 25540 3672 25596
rect 3672 25540 3676 25596
rect 3612 25536 3676 25540
rect 3692 25596 3756 25600
rect 3692 25540 3696 25596
rect 3696 25540 3752 25596
rect 3752 25540 3756 25596
rect 3692 25536 3756 25540
rect 3772 25596 3836 25600
rect 3772 25540 3776 25596
rect 3776 25540 3832 25596
rect 3832 25540 3836 25596
rect 3772 25536 3836 25540
rect 3852 25596 3916 25600
rect 3852 25540 3856 25596
rect 3856 25540 3912 25596
rect 3912 25540 3916 25596
rect 3852 25536 3916 25540
rect 5212 25596 5276 25600
rect 5212 25540 5216 25596
rect 5216 25540 5272 25596
rect 5272 25540 5276 25596
rect 5212 25536 5276 25540
rect 5292 25596 5356 25600
rect 5292 25540 5296 25596
rect 5296 25540 5352 25596
rect 5352 25540 5356 25596
rect 5292 25536 5356 25540
rect 5372 25596 5436 25600
rect 5372 25540 5376 25596
rect 5376 25540 5432 25596
rect 5432 25540 5436 25596
rect 5372 25536 5436 25540
rect 5452 25596 5516 25600
rect 5452 25540 5456 25596
rect 5456 25540 5512 25596
rect 5512 25540 5516 25596
rect 5452 25536 5516 25540
rect 6812 25596 6876 25600
rect 6812 25540 6816 25596
rect 6816 25540 6872 25596
rect 6872 25540 6876 25596
rect 6812 25536 6876 25540
rect 6892 25596 6956 25600
rect 6892 25540 6896 25596
rect 6896 25540 6952 25596
rect 6952 25540 6956 25596
rect 6892 25536 6956 25540
rect 6972 25596 7036 25600
rect 6972 25540 6976 25596
rect 6976 25540 7032 25596
rect 7032 25540 7036 25596
rect 6972 25536 7036 25540
rect 7052 25596 7116 25600
rect 7052 25540 7056 25596
rect 7056 25540 7112 25596
rect 7112 25540 7116 25596
rect 7052 25536 7116 25540
rect 8412 25596 8476 25600
rect 8412 25540 8416 25596
rect 8416 25540 8472 25596
rect 8472 25540 8476 25596
rect 8412 25536 8476 25540
rect 8492 25596 8556 25600
rect 8492 25540 8496 25596
rect 8496 25540 8552 25596
rect 8552 25540 8556 25596
rect 8492 25536 8556 25540
rect 8572 25596 8636 25600
rect 8572 25540 8576 25596
rect 8576 25540 8632 25596
rect 8632 25540 8636 25596
rect 8572 25536 8636 25540
rect 8652 25596 8716 25600
rect 8652 25540 8656 25596
rect 8656 25540 8712 25596
rect 8712 25540 8716 25596
rect 8652 25536 8716 25540
rect 2952 25052 3016 25056
rect 2952 24996 2956 25052
rect 2956 24996 3012 25052
rect 3012 24996 3016 25052
rect 2952 24992 3016 24996
rect 3032 25052 3096 25056
rect 3032 24996 3036 25052
rect 3036 24996 3092 25052
rect 3092 24996 3096 25052
rect 3032 24992 3096 24996
rect 3112 25052 3176 25056
rect 3112 24996 3116 25052
rect 3116 24996 3172 25052
rect 3172 24996 3176 25052
rect 3112 24992 3176 24996
rect 3192 25052 3256 25056
rect 3192 24996 3196 25052
rect 3196 24996 3252 25052
rect 3252 24996 3256 25052
rect 3192 24992 3256 24996
rect 4552 25052 4616 25056
rect 4552 24996 4556 25052
rect 4556 24996 4612 25052
rect 4612 24996 4616 25052
rect 4552 24992 4616 24996
rect 4632 25052 4696 25056
rect 4632 24996 4636 25052
rect 4636 24996 4692 25052
rect 4692 24996 4696 25052
rect 4632 24992 4696 24996
rect 4712 25052 4776 25056
rect 4712 24996 4716 25052
rect 4716 24996 4772 25052
rect 4772 24996 4776 25052
rect 4712 24992 4776 24996
rect 4792 25052 4856 25056
rect 4792 24996 4796 25052
rect 4796 24996 4852 25052
rect 4852 24996 4856 25052
rect 4792 24992 4856 24996
rect 6152 25052 6216 25056
rect 6152 24996 6156 25052
rect 6156 24996 6212 25052
rect 6212 24996 6216 25052
rect 6152 24992 6216 24996
rect 6232 25052 6296 25056
rect 6232 24996 6236 25052
rect 6236 24996 6292 25052
rect 6292 24996 6296 25052
rect 6232 24992 6296 24996
rect 6312 25052 6376 25056
rect 6312 24996 6316 25052
rect 6316 24996 6372 25052
rect 6372 24996 6376 25052
rect 6312 24992 6376 24996
rect 6392 25052 6456 25056
rect 6392 24996 6396 25052
rect 6396 24996 6452 25052
rect 6452 24996 6456 25052
rect 6392 24992 6456 24996
rect 7752 25052 7816 25056
rect 7752 24996 7756 25052
rect 7756 24996 7812 25052
rect 7812 24996 7816 25052
rect 7752 24992 7816 24996
rect 7832 25052 7896 25056
rect 7832 24996 7836 25052
rect 7836 24996 7892 25052
rect 7892 24996 7896 25052
rect 7832 24992 7896 24996
rect 7912 25052 7976 25056
rect 7912 24996 7916 25052
rect 7916 24996 7972 25052
rect 7972 24996 7976 25052
rect 7912 24992 7976 24996
rect 7992 25052 8056 25056
rect 7992 24996 7996 25052
rect 7996 24996 8052 25052
rect 8052 24996 8056 25052
rect 7992 24992 8056 24996
rect 9352 25052 9416 25056
rect 9352 24996 9356 25052
rect 9356 24996 9412 25052
rect 9412 24996 9416 25052
rect 9352 24992 9416 24996
rect 9432 25052 9496 25056
rect 9432 24996 9436 25052
rect 9436 24996 9492 25052
rect 9492 24996 9496 25052
rect 9432 24992 9496 24996
rect 9512 25052 9576 25056
rect 9512 24996 9516 25052
rect 9516 24996 9572 25052
rect 9572 24996 9576 25052
rect 9512 24992 9576 24996
rect 9592 25052 9656 25056
rect 9592 24996 9596 25052
rect 9596 24996 9652 25052
rect 9652 24996 9656 25052
rect 9592 24992 9656 24996
rect 3612 24508 3676 24512
rect 3612 24452 3616 24508
rect 3616 24452 3672 24508
rect 3672 24452 3676 24508
rect 3612 24448 3676 24452
rect 3692 24508 3756 24512
rect 3692 24452 3696 24508
rect 3696 24452 3752 24508
rect 3752 24452 3756 24508
rect 3692 24448 3756 24452
rect 3772 24508 3836 24512
rect 3772 24452 3776 24508
rect 3776 24452 3832 24508
rect 3832 24452 3836 24508
rect 3772 24448 3836 24452
rect 3852 24508 3916 24512
rect 3852 24452 3856 24508
rect 3856 24452 3912 24508
rect 3912 24452 3916 24508
rect 3852 24448 3916 24452
rect 5212 24508 5276 24512
rect 5212 24452 5216 24508
rect 5216 24452 5272 24508
rect 5272 24452 5276 24508
rect 5212 24448 5276 24452
rect 5292 24508 5356 24512
rect 5292 24452 5296 24508
rect 5296 24452 5352 24508
rect 5352 24452 5356 24508
rect 5292 24448 5356 24452
rect 5372 24508 5436 24512
rect 5372 24452 5376 24508
rect 5376 24452 5432 24508
rect 5432 24452 5436 24508
rect 5372 24448 5436 24452
rect 5452 24508 5516 24512
rect 5452 24452 5456 24508
rect 5456 24452 5512 24508
rect 5512 24452 5516 24508
rect 5452 24448 5516 24452
rect 6812 24508 6876 24512
rect 6812 24452 6816 24508
rect 6816 24452 6872 24508
rect 6872 24452 6876 24508
rect 6812 24448 6876 24452
rect 6892 24508 6956 24512
rect 6892 24452 6896 24508
rect 6896 24452 6952 24508
rect 6952 24452 6956 24508
rect 6892 24448 6956 24452
rect 6972 24508 7036 24512
rect 6972 24452 6976 24508
rect 6976 24452 7032 24508
rect 7032 24452 7036 24508
rect 6972 24448 7036 24452
rect 7052 24508 7116 24512
rect 7052 24452 7056 24508
rect 7056 24452 7112 24508
rect 7112 24452 7116 24508
rect 7052 24448 7116 24452
rect 8412 24508 8476 24512
rect 8412 24452 8416 24508
rect 8416 24452 8472 24508
rect 8472 24452 8476 24508
rect 8412 24448 8476 24452
rect 8492 24508 8556 24512
rect 8492 24452 8496 24508
rect 8496 24452 8552 24508
rect 8552 24452 8556 24508
rect 8492 24448 8556 24452
rect 8572 24508 8636 24512
rect 8572 24452 8576 24508
rect 8576 24452 8632 24508
rect 8632 24452 8636 24508
rect 8572 24448 8636 24452
rect 8652 24508 8716 24512
rect 8652 24452 8656 24508
rect 8656 24452 8712 24508
rect 8712 24452 8716 24508
rect 8652 24448 8716 24452
rect 2952 23964 3016 23968
rect 2952 23908 2956 23964
rect 2956 23908 3012 23964
rect 3012 23908 3016 23964
rect 2952 23904 3016 23908
rect 3032 23964 3096 23968
rect 3032 23908 3036 23964
rect 3036 23908 3092 23964
rect 3092 23908 3096 23964
rect 3032 23904 3096 23908
rect 3112 23964 3176 23968
rect 3112 23908 3116 23964
rect 3116 23908 3172 23964
rect 3172 23908 3176 23964
rect 3112 23904 3176 23908
rect 3192 23964 3256 23968
rect 3192 23908 3196 23964
rect 3196 23908 3252 23964
rect 3252 23908 3256 23964
rect 3192 23904 3256 23908
rect 4552 23964 4616 23968
rect 4552 23908 4556 23964
rect 4556 23908 4612 23964
rect 4612 23908 4616 23964
rect 4552 23904 4616 23908
rect 4632 23964 4696 23968
rect 4632 23908 4636 23964
rect 4636 23908 4692 23964
rect 4692 23908 4696 23964
rect 4632 23904 4696 23908
rect 4712 23964 4776 23968
rect 4712 23908 4716 23964
rect 4716 23908 4772 23964
rect 4772 23908 4776 23964
rect 4712 23904 4776 23908
rect 4792 23964 4856 23968
rect 4792 23908 4796 23964
rect 4796 23908 4852 23964
rect 4852 23908 4856 23964
rect 4792 23904 4856 23908
rect 6152 23964 6216 23968
rect 6152 23908 6156 23964
rect 6156 23908 6212 23964
rect 6212 23908 6216 23964
rect 6152 23904 6216 23908
rect 6232 23964 6296 23968
rect 6232 23908 6236 23964
rect 6236 23908 6292 23964
rect 6292 23908 6296 23964
rect 6232 23904 6296 23908
rect 6312 23964 6376 23968
rect 6312 23908 6316 23964
rect 6316 23908 6372 23964
rect 6372 23908 6376 23964
rect 6312 23904 6376 23908
rect 6392 23964 6456 23968
rect 6392 23908 6396 23964
rect 6396 23908 6452 23964
rect 6452 23908 6456 23964
rect 6392 23904 6456 23908
rect 7752 23964 7816 23968
rect 7752 23908 7756 23964
rect 7756 23908 7812 23964
rect 7812 23908 7816 23964
rect 7752 23904 7816 23908
rect 7832 23964 7896 23968
rect 7832 23908 7836 23964
rect 7836 23908 7892 23964
rect 7892 23908 7896 23964
rect 7832 23904 7896 23908
rect 7912 23964 7976 23968
rect 7912 23908 7916 23964
rect 7916 23908 7972 23964
rect 7972 23908 7976 23964
rect 7912 23904 7976 23908
rect 7992 23964 8056 23968
rect 7992 23908 7996 23964
rect 7996 23908 8052 23964
rect 8052 23908 8056 23964
rect 7992 23904 8056 23908
rect 9352 23964 9416 23968
rect 9352 23908 9356 23964
rect 9356 23908 9412 23964
rect 9412 23908 9416 23964
rect 9352 23904 9416 23908
rect 9432 23964 9496 23968
rect 9432 23908 9436 23964
rect 9436 23908 9492 23964
rect 9492 23908 9496 23964
rect 9432 23904 9496 23908
rect 9512 23964 9576 23968
rect 9512 23908 9516 23964
rect 9516 23908 9572 23964
rect 9572 23908 9576 23964
rect 9512 23904 9576 23908
rect 9592 23964 9656 23968
rect 9592 23908 9596 23964
rect 9596 23908 9652 23964
rect 9652 23908 9656 23964
rect 9592 23904 9656 23908
rect 3612 23420 3676 23424
rect 3612 23364 3616 23420
rect 3616 23364 3672 23420
rect 3672 23364 3676 23420
rect 3612 23360 3676 23364
rect 3692 23420 3756 23424
rect 3692 23364 3696 23420
rect 3696 23364 3752 23420
rect 3752 23364 3756 23420
rect 3692 23360 3756 23364
rect 3772 23420 3836 23424
rect 3772 23364 3776 23420
rect 3776 23364 3832 23420
rect 3832 23364 3836 23420
rect 3772 23360 3836 23364
rect 3852 23420 3916 23424
rect 3852 23364 3856 23420
rect 3856 23364 3912 23420
rect 3912 23364 3916 23420
rect 3852 23360 3916 23364
rect 5212 23420 5276 23424
rect 5212 23364 5216 23420
rect 5216 23364 5272 23420
rect 5272 23364 5276 23420
rect 5212 23360 5276 23364
rect 5292 23420 5356 23424
rect 5292 23364 5296 23420
rect 5296 23364 5352 23420
rect 5352 23364 5356 23420
rect 5292 23360 5356 23364
rect 5372 23420 5436 23424
rect 5372 23364 5376 23420
rect 5376 23364 5432 23420
rect 5432 23364 5436 23420
rect 5372 23360 5436 23364
rect 5452 23420 5516 23424
rect 5452 23364 5456 23420
rect 5456 23364 5512 23420
rect 5512 23364 5516 23420
rect 5452 23360 5516 23364
rect 6812 23420 6876 23424
rect 6812 23364 6816 23420
rect 6816 23364 6872 23420
rect 6872 23364 6876 23420
rect 6812 23360 6876 23364
rect 6892 23420 6956 23424
rect 6892 23364 6896 23420
rect 6896 23364 6952 23420
rect 6952 23364 6956 23420
rect 6892 23360 6956 23364
rect 6972 23420 7036 23424
rect 6972 23364 6976 23420
rect 6976 23364 7032 23420
rect 7032 23364 7036 23420
rect 6972 23360 7036 23364
rect 7052 23420 7116 23424
rect 7052 23364 7056 23420
rect 7056 23364 7112 23420
rect 7112 23364 7116 23420
rect 7052 23360 7116 23364
rect 8412 23420 8476 23424
rect 8412 23364 8416 23420
rect 8416 23364 8472 23420
rect 8472 23364 8476 23420
rect 8412 23360 8476 23364
rect 8492 23420 8556 23424
rect 8492 23364 8496 23420
rect 8496 23364 8552 23420
rect 8552 23364 8556 23420
rect 8492 23360 8556 23364
rect 8572 23420 8636 23424
rect 8572 23364 8576 23420
rect 8576 23364 8632 23420
rect 8632 23364 8636 23420
rect 8572 23360 8636 23364
rect 8652 23420 8716 23424
rect 8652 23364 8656 23420
rect 8656 23364 8712 23420
rect 8712 23364 8716 23420
rect 8652 23360 8716 23364
rect 2952 22876 3016 22880
rect 2952 22820 2956 22876
rect 2956 22820 3012 22876
rect 3012 22820 3016 22876
rect 2952 22816 3016 22820
rect 3032 22876 3096 22880
rect 3032 22820 3036 22876
rect 3036 22820 3092 22876
rect 3092 22820 3096 22876
rect 3032 22816 3096 22820
rect 3112 22876 3176 22880
rect 3112 22820 3116 22876
rect 3116 22820 3172 22876
rect 3172 22820 3176 22876
rect 3112 22816 3176 22820
rect 3192 22876 3256 22880
rect 3192 22820 3196 22876
rect 3196 22820 3252 22876
rect 3252 22820 3256 22876
rect 3192 22816 3256 22820
rect 4552 22876 4616 22880
rect 4552 22820 4556 22876
rect 4556 22820 4612 22876
rect 4612 22820 4616 22876
rect 4552 22816 4616 22820
rect 4632 22876 4696 22880
rect 4632 22820 4636 22876
rect 4636 22820 4692 22876
rect 4692 22820 4696 22876
rect 4632 22816 4696 22820
rect 4712 22876 4776 22880
rect 4712 22820 4716 22876
rect 4716 22820 4772 22876
rect 4772 22820 4776 22876
rect 4712 22816 4776 22820
rect 4792 22876 4856 22880
rect 4792 22820 4796 22876
rect 4796 22820 4852 22876
rect 4852 22820 4856 22876
rect 4792 22816 4856 22820
rect 6152 22876 6216 22880
rect 6152 22820 6156 22876
rect 6156 22820 6212 22876
rect 6212 22820 6216 22876
rect 6152 22816 6216 22820
rect 6232 22876 6296 22880
rect 6232 22820 6236 22876
rect 6236 22820 6292 22876
rect 6292 22820 6296 22876
rect 6232 22816 6296 22820
rect 6312 22876 6376 22880
rect 6312 22820 6316 22876
rect 6316 22820 6372 22876
rect 6372 22820 6376 22876
rect 6312 22816 6376 22820
rect 6392 22876 6456 22880
rect 6392 22820 6396 22876
rect 6396 22820 6452 22876
rect 6452 22820 6456 22876
rect 6392 22816 6456 22820
rect 7752 22876 7816 22880
rect 7752 22820 7756 22876
rect 7756 22820 7812 22876
rect 7812 22820 7816 22876
rect 7752 22816 7816 22820
rect 7832 22876 7896 22880
rect 7832 22820 7836 22876
rect 7836 22820 7892 22876
rect 7892 22820 7896 22876
rect 7832 22816 7896 22820
rect 7912 22876 7976 22880
rect 7912 22820 7916 22876
rect 7916 22820 7972 22876
rect 7972 22820 7976 22876
rect 7912 22816 7976 22820
rect 7992 22876 8056 22880
rect 7992 22820 7996 22876
rect 7996 22820 8052 22876
rect 8052 22820 8056 22876
rect 7992 22816 8056 22820
rect 9352 22876 9416 22880
rect 9352 22820 9356 22876
rect 9356 22820 9412 22876
rect 9412 22820 9416 22876
rect 9352 22816 9416 22820
rect 9432 22876 9496 22880
rect 9432 22820 9436 22876
rect 9436 22820 9492 22876
rect 9492 22820 9496 22876
rect 9432 22816 9496 22820
rect 9512 22876 9576 22880
rect 9512 22820 9516 22876
rect 9516 22820 9572 22876
rect 9572 22820 9576 22876
rect 9512 22816 9576 22820
rect 9592 22876 9656 22880
rect 9592 22820 9596 22876
rect 9596 22820 9652 22876
rect 9652 22820 9656 22876
rect 9592 22816 9656 22820
rect 3612 22332 3676 22336
rect 3612 22276 3616 22332
rect 3616 22276 3672 22332
rect 3672 22276 3676 22332
rect 3612 22272 3676 22276
rect 3692 22332 3756 22336
rect 3692 22276 3696 22332
rect 3696 22276 3752 22332
rect 3752 22276 3756 22332
rect 3692 22272 3756 22276
rect 3772 22332 3836 22336
rect 3772 22276 3776 22332
rect 3776 22276 3832 22332
rect 3832 22276 3836 22332
rect 3772 22272 3836 22276
rect 3852 22332 3916 22336
rect 3852 22276 3856 22332
rect 3856 22276 3912 22332
rect 3912 22276 3916 22332
rect 3852 22272 3916 22276
rect 5212 22332 5276 22336
rect 5212 22276 5216 22332
rect 5216 22276 5272 22332
rect 5272 22276 5276 22332
rect 5212 22272 5276 22276
rect 5292 22332 5356 22336
rect 5292 22276 5296 22332
rect 5296 22276 5352 22332
rect 5352 22276 5356 22332
rect 5292 22272 5356 22276
rect 5372 22332 5436 22336
rect 5372 22276 5376 22332
rect 5376 22276 5432 22332
rect 5432 22276 5436 22332
rect 5372 22272 5436 22276
rect 5452 22332 5516 22336
rect 5452 22276 5456 22332
rect 5456 22276 5512 22332
rect 5512 22276 5516 22332
rect 5452 22272 5516 22276
rect 6812 22332 6876 22336
rect 6812 22276 6816 22332
rect 6816 22276 6872 22332
rect 6872 22276 6876 22332
rect 6812 22272 6876 22276
rect 6892 22332 6956 22336
rect 6892 22276 6896 22332
rect 6896 22276 6952 22332
rect 6952 22276 6956 22332
rect 6892 22272 6956 22276
rect 6972 22332 7036 22336
rect 6972 22276 6976 22332
rect 6976 22276 7032 22332
rect 7032 22276 7036 22332
rect 6972 22272 7036 22276
rect 7052 22332 7116 22336
rect 7052 22276 7056 22332
rect 7056 22276 7112 22332
rect 7112 22276 7116 22332
rect 7052 22272 7116 22276
rect 8412 22332 8476 22336
rect 8412 22276 8416 22332
rect 8416 22276 8472 22332
rect 8472 22276 8476 22332
rect 8412 22272 8476 22276
rect 8492 22332 8556 22336
rect 8492 22276 8496 22332
rect 8496 22276 8552 22332
rect 8552 22276 8556 22332
rect 8492 22272 8556 22276
rect 8572 22332 8636 22336
rect 8572 22276 8576 22332
rect 8576 22276 8632 22332
rect 8632 22276 8636 22332
rect 8572 22272 8636 22276
rect 8652 22332 8716 22336
rect 8652 22276 8656 22332
rect 8656 22276 8712 22332
rect 8712 22276 8716 22332
rect 8652 22272 8716 22276
rect 2952 21788 3016 21792
rect 2952 21732 2956 21788
rect 2956 21732 3012 21788
rect 3012 21732 3016 21788
rect 2952 21728 3016 21732
rect 3032 21788 3096 21792
rect 3032 21732 3036 21788
rect 3036 21732 3092 21788
rect 3092 21732 3096 21788
rect 3032 21728 3096 21732
rect 3112 21788 3176 21792
rect 3112 21732 3116 21788
rect 3116 21732 3172 21788
rect 3172 21732 3176 21788
rect 3112 21728 3176 21732
rect 3192 21788 3256 21792
rect 3192 21732 3196 21788
rect 3196 21732 3252 21788
rect 3252 21732 3256 21788
rect 3192 21728 3256 21732
rect 4552 21788 4616 21792
rect 4552 21732 4556 21788
rect 4556 21732 4612 21788
rect 4612 21732 4616 21788
rect 4552 21728 4616 21732
rect 4632 21788 4696 21792
rect 4632 21732 4636 21788
rect 4636 21732 4692 21788
rect 4692 21732 4696 21788
rect 4632 21728 4696 21732
rect 4712 21788 4776 21792
rect 4712 21732 4716 21788
rect 4716 21732 4772 21788
rect 4772 21732 4776 21788
rect 4712 21728 4776 21732
rect 4792 21788 4856 21792
rect 4792 21732 4796 21788
rect 4796 21732 4852 21788
rect 4852 21732 4856 21788
rect 4792 21728 4856 21732
rect 6152 21788 6216 21792
rect 6152 21732 6156 21788
rect 6156 21732 6212 21788
rect 6212 21732 6216 21788
rect 6152 21728 6216 21732
rect 6232 21788 6296 21792
rect 6232 21732 6236 21788
rect 6236 21732 6292 21788
rect 6292 21732 6296 21788
rect 6232 21728 6296 21732
rect 6312 21788 6376 21792
rect 6312 21732 6316 21788
rect 6316 21732 6372 21788
rect 6372 21732 6376 21788
rect 6312 21728 6376 21732
rect 6392 21788 6456 21792
rect 6392 21732 6396 21788
rect 6396 21732 6452 21788
rect 6452 21732 6456 21788
rect 6392 21728 6456 21732
rect 7752 21788 7816 21792
rect 7752 21732 7756 21788
rect 7756 21732 7812 21788
rect 7812 21732 7816 21788
rect 7752 21728 7816 21732
rect 7832 21788 7896 21792
rect 7832 21732 7836 21788
rect 7836 21732 7892 21788
rect 7892 21732 7896 21788
rect 7832 21728 7896 21732
rect 7912 21788 7976 21792
rect 7912 21732 7916 21788
rect 7916 21732 7972 21788
rect 7972 21732 7976 21788
rect 7912 21728 7976 21732
rect 7992 21788 8056 21792
rect 7992 21732 7996 21788
rect 7996 21732 8052 21788
rect 8052 21732 8056 21788
rect 7992 21728 8056 21732
rect 9352 21788 9416 21792
rect 9352 21732 9356 21788
rect 9356 21732 9412 21788
rect 9412 21732 9416 21788
rect 9352 21728 9416 21732
rect 9432 21788 9496 21792
rect 9432 21732 9436 21788
rect 9436 21732 9492 21788
rect 9492 21732 9496 21788
rect 9432 21728 9496 21732
rect 9512 21788 9576 21792
rect 9512 21732 9516 21788
rect 9516 21732 9572 21788
rect 9572 21732 9576 21788
rect 9512 21728 9576 21732
rect 9592 21788 9656 21792
rect 9592 21732 9596 21788
rect 9596 21732 9652 21788
rect 9652 21732 9656 21788
rect 9592 21728 9656 21732
rect 3612 21244 3676 21248
rect 3612 21188 3616 21244
rect 3616 21188 3672 21244
rect 3672 21188 3676 21244
rect 3612 21184 3676 21188
rect 3692 21244 3756 21248
rect 3692 21188 3696 21244
rect 3696 21188 3752 21244
rect 3752 21188 3756 21244
rect 3692 21184 3756 21188
rect 3772 21244 3836 21248
rect 3772 21188 3776 21244
rect 3776 21188 3832 21244
rect 3832 21188 3836 21244
rect 3772 21184 3836 21188
rect 3852 21244 3916 21248
rect 3852 21188 3856 21244
rect 3856 21188 3912 21244
rect 3912 21188 3916 21244
rect 3852 21184 3916 21188
rect 5212 21244 5276 21248
rect 5212 21188 5216 21244
rect 5216 21188 5272 21244
rect 5272 21188 5276 21244
rect 5212 21184 5276 21188
rect 5292 21244 5356 21248
rect 5292 21188 5296 21244
rect 5296 21188 5352 21244
rect 5352 21188 5356 21244
rect 5292 21184 5356 21188
rect 5372 21244 5436 21248
rect 5372 21188 5376 21244
rect 5376 21188 5432 21244
rect 5432 21188 5436 21244
rect 5372 21184 5436 21188
rect 5452 21244 5516 21248
rect 5452 21188 5456 21244
rect 5456 21188 5512 21244
rect 5512 21188 5516 21244
rect 5452 21184 5516 21188
rect 6812 21244 6876 21248
rect 6812 21188 6816 21244
rect 6816 21188 6872 21244
rect 6872 21188 6876 21244
rect 6812 21184 6876 21188
rect 6892 21244 6956 21248
rect 6892 21188 6896 21244
rect 6896 21188 6952 21244
rect 6952 21188 6956 21244
rect 6892 21184 6956 21188
rect 6972 21244 7036 21248
rect 6972 21188 6976 21244
rect 6976 21188 7032 21244
rect 7032 21188 7036 21244
rect 6972 21184 7036 21188
rect 7052 21244 7116 21248
rect 7052 21188 7056 21244
rect 7056 21188 7112 21244
rect 7112 21188 7116 21244
rect 7052 21184 7116 21188
rect 8412 21244 8476 21248
rect 8412 21188 8416 21244
rect 8416 21188 8472 21244
rect 8472 21188 8476 21244
rect 8412 21184 8476 21188
rect 8492 21244 8556 21248
rect 8492 21188 8496 21244
rect 8496 21188 8552 21244
rect 8552 21188 8556 21244
rect 8492 21184 8556 21188
rect 8572 21244 8636 21248
rect 8572 21188 8576 21244
rect 8576 21188 8632 21244
rect 8632 21188 8636 21244
rect 8572 21184 8636 21188
rect 8652 21244 8716 21248
rect 8652 21188 8656 21244
rect 8656 21188 8712 21244
rect 8712 21188 8716 21244
rect 8652 21184 8716 21188
rect 2952 20700 3016 20704
rect 2952 20644 2956 20700
rect 2956 20644 3012 20700
rect 3012 20644 3016 20700
rect 2952 20640 3016 20644
rect 3032 20700 3096 20704
rect 3032 20644 3036 20700
rect 3036 20644 3092 20700
rect 3092 20644 3096 20700
rect 3032 20640 3096 20644
rect 3112 20700 3176 20704
rect 3112 20644 3116 20700
rect 3116 20644 3172 20700
rect 3172 20644 3176 20700
rect 3112 20640 3176 20644
rect 3192 20700 3256 20704
rect 3192 20644 3196 20700
rect 3196 20644 3252 20700
rect 3252 20644 3256 20700
rect 3192 20640 3256 20644
rect 4552 20700 4616 20704
rect 4552 20644 4556 20700
rect 4556 20644 4612 20700
rect 4612 20644 4616 20700
rect 4552 20640 4616 20644
rect 4632 20700 4696 20704
rect 4632 20644 4636 20700
rect 4636 20644 4692 20700
rect 4692 20644 4696 20700
rect 4632 20640 4696 20644
rect 4712 20700 4776 20704
rect 4712 20644 4716 20700
rect 4716 20644 4772 20700
rect 4772 20644 4776 20700
rect 4712 20640 4776 20644
rect 4792 20700 4856 20704
rect 4792 20644 4796 20700
rect 4796 20644 4852 20700
rect 4852 20644 4856 20700
rect 4792 20640 4856 20644
rect 6152 20700 6216 20704
rect 6152 20644 6156 20700
rect 6156 20644 6212 20700
rect 6212 20644 6216 20700
rect 6152 20640 6216 20644
rect 6232 20700 6296 20704
rect 6232 20644 6236 20700
rect 6236 20644 6292 20700
rect 6292 20644 6296 20700
rect 6232 20640 6296 20644
rect 6312 20700 6376 20704
rect 6312 20644 6316 20700
rect 6316 20644 6372 20700
rect 6372 20644 6376 20700
rect 6312 20640 6376 20644
rect 6392 20700 6456 20704
rect 6392 20644 6396 20700
rect 6396 20644 6452 20700
rect 6452 20644 6456 20700
rect 6392 20640 6456 20644
rect 7752 20700 7816 20704
rect 7752 20644 7756 20700
rect 7756 20644 7812 20700
rect 7812 20644 7816 20700
rect 7752 20640 7816 20644
rect 7832 20700 7896 20704
rect 7832 20644 7836 20700
rect 7836 20644 7892 20700
rect 7892 20644 7896 20700
rect 7832 20640 7896 20644
rect 7912 20700 7976 20704
rect 7912 20644 7916 20700
rect 7916 20644 7972 20700
rect 7972 20644 7976 20700
rect 7912 20640 7976 20644
rect 7992 20700 8056 20704
rect 7992 20644 7996 20700
rect 7996 20644 8052 20700
rect 8052 20644 8056 20700
rect 7992 20640 8056 20644
rect 9352 20700 9416 20704
rect 9352 20644 9356 20700
rect 9356 20644 9412 20700
rect 9412 20644 9416 20700
rect 9352 20640 9416 20644
rect 9432 20700 9496 20704
rect 9432 20644 9436 20700
rect 9436 20644 9492 20700
rect 9492 20644 9496 20700
rect 9432 20640 9496 20644
rect 9512 20700 9576 20704
rect 9512 20644 9516 20700
rect 9516 20644 9572 20700
rect 9572 20644 9576 20700
rect 9512 20640 9576 20644
rect 9592 20700 9656 20704
rect 9592 20644 9596 20700
rect 9596 20644 9652 20700
rect 9652 20644 9656 20700
rect 9592 20640 9656 20644
rect 3612 20156 3676 20160
rect 3612 20100 3616 20156
rect 3616 20100 3672 20156
rect 3672 20100 3676 20156
rect 3612 20096 3676 20100
rect 3692 20156 3756 20160
rect 3692 20100 3696 20156
rect 3696 20100 3752 20156
rect 3752 20100 3756 20156
rect 3692 20096 3756 20100
rect 3772 20156 3836 20160
rect 3772 20100 3776 20156
rect 3776 20100 3832 20156
rect 3832 20100 3836 20156
rect 3772 20096 3836 20100
rect 3852 20156 3916 20160
rect 3852 20100 3856 20156
rect 3856 20100 3912 20156
rect 3912 20100 3916 20156
rect 3852 20096 3916 20100
rect 5212 20156 5276 20160
rect 5212 20100 5216 20156
rect 5216 20100 5272 20156
rect 5272 20100 5276 20156
rect 5212 20096 5276 20100
rect 5292 20156 5356 20160
rect 5292 20100 5296 20156
rect 5296 20100 5352 20156
rect 5352 20100 5356 20156
rect 5292 20096 5356 20100
rect 5372 20156 5436 20160
rect 5372 20100 5376 20156
rect 5376 20100 5432 20156
rect 5432 20100 5436 20156
rect 5372 20096 5436 20100
rect 5452 20156 5516 20160
rect 5452 20100 5456 20156
rect 5456 20100 5512 20156
rect 5512 20100 5516 20156
rect 5452 20096 5516 20100
rect 6812 20156 6876 20160
rect 6812 20100 6816 20156
rect 6816 20100 6872 20156
rect 6872 20100 6876 20156
rect 6812 20096 6876 20100
rect 6892 20156 6956 20160
rect 6892 20100 6896 20156
rect 6896 20100 6952 20156
rect 6952 20100 6956 20156
rect 6892 20096 6956 20100
rect 6972 20156 7036 20160
rect 6972 20100 6976 20156
rect 6976 20100 7032 20156
rect 7032 20100 7036 20156
rect 6972 20096 7036 20100
rect 7052 20156 7116 20160
rect 7052 20100 7056 20156
rect 7056 20100 7112 20156
rect 7112 20100 7116 20156
rect 7052 20096 7116 20100
rect 8412 20156 8476 20160
rect 8412 20100 8416 20156
rect 8416 20100 8472 20156
rect 8472 20100 8476 20156
rect 8412 20096 8476 20100
rect 8492 20156 8556 20160
rect 8492 20100 8496 20156
rect 8496 20100 8552 20156
rect 8552 20100 8556 20156
rect 8492 20096 8556 20100
rect 8572 20156 8636 20160
rect 8572 20100 8576 20156
rect 8576 20100 8632 20156
rect 8632 20100 8636 20156
rect 8572 20096 8636 20100
rect 8652 20156 8716 20160
rect 8652 20100 8656 20156
rect 8656 20100 8712 20156
rect 8712 20100 8716 20156
rect 8652 20096 8716 20100
rect 2952 19612 3016 19616
rect 2952 19556 2956 19612
rect 2956 19556 3012 19612
rect 3012 19556 3016 19612
rect 2952 19552 3016 19556
rect 3032 19612 3096 19616
rect 3032 19556 3036 19612
rect 3036 19556 3092 19612
rect 3092 19556 3096 19612
rect 3032 19552 3096 19556
rect 3112 19612 3176 19616
rect 3112 19556 3116 19612
rect 3116 19556 3172 19612
rect 3172 19556 3176 19612
rect 3112 19552 3176 19556
rect 3192 19612 3256 19616
rect 3192 19556 3196 19612
rect 3196 19556 3252 19612
rect 3252 19556 3256 19612
rect 3192 19552 3256 19556
rect 4552 19612 4616 19616
rect 4552 19556 4556 19612
rect 4556 19556 4612 19612
rect 4612 19556 4616 19612
rect 4552 19552 4616 19556
rect 4632 19612 4696 19616
rect 4632 19556 4636 19612
rect 4636 19556 4692 19612
rect 4692 19556 4696 19612
rect 4632 19552 4696 19556
rect 4712 19612 4776 19616
rect 4712 19556 4716 19612
rect 4716 19556 4772 19612
rect 4772 19556 4776 19612
rect 4712 19552 4776 19556
rect 4792 19612 4856 19616
rect 4792 19556 4796 19612
rect 4796 19556 4852 19612
rect 4852 19556 4856 19612
rect 4792 19552 4856 19556
rect 6152 19612 6216 19616
rect 6152 19556 6156 19612
rect 6156 19556 6212 19612
rect 6212 19556 6216 19612
rect 6152 19552 6216 19556
rect 6232 19612 6296 19616
rect 6232 19556 6236 19612
rect 6236 19556 6292 19612
rect 6292 19556 6296 19612
rect 6232 19552 6296 19556
rect 6312 19612 6376 19616
rect 6312 19556 6316 19612
rect 6316 19556 6372 19612
rect 6372 19556 6376 19612
rect 6312 19552 6376 19556
rect 6392 19612 6456 19616
rect 6392 19556 6396 19612
rect 6396 19556 6452 19612
rect 6452 19556 6456 19612
rect 6392 19552 6456 19556
rect 7752 19612 7816 19616
rect 7752 19556 7756 19612
rect 7756 19556 7812 19612
rect 7812 19556 7816 19612
rect 7752 19552 7816 19556
rect 7832 19612 7896 19616
rect 7832 19556 7836 19612
rect 7836 19556 7892 19612
rect 7892 19556 7896 19612
rect 7832 19552 7896 19556
rect 7912 19612 7976 19616
rect 7912 19556 7916 19612
rect 7916 19556 7972 19612
rect 7972 19556 7976 19612
rect 7912 19552 7976 19556
rect 7992 19612 8056 19616
rect 7992 19556 7996 19612
rect 7996 19556 8052 19612
rect 8052 19556 8056 19612
rect 7992 19552 8056 19556
rect 9352 19612 9416 19616
rect 9352 19556 9356 19612
rect 9356 19556 9412 19612
rect 9412 19556 9416 19612
rect 9352 19552 9416 19556
rect 9432 19612 9496 19616
rect 9432 19556 9436 19612
rect 9436 19556 9492 19612
rect 9492 19556 9496 19612
rect 9432 19552 9496 19556
rect 9512 19612 9576 19616
rect 9512 19556 9516 19612
rect 9516 19556 9572 19612
rect 9572 19556 9576 19612
rect 9512 19552 9576 19556
rect 9592 19612 9656 19616
rect 9592 19556 9596 19612
rect 9596 19556 9652 19612
rect 9652 19556 9656 19612
rect 9592 19552 9656 19556
rect 3612 19068 3676 19072
rect 3612 19012 3616 19068
rect 3616 19012 3672 19068
rect 3672 19012 3676 19068
rect 3612 19008 3676 19012
rect 3692 19068 3756 19072
rect 3692 19012 3696 19068
rect 3696 19012 3752 19068
rect 3752 19012 3756 19068
rect 3692 19008 3756 19012
rect 3772 19068 3836 19072
rect 3772 19012 3776 19068
rect 3776 19012 3832 19068
rect 3832 19012 3836 19068
rect 3772 19008 3836 19012
rect 3852 19068 3916 19072
rect 3852 19012 3856 19068
rect 3856 19012 3912 19068
rect 3912 19012 3916 19068
rect 3852 19008 3916 19012
rect 5212 19068 5276 19072
rect 5212 19012 5216 19068
rect 5216 19012 5272 19068
rect 5272 19012 5276 19068
rect 5212 19008 5276 19012
rect 5292 19068 5356 19072
rect 5292 19012 5296 19068
rect 5296 19012 5352 19068
rect 5352 19012 5356 19068
rect 5292 19008 5356 19012
rect 5372 19068 5436 19072
rect 5372 19012 5376 19068
rect 5376 19012 5432 19068
rect 5432 19012 5436 19068
rect 5372 19008 5436 19012
rect 5452 19068 5516 19072
rect 5452 19012 5456 19068
rect 5456 19012 5512 19068
rect 5512 19012 5516 19068
rect 5452 19008 5516 19012
rect 6812 19068 6876 19072
rect 6812 19012 6816 19068
rect 6816 19012 6872 19068
rect 6872 19012 6876 19068
rect 6812 19008 6876 19012
rect 6892 19068 6956 19072
rect 6892 19012 6896 19068
rect 6896 19012 6952 19068
rect 6952 19012 6956 19068
rect 6892 19008 6956 19012
rect 6972 19068 7036 19072
rect 6972 19012 6976 19068
rect 6976 19012 7032 19068
rect 7032 19012 7036 19068
rect 6972 19008 7036 19012
rect 7052 19068 7116 19072
rect 7052 19012 7056 19068
rect 7056 19012 7112 19068
rect 7112 19012 7116 19068
rect 7052 19008 7116 19012
rect 8412 19068 8476 19072
rect 8412 19012 8416 19068
rect 8416 19012 8472 19068
rect 8472 19012 8476 19068
rect 8412 19008 8476 19012
rect 8492 19068 8556 19072
rect 8492 19012 8496 19068
rect 8496 19012 8552 19068
rect 8552 19012 8556 19068
rect 8492 19008 8556 19012
rect 8572 19068 8636 19072
rect 8572 19012 8576 19068
rect 8576 19012 8632 19068
rect 8632 19012 8636 19068
rect 8572 19008 8636 19012
rect 8652 19068 8716 19072
rect 8652 19012 8656 19068
rect 8656 19012 8712 19068
rect 8712 19012 8716 19068
rect 8652 19008 8716 19012
rect 2952 18524 3016 18528
rect 2952 18468 2956 18524
rect 2956 18468 3012 18524
rect 3012 18468 3016 18524
rect 2952 18464 3016 18468
rect 3032 18524 3096 18528
rect 3032 18468 3036 18524
rect 3036 18468 3092 18524
rect 3092 18468 3096 18524
rect 3032 18464 3096 18468
rect 3112 18524 3176 18528
rect 3112 18468 3116 18524
rect 3116 18468 3172 18524
rect 3172 18468 3176 18524
rect 3112 18464 3176 18468
rect 3192 18524 3256 18528
rect 3192 18468 3196 18524
rect 3196 18468 3252 18524
rect 3252 18468 3256 18524
rect 3192 18464 3256 18468
rect 4552 18524 4616 18528
rect 4552 18468 4556 18524
rect 4556 18468 4612 18524
rect 4612 18468 4616 18524
rect 4552 18464 4616 18468
rect 4632 18524 4696 18528
rect 4632 18468 4636 18524
rect 4636 18468 4692 18524
rect 4692 18468 4696 18524
rect 4632 18464 4696 18468
rect 4712 18524 4776 18528
rect 4712 18468 4716 18524
rect 4716 18468 4772 18524
rect 4772 18468 4776 18524
rect 4712 18464 4776 18468
rect 4792 18524 4856 18528
rect 4792 18468 4796 18524
rect 4796 18468 4852 18524
rect 4852 18468 4856 18524
rect 4792 18464 4856 18468
rect 6152 18524 6216 18528
rect 6152 18468 6156 18524
rect 6156 18468 6212 18524
rect 6212 18468 6216 18524
rect 6152 18464 6216 18468
rect 6232 18524 6296 18528
rect 6232 18468 6236 18524
rect 6236 18468 6292 18524
rect 6292 18468 6296 18524
rect 6232 18464 6296 18468
rect 6312 18524 6376 18528
rect 6312 18468 6316 18524
rect 6316 18468 6372 18524
rect 6372 18468 6376 18524
rect 6312 18464 6376 18468
rect 6392 18524 6456 18528
rect 6392 18468 6396 18524
rect 6396 18468 6452 18524
rect 6452 18468 6456 18524
rect 6392 18464 6456 18468
rect 7752 18524 7816 18528
rect 7752 18468 7756 18524
rect 7756 18468 7812 18524
rect 7812 18468 7816 18524
rect 7752 18464 7816 18468
rect 7832 18524 7896 18528
rect 7832 18468 7836 18524
rect 7836 18468 7892 18524
rect 7892 18468 7896 18524
rect 7832 18464 7896 18468
rect 7912 18524 7976 18528
rect 7912 18468 7916 18524
rect 7916 18468 7972 18524
rect 7972 18468 7976 18524
rect 7912 18464 7976 18468
rect 7992 18524 8056 18528
rect 7992 18468 7996 18524
rect 7996 18468 8052 18524
rect 8052 18468 8056 18524
rect 7992 18464 8056 18468
rect 9352 18524 9416 18528
rect 9352 18468 9356 18524
rect 9356 18468 9412 18524
rect 9412 18468 9416 18524
rect 9352 18464 9416 18468
rect 9432 18524 9496 18528
rect 9432 18468 9436 18524
rect 9436 18468 9492 18524
rect 9492 18468 9496 18524
rect 9432 18464 9496 18468
rect 9512 18524 9576 18528
rect 9512 18468 9516 18524
rect 9516 18468 9572 18524
rect 9572 18468 9576 18524
rect 9512 18464 9576 18468
rect 9592 18524 9656 18528
rect 9592 18468 9596 18524
rect 9596 18468 9652 18524
rect 9652 18468 9656 18524
rect 9592 18464 9656 18468
rect 3612 17980 3676 17984
rect 3612 17924 3616 17980
rect 3616 17924 3672 17980
rect 3672 17924 3676 17980
rect 3612 17920 3676 17924
rect 3692 17980 3756 17984
rect 3692 17924 3696 17980
rect 3696 17924 3752 17980
rect 3752 17924 3756 17980
rect 3692 17920 3756 17924
rect 3772 17980 3836 17984
rect 3772 17924 3776 17980
rect 3776 17924 3832 17980
rect 3832 17924 3836 17980
rect 3772 17920 3836 17924
rect 3852 17980 3916 17984
rect 3852 17924 3856 17980
rect 3856 17924 3912 17980
rect 3912 17924 3916 17980
rect 3852 17920 3916 17924
rect 5212 17980 5276 17984
rect 5212 17924 5216 17980
rect 5216 17924 5272 17980
rect 5272 17924 5276 17980
rect 5212 17920 5276 17924
rect 5292 17980 5356 17984
rect 5292 17924 5296 17980
rect 5296 17924 5352 17980
rect 5352 17924 5356 17980
rect 5292 17920 5356 17924
rect 5372 17980 5436 17984
rect 5372 17924 5376 17980
rect 5376 17924 5432 17980
rect 5432 17924 5436 17980
rect 5372 17920 5436 17924
rect 5452 17980 5516 17984
rect 5452 17924 5456 17980
rect 5456 17924 5512 17980
rect 5512 17924 5516 17980
rect 5452 17920 5516 17924
rect 6812 17980 6876 17984
rect 6812 17924 6816 17980
rect 6816 17924 6872 17980
rect 6872 17924 6876 17980
rect 6812 17920 6876 17924
rect 6892 17980 6956 17984
rect 6892 17924 6896 17980
rect 6896 17924 6952 17980
rect 6952 17924 6956 17980
rect 6892 17920 6956 17924
rect 6972 17980 7036 17984
rect 6972 17924 6976 17980
rect 6976 17924 7032 17980
rect 7032 17924 7036 17980
rect 6972 17920 7036 17924
rect 7052 17980 7116 17984
rect 7052 17924 7056 17980
rect 7056 17924 7112 17980
rect 7112 17924 7116 17980
rect 7052 17920 7116 17924
rect 8412 17980 8476 17984
rect 8412 17924 8416 17980
rect 8416 17924 8472 17980
rect 8472 17924 8476 17980
rect 8412 17920 8476 17924
rect 8492 17980 8556 17984
rect 8492 17924 8496 17980
rect 8496 17924 8552 17980
rect 8552 17924 8556 17980
rect 8492 17920 8556 17924
rect 8572 17980 8636 17984
rect 8572 17924 8576 17980
rect 8576 17924 8632 17980
rect 8632 17924 8636 17980
rect 8572 17920 8636 17924
rect 8652 17980 8716 17984
rect 8652 17924 8656 17980
rect 8656 17924 8712 17980
rect 8712 17924 8716 17980
rect 8652 17920 8716 17924
rect 2952 17436 3016 17440
rect 2952 17380 2956 17436
rect 2956 17380 3012 17436
rect 3012 17380 3016 17436
rect 2952 17376 3016 17380
rect 3032 17436 3096 17440
rect 3032 17380 3036 17436
rect 3036 17380 3092 17436
rect 3092 17380 3096 17436
rect 3032 17376 3096 17380
rect 3112 17436 3176 17440
rect 3112 17380 3116 17436
rect 3116 17380 3172 17436
rect 3172 17380 3176 17436
rect 3112 17376 3176 17380
rect 3192 17436 3256 17440
rect 3192 17380 3196 17436
rect 3196 17380 3252 17436
rect 3252 17380 3256 17436
rect 3192 17376 3256 17380
rect 4552 17436 4616 17440
rect 4552 17380 4556 17436
rect 4556 17380 4612 17436
rect 4612 17380 4616 17436
rect 4552 17376 4616 17380
rect 4632 17436 4696 17440
rect 4632 17380 4636 17436
rect 4636 17380 4692 17436
rect 4692 17380 4696 17436
rect 4632 17376 4696 17380
rect 4712 17436 4776 17440
rect 4712 17380 4716 17436
rect 4716 17380 4772 17436
rect 4772 17380 4776 17436
rect 4712 17376 4776 17380
rect 4792 17436 4856 17440
rect 4792 17380 4796 17436
rect 4796 17380 4852 17436
rect 4852 17380 4856 17436
rect 4792 17376 4856 17380
rect 6152 17436 6216 17440
rect 6152 17380 6156 17436
rect 6156 17380 6212 17436
rect 6212 17380 6216 17436
rect 6152 17376 6216 17380
rect 6232 17436 6296 17440
rect 6232 17380 6236 17436
rect 6236 17380 6292 17436
rect 6292 17380 6296 17436
rect 6232 17376 6296 17380
rect 6312 17436 6376 17440
rect 6312 17380 6316 17436
rect 6316 17380 6372 17436
rect 6372 17380 6376 17436
rect 6312 17376 6376 17380
rect 6392 17436 6456 17440
rect 6392 17380 6396 17436
rect 6396 17380 6452 17436
rect 6452 17380 6456 17436
rect 6392 17376 6456 17380
rect 7752 17436 7816 17440
rect 7752 17380 7756 17436
rect 7756 17380 7812 17436
rect 7812 17380 7816 17436
rect 7752 17376 7816 17380
rect 7832 17436 7896 17440
rect 7832 17380 7836 17436
rect 7836 17380 7892 17436
rect 7892 17380 7896 17436
rect 7832 17376 7896 17380
rect 7912 17436 7976 17440
rect 7912 17380 7916 17436
rect 7916 17380 7972 17436
rect 7972 17380 7976 17436
rect 7912 17376 7976 17380
rect 7992 17436 8056 17440
rect 7992 17380 7996 17436
rect 7996 17380 8052 17436
rect 8052 17380 8056 17436
rect 7992 17376 8056 17380
rect 9352 17436 9416 17440
rect 9352 17380 9356 17436
rect 9356 17380 9412 17436
rect 9412 17380 9416 17436
rect 9352 17376 9416 17380
rect 9432 17436 9496 17440
rect 9432 17380 9436 17436
rect 9436 17380 9492 17436
rect 9492 17380 9496 17436
rect 9432 17376 9496 17380
rect 9512 17436 9576 17440
rect 9512 17380 9516 17436
rect 9516 17380 9572 17436
rect 9572 17380 9576 17436
rect 9512 17376 9576 17380
rect 9592 17436 9656 17440
rect 9592 17380 9596 17436
rect 9596 17380 9652 17436
rect 9652 17380 9656 17436
rect 9592 17376 9656 17380
rect 3612 16892 3676 16896
rect 3612 16836 3616 16892
rect 3616 16836 3672 16892
rect 3672 16836 3676 16892
rect 3612 16832 3676 16836
rect 3692 16892 3756 16896
rect 3692 16836 3696 16892
rect 3696 16836 3752 16892
rect 3752 16836 3756 16892
rect 3692 16832 3756 16836
rect 3772 16892 3836 16896
rect 3772 16836 3776 16892
rect 3776 16836 3832 16892
rect 3832 16836 3836 16892
rect 3772 16832 3836 16836
rect 3852 16892 3916 16896
rect 3852 16836 3856 16892
rect 3856 16836 3912 16892
rect 3912 16836 3916 16892
rect 3852 16832 3916 16836
rect 5212 16892 5276 16896
rect 5212 16836 5216 16892
rect 5216 16836 5272 16892
rect 5272 16836 5276 16892
rect 5212 16832 5276 16836
rect 5292 16892 5356 16896
rect 5292 16836 5296 16892
rect 5296 16836 5352 16892
rect 5352 16836 5356 16892
rect 5292 16832 5356 16836
rect 5372 16892 5436 16896
rect 5372 16836 5376 16892
rect 5376 16836 5432 16892
rect 5432 16836 5436 16892
rect 5372 16832 5436 16836
rect 5452 16892 5516 16896
rect 5452 16836 5456 16892
rect 5456 16836 5512 16892
rect 5512 16836 5516 16892
rect 5452 16832 5516 16836
rect 6812 16892 6876 16896
rect 6812 16836 6816 16892
rect 6816 16836 6872 16892
rect 6872 16836 6876 16892
rect 6812 16832 6876 16836
rect 6892 16892 6956 16896
rect 6892 16836 6896 16892
rect 6896 16836 6952 16892
rect 6952 16836 6956 16892
rect 6892 16832 6956 16836
rect 6972 16892 7036 16896
rect 6972 16836 6976 16892
rect 6976 16836 7032 16892
rect 7032 16836 7036 16892
rect 6972 16832 7036 16836
rect 7052 16892 7116 16896
rect 7052 16836 7056 16892
rect 7056 16836 7112 16892
rect 7112 16836 7116 16892
rect 7052 16832 7116 16836
rect 8412 16892 8476 16896
rect 8412 16836 8416 16892
rect 8416 16836 8472 16892
rect 8472 16836 8476 16892
rect 8412 16832 8476 16836
rect 8492 16892 8556 16896
rect 8492 16836 8496 16892
rect 8496 16836 8552 16892
rect 8552 16836 8556 16892
rect 8492 16832 8556 16836
rect 8572 16892 8636 16896
rect 8572 16836 8576 16892
rect 8576 16836 8632 16892
rect 8632 16836 8636 16892
rect 8572 16832 8636 16836
rect 8652 16892 8716 16896
rect 8652 16836 8656 16892
rect 8656 16836 8712 16892
rect 8712 16836 8716 16892
rect 8652 16832 8716 16836
rect 2952 16348 3016 16352
rect 2952 16292 2956 16348
rect 2956 16292 3012 16348
rect 3012 16292 3016 16348
rect 2952 16288 3016 16292
rect 3032 16348 3096 16352
rect 3032 16292 3036 16348
rect 3036 16292 3092 16348
rect 3092 16292 3096 16348
rect 3032 16288 3096 16292
rect 3112 16348 3176 16352
rect 3112 16292 3116 16348
rect 3116 16292 3172 16348
rect 3172 16292 3176 16348
rect 3112 16288 3176 16292
rect 3192 16348 3256 16352
rect 3192 16292 3196 16348
rect 3196 16292 3252 16348
rect 3252 16292 3256 16348
rect 3192 16288 3256 16292
rect 4552 16348 4616 16352
rect 4552 16292 4556 16348
rect 4556 16292 4612 16348
rect 4612 16292 4616 16348
rect 4552 16288 4616 16292
rect 4632 16348 4696 16352
rect 4632 16292 4636 16348
rect 4636 16292 4692 16348
rect 4692 16292 4696 16348
rect 4632 16288 4696 16292
rect 4712 16348 4776 16352
rect 4712 16292 4716 16348
rect 4716 16292 4772 16348
rect 4772 16292 4776 16348
rect 4712 16288 4776 16292
rect 4792 16348 4856 16352
rect 4792 16292 4796 16348
rect 4796 16292 4852 16348
rect 4852 16292 4856 16348
rect 4792 16288 4856 16292
rect 6152 16348 6216 16352
rect 6152 16292 6156 16348
rect 6156 16292 6212 16348
rect 6212 16292 6216 16348
rect 6152 16288 6216 16292
rect 6232 16348 6296 16352
rect 6232 16292 6236 16348
rect 6236 16292 6292 16348
rect 6292 16292 6296 16348
rect 6232 16288 6296 16292
rect 6312 16348 6376 16352
rect 6312 16292 6316 16348
rect 6316 16292 6372 16348
rect 6372 16292 6376 16348
rect 6312 16288 6376 16292
rect 6392 16348 6456 16352
rect 6392 16292 6396 16348
rect 6396 16292 6452 16348
rect 6452 16292 6456 16348
rect 6392 16288 6456 16292
rect 7752 16348 7816 16352
rect 7752 16292 7756 16348
rect 7756 16292 7812 16348
rect 7812 16292 7816 16348
rect 7752 16288 7816 16292
rect 7832 16348 7896 16352
rect 7832 16292 7836 16348
rect 7836 16292 7892 16348
rect 7892 16292 7896 16348
rect 7832 16288 7896 16292
rect 7912 16348 7976 16352
rect 7912 16292 7916 16348
rect 7916 16292 7972 16348
rect 7972 16292 7976 16348
rect 7912 16288 7976 16292
rect 7992 16348 8056 16352
rect 7992 16292 7996 16348
rect 7996 16292 8052 16348
rect 8052 16292 8056 16348
rect 7992 16288 8056 16292
rect 9352 16348 9416 16352
rect 9352 16292 9356 16348
rect 9356 16292 9412 16348
rect 9412 16292 9416 16348
rect 9352 16288 9416 16292
rect 9432 16348 9496 16352
rect 9432 16292 9436 16348
rect 9436 16292 9492 16348
rect 9492 16292 9496 16348
rect 9432 16288 9496 16292
rect 9512 16348 9576 16352
rect 9512 16292 9516 16348
rect 9516 16292 9572 16348
rect 9572 16292 9576 16348
rect 9512 16288 9576 16292
rect 9592 16348 9656 16352
rect 9592 16292 9596 16348
rect 9596 16292 9652 16348
rect 9652 16292 9656 16348
rect 9592 16288 9656 16292
rect 3612 15804 3676 15808
rect 3612 15748 3616 15804
rect 3616 15748 3672 15804
rect 3672 15748 3676 15804
rect 3612 15744 3676 15748
rect 3692 15804 3756 15808
rect 3692 15748 3696 15804
rect 3696 15748 3752 15804
rect 3752 15748 3756 15804
rect 3692 15744 3756 15748
rect 3772 15804 3836 15808
rect 3772 15748 3776 15804
rect 3776 15748 3832 15804
rect 3832 15748 3836 15804
rect 3772 15744 3836 15748
rect 3852 15804 3916 15808
rect 3852 15748 3856 15804
rect 3856 15748 3912 15804
rect 3912 15748 3916 15804
rect 3852 15744 3916 15748
rect 5212 15804 5276 15808
rect 5212 15748 5216 15804
rect 5216 15748 5272 15804
rect 5272 15748 5276 15804
rect 5212 15744 5276 15748
rect 5292 15804 5356 15808
rect 5292 15748 5296 15804
rect 5296 15748 5352 15804
rect 5352 15748 5356 15804
rect 5292 15744 5356 15748
rect 5372 15804 5436 15808
rect 5372 15748 5376 15804
rect 5376 15748 5432 15804
rect 5432 15748 5436 15804
rect 5372 15744 5436 15748
rect 5452 15804 5516 15808
rect 5452 15748 5456 15804
rect 5456 15748 5512 15804
rect 5512 15748 5516 15804
rect 5452 15744 5516 15748
rect 6812 15804 6876 15808
rect 6812 15748 6816 15804
rect 6816 15748 6872 15804
rect 6872 15748 6876 15804
rect 6812 15744 6876 15748
rect 6892 15804 6956 15808
rect 6892 15748 6896 15804
rect 6896 15748 6952 15804
rect 6952 15748 6956 15804
rect 6892 15744 6956 15748
rect 6972 15804 7036 15808
rect 6972 15748 6976 15804
rect 6976 15748 7032 15804
rect 7032 15748 7036 15804
rect 6972 15744 7036 15748
rect 7052 15804 7116 15808
rect 7052 15748 7056 15804
rect 7056 15748 7112 15804
rect 7112 15748 7116 15804
rect 7052 15744 7116 15748
rect 8412 15804 8476 15808
rect 8412 15748 8416 15804
rect 8416 15748 8472 15804
rect 8472 15748 8476 15804
rect 8412 15744 8476 15748
rect 8492 15804 8556 15808
rect 8492 15748 8496 15804
rect 8496 15748 8552 15804
rect 8552 15748 8556 15804
rect 8492 15744 8556 15748
rect 8572 15804 8636 15808
rect 8572 15748 8576 15804
rect 8576 15748 8632 15804
rect 8632 15748 8636 15804
rect 8572 15744 8636 15748
rect 8652 15804 8716 15808
rect 8652 15748 8656 15804
rect 8656 15748 8712 15804
rect 8712 15748 8716 15804
rect 8652 15744 8716 15748
rect 2952 15260 3016 15264
rect 2952 15204 2956 15260
rect 2956 15204 3012 15260
rect 3012 15204 3016 15260
rect 2952 15200 3016 15204
rect 3032 15260 3096 15264
rect 3032 15204 3036 15260
rect 3036 15204 3092 15260
rect 3092 15204 3096 15260
rect 3032 15200 3096 15204
rect 3112 15260 3176 15264
rect 3112 15204 3116 15260
rect 3116 15204 3172 15260
rect 3172 15204 3176 15260
rect 3112 15200 3176 15204
rect 3192 15260 3256 15264
rect 3192 15204 3196 15260
rect 3196 15204 3252 15260
rect 3252 15204 3256 15260
rect 3192 15200 3256 15204
rect 4552 15260 4616 15264
rect 4552 15204 4556 15260
rect 4556 15204 4612 15260
rect 4612 15204 4616 15260
rect 4552 15200 4616 15204
rect 4632 15260 4696 15264
rect 4632 15204 4636 15260
rect 4636 15204 4692 15260
rect 4692 15204 4696 15260
rect 4632 15200 4696 15204
rect 4712 15260 4776 15264
rect 4712 15204 4716 15260
rect 4716 15204 4772 15260
rect 4772 15204 4776 15260
rect 4712 15200 4776 15204
rect 4792 15260 4856 15264
rect 4792 15204 4796 15260
rect 4796 15204 4852 15260
rect 4852 15204 4856 15260
rect 4792 15200 4856 15204
rect 6152 15260 6216 15264
rect 6152 15204 6156 15260
rect 6156 15204 6212 15260
rect 6212 15204 6216 15260
rect 6152 15200 6216 15204
rect 6232 15260 6296 15264
rect 6232 15204 6236 15260
rect 6236 15204 6292 15260
rect 6292 15204 6296 15260
rect 6232 15200 6296 15204
rect 6312 15260 6376 15264
rect 6312 15204 6316 15260
rect 6316 15204 6372 15260
rect 6372 15204 6376 15260
rect 6312 15200 6376 15204
rect 6392 15260 6456 15264
rect 6392 15204 6396 15260
rect 6396 15204 6452 15260
rect 6452 15204 6456 15260
rect 6392 15200 6456 15204
rect 7752 15260 7816 15264
rect 7752 15204 7756 15260
rect 7756 15204 7812 15260
rect 7812 15204 7816 15260
rect 7752 15200 7816 15204
rect 7832 15260 7896 15264
rect 7832 15204 7836 15260
rect 7836 15204 7892 15260
rect 7892 15204 7896 15260
rect 7832 15200 7896 15204
rect 7912 15260 7976 15264
rect 7912 15204 7916 15260
rect 7916 15204 7972 15260
rect 7972 15204 7976 15260
rect 7912 15200 7976 15204
rect 7992 15260 8056 15264
rect 7992 15204 7996 15260
rect 7996 15204 8052 15260
rect 8052 15204 8056 15260
rect 7992 15200 8056 15204
rect 9352 15260 9416 15264
rect 9352 15204 9356 15260
rect 9356 15204 9412 15260
rect 9412 15204 9416 15260
rect 9352 15200 9416 15204
rect 9432 15260 9496 15264
rect 9432 15204 9436 15260
rect 9436 15204 9492 15260
rect 9492 15204 9496 15260
rect 9432 15200 9496 15204
rect 9512 15260 9576 15264
rect 9512 15204 9516 15260
rect 9516 15204 9572 15260
rect 9572 15204 9576 15260
rect 9512 15200 9576 15204
rect 9592 15260 9656 15264
rect 9592 15204 9596 15260
rect 9596 15204 9652 15260
rect 9652 15204 9656 15260
rect 9592 15200 9656 15204
rect 3612 14716 3676 14720
rect 3612 14660 3616 14716
rect 3616 14660 3672 14716
rect 3672 14660 3676 14716
rect 3612 14656 3676 14660
rect 3692 14716 3756 14720
rect 3692 14660 3696 14716
rect 3696 14660 3752 14716
rect 3752 14660 3756 14716
rect 3692 14656 3756 14660
rect 3772 14716 3836 14720
rect 3772 14660 3776 14716
rect 3776 14660 3832 14716
rect 3832 14660 3836 14716
rect 3772 14656 3836 14660
rect 3852 14716 3916 14720
rect 3852 14660 3856 14716
rect 3856 14660 3912 14716
rect 3912 14660 3916 14716
rect 3852 14656 3916 14660
rect 5212 14716 5276 14720
rect 5212 14660 5216 14716
rect 5216 14660 5272 14716
rect 5272 14660 5276 14716
rect 5212 14656 5276 14660
rect 5292 14716 5356 14720
rect 5292 14660 5296 14716
rect 5296 14660 5352 14716
rect 5352 14660 5356 14716
rect 5292 14656 5356 14660
rect 5372 14716 5436 14720
rect 5372 14660 5376 14716
rect 5376 14660 5432 14716
rect 5432 14660 5436 14716
rect 5372 14656 5436 14660
rect 5452 14716 5516 14720
rect 5452 14660 5456 14716
rect 5456 14660 5512 14716
rect 5512 14660 5516 14716
rect 5452 14656 5516 14660
rect 6812 14716 6876 14720
rect 6812 14660 6816 14716
rect 6816 14660 6872 14716
rect 6872 14660 6876 14716
rect 6812 14656 6876 14660
rect 6892 14716 6956 14720
rect 6892 14660 6896 14716
rect 6896 14660 6952 14716
rect 6952 14660 6956 14716
rect 6892 14656 6956 14660
rect 6972 14716 7036 14720
rect 6972 14660 6976 14716
rect 6976 14660 7032 14716
rect 7032 14660 7036 14716
rect 6972 14656 7036 14660
rect 7052 14716 7116 14720
rect 7052 14660 7056 14716
rect 7056 14660 7112 14716
rect 7112 14660 7116 14716
rect 7052 14656 7116 14660
rect 8412 14716 8476 14720
rect 8412 14660 8416 14716
rect 8416 14660 8472 14716
rect 8472 14660 8476 14716
rect 8412 14656 8476 14660
rect 8492 14716 8556 14720
rect 8492 14660 8496 14716
rect 8496 14660 8552 14716
rect 8552 14660 8556 14716
rect 8492 14656 8556 14660
rect 8572 14716 8636 14720
rect 8572 14660 8576 14716
rect 8576 14660 8632 14716
rect 8632 14660 8636 14716
rect 8572 14656 8636 14660
rect 8652 14716 8716 14720
rect 8652 14660 8656 14716
rect 8656 14660 8712 14716
rect 8712 14660 8716 14716
rect 8652 14656 8716 14660
rect 2952 14172 3016 14176
rect 2952 14116 2956 14172
rect 2956 14116 3012 14172
rect 3012 14116 3016 14172
rect 2952 14112 3016 14116
rect 3032 14172 3096 14176
rect 3032 14116 3036 14172
rect 3036 14116 3092 14172
rect 3092 14116 3096 14172
rect 3032 14112 3096 14116
rect 3112 14172 3176 14176
rect 3112 14116 3116 14172
rect 3116 14116 3172 14172
rect 3172 14116 3176 14172
rect 3112 14112 3176 14116
rect 3192 14172 3256 14176
rect 3192 14116 3196 14172
rect 3196 14116 3252 14172
rect 3252 14116 3256 14172
rect 3192 14112 3256 14116
rect 4552 14172 4616 14176
rect 4552 14116 4556 14172
rect 4556 14116 4612 14172
rect 4612 14116 4616 14172
rect 4552 14112 4616 14116
rect 4632 14172 4696 14176
rect 4632 14116 4636 14172
rect 4636 14116 4692 14172
rect 4692 14116 4696 14172
rect 4632 14112 4696 14116
rect 4712 14172 4776 14176
rect 4712 14116 4716 14172
rect 4716 14116 4772 14172
rect 4772 14116 4776 14172
rect 4712 14112 4776 14116
rect 4792 14172 4856 14176
rect 4792 14116 4796 14172
rect 4796 14116 4852 14172
rect 4852 14116 4856 14172
rect 4792 14112 4856 14116
rect 6152 14172 6216 14176
rect 6152 14116 6156 14172
rect 6156 14116 6212 14172
rect 6212 14116 6216 14172
rect 6152 14112 6216 14116
rect 6232 14172 6296 14176
rect 6232 14116 6236 14172
rect 6236 14116 6292 14172
rect 6292 14116 6296 14172
rect 6232 14112 6296 14116
rect 6312 14172 6376 14176
rect 6312 14116 6316 14172
rect 6316 14116 6372 14172
rect 6372 14116 6376 14172
rect 6312 14112 6376 14116
rect 6392 14172 6456 14176
rect 6392 14116 6396 14172
rect 6396 14116 6452 14172
rect 6452 14116 6456 14172
rect 6392 14112 6456 14116
rect 7752 14172 7816 14176
rect 7752 14116 7756 14172
rect 7756 14116 7812 14172
rect 7812 14116 7816 14172
rect 7752 14112 7816 14116
rect 7832 14172 7896 14176
rect 7832 14116 7836 14172
rect 7836 14116 7892 14172
rect 7892 14116 7896 14172
rect 7832 14112 7896 14116
rect 7912 14172 7976 14176
rect 7912 14116 7916 14172
rect 7916 14116 7972 14172
rect 7972 14116 7976 14172
rect 7912 14112 7976 14116
rect 7992 14172 8056 14176
rect 7992 14116 7996 14172
rect 7996 14116 8052 14172
rect 8052 14116 8056 14172
rect 7992 14112 8056 14116
rect 9352 14172 9416 14176
rect 9352 14116 9356 14172
rect 9356 14116 9412 14172
rect 9412 14116 9416 14172
rect 9352 14112 9416 14116
rect 9432 14172 9496 14176
rect 9432 14116 9436 14172
rect 9436 14116 9492 14172
rect 9492 14116 9496 14172
rect 9432 14112 9496 14116
rect 9512 14172 9576 14176
rect 9512 14116 9516 14172
rect 9516 14116 9572 14172
rect 9572 14116 9576 14172
rect 9512 14112 9576 14116
rect 9592 14172 9656 14176
rect 9592 14116 9596 14172
rect 9596 14116 9652 14172
rect 9652 14116 9656 14172
rect 9592 14112 9656 14116
rect 3612 13628 3676 13632
rect 3612 13572 3616 13628
rect 3616 13572 3672 13628
rect 3672 13572 3676 13628
rect 3612 13568 3676 13572
rect 3692 13628 3756 13632
rect 3692 13572 3696 13628
rect 3696 13572 3752 13628
rect 3752 13572 3756 13628
rect 3692 13568 3756 13572
rect 3772 13628 3836 13632
rect 3772 13572 3776 13628
rect 3776 13572 3832 13628
rect 3832 13572 3836 13628
rect 3772 13568 3836 13572
rect 3852 13628 3916 13632
rect 3852 13572 3856 13628
rect 3856 13572 3912 13628
rect 3912 13572 3916 13628
rect 3852 13568 3916 13572
rect 5212 13628 5276 13632
rect 5212 13572 5216 13628
rect 5216 13572 5272 13628
rect 5272 13572 5276 13628
rect 5212 13568 5276 13572
rect 5292 13628 5356 13632
rect 5292 13572 5296 13628
rect 5296 13572 5352 13628
rect 5352 13572 5356 13628
rect 5292 13568 5356 13572
rect 5372 13628 5436 13632
rect 5372 13572 5376 13628
rect 5376 13572 5432 13628
rect 5432 13572 5436 13628
rect 5372 13568 5436 13572
rect 5452 13628 5516 13632
rect 5452 13572 5456 13628
rect 5456 13572 5512 13628
rect 5512 13572 5516 13628
rect 5452 13568 5516 13572
rect 6812 13628 6876 13632
rect 6812 13572 6816 13628
rect 6816 13572 6872 13628
rect 6872 13572 6876 13628
rect 6812 13568 6876 13572
rect 6892 13628 6956 13632
rect 6892 13572 6896 13628
rect 6896 13572 6952 13628
rect 6952 13572 6956 13628
rect 6892 13568 6956 13572
rect 6972 13628 7036 13632
rect 6972 13572 6976 13628
rect 6976 13572 7032 13628
rect 7032 13572 7036 13628
rect 6972 13568 7036 13572
rect 7052 13628 7116 13632
rect 7052 13572 7056 13628
rect 7056 13572 7112 13628
rect 7112 13572 7116 13628
rect 7052 13568 7116 13572
rect 8412 13628 8476 13632
rect 8412 13572 8416 13628
rect 8416 13572 8472 13628
rect 8472 13572 8476 13628
rect 8412 13568 8476 13572
rect 8492 13628 8556 13632
rect 8492 13572 8496 13628
rect 8496 13572 8552 13628
rect 8552 13572 8556 13628
rect 8492 13568 8556 13572
rect 8572 13628 8636 13632
rect 8572 13572 8576 13628
rect 8576 13572 8632 13628
rect 8632 13572 8636 13628
rect 8572 13568 8636 13572
rect 8652 13628 8716 13632
rect 8652 13572 8656 13628
rect 8656 13572 8712 13628
rect 8712 13572 8716 13628
rect 8652 13568 8716 13572
rect 2952 13084 3016 13088
rect 2952 13028 2956 13084
rect 2956 13028 3012 13084
rect 3012 13028 3016 13084
rect 2952 13024 3016 13028
rect 3032 13084 3096 13088
rect 3032 13028 3036 13084
rect 3036 13028 3092 13084
rect 3092 13028 3096 13084
rect 3032 13024 3096 13028
rect 3112 13084 3176 13088
rect 3112 13028 3116 13084
rect 3116 13028 3172 13084
rect 3172 13028 3176 13084
rect 3112 13024 3176 13028
rect 3192 13084 3256 13088
rect 3192 13028 3196 13084
rect 3196 13028 3252 13084
rect 3252 13028 3256 13084
rect 3192 13024 3256 13028
rect 4552 13084 4616 13088
rect 4552 13028 4556 13084
rect 4556 13028 4612 13084
rect 4612 13028 4616 13084
rect 4552 13024 4616 13028
rect 4632 13084 4696 13088
rect 4632 13028 4636 13084
rect 4636 13028 4692 13084
rect 4692 13028 4696 13084
rect 4632 13024 4696 13028
rect 4712 13084 4776 13088
rect 4712 13028 4716 13084
rect 4716 13028 4772 13084
rect 4772 13028 4776 13084
rect 4712 13024 4776 13028
rect 4792 13084 4856 13088
rect 4792 13028 4796 13084
rect 4796 13028 4852 13084
rect 4852 13028 4856 13084
rect 4792 13024 4856 13028
rect 6152 13084 6216 13088
rect 6152 13028 6156 13084
rect 6156 13028 6212 13084
rect 6212 13028 6216 13084
rect 6152 13024 6216 13028
rect 6232 13084 6296 13088
rect 6232 13028 6236 13084
rect 6236 13028 6292 13084
rect 6292 13028 6296 13084
rect 6232 13024 6296 13028
rect 6312 13084 6376 13088
rect 6312 13028 6316 13084
rect 6316 13028 6372 13084
rect 6372 13028 6376 13084
rect 6312 13024 6376 13028
rect 6392 13084 6456 13088
rect 6392 13028 6396 13084
rect 6396 13028 6452 13084
rect 6452 13028 6456 13084
rect 6392 13024 6456 13028
rect 7752 13084 7816 13088
rect 7752 13028 7756 13084
rect 7756 13028 7812 13084
rect 7812 13028 7816 13084
rect 7752 13024 7816 13028
rect 7832 13084 7896 13088
rect 7832 13028 7836 13084
rect 7836 13028 7892 13084
rect 7892 13028 7896 13084
rect 7832 13024 7896 13028
rect 7912 13084 7976 13088
rect 7912 13028 7916 13084
rect 7916 13028 7972 13084
rect 7972 13028 7976 13084
rect 7912 13024 7976 13028
rect 7992 13084 8056 13088
rect 7992 13028 7996 13084
rect 7996 13028 8052 13084
rect 8052 13028 8056 13084
rect 7992 13024 8056 13028
rect 9352 13084 9416 13088
rect 9352 13028 9356 13084
rect 9356 13028 9412 13084
rect 9412 13028 9416 13084
rect 9352 13024 9416 13028
rect 9432 13084 9496 13088
rect 9432 13028 9436 13084
rect 9436 13028 9492 13084
rect 9492 13028 9496 13084
rect 9432 13024 9496 13028
rect 9512 13084 9576 13088
rect 9512 13028 9516 13084
rect 9516 13028 9572 13084
rect 9572 13028 9576 13084
rect 9512 13024 9576 13028
rect 9592 13084 9656 13088
rect 9592 13028 9596 13084
rect 9596 13028 9652 13084
rect 9652 13028 9656 13084
rect 9592 13024 9656 13028
rect 3612 12540 3676 12544
rect 3612 12484 3616 12540
rect 3616 12484 3672 12540
rect 3672 12484 3676 12540
rect 3612 12480 3676 12484
rect 3692 12540 3756 12544
rect 3692 12484 3696 12540
rect 3696 12484 3752 12540
rect 3752 12484 3756 12540
rect 3692 12480 3756 12484
rect 3772 12540 3836 12544
rect 3772 12484 3776 12540
rect 3776 12484 3832 12540
rect 3832 12484 3836 12540
rect 3772 12480 3836 12484
rect 3852 12540 3916 12544
rect 3852 12484 3856 12540
rect 3856 12484 3912 12540
rect 3912 12484 3916 12540
rect 3852 12480 3916 12484
rect 5212 12540 5276 12544
rect 5212 12484 5216 12540
rect 5216 12484 5272 12540
rect 5272 12484 5276 12540
rect 5212 12480 5276 12484
rect 5292 12540 5356 12544
rect 5292 12484 5296 12540
rect 5296 12484 5352 12540
rect 5352 12484 5356 12540
rect 5292 12480 5356 12484
rect 5372 12540 5436 12544
rect 5372 12484 5376 12540
rect 5376 12484 5432 12540
rect 5432 12484 5436 12540
rect 5372 12480 5436 12484
rect 5452 12540 5516 12544
rect 5452 12484 5456 12540
rect 5456 12484 5512 12540
rect 5512 12484 5516 12540
rect 5452 12480 5516 12484
rect 6812 12540 6876 12544
rect 6812 12484 6816 12540
rect 6816 12484 6872 12540
rect 6872 12484 6876 12540
rect 6812 12480 6876 12484
rect 6892 12540 6956 12544
rect 6892 12484 6896 12540
rect 6896 12484 6952 12540
rect 6952 12484 6956 12540
rect 6892 12480 6956 12484
rect 6972 12540 7036 12544
rect 6972 12484 6976 12540
rect 6976 12484 7032 12540
rect 7032 12484 7036 12540
rect 6972 12480 7036 12484
rect 7052 12540 7116 12544
rect 7052 12484 7056 12540
rect 7056 12484 7112 12540
rect 7112 12484 7116 12540
rect 7052 12480 7116 12484
rect 8412 12540 8476 12544
rect 8412 12484 8416 12540
rect 8416 12484 8472 12540
rect 8472 12484 8476 12540
rect 8412 12480 8476 12484
rect 8492 12540 8556 12544
rect 8492 12484 8496 12540
rect 8496 12484 8552 12540
rect 8552 12484 8556 12540
rect 8492 12480 8556 12484
rect 8572 12540 8636 12544
rect 8572 12484 8576 12540
rect 8576 12484 8632 12540
rect 8632 12484 8636 12540
rect 8572 12480 8636 12484
rect 8652 12540 8716 12544
rect 8652 12484 8656 12540
rect 8656 12484 8712 12540
rect 8712 12484 8716 12540
rect 8652 12480 8716 12484
rect 2952 11996 3016 12000
rect 2952 11940 2956 11996
rect 2956 11940 3012 11996
rect 3012 11940 3016 11996
rect 2952 11936 3016 11940
rect 3032 11996 3096 12000
rect 3032 11940 3036 11996
rect 3036 11940 3092 11996
rect 3092 11940 3096 11996
rect 3032 11936 3096 11940
rect 3112 11996 3176 12000
rect 3112 11940 3116 11996
rect 3116 11940 3172 11996
rect 3172 11940 3176 11996
rect 3112 11936 3176 11940
rect 3192 11996 3256 12000
rect 3192 11940 3196 11996
rect 3196 11940 3252 11996
rect 3252 11940 3256 11996
rect 3192 11936 3256 11940
rect 4552 11996 4616 12000
rect 4552 11940 4556 11996
rect 4556 11940 4612 11996
rect 4612 11940 4616 11996
rect 4552 11936 4616 11940
rect 4632 11996 4696 12000
rect 4632 11940 4636 11996
rect 4636 11940 4692 11996
rect 4692 11940 4696 11996
rect 4632 11936 4696 11940
rect 4712 11996 4776 12000
rect 4712 11940 4716 11996
rect 4716 11940 4772 11996
rect 4772 11940 4776 11996
rect 4712 11936 4776 11940
rect 4792 11996 4856 12000
rect 4792 11940 4796 11996
rect 4796 11940 4852 11996
rect 4852 11940 4856 11996
rect 4792 11936 4856 11940
rect 6152 11996 6216 12000
rect 6152 11940 6156 11996
rect 6156 11940 6212 11996
rect 6212 11940 6216 11996
rect 6152 11936 6216 11940
rect 6232 11996 6296 12000
rect 6232 11940 6236 11996
rect 6236 11940 6292 11996
rect 6292 11940 6296 11996
rect 6232 11936 6296 11940
rect 6312 11996 6376 12000
rect 6312 11940 6316 11996
rect 6316 11940 6372 11996
rect 6372 11940 6376 11996
rect 6312 11936 6376 11940
rect 6392 11996 6456 12000
rect 6392 11940 6396 11996
rect 6396 11940 6452 11996
rect 6452 11940 6456 11996
rect 6392 11936 6456 11940
rect 7752 11996 7816 12000
rect 7752 11940 7756 11996
rect 7756 11940 7812 11996
rect 7812 11940 7816 11996
rect 7752 11936 7816 11940
rect 7832 11996 7896 12000
rect 7832 11940 7836 11996
rect 7836 11940 7892 11996
rect 7892 11940 7896 11996
rect 7832 11936 7896 11940
rect 7912 11996 7976 12000
rect 7912 11940 7916 11996
rect 7916 11940 7972 11996
rect 7972 11940 7976 11996
rect 7912 11936 7976 11940
rect 7992 11996 8056 12000
rect 7992 11940 7996 11996
rect 7996 11940 8052 11996
rect 8052 11940 8056 11996
rect 7992 11936 8056 11940
rect 9352 11996 9416 12000
rect 9352 11940 9356 11996
rect 9356 11940 9412 11996
rect 9412 11940 9416 11996
rect 9352 11936 9416 11940
rect 9432 11996 9496 12000
rect 9432 11940 9436 11996
rect 9436 11940 9492 11996
rect 9492 11940 9496 11996
rect 9432 11936 9496 11940
rect 9512 11996 9576 12000
rect 9512 11940 9516 11996
rect 9516 11940 9572 11996
rect 9572 11940 9576 11996
rect 9512 11936 9576 11940
rect 9592 11996 9656 12000
rect 9592 11940 9596 11996
rect 9596 11940 9652 11996
rect 9652 11940 9656 11996
rect 9592 11936 9656 11940
rect 3612 11452 3676 11456
rect 3612 11396 3616 11452
rect 3616 11396 3672 11452
rect 3672 11396 3676 11452
rect 3612 11392 3676 11396
rect 3692 11452 3756 11456
rect 3692 11396 3696 11452
rect 3696 11396 3752 11452
rect 3752 11396 3756 11452
rect 3692 11392 3756 11396
rect 3772 11452 3836 11456
rect 3772 11396 3776 11452
rect 3776 11396 3832 11452
rect 3832 11396 3836 11452
rect 3772 11392 3836 11396
rect 3852 11452 3916 11456
rect 3852 11396 3856 11452
rect 3856 11396 3912 11452
rect 3912 11396 3916 11452
rect 3852 11392 3916 11396
rect 5212 11452 5276 11456
rect 5212 11396 5216 11452
rect 5216 11396 5272 11452
rect 5272 11396 5276 11452
rect 5212 11392 5276 11396
rect 5292 11452 5356 11456
rect 5292 11396 5296 11452
rect 5296 11396 5352 11452
rect 5352 11396 5356 11452
rect 5292 11392 5356 11396
rect 5372 11452 5436 11456
rect 5372 11396 5376 11452
rect 5376 11396 5432 11452
rect 5432 11396 5436 11452
rect 5372 11392 5436 11396
rect 5452 11452 5516 11456
rect 5452 11396 5456 11452
rect 5456 11396 5512 11452
rect 5512 11396 5516 11452
rect 5452 11392 5516 11396
rect 6812 11452 6876 11456
rect 6812 11396 6816 11452
rect 6816 11396 6872 11452
rect 6872 11396 6876 11452
rect 6812 11392 6876 11396
rect 6892 11452 6956 11456
rect 6892 11396 6896 11452
rect 6896 11396 6952 11452
rect 6952 11396 6956 11452
rect 6892 11392 6956 11396
rect 6972 11452 7036 11456
rect 6972 11396 6976 11452
rect 6976 11396 7032 11452
rect 7032 11396 7036 11452
rect 6972 11392 7036 11396
rect 7052 11452 7116 11456
rect 7052 11396 7056 11452
rect 7056 11396 7112 11452
rect 7112 11396 7116 11452
rect 7052 11392 7116 11396
rect 8412 11452 8476 11456
rect 8412 11396 8416 11452
rect 8416 11396 8472 11452
rect 8472 11396 8476 11452
rect 8412 11392 8476 11396
rect 8492 11452 8556 11456
rect 8492 11396 8496 11452
rect 8496 11396 8552 11452
rect 8552 11396 8556 11452
rect 8492 11392 8556 11396
rect 8572 11452 8636 11456
rect 8572 11396 8576 11452
rect 8576 11396 8632 11452
rect 8632 11396 8636 11452
rect 8572 11392 8636 11396
rect 8652 11452 8716 11456
rect 8652 11396 8656 11452
rect 8656 11396 8712 11452
rect 8712 11396 8716 11452
rect 8652 11392 8716 11396
rect 2952 10908 3016 10912
rect 2952 10852 2956 10908
rect 2956 10852 3012 10908
rect 3012 10852 3016 10908
rect 2952 10848 3016 10852
rect 3032 10908 3096 10912
rect 3032 10852 3036 10908
rect 3036 10852 3092 10908
rect 3092 10852 3096 10908
rect 3032 10848 3096 10852
rect 3112 10908 3176 10912
rect 3112 10852 3116 10908
rect 3116 10852 3172 10908
rect 3172 10852 3176 10908
rect 3112 10848 3176 10852
rect 3192 10908 3256 10912
rect 3192 10852 3196 10908
rect 3196 10852 3252 10908
rect 3252 10852 3256 10908
rect 3192 10848 3256 10852
rect 4552 10908 4616 10912
rect 4552 10852 4556 10908
rect 4556 10852 4612 10908
rect 4612 10852 4616 10908
rect 4552 10848 4616 10852
rect 4632 10908 4696 10912
rect 4632 10852 4636 10908
rect 4636 10852 4692 10908
rect 4692 10852 4696 10908
rect 4632 10848 4696 10852
rect 4712 10908 4776 10912
rect 4712 10852 4716 10908
rect 4716 10852 4772 10908
rect 4772 10852 4776 10908
rect 4712 10848 4776 10852
rect 4792 10908 4856 10912
rect 4792 10852 4796 10908
rect 4796 10852 4852 10908
rect 4852 10852 4856 10908
rect 4792 10848 4856 10852
rect 6152 10908 6216 10912
rect 6152 10852 6156 10908
rect 6156 10852 6212 10908
rect 6212 10852 6216 10908
rect 6152 10848 6216 10852
rect 6232 10908 6296 10912
rect 6232 10852 6236 10908
rect 6236 10852 6292 10908
rect 6292 10852 6296 10908
rect 6232 10848 6296 10852
rect 6312 10908 6376 10912
rect 6312 10852 6316 10908
rect 6316 10852 6372 10908
rect 6372 10852 6376 10908
rect 6312 10848 6376 10852
rect 6392 10908 6456 10912
rect 6392 10852 6396 10908
rect 6396 10852 6452 10908
rect 6452 10852 6456 10908
rect 6392 10848 6456 10852
rect 7752 10908 7816 10912
rect 7752 10852 7756 10908
rect 7756 10852 7812 10908
rect 7812 10852 7816 10908
rect 7752 10848 7816 10852
rect 7832 10908 7896 10912
rect 7832 10852 7836 10908
rect 7836 10852 7892 10908
rect 7892 10852 7896 10908
rect 7832 10848 7896 10852
rect 7912 10908 7976 10912
rect 7912 10852 7916 10908
rect 7916 10852 7972 10908
rect 7972 10852 7976 10908
rect 7912 10848 7976 10852
rect 7992 10908 8056 10912
rect 7992 10852 7996 10908
rect 7996 10852 8052 10908
rect 8052 10852 8056 10908
rect 7992 10848 8056 10852
rect 9352 10908 9416 10912
rect 9352 10852 9356 10908
rect 9356 10852 9412 10908
rect 9412 10852 9416 10908
rect 9352 10848 9416 10852
rect 9432 10908 9496 10912
rect 9432 10852 9436 10908
rect 9436 10852 9492 10908
rect 9492 10852 9496 10908
rect 9432 10848 9496 10852
rect 9512 10908 9576 10912
rect 9512 10852 9516 10908
rect 9516 10852 9572 10908
rect 9572 10852 9576 10908
rect 9512 10848 9576 10852
rect 9592 10908 9656 10912
rect 9592 10852 9596 10908
rect 9596 10852 9652 10908
rect 9652 10852 9656 10908
rect 9592 10848 9656 10852
rect 3612 10364 3676 10368
rect 3612 10308 3616 10364
rect 3616 10308 3672 10364
rect 3672 10308 3676 10364
rect 3612 10304 3676 10308
rect 3692 10364 3756 10368
rect 3692 10308 3696 10364
rect 3696 10308 3752 10364
rect 3752 10308 3756 10364
rect 3692 10304 3756 10308
rect 3772 10364 3836 10368
rect 3772 10308 3776 10364
rect 3776 10308 3832 10364
rect 3832 10308 3836 10364
rect 3772 10304 3836 10308
rect 3852 10364 3916 10368
rect 3852 10308 3856 10364
rect 3856 10308 3912 10364
rect 3912 10308 3916 10364
rect 3852 10304 3916 10308
rect 5212 10364 5276 10368
rect 5212 10308 5216 10364
rect 5216 10308 5272 10364
rect 5272 10308 5276 10364
rect 5212 10304 5276 10308
rect 5292 10364 5356 10368
rect 5292 10308 5296 10364
rect 5296 10308 5352 10364
rect 5352 10308 5356 10364
rect 5292 10304 5356 10308
rect 5372 10364 5436 10368
rect 5372 10308 5376 10364
rect 5376 10308 5432 10364
rect 5432 10308 5436 10364
rect 5372 10304 5436 10308
rect 5452 10364 5516 10368
rect 5452 10308 5456 10364
rect 5456 10308 5512 10364
rect 5512 10308 5516 10364
rect 5452 10304 5516 10308
rect 6812 10364 6876 10368
rect 6812 10308 6816 10364
rect 6816 10308 6872 10364
rect 6872 10308 6876 10364
rect 6812 10304 6876 10308
rect 6892 10364 6956 10368
rect 6892 10308 6896 10364
rect 6896 10308 6952 10364
rect 6952 10308 6956 10364
rect 6892 10304 6956 10308
rect 6972 10364 7036 10368
rect 6972 10308 6976 10364
rect 6976 10308 7032 10364
rect 7032 10308 7036 10364
rect 6972 10304 7036 10308
rect 7052 10364 7116 10368
rect 7052 10308 7056 10364
rect 7056 10308 7112 10364
rect 7112 10308 7116 10364
rect 7052 10304 7116 10308
rect 8412 10364 8476 10368
rect 8412 10308 8416 10364
rect 8416 10308 8472 10364
rect 8472 10308 8476 10364
rect 8412 10304 8476 10308
rect 8492 10364 8556 10368
rect 8492 10308 8496 10364
rect 8496 10308 8552 10364
rect 8552 10308 8556 10364
rect 8492 10304 8556 10308
rect 8572 10364 8636 10368
rect 8572 10308 8576 10364
rect 8576 10308 8632 10364
rect 8632 10308 8636 10364
rect 8572 10304 8636 10308
rect 8652 10364 8716 10368
rect 8652 10308 8656 10364
rect 8656 10308 8712 10364
rect 8712 10308 8716 10364
rect 8652 10304 8716 10308
rect 2952 9820 3016 9824
rect 2952 9764 2956 9820
rect 2956 9764 3012 9820
rect 3012 9764 3016 9820
rect 2952 9760 3016 9764
rect 3032 9820 3096 9824
rect 3032 9764 3036 9820
rect 3036 9764 3092 9820
rect 3092 9764 3096 9820
rect 3032 9760 3096 9764
rect 3112 9820 3176 9824
rect 3112 9764 3116 9820
rect 3116 9764 3172 9820
rect 3172 9764 3176 9820
rect 3112 9760 3176 9764
rect 3192 9820 3256 9824
rect 3192 9764 3196 9820
rect 3196 9764 3252 9820
rect 3252 9764 3256 9820
rect 3192 9760 3256 9764
rect 4552 9820 4616 9824
rect 4552 9764 4556 9820
rect 4556 9764 4612 9820
rect 4612 9764 4616 9820
rect 4552 9760 4616 9764
rect 4632 9820 4696 9824
rect 4632 9764 4636 9820
rect 4636 9764 4692 9820
rect 4692 9764 4696 9820
rect 4632 9760 4696 9764
rect 4712 9820 4776 9824
rect 4712 9764 4716 9820
rect 4716 9764 4772 9820
rect 4772 9764 4776 9820
rect 4712 9760 4776 9764
rect 4792 9820 4856 9824
rect 4792 9764 4796 9820
rect 4796 9764 4852 9820
rect 4852 9764 4856 9820
rect 4792 9760 4856 9764
rect 6152 9820 6216 9824
rect 6152 9764 6156 9820
rect 6156 9764 6212 9820
rect 6212 9764 6216 9820
rect 6152 9760 6216 9764
rect 6232 9820 6296 9824
rect 6232 9764 6236 9820
rect 6236 9764 6292 9820
rect 6292 9764 6296 9820
rect 6232 9760 6296 9764
rect 6312 9820 6376 9824
rect 6312 9764 6316 9820
rect 6316 9764 6372 9820
rect 6372 9764 6376 9820
rect 6312 9760 6376 9764
rect 6392 9820 6456 9824
rect 6392 9764 6396 9820
rect 6396 9764 6452 9820
rect 6452 9764 6456 9820
rect 6392 9760 6456 9764
rect 7752 9820 7816 9824
rect 7752 9764 7756 9820
rect 7756 9764 7812 9820
rect 7812 9764 7816 9820
rect 7752 9760 7816 9764
rect 7832 9820 7896 9824
rect 7832 9764 7836 9820
rect 7836 9764 7892 9820
rect 7892 9764 7896 9820
rect 7832 9760 7896 9764
rect 7912 9820 7976 9824
rect 7912 9764 7916 9820
rect 7916 9764 7972 9820
rect 7972 9764 7976 9820
rect 7912 9760 7976 9764
rect 7992 9820 8056 9824
rect 7992 9764 7996 9820
rect 7996 9764 8052 9820
rect 8052 9764 8056 9820
rect 7992 9760 8056 9764
rect 9352 9820 9416 9824
rect 9352 9764 9356 9820
rect 9356 9764 9412 9820
rect 9412 9764 9416 9820
rect 9352 9760 9416 9764
rect 9432 9820 9496 9824
rect 9432 9764 9436 9820
rect 9436 9764 9492 9820
rect 9492 9764 9496 9820
rect 9432 9760 9496 9764
rect 9512 9820 9576 9824
rect 9512 9764 9516 9820
rect 9516 9764 9572 9820
rect 9572 9764 9576 9820
rect 9512 9760 9576 9764
rect 9592 9820 9656 9824
rect 9592 9764 9596 9820
rect 9596 9764 9652 9820
rect 9652 9764 9656 9820
rect 9592 9760 9656 9764
rect 3612 9276 3676 9280
rect 3612 9220 3616 9276
rect 3616 9220 3672 9276
rect 3672 9220 3676 9276
rect 3612 9216 3676 9220
rect 3692 9276 3756 9280
rect 3692 9220 3696 9276
rect 3696 9220 3752 9276
rect 3752 9220 3756 9276
rect 3692 9216 3756 9220
rect 3772 9276 3836 9280
rect 3772 9220 3776 9276
rect 3776 9220 3832 9276
rect 3832 9220 3836 9276
rect 3772 9216 3836 9220
rect 3852 9276 3916 9280
rect 3852 9220 3856 9276
rect 3856 9220 3912 9276
rect 3912 9220 3916 9276
rect 3852 9216 3916 9220
rect 5212 9276 5276 9280
rect 5212 9220 5216 9276
rect 5216 9220 5272 9276
rect 5272 9220 5276 9276
rect 5212 9216 5276 9220
rect 5292 9276 5356 9280
rect 5292 9220 5296 9276
rect 5296 9220 5352 9276
rect 5352 9220 5356 9276
rect 5292 9216 5356 9220
rect 5372 9276 5436 9280
rect 5372 9220 5376 9276
rect 5376 9220 5432 9276
rect 5432 9220 5436 9276
rect 5372 9216 5436 9220
rect 5452 9276 5516 9280
rect 5452 9220 5456 9276
rect 5456 9220 5512 9276
rect 5512 9220 5516 9276
rect 5452 9216 5516 9220
rect 6812 9276 6876 9280
rect 6812 9220 6816 9276
rect 6816 9220 6872 9276
rect 6872 9220 6876 9276
rect 6812 9216 6876 9220
rect 6892 9276 6956 9280
rect 6892 9220 6896 9276
rect 6896 9220 6952 9276
rect 6952 9220 6956 9276
rect 6892 9216 6956 9220
rect 6972 9276 7036 9280
rect 6972 9220 6976 9276
rect 6976 9220 7032 9276
rect 7032 9220 7036 9276
rect 6972 9216 7036 9220
rect 7052 9276 7116 9280
rect 7052 9220 7056 9276
rect 7056 9220 7112 9276
rect 7112 9220 7116 9276
rect 7052 9216 7116 9220
rect 8412 9276 8476 9280
rect 8412 9220 8416 9276
rect 8416 9220 8472 9276
rect 8472 9220 8476 9276
rect 8412 9216 8476 9220
rect 8492 9276 8556 9280
rect 8492 9220 8496 9276
rect 8496 9220 8552 9276
rect 8552 9220 8556 9276
rect 8492 9216 8556 9220
rect 8572 9276 8636 9280
rect 8572 9220 8576 9276
rect 8576 9220 8632 9276
rect 8632 9220 8636 9276
rect 8572 9216 8636 9220
rect 8652 9276 8716 9280
rect 8652 9220 8656 9276
rect 8656 9220 8712 9276
rect 8712 9220 8716 9276
rect 8652 9216 8716 9220
rect 2952 8732 3016 8736
rect 2952 8676 2956 8732
rect 2956 8676 3012 8732
rect 3012 8676 3016 8732
rect 2952 8672 3016 8676
rect 3032 8732 3096 8736
rect 3032 8676 3036 8732
rect 3036 8676 3092 8732
rect 3092 8676 3096 8732
rect 3032 8672 3096 8676
rect 3112 8732 3176 8736
rect 3112 8676 3116 8732
rect 3116 8676 3172 8732
rect 3172 8676 3176 8732
rect 3112 8672 3176 8676
rect 3192 8732 3256 8736
rect 3192 8676 3196 8732
rect 3196 8676 3252 8732
rect 3252 8676 3256 8732
rect 3192 8672 3256 8676
rect 4552 8732 4616 8736
rect 4552 8676 4556 8732
rect 4556 8676 4612 8732
rect 4612 8676 4616 8732
rect 4552 8672 4616 8676
rect 4632 8732 4696 8736
rect 4632 8676 4636 8732
rect 4636 8676 4692 8732
rect 4692 8676 4696 8732
rect 4632 8672 4696 8676
rect 4712 8732 4776 8736
rect 4712 8676 4716 8732
rect 4716 8676 4772 8732
rect 4772 8676 4776 8732
rect 4712 8672 4776 8676
rect 4792 8732 4856 8736
rect 4792 8676 4796 8732
rect 4796 8676 4852 8732
rect 4852 8676 4856 8732
rect 4792 8672 4856 8676
rect 6152 8732 6216 8736
rect 6152 8676 6156 8732
rect 6156 8676 6212 8732
rect 6212 8676 6216 8732
rect 6152 8672 6216 8676
rect 6232 8732 6296 8736
rect 6232 8676 6236 8732
rect 6236 8676 6292 8732
rect 6292 8676 6296 8732
rect 6232 8672 6296 8676
rect 6312 8732 6376 8736
rect 6312 8676 6316 8732
rect 6316 8676 6372 8732
rect 6372 8676 6376 8732
rect 6312 8672 6376 8676
rect 6392 8732 6456 8736
rect 6392 8676 6396 8732
rect 6396 8676 6452 8732
rect 6452 8676 6456 8732
rect 6392 8672 6456 8676
rect 7752 8732 7816 8736
rect 7752 8676 7756 8732
rect 7756 8676 7812 8732
rect 7812 8676 7816 8732
rect 7752 8672 7816 8676
rect 7832 8732 7896 8736
rect 7832 8676 7836 8732
rect 7836 8676 7892 8732
rect 7892 8676 7896 8732
rect 7832 8672 7896 8676
rect 7912 8732 7976 8736
rect 7912 8676 7916 8732
rect 7916 8676 7972 8732
rect 7972 8676 7976 8732
rect 7912 8672 7976 8676
rect 7992 8732 8056 8736
rect 7992 8676 7996 8732
rect 7996 8676 8052 8732
rect 8052 8676 8056 8732
rect 7992 8672 8056 8676
rect 9352 8732 9416 8736
rect 9352 8676 9356 8732
rect 9356 8676 9412 8732
rect 9412 8676 9416 8732
rect 9352 8672 9416 8676
rect 9432 8732 9496 8736
rect 9432 8676 9436 8732
rect 9436 8676 9492 8732
rect 9492 8676 9496 8732
rect 9432 8672 9496 8676
rect 9512 8732 9576 8736
rect 9512 8676 9516 8732
rect 9516 8676 9572 8732
rect 9572 8676 9576 8732
rect 9512 8672 9576 8676
rect 9592 8732 9656 8736
rect 9592 8676 9596 8732
rect 9596 8676 9652 8732
rect 9652 8676 9656 8732
rect 9592 8672 9656 8676
rect 3612 8188 3676 8192
rect 3612 8132 3616 8188
rect 3616 8132 3672 8188
rect 3672 8132 3676 8188
rect 3612 8128 3676 8132
rect 3692 8188 3756 8192
rect 3692 8132 3696 8188
rect 3696 8132 3752 8188
rect 3752 8132 3756 8188
rect 3692 8128 3756 8132
rect 3772 8188 3836 8192
rect 3772 8132 3776 8188
rect 3776 8132 3832 8188
rect 3832 8132 3836 8188
rect 3772 8128 3836 8132
rect 3852 8188 3916 8192
rect 3852 8132 3856 8188
rect 3856 8132 3912 8188
rect 3912 8132 3916 8188
rect 3852 8128 3916 8132
rect 5212 8188 5276 8192
rect 5212 8132 5216 8188
rect 5216 8132 5272 8188
rect 5272 8132 5276 8188
rect 5212 8128 5276 8132
rect 5292 8188 5356 8192
rect 5292 8132 5296 8188
rect 5296 8132 5352 8188
rect 5352 8132 5356 8188
rect 5292 8128 5356 8132
rect 5372 8188 5436 8192
rect 5372 8132 5376 8188
rect 5376 8132 5432 8188
rect 5432 8132 5436 8188
rect 5372 8128 5436 8132
rect 5452 8188 5516 8192
rect 5452 8132 5456 8188
rect 5456 8132 5512 8188
rect 5512 8132 5516 8188
rect 5452 8128 5516 8132
rect 6812 8188 6876 8192
rect 6812 8132 6816 8188
rect 6816 8132 6872 8188
rect 6872 8132 6876 8188
rect 6812 8128 6876 8132
rect 6892 8188 6956 8192
rect 6892 8132 6896 8188
rect 6896 8132 6952 8188
rect 6952 8132 6956 8188
rect 6892 8128 6956 8132
rect 6972 8188 7036 8192
rect 6972 8132 6976 8188
rect 6976 8132 7032 8188
rect 7032 8132 7036 8188
rect 6972 8128 7036 8132
rect 7052 8188 7116 8192
rect 7052 8132 7056 8188
rect 7056 8132 7112 8188
rect 7112 8132 7116 8188
rect 7052 8128 7116 8132
rect 8412 8188 8476 8192
rect 8412 8132 8416 8188
rect 8416 8132 8472 8188
rect 8472 8132 8476 8188
rect 8412 8128 8476 8132
rect 8492 8188 8556 8192
rect 8492 8132 8496 8188
rect 8496 8132 8552 8188
rect 8552 8132 8556 8188
rect 8492 8128 8556 8132
rect 8572 8188 8636 8192
rect 8572 8132 8576 8188
rect 8576 8132 8632 8188
rect 8632 8132 8636 8188
rect 8572 8128 8636 8132
rect 8652 8188 8716 8192
rect 8652 8132 8656 8188
rect 8656 8132 8712 8188
rect 8712 8132 8716 8188
rect 8652 8128 8716 8132
rect 2952 7644 3016 7648
rect 2952 7588 2956 7644
rect 2956 7588 3012 7644
rect 3012 7588 3016 7644
rect 2952 7584 3016 7588
rect 3032 7644 3096 7648
rect 3032 7588 3036 7644
rect 3036 7588 3092 7644
rect 3092 7588 3096 7644
rect 3032 7584 3096 7588
rect 3112 7644 3176 7648
rect 3112 7588 3116 7644
rect 3116 7588 3172 7644
rect 3172 7588 3176 7644
rect 3112 7584 3176 7588
rect 3192 7644 3256 7648
rect 3192 7588 3196 7644
rect 3196 7588 3252 7644
rect 3252 7588 3256 7644
rect 3192 7584 3256 7588
rect 4552 7644 4616 7648
rect 4552 7588 4556 7644
rect 4556 7588 4612 7644
rect 4612 7588 4616 7644
rect 4552 7584 4616 7588
rect 4632 7644 4696 7648
rect 4632 7588 4636 7644
rect 4636 7588 4692 7644
rect 4692 7588 4696 7644
rect 4632 7584 4696 7588
rect 4712 7644 4776 7648
rect 4712 7588 4716 7644
rect 4716 7588 4772 7644
rect 4772 7588 4776 7644
rect 4712 7584 4776 7588
rect 4792 7644 4856 7648
rect 4792 7588 4796 7644
rect 4796 7588 4852 7644
rect 4852 7588 4856 7644
rect 4792 7584 4856 7588
rect 6152 7644 6216 7648
rect 6152 7588 6156 7644
rect 6156 7588 6212 7644
rect 6212 7588 6216 7644
rect 6152 7584 6216 7588
rect 6232 7644 6296 7648
rect 6232 7588 6236 7644
rect 6236 7588 6292 7644
rect 6292 7588 6296 7644
rect 6232 7584 6296 7588
rect 6312 7644 6376 7648
rect 6312 7588 6316 7644
rect 6316 7588 6372 7644
rect 6372 7588 6376 7644
rect 6312 7584 6376 7588
rect 6392 7644 6456 7648
rect 6392 7588 6396 7644
rect 6396 7588 6452 7644
rect 6452 7588 6456 7644
rect 6392 7584 6456 7588
rect 7752 7644 7816 7648
rect 7752 7588 7756 7644
rect 7756 7588 7812 7644
rect 7812 7588 7816 7644
rect 7752 7584 7816 7588
rect 7832 7644 7896 7648
rect 7832 7588 7836 7644
rect 7836 7588 7892 7644
rect 7892 7588 7896 7644
rect 7832 7584 7896 7588
rect 7912 7644 7976 7648
rect 7912 7588 7916 7644
rect 7916 7588 7972 7644
rect 7972 7588 7976 7644
rect 7912 7584 7976 7588
rect 7992 7644 8056 7648
rect 7992 7588 7996 7644
rect 7996 7588 8052 7644
rect 8052 7588 8056 7644
rect 7992 7584 8056 7588
rect 9352 7644 9416 7648
rect 9352 7588 9356 7644
rect 9356 7588 9412 7644
rect 9412 7588 9416 7644
rect 9352 7584 9416 7588
rect 9432 7644 9496 7648
rect 9432 7588 9436 7644
rect 9436 7588 9492 7644
rect 9492 7588 9496 7644
rect 9432 7584 9496 7588
rect 9512 7644 9576 7648
rect 9512 7588 9516 7644
rect 9516 7588 9572 7644
rect 9572 7588 9576 7644
rect 9512 7584 9576 7588
rect 9592 7644 9656 7648
rect 9592 7588 9596 7644
rect 9596 7588 9652 7644
rect 9652 7588 9656 7644
rect 9592 7584 9656 7588
rect 3612 7100 3676 7104
rect 3612 7044 3616 7100
rect 3616 7044 3672 7100
rect 3672 7044 3676 7100
rect 3612 7040 3676 7044
rect 3692 7100 3756 7104
rect 3692 7044 3696 7100
rect 3696 7044 3752 7100
rect 3752 7044 3756 7100
rect 3692 7040 3756 7044
rect 3772 7100 3836 7104
rect 3772 7044 3776 7100
rect 3776 7044 3832 7100
rect 3832 7044 3836 7100
rect 3772 7040 3836 7044
rect 3852 7100 3916 7104
rect 3852 7044 3856 7100
rect 3856 7044 3912 7100
rect 3912 7044 3916 7100
rect 3852 7040 3916 7044
rect 5212 7100 5276 7104
rect 5212 7044 5216 7100
rect 5216 7044 5272 7100
rect 5272 7044 5276 7100
rect 5212 7040 5276 7044
rect 5292 7100 5356 7104
rect 5292 7044 5296 7100
rect 5296 7044 5352 7100
rect 5352 7044 5356 7100
rect 5292 7040 5356 7044
rect 5372 7100 5436 7104
rect 5372 7044 5376 7100
rect 5376 7044 5432 7100
rect 5432 7044 5436 7100
rect 5372 7040 5436 7044
rect 5452 7100 5516 7104
rect 5452 7044 5456 7100
rect 5456 7044 5512 7100
rect 5512 7044 5516 7100
rect 5452 7040 5516 7044
rect 6812 7100 6876 7104
rect 6812 7044 6816 7100
rect 6816 7044 6872 7100
rect 6872 7044 6876 7100
rect 6812 7040 6876 7044
rect 6892 7100 6956 7104
rect 6892 7044 6896 7100
rect 6896 7044 6952 7100
rect 6952 7044 6956 7100
rect 6892 7040 6956 7044
rect 6972 7100 7036 7104
rect 6972 7044 6976 7100
rect 6976 7044 7032 7100
rect 7032 7044 7036 7100
rect 6972 7040 7036 7044
rect 7052 7100 7116 7104
rect 7052 7044 7056 7100
rect 7056 7044 7112 7100
rect 7112 7044 7116 7100
rect 7052 7040 7116 7044
rect 8412 7100 8476 7104
rect 8412 7044 8416 7100
rect 8416 7044 8472 7100
rect 8472 7044 8476 7100
rect 8412 7040 8476 7044
rect 8492 7100 8556 7104
rect 8492 7044 8496 7100
rect 8496 7044 8552 7100
rect 8552 7044 8556 7100
rect 8492 7040 8556 7044
rect 8572 7100 8636 7104
rect 8572 7044 8576 7100
rect 8576 7044 8632 7100
rect 8632 7044 8636 7100
rect 8572 7040 8636 7044
rect 8652 7100 8716 7104
rect 8652 7044 8656 7100
rect 8656 7044 8712 7100
rect 8712 7044 8716 7100
rect 8652 7040 8716 7044
rect 2952 6556 3016 6560
rect 2952 6500 2956 6556
rect 2956 6500 3012 6556
rect 3012 6500 3016 6556
rect 2952 6496 3016 6500
rect 3032 6556 3096 6560
rect 3032 6500 3036 6556
rect 3036 6500 3092 6556
rect 3092 6500 3096 6556
rect 3032 6496 3096 6500
rect 3112 6556 3176 6560
rect 3112 6500 3116 6556
rect 3116 6500 3172 6556
rect 3172 6500 3176 6556
rect 3112 6496 3176 6500
rect 3192 6556 3256 6560
rect 3192 6500 3196 6556
rect 3196 6500 3252 6556
rect 3252 6500 3256 6556
rect 3192 6496 3256 6500
rect 4552 6556 4616 6560
rect 4552 6500 4556 6556
rect 4556 6500 4612 6556
rect 4612 6500 4616 6556
rect 4552 6496 4616 6500
rect 4632 6556 4696 6560
rect 4632 6500 4636 6556
rect 4636 6500 4692 6556
rect 4692 6500 4696 6556
rect 4632 6496 4696 6500
rect 4712 6556 4776 6560
rect 4712 6500 4716 6556
rect 4716 6500 4772 6556
rect 4772 6500 4776 6556
rect 4712 6496 4776 6500
rect 4792 6556 4856 6560
rect 4792 6500 4796 6556
rect 4796 6500 4852 6556
rect 4852 6500 4856 6556
rect 4792 6496 4856 6500
rect 6152 6556 6216 6560
rect 6152 6500 6156 6556
rect 6156 6500 6212 6556
rect 6212 6500 6216 6556
rect 6152 6496 6216 6500
rect 6232 6556 6296 6560
rect 6232 6500 6236 6556
rect 6236 6500 6292 6556
rect 6292 6500 6296 6556
rect 6232 6496 6296 6500
rect 6312 6556 6376 6560
rect 6312 6500 6316 6556
rect 6316 6500 6372 6556
rect 6372 6500 6376 6556
rect 6312 6496 6376 6500
rect 6392 6556 6456 6560
rect 6392 6500 6396 6556
rect 6396 6500 6452 6556
rect 6452 6500 6456 6556
rect 6392 6496 6456 6500
rect 7752 6556 7816 6560
rect 7752 6500 7756 6556
rect 7756 6500 7812 6556
rect 7812 6500 7816 6556
rect 7752 6496 7816 6500
rect 7832 6556 7896 6560
rect 7832 6500 7836 6556
rect 7836 6500 7892 6556
rect 7892 6500 7896 6556
rect 7832 6496 7896 6500
rect 7912 6556 7976 6560
rect 7912 6500 7916 6556
rect 7916 6500 7972 6556
rect 7972 6500 7976 6556
rect 7912 6496 7976 6500
rect 7992 6556 8056 6560
rect 7992 6500 7996 6556
rect 7996 6500 8052 6556
rect 8052 6500 8056 6556
rect 7992 6496 8056 6500
rect 9352 6556 9416 6560
rect 9352 6500 9356 6556
rect 9356 6500 9412 6556
rect 9412 6500 9416 6556
rect 9352 6496 9416 6500
rect 9432 6556 9496 6560
rect 9432 6500 9436 6556
rect 9436 6500 9492 6556
rect 9492 6500 9496 6556
rect 9432 6496 9496 6500
rect 9512 6556 9576 6560
rect 9512 6500 9516 6556
rect 9516 6500 9572 6556
rect 9572 6500 9576 6556
rect 9512 6496 9576 6500
rect 9592 6556 9656 6560
rect 9592 6500 9596 6556
rect 9596 6500 9652 6556
rect 9652 6500 9656 6556
rect 9592 6496 9656 6500
rect 3612 6012 3676 6016
rect 3612 5956 3616 6012
rect 3616 5956 3672 6012
rect 3672 5956 3676 6012
rect 3612 5952 3676 5956
rect 3692 6012 3756 6016
rect 3692 5956 3696 6012
rect 3696 5956 3752 6012
rect 3752 5956 3756 6012
rect 3692 5952 3756 5956
rect 3772 6012 3836 6016
rect 3772 5956 3776 6012
rect 3776 5956 3832 6012
rect 3832 5956 3836 6012
rect 3772 5952 3836 5956
rect 3852 6012 3916 6016
rect 3852 5956 3856 6012
rect 3856 5956 3912 6012
rect 3912 5956 3916 6012
rect 3852 5952 3916 5956
rect 5212 6012 5276 6016
rect 5212 5956 5216 6012
rect 5216 5956 5272 6012
rect 5272 5956 5276 6012
rect 5212 5952 5276 5956
rect 5292 6012 5356 6016
rect 5292 5956 5296 6012
rect 5296 5956 5352 6012
rect 5352 5956 5356 6012
rect 5292 5952 5356 5956
rect 5372 6012 5436 6016
rect 5372 5956 5376 6012
rect 5376 5956 5432 6012
rect 5432 5956 5436 6012
rect 5372 5952 5436 5956
rect 5452 6012 5516 6016
rect 5452 5956 5456 6012
rect 5456 5956 5512 6012
rect 5512 5956 5516 6012
rect 5452 5952 5516 5956
rect 6812 6012 6876 6016
rect 6812 5956 6816 6012
rect 6816 5956 6872 6012
rect 6872 5956 6876 6012
rect 6812 5952 6876 5956
rect 6892 6012 6956 6016
rect 6892 5956 6896 6012
rect 6896 5956 6952 6012
rect 6952 5956 6956 6012
rect 6892 5952 6956 5956
rect 6972 6012 7036 6016
rect 6972 5956 6976 6012
rect 6976 5956 7032 6012
rect 7032 5956 7036 6012
rect 6972 5952 7036 5956
rect 7052 6012 7116 6016
rect 7052 5956 7056 6012
rect 7056 5956 7112 6012
rect 7112 5956 7116 6012
rect 7052 5952 7116 5956
rect 8412 6012 8476 6016
rect 8412 5956 8416 6012
rect 8416 5956 8472 6012
rect 8472 5956 8476 6012
rect 8412 5952 8476 5956
rect 8492 6012 8556 6016
rect 8492 5956 8496 6012
rect 8496 5956 8552 6012
rect 8552 5956 8556 6012
rect 8492 5952 8556 5956
rect 8572 6012 8636 6016
rect 8572 5956 8576 6012
rect 8576 5956 8632 6012
rect 8632 5956 8636 6012
rect 8572 5952 8636 5956
rect 8652 6012 8716 6016
rect 8652 5956 8656 6012
rect 8656 5956 8712 6012
rect 8712 5956 8716 6012
rect 8652 5952 8716 5956
rect 2952 5468 3016 5472
rect 2952 5412 2956 5468
rect 2956 5412 3012 5468
rect 3012 5412 3016 5468
rect 2952 5408 3016 5412
rect 3032 5468 3096 5472
rect 3032 5412 3036 5468
rect 3036 5412 3092 5468
rect 3092 5412 3096 5468
rect 3032 5408 3096 5412
rect 3112 5468 3176 5472
rect 3112 5412 3116 5468
rect 3116 5412 3172 5468
rect 3172 5412 3176 5468
rect 3112 5408 3176 5412
rect 3192 5468 3256 5472
rect 3192 5412 3196 5468
rect 3196 5412 3252 5468
rect 3252 5412 3256 5468
rect 3192 5408 3256 5412
rect 4552 5468 4616 5472
rect 4552 5412 4556 5468
rect 4556 5412 4612 5468
rect 4612 5412 4616 5468
rect 4552 5408 4616 5412
rect 4632 5468 4696 5472
rect 4632 5412 4636 5468
rect 4636 5412 4692 5468
rect 4692 5412 4696 5468
rect 4632 5408 4696 5412
rect 4712 5468 4776 5472
rect 4712 5412 4716 5468
rect 4716 5412 4772 5468
rect 4772 5412 4776 5468
rect 4712 5408 4776 5412
rect 4792 5468 4856 5472
rect 4792 5412 4796 5468
rect 4796 5412 4852 5468
rect 4852 5412 4856 5468
rect 4792 5408 4856 5412
rect 6152 5468 6216 5472
rect 6152 5412 6156 5468
rect 6156 5412 6212 5468
rect 6212 5412 6216 5468
rect 6152 5408 6216 5412
rect 6232 5468 6296 5472
rect 6232 5412 6236 5468
rect 6236 5412 6292 5468
rect 6292 5412 6296 5468
rect 6232 5408 6296 5412
rect 6312 5468 6376 5472
rect 6312 5412 6316 5468
rect 6316 5412 6372 5468
rect 6372 5412 6376 5468
rect 6312 5408 6376 5412
rect 6392 5468 6456 5472
rect 6392 5412 6396 5468
rect 6396 5412 6452 5468
rect 6452 5412 6456 5468
rect 6392 5408 6456 5412
rect 7752 5468 7816 5472
rect 7752 5412 7756 5468
rect 7756 5412 7812 5468
rect 7812 5412 7816 5468
rect 7752 5408 7816 5412
rect 7832 5468 7896 5472
rect 7832 5412 7836 5468
rect 7836 5412 7892 5468
rect 7892 5412 7896 5468
rect 7832 5408 7896 5412
rect 7912 5468 7976 5472
rect 7912 5412 7916 5468
rect 7916 5412 7972 5468
rect 7972 5412 7976 5468
rect 7912 5408 7976 5412
rect 7992 5468 8056 5472
rect 7992 5412 7996 5468
rect 7996 5412 8052 5468
rect 8052 5412 8056 5468
rect 7992 5408 8056 5412
rect 9352 5468 9416 5472
rect 9352 5412 9356 5468
rect 9356 5412 9412 5468
rect 9412 5412 9416 5468
rect 9352 5408 9416 5412
rect 9432 5468 9496 5472
rect 9432 5412 9436 5468
rect 9436 5412 9492 5468
rect 9492 5412 9496 5468
rect 9432 5408 9496 5412
rect 9512 5468 9576 5472
rect 9512 5412 9516 5468
rect 9516 5412 9572 5468
rect 9572 5412 9576 5468
rect 9512 5408 9576 5412
rect 9592 5468 9656 5472
rect 9592 5412 9596 5468
rect 9596 5412 9652 5468
rect 9652 5412 9656 5468
rect 9592 5408 9656 5412
rect 3612 4924 3676 4928
rect 3612 4868 3616 4924
rect 3616 4868 3672 4924
rect 3672 4868 3676 4924
rect 3612 4864 3676 4868
rect 3692 4924 3756 4928
rect 3692 4868 3696 4924
rect 3696 4868 3752 4924
rect 3752 4868 3756 4924
rect 3692 4864 3756 4868
rect 3772 4924 3836 4928
rect 3772 4868 3776 4924
rect 3776 4868 3832 4924
rect 3832 4868 3836 4924
rect 3772 4864 3836 4868
rect 3852 4924 3916 4928
rect 3852 4868 3856 4924
rect 3856 4868 3912 4924
rect 3912 4868 3916 4924
rect 3852 4864 3916 4868
rect 5212 4924 5276 4928
rect 5212 4868 5216 4924
rect 5216 4868 5272 4924
rect 5272 4868 5276 4924
rect 5212 4864 5276 4868
rect 5292 4924 5356 4928
rect 5292 4868 5296 4924
rect 5296 4868 5352 4924
rect 5352 4868 5356 4924
rect 5292 4864 5356 4868
rect 5372 4924 5436 4928
rect 5372 4868 5376 4924
rect 5376 4868 5432 4924
rect 5432 4868 5436 4924
rect 5372 4864 5436 4868
rect 5452 4924 5516 4928
rect 5452 4868 5456 4924
rect 5456 4868 5512 4924
rect 5512 4868 5516 4924
rect 5452 4864 5516 4868
rect 6812 4924 6876 4928
rect 6812 4868 6816 4924
rect 6816 4868 6872 4924
rect 6872 4868 6876 4924
rect 6812 4864 6876 4868
rect 6892 4924 6956 4928
rect 6892 4868 6896 4924
rect 6896 4868 6952 4924
rect 6952 4868 6956 4924
rect 6892 4864 6956 4868
rect 6972 4924 7036 4928
rect 6972 4868 6976 4924
rect 6976 4868 7032 4924
rect 7032 4868 7036 4924
rect 6972 4864 7036 4868
rect 7052 4924 7116 4928
rect 7052 4868 7056 4924
rect 7056 4868 7112 4924
rect 7112 4868 7116 4924
rect 7052 4864 7116 4868
rect 8412 4924 8476 4928
rect 8412 4868 8416 4924
rect 8416 4868 8472 4924
rect 8472 4868 8476 4924
rect 8412 4864 8476 4868
rect 8492 4924 8556 4928
rect 8492 4868 8496 4924
rect 8496 4868 8552 4924
rect 8552 4868 8556 4924
rect 8492 4864 8556 4868
rect 8572 4924 8636 4928
rect 8572 4868 8576 4924
rect 8576 4868 8632 4924
rect 8632 4868 8636 4924
rect 8572 4864 8636 4868
rect 8652 4924 8716 4928
rect 8652 4868 8656 4924
rect 8656 4868 8712 4924
rect 8712 4868 8716 4924
rect 8652 4864 8716 4868
rect 2952 4380 3016 4384
rect 2952 4324 2956 4380
rect 2956 4324 3012 4380
rect 3012 4324 3016 4380
rect 2952 4320 3016 4324
rect 3032 4380 3096 4384
rect 3032 4324 3036 4380
rect 3036 4324 3092 4380
rect 3092 4324 3096 4380
rect 3032 4320 3096 4324
rect 3112 4380 3176 4384
rect 3112 4324 3116 4380
rect 3116 4324 3172 4380
rect 3172 4324 3176 4380
rect 3112 4320 3176 4324
rect 3192 4380 3256 4384
rect 3192 4324 3196 4380
rect 3196 4324 3252 4380
rect 3252 4324 3256 4380
rect 3192 4320 3256 4324
rect 4552 4380 4616 4384
rect 4552 4324 4556 4380
rect 4556 4324 4612 4380
rect 4612 4324 4616 4380
rect 4552 4320 4616 4324
rect 4632 4380 4696 4384
rect 4632 4324 4636 4380
rect 4636 4324 4692 4380
rect 4692 4324 4696 4380
rect 4632 4320 4696 4324
rect 4712 4380 4776 4384
rect 4712 4324 4716 4380
rect 4716 4324 4772 4380
rect 4772 4324 4776 4380
rect 4712 4320 4776 4324
rect 4792 4380 4856 4384
rect 4792 4324 4796 4380
rect 4796 4324 4852 4380
rect 4852 4324 4856 4380
rect 4792 4320 4856 4324
rect 6152 4380 6216 4384
rect 6152 4324 6156 4380
rect 6156 4324 6212 4380
rect 6212 4324 6216 4380
rect 6152 4320 6216 4324
rect 6232 4380 6296 4384
rect 6232 4324 6236 4380
rect 6236 4324 6292 4380
rect 6292 4324 6296 4380
rect 6232 4320 6296 4324
rect 6312 4380 6376 4384
rect 6312 4324 6316 4380
rect 6316 4324 6372 4380
rect 6372 4324 6376 4380
rect 6312 4320 6376 4324
rect 6392 4380 6456 4384
rect 6392 4324 6396 4380
rect 6396 4324 6452 4380
rect 6452 4324 6456 4380
rect 6392 4320 6456 4324
rect 7752 4380 7816 4384
rect 7752 4324 7756 4380
rect 7756 4324 7812 4380
rect 7812 4324 7816 4380
rect 7752 4320 7816 4324
rect 7832 4380 7896 4384
rect 7832 4324 7836 4380
rect 7836 4324 7892 4380
rect 7892 4324 7896 4380
rect 7832 4320 7896 4324
rect 7912 4380 7976 4384
rect 7912 4324 7916 4380
rect 7916 4324 7972 4380
rect 7972 4324 7976 4380
rect 7912 4320 7976 4324
rect 7992 4380 8056 4384
rect 7992 4324 7996 4380
rect 7996 4324 8052 4380
rect 8052 4324 8056 4380
rect 7992 4320 8056 4324
rect 9352 4380 9416 4384
rect 9352 4324 9356 4380
rect 9356 4324 9412 4380
rect 9412 4324 9416 4380
rect 9352 4320 9416 4324
rect 9432 4380 9496 4384
rect 9432 4324 9436 4380
rect 9436 4324 9492 4380
rect 9492 4324 9496 4380
rect 9432 4320 9496 4324
rect 9512 4380 9576 4384
rect 9512 4324 9516 4380
rect 9516 4324 9572 4380
rect 9572 4324 9576 4380
rect 9512 4320 9576 4324
rect 9592 4380 9656 4384
rect 9592 4324 9596 4380
rect 9596 4324 9652 4380
rect 9652 4324 9656 4380
rect 9592 4320 9656 4324
rect 17854 3904 17918 3908
rect 17854 3848 17866 3904
rect 17866 3848 17918 3904
rect 17854 3844 17918 3848
rect 39206 3904 39270 3908
rect 39206 3848 39210 3904
rect 39210 3848 39266 3904
rect 39266 3848 39270 3904
rect 39206 3844 39270 3848
rect 40294 3904 40358 3908
rect 40294 3848 40314 3904
rect 40314 3848 40358 3904
rect 40294 3844 40358 3848
rect 45054 3904 45118 3908
rect 45054 3848 45062 3904
rect 45062 3848 45118 3904
rect 45054 3844 45118 3848
rect 46142 3904 46206 3908
rect 46142 3848 46166 3904
rect 46166 3848 46206 3904
rect 46142 3844 46206 3848
rect 50902 3904 50966 3908
rect 50902 3848 50950 3904
rect 50950 3848 50966 3904
rect 50902 3844 50966 3848
rect 54438 3904 54502 3908
rect 54438 3848 54446 3904
rect 54446 3848 54502 3904
rect 54438 3844 54502 3848
rect 93900 3844 93964 3908
rect 94966 3844 95030 3908
rect 3612 3836 3676 3840
rect 3612 3780 3616 3836
rect 3616 3780 3672 3836
rect 3672 3780 3676 3836
rect 3612 3776 3676 3780
rect 3692 3836 3756 3840
rect 3692 3780 3696 3836
rect 3696 3780 3752 3836
rect 3752 3780 3756 3836
rect 3692 3776 3756 3780
rect 3772 3836 3836 3840
rect 3772 3780 3776 3836
rect 3776 3780 3832 3836
rect 3832 3780 3836 3836
rect 3772 3776 3836 3780
rect 3852 3836 3916 3840
rect 3852 3780 3856 3836
rect 3856 3780 3912 3836
rect 3912 3780 3916 3836
rect 3852 3776 3916 3780
rect 5212 3836 5276 3840
rect 5212 3780 5216 3836
rect 5216 3780 5272 3836
rect 5272 3780 5276 3836
rect 5212 3776 5276 3780
rect 5292 3836 5356 3840
rect 5292 3780 5296 3836
rect 5296 3780 5352 3836
rect 5352 3780 5356 3836
rect 5292 3776 5356 3780
rect 5372 3836 5436 3840
rect 5372 3780 5376 3836
rect 5376 3780 5432 3836
rect 5432 3780 5436 3836
rect 5372 3776 5436 3780
rect 5452 3836 5516 3840
rect 5452 3780 5456 3836
rect 5456 3780 5512 3836
rect 5512 3780 5516 3836
rect 5452 3776 5516 3780
rect 6812 3836 6876 3840
rect 6812 3780 6816 3836
rect 6816 3780 6872 3836
rect 6872 3780 6876 3836
rect 6812 3776 6876 3780
rect 6892 3836 6956 3840
rect 6892 3780 6896 3836
rect 6896 3780 6952 3836
rect 6952 3780 6956 3836
rect 6892 3776 6956 3780
rect 6972 3836 7036 3840
rect 6972 3780 6976 3836
rect 6976 3780 7032 3836
rect 7032 3780 7036 3836
rect 6972 3776 7036 3780
rect 7052 3836 7116 3840
rect 7052 3780 7056 3836
rect 7056 3780 7112 3836
rect 7112 3780 7116 3836
rect 7052 3776 7116 3780
rect 8412 3836 8476 3840
rect 8412 3780 8416 3836
rect 8416 3780 8472 3836
rect 8472 3780 8476 3836
rect 8412 3776 8476 3780
rect 8492 3836 8556 3840
rect 8492 3780 8496 3836
rect 8496 3780 8552 3836
rect 8552 3780 8556 3836
rect 8492 3776 8556 3780
rect 8572 3836 8636 3840
rect 8572 3780 8576 3836
rect 8576 3780 8632 3836
rect 8632 3780 8636 3836
rect 8572 3776 8636 3780
rect 8652 3836 8716 3840
rect 8652 3780 8656 3836
rect 8656 3780 8712 3836
rect 8712 3780 8716 3836
rect 8652 3776 8716 3780
rect 28734 3768 28798 3772
rect 28734 3712 28778 3768
rect 28778 3712 28798 3768
rect 28734 3708 28798 3712
rect 29822 3768 29886 3772
rect 29822 3712 29826 3768
rect 29826 3712 29882 3768
rect 29882 3712 29886 3768
rect 29822 3708 29886 3712
rect 47502 3768 47566 3772
rect 47502 3712 47546 3768
rect 47546 3712 47566 3768
rect 47502 3708 47566 3712
rect 2952 3292 3016 3296
rect 2952 3236 2956 3292
rect 2956 3236 3012 3292
rect 3012 3236 3016 3292
rect 2952 3232 3016 3236
rect 3032 3292 3096 3296
rect 3032 3236 3036 3292
rect 3036 3236 3092 3292
rect 3092 3236 3096 3292
rect 3032 3232 3096 3236
rect 3112 3292 3176 3296
rect 3112 3236 3116 3292
rect 3116 3236 3172 3292
rect 3172 3236 3176 3292
rect 3112 3232 3176 3236
rect 3192 3292 3256 3296
rect 3192 3236 3196 3292
rect 3196 3236 3252 3292
rect 3252 3236 3256 3292
rect 3192 3232 3256 3236
rect 4552 3292 4616 3296
rect 4552 3236 4556 3292
rect 4556 3236 4612 3292
rect 4612 3236 4616 3292
rect 4552 3232 4616 3236
rect 4632 3292 4696 3296
rect 4632 3236 4636 3292
rect 4636 3236 4692 3292
rect 4692 3236 4696 3292
rect 4632 3232 4696 3236
rect 4712 3292 4776 3296
rect 4712 3236 4716 3292
rect 4716 3236 4772 3292
rect 4772 3236 4776 3292
rect 4712 3232 4776 3236
rect 4792 3292 4856 3296
rect 4792 3236 4796 3292
rect 4796 3236 4852 3292
rect 4852 3236 4856 3292
rect 4792 3232 4856 3236
rect 6152 3292 6216 3296
rect 6152 3236 6156 3292
rect 6156 3236 6212 3292
rect 6212 3236 6216 3292
rect 6152 3232 6216 3236
rect 6232 3292 6296 3296
rect 6232 3236 6236 3292
rect 6236 3236 6292 3292
rect 6292 3236 6296 3292
rect 6232 3232 6296 3236
rect 6312 3292 6376 3296
rect 6312 3236 6316 3292
rect 6316 3236 6372 3292
rect 6372 3236 6376 3292
rect 6312 3232 6376 3236
rect 6392 3292 6456 3296
rect 6392 3236 6396 3292
rect 6396 3236 6452 3292
rect 6452 3236 6456 3292
rect 6392 3232 6456 3236
rect 7752 3292 7816 3296
rect 7752 3236 7756 3292
rect 7756 3236 7812 3292
rect 7812 3236 7816 3292
rect 7752 3232 7816 3236
rect 7832 3292 7896 3296
rect 7832 3236 7836 3292
rect 7836 3236 7892 3292
rect 7892 3236 7896 3292
rect 7832 3232 7896 3236
rect 7912 3292 7976 3296
rect 7912 3236 7916 3292
rect 7916 3236 7972 3292
rect 7972 3236 7976 3292
rect 7912 3232 7976 3236
rect 7992 3292 8056 3296
rect 7992 3236 7996 3292
rect 7996 3236 8052 3292
rect 8052 3236 8056 3292
rect 7992 3232 8056 3236
rect 9352 3292 9416 3296
rect 9352 3236 9356 3292
rect 9356 3236 9412 3292
rect 9412 3236 9416 3292
rect 9352 3232 9416 3236
rect 9432 3292 9496 3296
rect 9432 3236 9436 3292
rect 9436 3236 9492 3292
rect 9492 3236 9496 3292
rect 9432 3232 9496 3236
rect 9512 3292 9576 3296
rect 9512 3236 9516 3292
rect 9516 3236 9572 3292
rect 9572 3236 9576 3292
rect 9512 3232 9576 3236
rect 9592 3292 9656 3296
rect 9592 3236 9596 3292
rect 9596 3236 9652 3292
rect 9652 3236 9656 3292
rect 9592 3232 9656 3236
rect 3612 2748 3676 2752
rect 3612 2692 3616 2748
rect 3616 2692 3672 2748
rect 3672 2692 3676 2748
rect 3612 2688 3676 2692
rect 3692 2748 3756 2752
rect 3692 2692 3696 2748
rect 3696 2692 3752 2748
rect 3752 2692 3756 2748
rect 3692 2688 3756 2692
rect 3772 2748 3836 2752
rect 3772 2692 3776 2748
rect 3776 2692 3832 2748
rect 3832 2692 3836 2748
rect 3772 2688 3836 2692
rect 3852 2748 3916 2752
rect 3852 2692 3856 2748
rect 3856 2692 3912 2748
rect 3912 2692 3916 2748
rect 3852 2688 3916 2692
rect 5212 2748 5276 2752
rect 5212 2692 5216 2748
rect 5216 2692 5272 2748
rect 5272 2692 5276 2748
rect 5212 2688 5276 2692
rect 5292 2748 5356 2752
rect 5292 2692 5296 2748
rect 5296 2692 5352 2748
rect 5352 2692 5356 2748
rect 5292 2688 5356 2692
rect 5372 2748 5436 2752
rect 5372 2692 5376 2748
rect 5376 2692 5432 2748
rect 5432 2692 5436 2748
rect 5372 2688 5436 2692
rect 5452 2748 5516 2752
rect 5452 2692 5456 2748
rect 5456 2692 5512 2748
rect 5512 2692 5516 2748
rect 5452 2688 5516 2692
rect 6812 2748 6876 2752
rect 6812 2692 6816 2748
rect 6816 2692 6872 2748
rect 6872 2692 6876 2748
rect 6812 2688 6876 2692
rect 6892 2748 6956 2752
rect 6892 2692 6896 2748
rect 6896 2692 6952 2748
rect 6952 2692 6956 2748
rect 6892 2688 6956 2692
rect 6972 2748 7036 2752
rect 6972 2692 6976 2748
rect 6976 2692 7032 2748
rect 7032 2692 7036 2748
rect 6972 2688 7036 2692
rect 7052 2748 7116 2752
rect 7052 2692 7056 2748
rect 7056 2692 7112 2748
rect 7112 2692 7116 2748
rect 7052 2688 7116 2692
rect 8412 2748 8476 2752
rect 8412 2692 8416 2748
rect 8416 2692 8472 2748
rect 8472 2692 8476 2748
rect 8412 2688 8476 2692
rect 8492 2748 8556 2752
rect 8492 2692 8496 2748
rect 8496 2692 8552 2748
rect 8552 2692 8556 2748
rect 8492 2688 8556 2692
rect 8572 2748 8636 2752
rect 8572 2692 8576 2748
rect 8576 2692 8632 2748
rect 8632 2692 8636 2748
rect 8572 2688 8636 2692
rect 8652 2748 8716 2752
rect 8652 2692 8656 2748
rect 8656 2692 8712 2748
rect 8712 2692 8716 2748
rect 8652 2688 8716 2692
rect 11836 2620 11900 2684
rect 35572 2620 35636 2684
rect 37044 2680 37108 2684
rect 37044 2624 37058 2680
rect 37058 2624 37108 2680
rect 37044 2620 37108 2624
rect 49740 2680 49804 2684
rect 49740 2624 49754 2680
rect 49754 2624 49804 2680
rect 49740 2620 49804 2624
rect 55444 2680 55508 2684
rect 55444 2624 55458 2680
rect 55458 2624 55508 2680
rect 55444 2620 55508 2624
rect 58020 2680 58084 2684
rect 58020 2624 58034 2680
rect 58034 2624 58084 2680
rect 58020 2620 58084 2624
rect 94820 2484 94884 2548
rect 95004 2544 95068 2548
rect 95004 2488 95018 2544
rect 95018 2488 95068 2544
rect 95004 2484 95068 2488
rect 32076 2408 32140 2412
rect 32076 2352 32090 2408
rect 32090 2352 32140 2408
rect 32076 2348 32140 2352
rect 42748 2408 42812 2412
rect 42748 2352 42798 2408
rect 42798 2352 42812 2408
rect 42748 2348 42812 2352
rect 43852 2408 43916 2412
rect 43852 2352 43866 2408
rect 43866 2352 43916 2408
rect 43852 2348 43916 2352
rect 48636 2408 48700 2412
rect 48636 2352 48650 2408
rect 48650 2352 48700 2408
rect 48636 2348 48700 2352
rect 2952 2204 3016 2208
rect 2952 2148 2956 2204
rect 2956 2148 3012 2204
rect 3012 2148 3016 2204
rect 2952 2144 3016 2148
rect 3032 2204 3096 2208
rect 3032 2148 3036 2204
rect 3036 2148 3092 2204
rect 3092 2148 3096 2204
rect 3032 2144 3096 2148
rect 3112 2204 3176 2208
rect 3112 2148 3116 2204
rect 3116 2148 3172 2204
rect 3172 2148 3176 2204
rect 3112 2144 3176 2148
rect 3192 2204 3256 2208
rect 3192 2148 3196 2204
rect 3196 2148 3252 2204
rect 3252 2148 3256 2204
rect 3192 2144 3256 2148
rect 4552 2204 4616 2208
rect 4552 2148 4556 2204
rect 4556 2148 4612 2204
rect 4612 2148 4616 2204
rect 4552 2144 4616 2148
rect 4632 2204 4696 2208
rect 4632 2148 4636 2204
rect 4636 2148 4692 2204
rect 4692 2148 4696 2204
rect 4632 2144 4696 2148
rect 4712 2204 4776 2208
rect 4712 2148 4716 2204
rect 4716 2148 4772 2204
rect 4772 2148 4776 2204
rect 4712 2144 4776 2148
rect 4792 2204 4856 2208
rect 4792 2148 4796 2204
rect 4796 2148 4852 2204
rect 4852 2148 4856 2204
rect 4792 2144 4856 2148
rect 6152 2204 6216 2208
rect 6152 2148 6156 2204
rect 6156 2148 6212 2204
rect 6212 2148 6216 2204
rect 6152 2144 6216 2148
rect 6232 2204 6296 2208
rect 6232 2148 6236 2204
rect 6236 2148 6292 2204
rect 6292 2148 6296 2204
rect 6232 2144 6296 2148
rect 6312 2204 6376 2208
rect 6312 2148 6316 2204
rect 6316 2148 6372 2204
rect 6372 2148 6376 2204
rect 6312 2144 6376 2148
rect 6392 2204 6456 2208
rect 6392 2148 6396 2204
rect 6396 2148 6452 2204
rect 6452 2148 6456 2204
rect 6392 2144 6456 2148
rect 7752 2204 7816 2208
rect 7752 2148 7756 2204
rect 7756 2148 7812 2204
rect 7812 2148 7816 2204
rect 7752 2144 7816 2148
rect 7832 2204 7896 2208
rect 7832 2148 7836 2204
rect 7836 2148 7892 2204
rect 7892 2148 7896 2204
rect 7832 2144 7896 2148
rect 7912 2204 7976 2208
rect 7912 2148 7916 2204
rect 7916 2148 7972 2204
rect 7972 2148 7976 2204
rect 7912 2144 7976 2148
rect 7992 2204 8056 2208
rect 7992 2148 7996 2204
rect 7996 2148 8052 2204
rect 8052 2148 8056 2204
rect 7992 2144 8056 2148
rect 9352 2204 9416 2208
rect 9352 2148 9356 2204
rect 9356 2148 9412 2204
rect 9412 2148 9416 2204
rect 9352 2144 9416 2148
rect 9432 2204 9496 2208
rect 9432 2148 9436 2204
rect 9436 2148 9492 2204
rect 9492 2148 9496 2204
rect 9432 2144 9496 2148
rect 9512 2204 9576 2208
rect 9512 2148 9516 2204
rect 9516 2148 9572 2204
rect 9572 2148 9576 2204
rect 9512 2144 9576 2148
rect 9592 2204 9656 2208
rect 9592 2148 9596 2204
rect 9596 2148 9652 2204
rect 9652 2148 9656 2204
rect 9592 2144 9656 2148
rect 11652 2076 11716 2140
rect 94636 1940 94700 2004
rect 3612 1660 3676 1664
rect 3612 1604 3616 1660
rect 3616 1604 3672 1660
rect 3672 1604 3676 1660
rect 3612 1600 3676 1604
rect 3692 1660 3756 1664
rect 3692 1604 3696 1660
rect 3696 1604 3752 1660
rect 3752 1604 3756 1660
rect 3692 1600 3756 1604
rect 3772 1660 3836 1664
rect 3772 1604 3776 1660
rect 3776 1604 3832 1660
rect 3832 1604 3836 1660
rect 3772 1600 3836 1604
rect 3852 1660 3916 1664
rect 3852 1604 3856 1660
rect 3856 1604 3912 1660
rect 3912 1604 3916 1660
rect 3852 1600 3916 1604
rect 5212 1660 5276 1664
rect 5212 1604 5216 1660
rect 5216 1604 5272 1660
rect 5272 1604 5276 1660
rect 5212 1600 5276 1604
rect 5292 1660 5356 1664
rect 5292 1604 5296 1660
rect 5296 1604 5352 1660
rect 5352 1604 5356 1660
rect 5292 1600 5356 1604
rect 5372 1660 5436 1664
rect 5372 1604 5376 1660
rect 5376 1604 5432 1660
rect 5432 1604 5436 1660
rect 5372 1600 5436 1604
rect 5452 1660 5516 1664
rect 5452 1604 5456 1660
rect 5456 1604 5512 1660
rect 5512 1604 5516 1660
rect 5452 1600 5516 1604
rect 6812 1660 6876 1664
rect 6812 1604 6816 1660
rect 6816 1604 6872 1660
rect 6872 1604 6876 1660
rect 6812 1600 6876 1604
rect 6892 1660 6956 1664
rect 6892 1604 6896 1660
rect 6896 1604 6952 1660
rect 6952 1604 6956 1660
rect 6892 1600 6956 1604
rect 6972 1660 7036 1664
rect 6972 1604 6976 1660
rect 6976 1604 7032 1660
rect 7032 1604 7036 1660
rect 6972 1600 7036 1604
rect 7052 1660 7116 1664
rect 7052 1604 7056 1660
rect 7056 1604 7112 1660
rect 7112 1604 7116 1660
rect 7052 1600 7116 1604
rect 8412 1660 8476 1664
rect 8412 1604 8416 1660
rect 8416 1604 8472 1660
rect 8472 1604 8476 1660
rect 8412 1600 8476 1604
rect 8492 1660 8556 1664
rect 8492 1604 8496 1660
rect 8496 1604 8552 1660
rect 8552 1604 8556 1660
rect 8492 1600 8556 1604
rect 8572 1660 8636 1664
rect 8572 1604 8576 1660
rect 8576 1604 8632 1660
rect 8632 1604 8636 1660
rect 8572 1600 8636 1604
rect 8652 1660 8716 1664
rect 8652 1604 8656 1660
rect 8656 1604 8712 1660
rect 8712 1604 8716 1660
rect 8652 1600 8716 1604
rect 10012 1660 10076 1664
rect 10012 1604 10016 1660
rect 10016 1604 10072 1660
rect 10072 1604 10076 1660
rect 10012 1600 10076 1604
rect 10092 1660 10156 1664
rect 10092 1604 10096 1660
rect 10096 1604 10152 1660
rect 10152 1604 10156 1660
rect 10092 1600 10156 1604
rect 10172 1660 10236 1664
rect 10172 1604 10176 1660
rect 10176 1604 10232 1660
rect 10232 1604 10236 1660
rect 10172 1600 10236 1604
rect 10252 1660 10316 1664
rect 10252 1604 10256 1660
rect 10256 1604 10312 1660
rect 10312 1604 10316 1660
rect 10252 1600 10316 1604
rect 11612 1660 11676 1664
rect 11612 1604 11616 1660
rect 11616 1604 11672 1660
rect 11672 1604 11676 1660
rect 11612 1600 11676 1604
rect 11692 1660 11756 1664
rect 11692 1604 11696 1660
rect 11696 1604 11752 1660
rect 11752 1604 11756 1660
rect 11692 1600 11756 1604
rect 11772 1660 11836 1664
rect 11772 1604 11776 1660
rect 11776 1604 11832 1660
rect 11832 1604 11836 1660
rect 11772 1600 11836 1604
rect 11852 1660 11916 1664
rect 11852 1604 11856 1660
rect 11856 1604 11912 1660
rect 11912 1604 11916 1660
rect 11852 1600 11916 1604
rect 13212 1660 13276 1664
rect 13212 1604 13216 1660
rect 13216 1604 13272 1660
rect 13272 1604 13276 1660
rect 13212 1600 13276 1604
rect 13292 1660 13356 1664
rect 13292 1604 13296 1660
rect 13296 1604 13352 1660
rect 13352 1604 13356 1660
rect 13292 1600 13356 1604
rect 13372 1660 13436 1664
rect 13372 1604 13376 1660
rect 13376 1604 13432 1660
rect 13432 1604 13436 1660
rect 13372 1600 13436 1604
rect 13452 1660 13516 1664
rect 13452 1604 13456 1660
rect 13456 1604 13512 1660
rect 13512 1604 13516 1660
rect 13452 1600 13516 1604
rect 14812 1660 14876 1664
rect 14812 1604 14816 1660
rect 14816 1604 14872 1660
rect 14872 1604 14876 1660
rect 14812 1600 14876 1604
rect 14892 1660 14956 1664
rect 14892 1604 14896 1660
rect 14896 1604 14952 1660
rect 14952 1604 14956 1660
rect 14892 1600 14956 1604
rect 14972 1660 15036 1664
rect 14972 1604 14976 1660
rect 14976 1604 15032 1660
rect 15032 1604 15036 1660
rect 14972 1600 15036 1604
rect 15052 1660 15116 1664
rect 15052 1604 15056 1660
rect 15056 1604 15112 1660
rect 15112 1604 15116 1660
rect 15052 1600 15116 1604
rect 16412 1660 16476 1664
rect 16412 1604 16416 1660
rect 16416 1604 16472 1660
rect 16472 1604 16476 1660
rect 16412 1600 16476 1604
rect 16492 1660 16556 1664
rect 16492 1604 16496 1660
rect 16496 1604 16552 1660
rect 16552 1604 16556 1660
rect 16492 1600 16556 1604
rect 16572 1660 16636 1664
rect 16572 1604 16576 1660
rect 16576 1604 16632 1660
rect 16632 1604 16636 1660
rect 16572 1600 16636 1604
rect 16652 1660 16716 1664
rect 16652 1604 16656 1660
rect 16656 1604 16712 1660
rect 16712 1604 16716 1660
rect 16652 1600 16716 1604
rect 18012 1660 18076 1664
rect 18012 1604 18016 1660
rect 18016 1604 18072 1660
rect 18072 1604 18076 1660
rect 18012 1600 18076 1604
rect 18092 1660 18156 1664
rect 18092 1604 18096 1660
rect 18096 1604 18152 1660
rect 18152 1604 18156 1660
rect 18092 1600 18156 1604
rect 18172 1660 18236 1664
rect 18172 1604 18176 1660
rect 18176 1604 18232 1660
rect 18232 1604 18236 1660
rect 18172 1600 18236 1604
rect 18252 1660 18316 1664
rect 18252 1604 18256 1660
rect 18256 1604 18312 1660
rect 18312 1604 18316 1660
rect 18252 1600 18316 1604
rect 19612 1660 19676 1664
rect 19612 1604 19616 1660
rect 19616 1604 19672 1660
rect 19672 1604 19676 1660
rect 19612 1600 19676 1604
rect 19692 1660 19756 1664
rect 19692 1604 19696 1660
rect 19696 1604 19752 1660
rect 19752 1604 19756 1660
rect 19692 1600 19756 1604
rect 19772 1660 19836 1664
rect 19772 1604 19776 1660
rect 19776 1604 19832 1660
rect 19832 1604 19836 1660
rect 19772 1600 19836 1604
rect 19852 1660 19916 1664
rect 19852 1604 19856 1660
rect 19856 1604 19912 1660
rect 19912 1604 19916 1660
rect 19852 1600 19916 1604
rect 21212 1660 21276 1664
rect 21212 1604 21216 1660
rect 21216 1604 21272 1660
rect 21272 1604 21276 1660
rect 21212 1600 21276 1604
rect 21292 1660 21356 1664
rect 21292 1604 21296 1660
rect 21296 1604 21352 1660
rect 21352 1604 21356 1660
rect 21292 1600 21356 1604
rect 21372 1660 21436 1664
rect 21372 1604 21376 1660
rect 21376 1604 21432 1660
rect 21432 1604 21436 1660
rect 21372 1600 21436 1604
rect 21452 1660 21516 1664
rect 21452 1604 21456 1660
rect 21456 1604 21512 1660
rect 21512 1604 21516 1660
rect 21452 1600 21516 1604
rect 22812 1660 22876 1664
rect 22812 1604 22816 1660
rect 22816 1604 22872 1660
rect 22872 1604 22876 1660
rect 22812 1600 22876 1604
rect 22892 1660 22956 1664
rect 22892 1604 22896 1660
rect 22896 1604 22952 1660
rect 22952 1604 22956 1660
rect 22892 1600 22956 1604
rect 22972 1660 23036 1664
rect 22972 1604 22976 1660
rect 22976 1604 23032 1660
rect 23032 1604 23036 1660
rect 22972 1600 23036 1604
rect 23052 1660 23116 1664
rect 23052 1604 23056 1660
rect 23056 1604 23112 1660
rect 23112 1604 23116 1660
rect 23052 1600 23116 1604
rect 24412 1660 24476 1664
rect 24412 1604 24416 1660
rect 24416 1604 24472 1660
rect 24472 1604 24476 1660
rect 24412 1600 24476 1604
rect 24492 1660 24556 1664
rect 24492 1604 24496 1660
rect 24496 1604 24552 1660
rect 24552 1604 24556 1660
rect 24492 1600 24556 1604
rect 24572 1660 24636 1664
rect 24572 1604 24576 1660
rect 24576 1604 24632 1660
rect 24632 1604 24636 1660
rect 24572 1600 24636 1604
rect 24652 1660 24716 1664
rect 24652 1604 24656 1660
rect 24656 1604 24712 1660
rect 24712 1604 24716 1660
rect 24652 1600 24716 1604
rect 26012 1660 26076 1664
rect 26012 1604 26016 1660
rect 26016 1604 26072 1660
rect 26072 1604 26076 1660
rect 26012 1600 26076 1604
rect 26092 1660 26156 1664
rect 26092 1604 26096 1660
rect 26096 1604 26152 1660
rect 26152 1604 26156 1660
rect 26092 1600 26156 1604
rect 26172 1660 26236 1664
rect 26172 1604 26176 1660
rect 26176 1604 26232 1660
rect 26232 1604 26236 1660
rect 26172 1600 26236 1604
rect 26252 1660 26316 1664
rect 26252 1604 26256 1660
rect 26256 1604 26312 1660
rect 26312 1604 26316 1660
rect 26252 1600 26316 1604
rect 27612 1660 27676 1664
rect 27612 1604 27616 1660
rect 27616 1604 27672 1660
rect 27672 1604 27676 1660
rect 27612 1600 27676 1604
rect 27692 1660 27756 1664
rect 27692 1604 27696 1660
rect 27696 1604 27752 1660
rect 27752 1604 27756 1660
rect 27692 1600 27756 1604
rect 27772 1660 27836 1664
rect 27772 1604 27776 1660
rect 27776 1604 27832 1660
rect 27832 1604 27836 1660
rect 27772 1600 27836 1604
rect 27852 1660 27916 1664
rect 27852 1604 27856 1660
rect 27856 1604 27912 1660
rect 27912 1604 27916 1660
rect 27852 1600 27916 1604
rect 29212 1660 29276 1664
rect 29212 1604 29216 1660
rect 29216 1604 29272 1660
rect 29272 1604 29276 1660
rect 29212 1600 29276 1604
rect 29292 1660 29356 1664
rect 29292 1604 29296 1660
rect 29296 1604 29352 1660
rect 29352 1604 29356 1660
rect 29292 1600 29356 1604
rect 29372 1660 29436 1664
rect 29372 1604 29376 1660
rect 29376 1604 29432 1660
rect 29432 1604 29436 1660
rect 29372 1600 29436 1604
rect 29452 1660 29516 1664
rect 29452 1604 29456 1660
rect 29456 1604 29512 1660
rect 29512 1604 29516 1660
rect 29452 1600 29516 1604
rect 30812 1660 30876 1664
rect 30812 1604 30816 1660
rect 30816 1604 30872 1660
rect 30872 1604 30876 1660
rect 30812 1600 30876 1604
rect 30892 1660 30956 1664
rect 30892 1604 30896 1660
rect 30896 1604 30952 1660
rect 30952 1604 30956 1660
rect 30892 1600 30956 1604
rect 30972 1660 31036 1664
rect 30972 1604 30976 1660
rect 30976 1604 31032 1660
rect 31032 1604 31036 1660
rect 30972 1600 31036 1604
rect 31052 1660 31116 1664
rect 31052 1604 31056 1660
rect 31056 1604 31112 1660
rect 31112 1604 31116 1660
rect 31052 1600 31116 1604
rect 32412 1660 32476 1664
rect 32412 1604 32416 1660
rect 32416 1604 32472 1660
rect 32472 1604 32476 1660
rect 32412 1600 32476 1604
rect 32492 1660 32556 1664
rect 32492 1604 32496 1660
rect 32496 1604 32552 1660
rect 32552 1604 32556 1660
rect 32492 1600 32556 1604
rect 32572 1660 32636 1664
rect 32572 1604 32576 1660
rect 32576 1604 32632 1660
rect 32632 1604 32636 1660
rect 32572 1600 32636 1604
rect 32652 1660 32716 1664
rect 32652 1604 32656 1660
rect 32656 1604 32712 1660
rect 32712 1604 32716 1660
rect 32652 1600 32716 1604
rect 34012 1660 34076 1664
rect 34012 1604 34016 1660
rect 34016 1604 34072 1660
rect 34072 1604 34076 1660
rect 34012 1600 34076 1604
rect 34092 1660 34156 1664
rect 34092 1604 34096 1660
rect 34096 1604 34152 1660
rect 34152 1604 34156 1660
rect 34092 1600 34156 1604
rect 34172 1660 34236 1664
rect 34172 1604 34176 1660
rect 34176 1604 34232 1660
rect 34232 1604 34236 1660
rect 34172 1600 34236 1604
rect 34252 1660 34316 1664
rect 34252 1604 34256 1660
rect 34256 1604 34312 1660
rect 34312 1604 34316 1660
rect 34252 1600 34316 1604
rect 35612 1660 35676 1664
rect 35612 1604 35616 1660
rect 35616 1604 35672 1660
rect 35672 1604 35676 1660
rect 35612 1600 35676 1604
rect 35692 1660 35756 1664
rect 35692 1604 35696 1660
rect 35696 1604 35752 1660
rect 35752 1604 35756 1660
rect 35692 1600 35756 1604
rect 35772 1660 35836 1664
rect 35772 1604 35776 1660
rect 35776 1604 35832 1660
rect 35832 1604 35836 1660
rect 35772 1600 35836 1604
rect 35852 1660 35916 1664
rect 35852 1604 35856 1660
rect 35856 1604 35912 1660
rect 35912 1604 35916 1660
rect 35852 1600 35916 1604
rect 37212 1660 37276 1664
rect 37212 1604 37216 1660
rect 37216 1604 37272 1660
rect 37272 1604 37276 1660
rect 37212 1600 37276 1604
rect 37292 1660 37356 1664
rect 37292 1604 37296 1660
rect 37296 1604 37352 1660
rect 37352 1604 37356 1660
rect 37292 1600 37356 1604
rect 37372 1660 37436 1664
rect 37372 1604 37376 1660
rect 37376 1604 37432 1660
rect 37432 1604 37436 1660
rect 37372 1600 37436 1604
rect 37452 1660 37516 1664
rect 37452 1604 37456 1660
rect 37456 1604 37512 1660
rect 37512 1604 37516 1660
rect 37452 1600 37516 1604
rect 38812 1660 38876 1664
rect 38812 1604 38816 1660
rect 38816 1604 38872 1660
rect 38872 1604 38876 1660
rect 38812 1600 38876 1604
rect 38892 1660 38956 1664
rect 38892 1604 38896 1660
rect 38896 1604 38952 1660
rect 38952 1604 38956 1660
rect 38892 1600 38956 1604
rect 38972 1660 39036 1664
rect 38972 1604 38976 1660
rect 38976 1604 39032 1660
rect 39032 1604 39036 1660
rect 38972 1600 39036 1604
rect 39052 1660 39116 1664
rect 39052 1604 39056 1660
rect 39056 1604 39112 1660
rect 39112 1604 39116 1660
rect 39052 1600 39116 1604
rect 40412 1660 40476 1664
rect 40412 1604 40416 1660
rect 40416 1604 40472 1660
rect 40472 1604 40476 1660
rect 40412 1600 40476 1604
rect 40492 1660 40556 1664
rect 40492 1604 40496 1660
rect 40496 1604 40552 1660
rect 40552 1604 40556 1660
rect 40492 1600 40556 1604
rect 40572 1660 40636 1664
rect 40572 1604 40576 1660
rect 40576 1604 40632 1660
rect 40632 1604 40636 1660
rect 40572 1600 40636 1604
rect 40652 1660 40716 1664
rect 40652 1604 40656 1660
rect 40656 1604 40712 1660
rect 40712 1604 40716 1660
rect 40652 1600 40716 1604
rect 42012 1660 42076 1664
rect 42012 1604 42016 1660
rect 42016 1604 42072 1660
rect 42072 1604 42076 1660
rect 42012 1600 42076 1604
rect 42092 1660 42156 1664
rect 42092 1604 42096 1660
rect 42096 1604 42152 1660
rect 42152 1604 42156 1660
rect 42092 1600 42156 1604
rect 42172 1660 42236 1664
rect 42172 1604 42176 1660
rect 42176 1604 42232 1660
rect 42232 1604 42236 1660
rect 42172 1600 42236 1604
rect 42252 1660 42316 1664
rect 42252 1604 42256 1660
rect 42256 1604 42312 1660
rect 42312 1604 42316 1660
rect 42252 1600 42316 1604
rect 43612 1660 43676 1664
rect 43612 1604 43616 1660
rect 43616 1604 43672 1660
rect 43672 1604 43676 1660
rect 43612 1600 43676 1604
rect 43692 1660 43756 1664
rect 43692 1604 43696 1660
rect 43696 1604 43752 1660
rect 43752 1604 43756 1660
rect 43692 1600 43756 1604
rect 43772 1660 43836 1664
rect 43772 1604 43776 1660
rect 43776 1604 43832 1660
rect 43832 1604 43836 1660
rect 43772 1600 43836 1604
rect 43852 1660 43916 1664
rect 43852 1604 43856 1660
rect 43856 1604 43912 1660
rect 43912 1604 43916 1660
rect 43852 1600 43916 1604
rect 45212 1660 45276 1664
rect 45212 1604 45216 1660
rect 45216 1604 45272 1660
rect 45272 1604 45276 1660
rect 45212 1600 45276 1604
rect 45292 1660 45356 1664
rect 45292 1604 45296 1660
rect 45296 1604 45352 1660
rect 45352 1604 45356 1660
rect 45292 1600 45356 1604
rect 45372 1660 45436 1664
rect 45372 1604 45376 1660
rect 45376 1604 45432 1660
rect 45432 1604 45436 1660
rect 45372 1600 45436 1604
rect 45452 1660 45516 1664
rect 45452 1604 45456 1660
rect 45456 1604 45512 1660
rect 45512 1604 45516 1660
rect 45452 1600 45516 1604
rect 46812 1660 46876 1664
rect 46812 1604 46816 1660
rect 46816 1604 46872 1660
rect 46872 1604 46876 1660
rect 46812 1600 46876 1604
rect 46892 1660 46956 1664
rect 46892 1604 46896 1660
rect 46896 1604 46952 1660
rect 46952 1604 46956 1660
rect 46892 1600 46956 1604
rect 46972 1660 47036 1664
rect 46972 1604 46976 1660
rect 46976 1604 47032 1660
rect 47032 1604 47036 1660
rect 46972 1600 47036 1604
rect 47052 1660 47116 1664
rect 47052 1604 47056 1660
rect 47056 1604 47112 1660
rect 47112 1604 47116 1660
rect 47052 1600 47116 1604
rect 48412 1660 48476 1664
rect 48412 1604 48416 1660
rect 48416 1604 48472 1660
rect 48472 1604 48476 1660
rect 48412 1600 48476 1604
rect 48492 1660 48556 1664
rect 48492 1604 48496 1660
rect 48496 1604 48552 1660
rect 48552 1604 48556 1660
rect 48492 1600 48556 1604
rect 48572 1660 48636 1664
rect 48572 1604 48576 1660
rect 48576 1604 48632 1660
rect 48632 1604 48636 1660
rect 48572 1600 48636 1604
rect 48652 1660 48716 1664
rect 48652 1604 48656 1660
rect 48656 1604 48712 1660
rect 48712 1604 48716 1660
rect 48652 1600 48716 1604
rect 50012 1660 50076 1664
rect 50012 1604 50016 1660
rect 50016 1604 50072 1660
rect 50072 1604 50076 1660
rect 50012 1600 50076 1604
rect 50092 1660 50156 1664
rect 50092 1604 50096 1660
rect 50096 1604 50152 1660
rect 50152 1604 50156 1660
rect 50092 1600 50156 1604
rect 50172 1660 50236 1664
rect 50172 1604 50176 1660
rect 50176 1604 50232 1660
rect 50232 1604 50236 1660
rect 50172 1600 50236 1604
rect 50252 1660 50316 1664
rect 50252 1604 50256 1660
rect 50256 1604 50312 1660
rect 50312 1604 50316 1660
rect 50252 1600 50316 1604
rect 51612 1660 51676 1664
rect 51612 1604 51616 1660
rect 51616 1604 51672 1660
rect 51672 1604 51676 1660
rect 51612 1600 51676 1604
rect 51692 1660 51756 1664
rect 51692 1604 51696 1660
rect 51696 1604 51752 1660
rect 51752 1604 51756 1660
rect 51692 1600 51756 1604
rect 51772 1660 51836 1664
rect 51772 1604 51776 1660
rect 51776 1604 51832 1660
rect 51832 1604 51836 1660
rect 51772 1600 51836 1604
rect 51852 1660 51916 1664
rect 51852 1604 51856 1660
rect 51856 1604 51912 1660
rect 51912 1604 51916 1660
rect 51852 1600 51916 1604
rect 53212 1660 53276 1664
rect 53212 1604 53216 1660
rect 53216 1604 53272 1660
rect 53272 1604 53276 1660
rect 53212 1600 53276 1604
rect 53292 1660 53356 1664
rect 53292 1604 53296 1660
rect 53296 1604 53352 1660
rect 53352 1604 53356 1660
rect 53292 1600 53356 1604
rect 53372 1660 53436 1664
rect 53372 1604 53376 1660
rect 53376 1604 53432 1660
rect 53432 1604 53436 1660
rect 53372 1600 53436 1604
rect 53452 1660 53516 1664
rect 53452 1604 53456 1660
rect 53456 1604 53512 1660
rect 53512 1604 53516 1660
rect 53452 1600 53516 1604
rect 54812 1660 54876 1664
rect 54812 1604 54816 1660
rect 54816 1604 54872 1660
rect 54872 1604 54876 1660
rect 54812 1600 54876 1604
rect 54892 1660 54956 1664
rect 54892 1604 54896 1660
rect 54896 1604 54952 1660
rect 54952 1604 54956 1660
rect 54892 1600 54956 1604
rect 54972 1660 55036 1664
rect 54972 1604 54976 1660
rect 54976 1604 55032 1660
rect 55032 1604 55036 1660
rect 54972 1600 55036 1604
rect 55052 1660 55116 1664
rect 55052 1604 55056 1660
rect 55056 1604 55112 1660
rect 55112 1604 55116 1660
rect 55052 1600 55116 1604
rect 56412 1660 56476 1664
rect 56412 1604 56416 1660
rect 56416 1604 56472 1660
rect 56472 1604 56476 1660
rect 56412 1600 56476 1604
rect 56492 1660 56556 1664
rect 56492 1604 56496 1660
rect 56496 1604 56552 1660
rect 56552 1604 56556 1660
rect 56492 1600 56556 1604
rect 56572 1660 56636 1664
rect 56572 1604 56576 1660
rect 56576 1604 56632 1660
rect 56632 1604 56636 1660
rect 56572 1600 56636 1604
rect 56652 1660 56716 1664
rect 56652 1604 56656 1660
rect 56656 1604 56712 1660
rect 56712 1604 56716 1660
rect 56652 1600 56716 1604
rect 58012 1660 58076 1664
rect 58012 1604 58016 1660
rect 58016 1604 58072 1660
rect 58072 1604 58076 1660
rect 58012 1600 58076 1604
rect 58092 1660 58156 1664
rect 58092 1604 58096 1660
rect 58096 1604 58152 1660
rect 58152 1604 58156 1660
rect 58092 1600 58156 1604
rect 58172 1660 58236 1664
rect 58172 1604 58176 1660
rect 58176 1604 58232 1660
rect 58232 1604 58236 1660
rect 58172 1600 58236 1604
rect 58252 1660 58316 1664
rect 58252 1604 58256 1660
rect 58256 1604 58312 1660
rect 58312 1604 58316 1660
rect 58252 1600 58316 1604
rect 59612 1660 59676 1664
rect 59612 1604 59616 1660
rect 59616 1604 59672 1660
rect 59672 1604 59676 1660
rect 59612 1600 59676 1604
rect 59692 1660 59756 1664
rect 59692 1604 59696 1660
rect 59696 1604 59752 1660
rect 59752 1604 59756 1660
rect 59692 1600 59756 1604
rect 59772 1660 59836 1664
rect 59772 1604 59776 1660
rect 59776 1604 59832 1660
rect 59832 1604 59836 1660
rect 59772 1600 59836 1604
rect 59852 1660 59916 1664
rect 59852 1604 59856 1660
rect 59856 1604 59912 1660
rect 59912 1604 59916 1660
rect 59852 1600 59916 1604
rect 61212 1660 61276 1664
rect 61212 1604 61216 1660
rect 61216 1604 61272 1660
rect 61272 1604 61276 1660
rect 61212 1600 61276 1604
rect 61292 1660 61356 1664
rect 61292 1604 61296 1660
rect 61296 1604 61352 1660
rect 61352 1604 61356 1660
rect 61292 1600 61356 1604
rect 61372 1660 61436 1664
rect 61372 1604 61376 1660
rect 61376 1604 61432 1660
rect 61432 1604 61436 1660
rect 61372 1600 61436 1604
rect 61452 1660 61516 1664
rect 61452 1604 61456 1660
rect 61456 1604 61512 1660
rect 61512 1604 61516 1660
rect 61452 1600 61516 1604
rect 62812 1660 62876 1664
rect 62812 1604 62816 1660
rect 62816 1604 62872 1660
rect 62872 1604 62876 1660
rect 62812 1600 62876 1604
rect 62892 1660 62956 1664
rect 62892 1604 62896 1660
rect 62896 1604 62952 1660
rect 62952 1604 62956 1660
rect 62892 1600 62956 1604
rect 62972 1660 63036 1664
rect 62972 1604 62976 1660
rect 62976 1604 63032 1660
rect 63032 1604 63036 1660
rect 62972 1600 63036 1604
rect 63052 1660 63116 1664
rect 63052 1604 63056 1660
rect 63056 1604 63112 1660
rect 63112 1604 63116 1660
rect 63052 1600 63116 1604
rect 64412 1660 64476 1664
rect 64412 1604 64416 1660
rect 64416 1604 64472 1660
rect 64472 1604 64476 1660
rect 64412 1600 64476 1604
rect 64492 1660 64556 1664
rect 64492 1604 64496 1660
rect 64496 1604 64552 1660
rect 64552 1604 64556 1660
rect 64492 1600 64556 1604
rect 64572 1660 64636 1664
rect 64572 1604 64576 1660
rect 64576 1604 64632 1660
rect 64632 1604 64636 1660
rect 64572 1600 64636 1604
rect 64652 1660 64716 1664
rect 64652 1604 64656 1660
rect 64656 1604 64712 1660
rect 64712 1604 64716 1660
rect 64652 1600 64716 1604
rect 66012 1660 66076 1664
rect 66012 1604 66016 1660
rect 66016 1604 66072 1660
rect 66072 1604 66076 1660
rect 66012 1600 66076 1604
rect 66092 1660 66156 1664
rect 66092 1604 66096 1660
rect 66096 1604 66152 1660
rect 66152 1604 66156 1660
rect 66092 1600 66156 1604
rect 66172 1660 66236 1664
rect 66172 1604 66176 1660
rect 66176 1604 66232 1660
rect 66232 1604 66236 1660
rect 66172 1600 66236 1604
rect 66252 1660 66316 1664
rect 66252 1604 66256 1660
rect 66256 1604 66312 1660
rect 66312 1604 66316 1660
rect 66252 1600 66316 1604
rect 67612 1660 67676 1664
rect 67612 1604 67616 1660
rect 67616 1604 67672 1660
rect 67672 1604 67676 1660
rect 67612 1600 67676 1604
rect 67692 1660 67756 1664
rect 67692 1604 67696 1660
rect 67696 1604 67752 1660
rect 67752 1604 67756 1660
rect 67692 1600 67756 1604
rect 67772 1660 67836 1664
rect 67772 1604 67776 1660
rect 67776 1604 67832 1660
rect 67832 1604 67836 1660
rect 67772 1600 67836 1604
rect 67852 1660 67916 1664
rect 67852 1604 67856 1660
rect 67856 1604 67912 1660
rect 67912 1604 67916 1660
rect 67852 1600 67916 1604
rect 69212 1660 69276 1664
rect 69212 1604 69216 1660
rect 69216 1604 69272 1660
rect 69272 1604 69276 1660
rect 69212 1600 69276 1604
rect 69292 1660 69356 1664
rect 69292 1604 69296 1660
rect 69296 1604 69352 1660
rect 69352 1604 69356 1660
rect 69292 1600 69356 1604
rect 69372 1660 69436 1664
rect 69372 1604 69376 1660
rect 69376 1604 69432 1660
rect 69432 1604 69436 1660
rect 69372 1600 69436 1604
rect 69452 1660 69516 1664
rect 69452 1604 69456 1660
rect 69456 1604 69512 1660
rect 69512 1604 69516 1660
rect 69452 1600 69516 1604
rect 70812 1660 70876 1664
rect 70812 1604 70816 1660
rect 70816 1604 70872 1660
rect 70872 1604 70876 1660
rect 70812 1600 70876 1604
rect 70892 1660 70956 1664
rect 70892 1604 70896 1660
rect 70896 1604 70952 1660
rect 70952 1604 70956 1660
rect 70892 1600 70956 1604
rect 70972 1660 71036 1664
rect 70972 1604 70976 1660
rect 70976 1604 71032 1660
rect 71032 1604 71036 1660
rect 70972 1600 71036 1604
rect 71052 1660 71116 1664
rect 71052 1604 71056 1660
rect 71056 1604 71112 1660
rect 71112 1604 71116 1660
rect 71052 1600 71116 1604
rect 72412 1660 72476 1664
rect 72412 1604 72416 1660
rect 72416 1604 72472 1660
rect 72472 1604 72476 1660
rect 72412 1600 72476 1604
rect 72492 1660 72556 1664
rect 72492 1604 72496 1660
rect 72496 1604 72552 1660
rect 72552 1604 72556 1660
rect 72492 1600 72556 1604
rect 72572 1660 72636 1664
rect 72572 1604 72576 1660
rect 72576 1604 72632 1660
rect 72632 1604 72636 1660
rect 72572 1600 72636 1604
rect 72652 1660 72716 1664
rect 72652 1604 72656 1660
rect 72656 1604 72712 1660
rect 72712 1604 72716 1660
rect 72652 1600 72716 1604
rect 74012 1660 74076 1664
rect 74012 1604 74016 1660
rect 74016 1604 74072 1660
rect 74072 1604 74076 1660
rect 74012 1600 74076 1604
rect 74092 1660 74156 1664
rect 74092 1604 74096 1660
rect 74096 1604 74152 1660
rect 74152 1604 74156 1660
rect 74092 1600 74156 1604
rect 74172 1660 74236 1664
rect 74172 1604 74176 1660
rect 74176 1604 74232 1660
rect 74232 1604 74236 1660
rect 74172 1600 74236 1604
rect 74252 1660 74316 1664
rect 74252 1604 74256 1660
rect 74256 1604 74312 1660
rect 74312 1604 74316 1660
rect 74252 1600 74316 1604
rect 75612 1660 75676 1664
rect 75612 1604 75616 1660
rect 75616 1604 75672 1660
rect 75672 1604 75676 1660
rect 75612 1600 75676 1604
rect 75692 1660 75756 1664
rect 75692 1604 75696 1660
rect 75696 1604 75752 1660
rect 75752 1604 75756 1660
rect 75692 1600 75756 1604
rect 75772 1660 75836 1664
rect 75772 1604 75776 1660
rect 75776 1604 75832 1660
rect 75832 1604 75836 1660
rect 75772 1600 75836 1604
rect 75852 1660 75916 1664
rect 75852 1604 75856 1660
rect 75856 1604 75912 1660
rect 75912 1604 75916 1660
rect 75852 1600 75916 1604
rect 77212 1660 77276 1664
rect 77212 1604 77216 1660
rect 77216 1604 77272 1660
rect 77272 1604 77276 1660
rect 77212 1600 77276 1604
rect 77292 1660 77356 1664
rect 77292 1604 77296 1660
rect 77296 1604 77352 1660
rect 77352 1604 77356 1660
rect 77292 1600 77356 1604
rect 77372 1660 77436 1664
rect 77372 1604 77376 1660
rect 77376 1604 77432 1660
rect 77432 1604 77436 1660
rect 77372 1600 77436 1604
rect 77452 1660 77516 1664
rect 77452 1604 77456 1660
rect 77456 1604 77512 1660
rect 77512 1604 77516 1660
rect 77452 1600 77516 1604
rect 78812 1660 78876 1664
rect 78812 1604 78816 1660
rect 78816 1604 78872 1660
rect 78872 1604 78876 1660
rect 78812 1600 78876 1604
rect 78892 1660 78956 1664
rect 78892 1604 78896 1660
rect 78896 1604 78952 1660
rect 78952 1604 78956 1660
rect 78892 1600 78956 1604
rect 78972 1660 79036 1664
rect 78972 1604 78976 1660
rect 78976 1604 79032 1660
rect 79032 1604 79036 1660
rect 78972 1600 79036 1604
rect 79052 1660 79116 1664
rect 79052 1604 79056 1660
rect 79056 1604 79112 1660
rect 79112 1604 79116 1660
rect 79052 1600 79116 1604
rect 80412 1660 80476 1664
rect 80412 1604 80416 1660
rect 80416 1604 80472 1660
rect 80472 1604 80476 1660
rect 80412 1600 80476 1604
rect 80492 1660 80556 1664
rect 80492 1604 80496 1660
rect 80496 1604 80552 1660
rect 80552 1604 80556 1660
rect 80492 1600 80556 1604
rect 80572 1660 80636 1664
rect 80572 1604 80576 1660
rect 80576 1604 80632 1660
rect 80632 1604 80636 1660
rect 80572 1600 80636 1604
rect 80652 1660 80716 1664
rect 80652 1604 80656 1660
rect 80656 1604 80712 1660
rect 80712 1604 80716 1660
rect 80652 1600 80716 1604
rect 82012 1660 82076 1664
rect 82012 1604 82016 1660
rect 82016 1604 82072 1660
rect 82072 1604 82076 1660
rect 82012 1600 82076 1604
rect 82092 1660 82156 1664
rect 82092 1604 82096 1660
rect 82096 1604 82152 1660
rect 82152 1604 82156 1660
rect 82092 1600 82156 1604
rect 82172 1660 82236 1664
rect 82172 1604 82176 1660
rect 82176 1604 82232 1660
rect 82232 1604 82236 1660
rect 82172 1600 82236 1604
rect 82252 1660 82316 1664
rect 82252 1604 82256 1660
rect 82256 1604 82312 1660
rect 82312 1604 82316 1660
rect 82252 1600 82316 1604
rect 83612 1660 83676 1664
rect 83612 1604 83616 1660
rect 83616 1604 83672 1660
rect 83672 1604 83676 1660
rect 83612 1600 83676 1604
rect 83692 1660 83756 1664
rect 83692 1604 83696 1660
rect 83696 1604 83752 1660
rect 83752 1604 83756 1660
rect 83692 1600 83756 1604
rect 83772 1660 83836 1664
rect 83772 1604 83776 1660
rect 83776 1604 83832 1660
rect 83832 1604 83836 1660
rect 83772 1600 83836 1604
rect 83852 1660 83916 1664
rect 83852 1604 83856 1660
rect 83856 1604 83912 1660
rect 83912 1604 83916 1660
rect 83852 1600 83916 1604
rect 85212 1660 85276 1664
rect 85212 1604 85216 1660
rect 85216 1604 85272 1660
rect 85272 1604 85276 1660
rect 85212 1600 85276 1604
rect 85292 1660 85356 1664
rect 85292 1604 85296 1660
rect 85296 1604 85352 1660
rect 85352 1604 85356 1660
rect 85292 1600 85356 1604
rect 85372 1660 85436 1664
rect 85372 1604 85376 1660
rect 85376 1604 85432 1660
rect 85432 1604 85436 1660
rect 85372 1600 85436 1604
rect 85452 1660 85516 1664
rect 85452 1604 85456 1660
rect 85456 1604 85512 1660
rect 85512 1604 85516 1660
rect 85452 1600 85516 1604
rect 86812 1660 86876 1664
rect 86812 1604 86816 1660
rect 86816 1604 86872 1660
rect 86872 1604 86876 1660
rect 86812 1600 86876 1604
rect 86892 1660 86956 1664
rect 86892 1604 86896 1660
rect 86896 1604 86952 1660
rect 86952 1604 86956 1660
rect 86892 1600 86956 1604
rect 86972 1660 87036 1664
rect 86972 1604 86976 1660
rect 86976 1604 87032 1660
rect 87032 1604 87036 1660
rect 86972 1600 87036 1604
rect 87052 1660 87116 1664
rect 87052 1604 87056 1660
rect 87056 1604 87112 1660
rect 87112 1604 87116 1660
rect 87052 1600 87116 1604
rect 88412 1660 88476 1664
rect 88412 1604 88416 1660
rect 88416 1604 88472 1660
rect 88472 1604 88476 1660
rect 88412 1600 88476 1604
rect 88492 1660 88556 1664
rect 88492 1604 88496 1660
rect 88496 1604 88552 1660
rect 88552 1604 88556 1660
rect 88492 1600 88556 1604
rect 88572 1660 88636 1664
rect 88572 1604 88576 1660
rect 88576 1604 88632 1660
rect 88632 1604 88636 1660
rect 88572 1600 88636 1604
rect 88652 1660 88716 1664
rect 88652 1604 88656 1660
rect 88656 1604 88712 1660
rect 88712 1604 88716 1660
rect 88652 1600 88716 1604
rect 90012 1660 90076 1664
rect 90012 1604 90016 1660
rect 90016 1604 90072 1660
rect 90072 1604 90076 1660
rect 90012 1600 90076 1604
rect 90092 1660 90156 1664
rect 90092 1604 90096 1660
rect 90096 1604 90152 1660
rect 90152 1604 90156 1660
rect 90092 1600 90156 1604
rect 90172 1660 90236 1664
rect 90172 1604 90176 1660
rect 90176 1604 90232 1660
rect 90232 1604 90236 1660
rect 90172 1600 90236 1604
rect 90252 1660 90316 1664
rect 90252 1604 90256 1660
rect 90256 1604 90312 1660
rect 90312 1604 90316 1660
rect 90252 1600 90316 1604
rect 91612 1660 91676 1664
rect 91612 1604 91616 1660
rect 91616 1604 91672 1660
rect 91672 1604 91676 1660
rect 91612 1600 91676 1604
rect 91692 1660 91756 1664
rect 91692 1604 91696 1660
rect 91696 1604 91752 1660
rect 91752 1604 91756 1660
rect 91692 1600 91756 1604
rect 91772 1660 91836 1664
rect 91772 1604 91776 1660
rect 91776 1604 91832 1660
rect 91832 1604 91836 1660
rect 91772 1600 91836 1604
rect 91852 1660 91916 1664
rect 91852 1604 91856 1660
rect 91856 1604 91912 1660
rect 91912 1604 91916 1660
rect 91852 1600 91916 1604
rect 93212 1660 93276 1664
rect 93212 1604 93216 1660
rect 93216 1604 93272 1660
rect 93272 1604 93276 1660
rect 93212 1600 93276 1604
rect 93292 1660 93356 1664
rect 93292 1604 93296 1660
rect 93296 1604 93352 1660
rect 93352 1604 93356 1660
rect 93292 1600 93356 1604
rect 93372 1660 93436 1664
rect 93372 1604 93376 1660
rect 93376 1604 93432 1660
rect 93432 1604 93436 1660
rect 93372 1600 93436 1604
rect 93452 1660 93516 1664
rect 93452 1604 93456 1660
rect 93456 1604 93512 1660
rect 93512 1604 93516 1660
rect 93452 1600 93516 1604
rect 94812 1660 94876 1664
rect 94812 1604 94816 1660
rect 94816 1604 94872 1660
rect 94872 1604 94876 1660
rect 94812 1600 94876 1604
rect 94892 1660 94956 1664
rect 94892 1604 94896 1660
rect 94896 1604 94952 1660
rect 94952 1604 94956 1660
rect 94892 1600 94956 1604
rect 94972 1660 95036 1664
rect 94972 1604 94976 1660
rect 94976 1604 95032 1660
rect 95032 1604 95036 1660
rect 94972 1600 95036 1604
rect 95052 1660 95116 1664
rect 95052 1604 95056 1660
rect 95056 1604 95112 1660
rect 95112 1604 95116 1660
rect 95052 1600 95116 1604
rect 96412 1660 96476 1664
rect 96412 1604 96416 1660
rect 96416 1604 96472 1660
rect 96472 1604 96476 1660
rect 96412 1600 96476 1604
rect 96492 1660 96556 1664
rect 96492 1604 96496 1660
rect 96496 1604 96552 1660
rect 96552 1604 96556 1660
rect 96492 1600 96556 1604
rect 96572 1660 96636 1664
rect 96572 1604 96576 1660
rect 96576 1604 96632 1660
rect 96632 1604 96636 1660
rect 96572 1600 96636 1604
rect 96652 1660 96716 1664
rect 96652 1604 96656 1660
rect 96656 1604 96712 1660
rect 96712 1604 96716 1660
rect 96652 1600 96716 1604
rect 98012 1660 98076 1664
rect 98012 1604 98016 1660
rect 98016 1604 98072 1660
rect 98072 1604 98076 1660
rect 98012 1600 98076 1604
rect 98092 1660 98156 1664
rect 98092 1604 98096 1660
rect 98096 1604 98152 1660
rect 98152 1604 98156 1660
rect 98092 1600 98156 1604
rect 98172 1660 98236 1664
rect 98172 1604 98176 1660
rect 98176 1604 98232 1660
rect 98232 1604 98236 1660
rect 98172 1600 98236 1604
rect 98252 1660 98316 1664
rect 98252 1604 98256 1660
rect 98256 1604 98312 1660
rect 98312 1604 98316 1660
rect 98252 1600 98316 1604
rect 99612 1660 99676 1664
rect 99612 1604 99616 1660
rect 99616 1604 99672 1660
rect 99672 1604 99676 1660
rect 99612 1600 99676 1604
rect 99692 1660 99756 1664
rect 99692 1604 99696 1660
rect 99696 1604 99752 1660
rect 99752 1604 99756 1660
rect 99692 1600 99756 1604
rect 99772 1660 99836 1664
rect 99772 1604 99776 1660
rect 99776 1604 99832 1660
rect 99832 1604 99836 1660
rect 99772 1600 99836 1604
rect 99852 1660 99916 1664
rect 99852 1604 99856 1660
rect 99856 1604 99912 1660
rect 99912 1604 99916 1660
rect 99852 1600 99916 1604
rect 101212 1660 101276 1664
rect 101212 1604 101216 1660
rect 101216 1604 101272 1660
rect 101272 1604 101276 1660
rect 101212 1600 101276 1604
rect 101292 1660 101356 1664
rect 101292 1604 101296 1660
rect 101296 1604 101352 1660
rect 101352 1604 101356 1660
rect 101292 1600 101356 1604
rect 101372 1660 101436 1664
rect 101372 1604 101376 1660
rect 101376 1604 101432 1660
rect 101432 1604 101436 1660
rect 101372 1600 101436 1604
rect 101452 1660 101516 1664
rect 101452 1604 101456 1660
rect 101456 1604 101512 1660
rect 101512 1604 101516 1660
rect 101452 1600 101516 1604
rect 102812 1660 102876 1664
rect 102812 1604 102816 1660
rect 102816 1604 102872 1660
rect 102872 1604 102876 1660
rect 102812 1600 102876 1604
rect 102892 1660 102956 1664
rect 102892 1604 102896 1660
rect 102896 1604 102952 1660
rect 102952 1604 102956 1660
rect 102892 1600 102956 1604
rect 102972 1660 103036 1664
rect 102972 1604 102976 1660
rect 102976 1604 103032 1660
rect 103032 1604 103036 1660
rect 102972 1600 103036 1604
rect 103052 1660 103116 1664
rect 103052 1604 103056 1660
rect 103056 1604 103112 1660
rect 103112 1604 103116 1660
rect 103052 1600 103116 1604
rect 104412 1660 104476 1664
rect 104412 1604 104416 1660
rect 104416 1604 104472 1660
rect 104472 1604 104476 1660
rect 104412 1600 104476 1604
rect 104492 1660 104556 1664
rect 104492 1604 104496 1660
rect 104496 1604 104552 1660
rect 104552 1604 104556 1660
rect 104492 1600 104556 1604
rect 104572 1660 104636 1664
rect 104572 1604 104576 1660
rect 104576 1604 104632 1660
rect 104632 1604 104636 1660
rect 104572 1600 104636 1604
rect 104652 1660 104716 1664
rect 104652 1604 104656 1660
rect 104656 1604 104712 1660
rect 104712 1604 104716 1660
rect 104652 1600 104716 1604
rect 106012 1660 106076 1664
rect 106012 1604 106016 1660
rect 106016 1604 106072 1660
rect 106072 1604 106076 1660
rect 106012 1600 106076 1604
rect 106092 1660 106156 1664
rect 106092 1604 106096 1660
rect 106096 1604 106152 1660
rect 106152 1604 106156 1660
rect 106092 1600 106156 1604
rect 106172 1660 106236 1664
rect 106172 1604 106176 1660
rect 106176 1604 106232 1660
rect 106232 1604 106236 1660
rect 106172 1600 106236 1604
rect 106252 1660 106316 1664
rect 106252 1604 106256 1660
rect 106256 1604 106312 1660
rect 106312 1604 106316 1660
rect 106252 1600 106316 1604
rect 107612 1660 107676 1664
rect 107612 1604 107616 1660
rect 107616 1604 107672 1660
rect 107672 1604 107676 1660
rect 107612 1600 107676 1604
rect 107692 1660 107756 1664
rect 107692 1604 107696 1660
rect 107696 1604 107752 1660
rect 107752 1604 107756 1660
rect 107692 1600 107756 1604
rect 107772 1660 107836 1664
rect 107772 1604 107776 1660
rect 107776 1604 107832 1660
rect 107832 1604 107836 1660
rect 107772 1600 107836 1604
rect 107852 1660 107916 1664
rect 107852 1604 107856 1660
rect 107856 1604 107912 1660
rect 107912 1604 107916 1660
rect 107852 1600 107916 1604
rect 31340 1260 31404 1324
rect 33180 1320 33244 1324
rect 33180 1264 33230 1320
rect 33230 1264 33244 1320
rect 33180 1260 33244 1264
rect 34468 1320 34532 1324
rect 34468 1264 34518 1320
rect 34518 1264 34532 1320
rect 34468 1260 34532 1264
rect 37964 1260 38028 1324
rect 56916 1260 56980 1324
rect 58756 1260 58820 1324
rect 60228 1260 60292 1324
rect 60964 1320 61028 1324
rect 60964 1264 60978 1320
rect 60978 1264 61028 1320
rect 60964 1260 61028 1264
rect 62620 1260 62684 1324
rect 63540 1320 63604 1324
rect 63540 1264 63554 1320
rect 63554 1264 63604 1320
rect 63540 1260 63604 1264
rect 65012 1260 65076 1324
rect 65748 1260 65812 1324
rect 67404 1260 67468 1324
rect 68324 1260 68388 1324
rect 69612 1260 69676 1324
rect 2952 1116 3016 1120
rect 2952 1060 2956 1116
rect 2956 1060 3012 1116
rect 3012 1060 3016 1116
rect 2952 1056 3016 1060
rect 3032 1116 3096 1120
rect 3032 1060 3036 1116
rect 3036 1060 3092 1116
rect 3092 1060 3096 1116
rect 3032 1056 3096 1060
rect 3112 1116 3176 1120
rect 3112 1060 3116 1116
rect 3116 1060 3172 1116
rect 3172 1060 3176 1116
rect 3112 1056 3176 1060
rect 3192 1116 3256 1120
rect 3192 1060 3196 1116
rect 3196 1060 3252 1116
rect 3252 1060 3256 1116
rect 3192 1056 3256 1060
rect 4552 1116 4616 1120
rect 4552 1060 4556 1116
rect 4556 1060 4612 1116
rect 4612 1060 4616 1116
rect 4552 1056 4616 1060
rect 4632 1116 4696 1120
rect 4632 1060 4636 1116
rect 4636 1060 4692 1116
rect 4692 1060 4696 1116
rect 4632 1056 4696 1060
rect 4712 1116 4776 1120
rect 4712 1060 4716 1116
rect 4716 1060 4772 1116
rect 4772 1060 4776 1116
rect 4712 1056 4776 1060
rect 4792 1116 4856 1120
rect 4792 1060 4796 1116
rect 4796 1060 4852 1116
rect 4852 1060 4856 1116
rect 4792 1056 4856 1060
rect 6152 1116 6216 1120
rect 6152 1060 6156 1116
rect 6156 1060 6212 1116
rect 6212 1060 6216 1116
rect 6152 1056 6216 1060
rect 6232 1116 6296 1120
rect 6232 1060 6236 1116
rect 6236 1060 6292 1116
rect 6292 1060 6296 1116
rect 6232 1056 6296 1060
rect 6312 1116 6376 1120
rect 6312 1060 6316 1116
rect 6316 1060 6372 1116
rect 6372 1060 6376 1116
rect 6312 1056 6376 1060
rect 6392 1116 6456 1120
rect 6392 1060 6396 1116
rect 6396 1060 6452 1116
rect 6452 1060 6456 1116
rect 6392 1056 6456 1060
rect 7752 1116 7816 1120
rect 7752 1060 7756 1116
rect 7756 1060 7812 1116
rect 7812 1060 7816 1116
rect 7752 1056 7816 1060
rect 7832 1116 7896 1120
rect 7832 1060 7836 1116
rect 7836 1060 7892 1116
rect 7892 1060 7896 1116
rect 7832 1056 7896 1060
rect 7912 1116 7976 1120
rect 7912 1060 7916 1116
rect 7916 1060 7972 1116
rect 7972 1060 7976 1116
rect 7912 1056 7976 1060
rect 7992 1116 8056 1120
rect 7992 1060 7996 1116
rect 7996 1060 8052 1116
rect 8052 1060 8056 1116
rect 7992 1056 8056 1060
rect 9352 1116 9416 1120
rect 9352 1060 9356 1116
rect 9356 1060 9412 1116
rect 9412 1060 9416 1116
rect 9352 1056 9416 1060
rect 9432 1116 9496 1120
rect 9432 1060 9436 1116
rect 9436 1060 9492 1116
rect 9492 1060 9496 1116
rect 9432 1056 9496 1060
rect 9512 1116 9576 1120
rect 9512 1060 9516 1116
rect 9516 1060 9572 1116
rect 9572 1060 9576 1116
rect 9512 1056 9576 1060
rect 9592 1116 9656 1120
rect 9592 1060 9596 1116
rect 9596 1060 9652 1116
rect 9652 1060 9656 1116
rect 9592 1056 9656 1060
rect 10952 1116 11016 1120
rect 10952 1060 10956 1116
rect 10956 1060 11012 1116
rect 11012 1060 11016 1116
rect 10952 1056 11016 1060
rect 11032 1116 11096 1120
rect 11032 1060 11036 1116
rect 11036 1060 11092 1116
rect 11092 1060 11096 1116
rect 11032 1056 11096 1060
rect 11112 1116 11176 1120
rect 11112 1060 11116 1116
rect 11116 1060 11172 1116
rect 11172 1060 11176 1116
rect 11112 1056 11176 1060
rect 11192 1116 11256 1120
rect 11192 1060 11196 1116
rect 11196 1060 11252 1116
rect 11252 1060 11256 1116
rect 11192 1056 11256 1060
rect 12552 1116 12616 1120
rect 12552 1060 12556 1116
rect 12556 1060 12612 1116
rect 12612 1060 12616 1116
rect 12552 1056 12616 1060
rect 12632 1116 12696 1120
rect 12632 1060 12636 1116
rect 12636 1060 12692 1116
rect 12692 1060 12696 1116
rect 12632 1056 12696 1060
rect 12712 1116 12776 1120
rect 12712 1060 12716 1116
rect 12716 1060 12772 1116
rect 12772 1060 12776 1116
rect 12712 1056 12776 1060
rect 12792 1116 12856 1120
rect 12792 1060 12796 1116
rect 12796 1060 12852 1116
rect 12852 1060 12856 1116
rect 12792 1056 12856 1060
rect 14152 1116 14216 1120
rect 14152 1060 14156 1116
rect 14156 1060 14212 1116
rect 14212 1060 14216 1116
rect 14152 1056 14216 1060
rect 14232 1116 14296 1120
rect 14232 1060 14236 1116
rect 14236 1060 14292 1116
rect 14292 1060 14296 1116
rect 14232 1056 14296 1060
rect 14312 1116 14376 1120
rect 14312 1060 14316 1116
rect 14316 1060 14372 1116
rect 14372 1060 14376 1116
rect 14312 1056 14376 1060
rect 14392 1116 14456 1120
rect 14392 1060 14396 1116
rect 14396 1060 14452 1116
rect 14452 1060 14456 1116
rect 14392 1056 14456 1060
rect 15752 1116 15816 1120
rect 15752 1060 15756 1116
rect 15756 1060 15812 1116
rect 15812 1060 15816 1116
rect 15752 1056 15816 1060
rect 15832 1116 15896 1120
rect 15832 1060 15836 1116
rect 15836 1060 15892 1116
rect 15892 1060 15896 1116
rect 15832 1056 15896 1060
rect 15912 1116 15976 1120
rect 15912 1060 15916 1116
rect 15916 1060 15972 1116
rect 15972 1060 15976 1116
rect 15912 1056 15976 1060
rect 15992 1116 16056 1120
rect 15992 1060 15996 1116
rect 15996 1060 16052 1116
rect 16052 1060 16056 1116
rect 15992 1056 16056 1060
rect 17352 1116 17416 1120
rect 17352 1060 17356 1116
rect 17356 1060 17412 1116
rect 17412 1060 17416 1116
rect 17352 1056 17416 1060
rect 17432 1116 17496 1120
rect 17432 1060 17436 1116
rect 17436 1060 17492 1116
rect 17492 1060 17496 1116
rect 17432 1056 17496 1060
rect 17512 1116 17576 1120
rect 17512 1060 17516 1116
rect 17516 1060 17572 1116
rect 17572 1060 17576 1116
rect 17512 1056 17576 1060
rect 17592 1116 17656 1120
rect 17592 1060 17596 1116
rect 17596 1060 17652 1116
rect 17652 1060 17656 1116
rect 17592 1056 17656 1060
rect 18952 1116 19016 1120
rect 18952 1060 18956 1116
rect 18956 1060 19012 1116
rect 19012 1060 19016 1116
rect 18952 1056 19016 1060
rect 19032 1116 19096 1120
rect 19032 1060 19036 1116
rect 19036 1060 19092 1116
rect 19092 1060 19096 1116
rect 19032 1056 19096 1060
rect 19112 1116 19176 1120
rect 19112 1060 19116 1116
rect 19116 1060 19172 1116
rect 19172 1060 19176 1116
rect 19112 1056 19176 1060
rect 19192 1116 19256 1120
rect 19192 1060 19196 1116
rect 19196 1060 19252 1116
rect 19252 1060 19256 1116
rect 19192 1056 19256 1060
rect 20552 1116 20616 1120
rect 20552 1060 20556 1116
rect 20556 1060 20612 1116
rect 20612 1060 20616 1116
rect 20552 1056 20616 1060
rect 20632 1116 20696 1120
rect 20632 1060 20636 1116
rect 20636 1060 20692 1116
rect 20692 1060 20696 1116
rect 20632 1056 20696 1060
rect 20712 1116 20776 1120
rect 20712 1060 20716 1116
rect 20716 1060 20772 1116
rect 20772 1060 20776 1116
rect 20712 1056 20776 1060
rect 20792 1116 20856 1120
rect 20792 1060 20796 1116
rect 20796 1060 20852 1116
rect 20852 1060 20856 1116
rect 20792 1056 20856 1060
rect 22152 1116 22216 1120
rect 22152 1060 22156 1116
rect 22156 1060 22212 1116
rect 22212 1060 22216 1116
rect 22152 1056 22216 1060
rect 22232 1116 22296 1120
rect 22232 1060 22236 1116
rect 22236 1060 22292 1116
rect 22292 1060 22296 1116
rect 22232 1056 22296 1060
rect 22312 1116 22376 1120
rect 22312 1060 22316 1116
rect 22316 1060 22372 1116
rect 22372 1060 22376 1116
rect 22312 1056 22376 1060
rect 22392 1116 22456 1120
rect 22392 1060 22396 1116
rect 22396 1060 22452 1116
rect 22452 1060 22456 1116
rect 22392 1056 22456 1060
rect 23752 1116 23816 1120
rect 23752 1060 23756 1116
rect 23756 1060 23812 1116
rect 23812 1060 23816 1116
rect 23752 1056 23816 1060
rect 23832 1116 23896 1120
rect 23832 1060 23836 1116
rect 23836 1060 23892 1116
rect 23892 1060 23896 1116
rect 23832 1056 23896 1060
rect 23912 1116 23976 1120
rect 23912 1060 23916 1116
rect 23916 1060 23972 1116
rect 23972 1060 23976 1116
rect 23912 1056 23976 1060
rect 23992 1116 24056 1120
rect 23992 1060 23996 1116
rect 23996 1060 24052 1116
rect 24052 1060 24056 1116
rect 23992 1056 24056 1060
rect 25352 1116 25416 1120
rect 25352 1060 25356 1116
rect 25356 1060 25412 1116
rect 25412 1060 25416 1116
rect 25352 1056 25416 1060
rect 25432 1116 25496 1120
rect 25432 1060 25436 1116
rect 25436 1060 25492 1116
rect 25492 1060 25496 1116
rect 25432 1056 25496 1060
rect 25512 1116 25576 1120
rect 25512 1060 25516 1116
rect 25516 1060 25572 1116
rect 25572 1060 25576 1116
rect 25512 1056 25576 1060
rect 25592 1116 25656 1120
rect 25592 1060 25596 1116
rect 25596 1060 25652 1116
rect 25652 1060 25656 1116
rect 25592 1056 25656 1060
rect 26952 1116 27016 1120
rect 26952 1060 26956 1116
rect 26956 1060 27012 1116
rect 27012 1060 27016 1116
rect 26952 1056 27016 1060
rect 27032 1116 27096 1120
rect 27032 1060 27036 1116
rect 27036 1060 27092 1116
rect 27092 1060 27096 1116
rect 27032 1056 27096 1060
rect 27112 1116 27176 1120
rect 27112 1060 27116 1116
rect 27116 1060 27172 1116
rect 27172 1060 27176 1116
rect 27112 1056 27176 1060
rect 27192 1116 27256 1120
rect 27192 1060 27196 1116
rect 27196 1060 27252 1116
rect 27252 1060 27256 1116
rect 27192 1056 27256 1060
rect 28552 1116 28616 1120
rect 28552 1060 28556 1116
rect 28556 1060 28612 1116
rect 28612 1060 28616 1116
rect 28552 1056 28616 1060
rect 28632 1116 28696 1120
rect 28632 1060 28636 1116
rect 28636 1060 28692 1116
rect 28692 1060 28696 1116
rect 28632 1056 28696 1060
rect 28712 1116 28776 1120
rect 28712 1060 28716 1116
rect 28716 1060 28772 1116
rect 28772 1060 28776 1116
rect 28712 1056 28776 1060
rect 28792 1116 28856 1120
rect 28792 1060 28796 1116
rect 28796 1060 28852 1116
rect 28852 1060 28856 1116
rect 28792 1056 28856 1060
rect 30152 1116 30216 1120
rect 30152 1060 30156 1116
rect 30156 1060 30212 1116
rect 30212 1060 30216 1116
rect 30152 1056 30216 1060
rect 30232 1116 30296 1120
rect 30232 1060 30236 1116
rect 30236 1060 30292 1116
rect 30292 1060 30296 1116
rect 30232 1056 30296 1060
rect 30312 1116 30376 1120
rect 30312 1060 30316 1116
rect 30316 1060 30372 1116
rect 30372 1060 30376 1116
rect 30312 1056 30376 1060
rect 30392 1116 30456 1120
rect 30392 1060 30396 1116
rect 30396 1060 30452 1116
rect 30452 1060 30456 1116
rect 30392 1056 30456 1060
rect 31752 1116 31816 1120
rect 31752 1060 31756 1116
rect 31756 1060 31812 1116
rect 31812 1060 31816 1116
rect 31752 1056 31816 1060
rect 31832 1116 31896 1120
rect 31832 1060 31836 1116
rect 31836 1060 31892 1116
rect 31892 1060 31896 1116
rect 31832 1056 31896 1060
rect 31912 1116 31976 1120
rect 31912 1060 31916 1116
rect 31916 1060 31972 1116
rect 31972 1060 31976 1116
rect 31912 1056 31976 1060
rect 31992 1116 32056 1120
rect 31992 1060 31996 1116
rect 31996 1060 32052 1116
rect 32052 1060 32056 1116
rect 31992 1056 32056 1060
rect 33352 1116 33416 1120
rect 33352 1060 33356 1116
rect 33356 1060 33412 1116
rect 33412 1060 33416 1116
rect 33352 1056 33416 1060
rect 33432 1116 33496 1120
rect 33432 1060 33436 1116
rect 33436 1060 33492 1116
rect 33492 1060 33496 1116
rect 33432 1056 33496 1060
rect 33512 1116 33576 1120
rect 33512 1060 33516 1116
rect 33516 1060 33572 1116
rect 33572 1060 33576 1116
rect 33512 1056 33576 1060
rect 33592 1116 33656 1120
rect 33592 1060 33596 1116
rect 33596 1060 33652 1116
rect 33652 1060 33656 1116
rect 33592 1056 33656 1060
rect 34952 1116 35016 1120
rect 34952 1060 34956 1116
rect 34956 1060 35012 1116
rect 35012 1060 35016 1116
rect 34952 1056 35016 1060
rect 35032 1116 35096 1120
rect 35032 1060 35036 1116
rect 35036 1060 35092 1116
rect 35092 1060 35096 1116
rect 35032 1056 35096 1060
rect 35112 1116 35176 1120
rect 35112 1060 35116 1116
rect 35116 1060 35172 1116
rect 35172 1060 35176 1116
rect 35112 1056 35176 1060
rect 35192 1116 35256 1120
rect 35192 1060 35196 1116
rect 35196 1060 35252 1116
rect 35252 1060 35256 1116
rect 35192 1056 35256 1060
rect 36552 1116 36616 1120
rect 36552 1060 36556 1116
rect 36556 1060 36612 1116
rect 36612 1060 36616 1116
rect 36552 1056 36616 1060
rect 36632 1116 36696 1120
rect 36632 1060 36636 1116
rect 36636 1060 36692 1116
rect 36692 1060 36696 1116
rect 36632 1056 36696 1060
rect 36712 1116 36776 1120
rect 36712 1060 36716 1116
rect 36716 1060 36772 1116
rect 36772 1060 36776 1116
rect 36712 1056 36776 1060
rect 36792 1116 36856 1120
rect 36792 1060 36796 1116
rect 36796 1060 36852 1116
rect 36852 1060 36856 1116
rect 36792 1056 36856 1060
rect 38152 1116 38216 1120
rect 38152 1060 38156 1116
rect 38156 1060 38212 1116
rect 38212 1060 38216 1116
rect 38152 1056 38216 1060
rect 38232 1116 38296 1120
rect 38232 1060 38236 1116
rect 38236 1060 38292 1116
rect 38292 1060 38296 1116
rect 38232 1056 38296 1060
rect 38312 1116 38376 1120
rect 38312 1060 38316 1116
rect 38316 1060 38372 1116
rect 38372 1060 38376 1116
rect 38312 1056 38376 1060
rect 38392 1116 38456 1120
rect 38392 1060 38396 1116
rect 38396 1060 38452 1116
rect 38452 1060 38456 1116
rect 38392 1056 38456 1060
rect 39752 1116 39816 1120
rect 39752 1060 39756 1116
rect 39756 1060 39812 1116
rect 39812 1060 39816 1116
rect 39752 1056 39816 1060
rect 39832 1116 39896 1120
rect 39832 1060 39836 1116
rect 39836 1060 39892 1116
rect 39892 1060 39896 1116
rect 39832 1056 39896 1060
rect 39912 1116 39976 1120
rect 39912 1060 39916 1116
rect 39916 1060 39972 1116
rect 39972 1060 39976 1116
rect 39912 1056 39976 1060
rect 39992 1116 40056 1120
rect 39992 1060 39996 1116
rect 39996 1060 40052 1116
rect 40052 1060 40056 1116
rect 39992 1056 40056 1060
rect 41352 1116 41416 1120
rect 41352 1060 41356 1116
rect 41356 1060 41412 1116
rect 41412 1060 41416 1116
rect 41352 1056 41416 1060
rect 41432 1116 41496 1120
rect 41432 1060 41436 1116
rect 41436 1060 41492 1116
rect 41492 1060 41496 1116
rect 41432 1056 41496 1060
rect 41512 1116 41576 1120
rect 41512 1060 41516 1116
rect 41516 1060 41572 1116
rect 41572 1060 41576 1116
rect 41512 1056 41576 1060
rect 41592 1116 41656 1120
rect 41592 1060 41596 1116
rect 41596 1060 41652 1116
rect 41652 1060 41656 1116
rect 41592 1056 41656 1060
rect 42952 1116 43016 1120
rect 42952 1060 42956 1116
rect 42956 1060 43012 1116
rect 43012 1060 43016 1116
rect 42952 1056 43016 1060
rect 43032 1116 43096 1120
rect 43032 1060 43036 1116
rect 43036 1060 43092 1116
rect 43092 1060 43096 1116
rect 43032 1056 43096 1060
rect 43112 1116 43176 1120
rect 43112 1060 43116 1116
rect 43116 1060 43172 1116
rect 43172 1060 43176 1116
rect 43112 1056 43176 1060
rect 43192 1116 43256 1120
rect 43192 1060 43196 1116
rect 43196 1060 43252 1116
rect 43252 1060 43256 1116
rect 43192 1056 43256 1060
rect 44552 1116 44616 1120
rect 44552 1060 44556 1116
rect 44556 1060 44612 1116
rect 44612 1060 44616 1116
rect 44552 1056 44616 1060
rect 44632 1116 44696 1120
rect 44632 1060 44636 1116
rect 44636 1060 44692 1116
rect 44692 1060 44696 1116
rect 44632 1056 44696 1060
rect 44712 1116 44776 1120
rect 44712 1060 44716 1116
rect 44716 1060 44772 1116
rect 44772 1060 44776 1116
rect 44712 1056 44776 1060
rect 44792 1116 44856 1120
rect 44792 1060 44796 1116
rect 44796 1060 44852 1116
rect 44852 1060 44856 1116
rect 44792 1056 44856 1060
rect 46152 1116 46216 1120
rect 46152 1060 46156 1116
rect 46156 1060 46212 1116
rect 46212 1060 46216 1116
rect 46152 1056 46216 1060
rect 46232 1116 46296 1120
rect 46232 1060 46236 1116
rect 46236 1060 46292 1116
rect 46292 1060 46296 1116
rect 46232 1056 46296 1060
rect 46312 1116 46376 1120
rect 46312 1060 46316 1116
rect 46316 1060 46372 1116
rect 46372 1060 46376 1116
rect 46312 1056 46376 1060
rect 46392 1116 46456 1120
rect 46392 1060 46396 1116
rect 46396 1060 46452 1116
rect 46452 1060 46456 1116
rect 46392 1056 46456 1060
rect 47752 1116 47816 1120
rect 47752 1060 47756 1116
rect 47756 1060 47812 1116
rect 47812 1060 47816 1116
rect 47752 1056 47816 1060
rect 47832 1116 47896 1120
rect 47832 1060 47836 1116
rect 47836 1060 47892 1116
rect 47892 1060 47896 1116
rect 47832 1056 47896 1060
rect 47912 1116 47976 1120
rect 47912 1060 47916 1116
rect 47916 1060 47972 1116
rect 47972 1060 47976 1116
rect 47912 1056 47976 1060
rect 47992 1116 48056 1120
rect 47992 1060 47996 1116
rect 47996 1060 48052 1116
rect 48052 1060 48056 1116
rect 47992 1056 48056 1060
rect 49352 1116 49416 1120
rect 49352 1060 49356 1116
rect 49356 1060 49412 1116
rect 49412 1060 49416 1116
rect 49352 1056 49416 1060
rect 49432 1116 49496 1120
rect 49432 1060 49436 1116
rect 49436 1060 49492 1116
rect 49492 1060 49496 1116
rect 49432 1056 49496 1060
rect 49512 1116 49576 1120
rect 49512 1060 49516 1116
rect 49516 1060 49572 1116
rect 49572 1060 49576 1116
rect 49512 1056 49576 1060
rect 49592 1116 49656 1120
rect 49592 1060 49596 1116
rect 49596 1060 49652 1116
rect 49652 1060 49656 1116
rect 49592 1056 49656 1060
rect 50952 1116 51016 1120
rect 50952 1060 50956 1116
rect 50956 1060 51012 1116
rect 51012 1060 51016 1116
rect 50952 1056 51016 1060
rect 51032 1116 51096 1120
rect 51032 1060 51036 1116
rect 51036 1060 51092 1116
rect 51092 1060 51096 1116
rect 51032 1056 51096 1060
rect 51112 1116 51176 1120
rect 51112 1060 51116 1116
rect 51116 1060 51172 1116
rect 51172 1060 51176 1116
rect 51112 1056 51176 1060
rect 51192 1116 51256 1120
rect 51192 1060 51196 1116
rect 51196 1060 51252 1116
rect 51252 1060 51256 1116
rect 51192 1056 51256 1060
rect 52552 1116 52616 1120
rect 52552 1060 52556 1116
rect 52556 1060 52612 1116
rect 52612 1060 52616 1116
rect 52552 1056 52616 1060
rect 52632 1116 52696 1120
rect 52632 1060 52636 1116
rect 52636 1060 52692 1116
rect 52692 1060 52696 1116
rect 52632 1056 52696 1060
rect 52712 1116 52776 1120
rect 52712 1060 52716 1116
rect 52716 1060 52772 1116
rect 52772 1060 52776 1116
rect 52712 1056 52776 1060
rect 52792 1116 52856 1120
rect 52792 1060 52796 1116
rect 52796 1060 52852 1116
rect 52852 1060 52856 1116
rect 52792 1056 52856 1060
rect 54152 1116 54216 1120
rect 54152 1060 54156 1116
rect 54156 1060 54212 1116
rect 54212 1060 54216 1116
rect 54152 1056 54216 1060
rect 54232 1116 54296 1120
rect 54232 1060 54236 1116
rect 54236 1060 54292 1116
rect 54292 1060 54296 1116
rect 54232 1056 54296 1060
rect 54312 1116 54376 1120
rect 54312 1060 54316 1116
rect 54316 1060 54372 1116
rect 54372 1060 54376 1116
rect 54312 1056 54376 1060
rect 54392 1116 54456 1120
rect 54392 1060 54396 1116
rect 54396 1060 54452 1116
rect 54452 1060 54456 1116
rect 54392 1056 54456 1060
rect 55752 1116 55816 1120
rect 55752 1060 55756 1116
rect 55756 1060 55812 1116
rect 55812 1060 55816 1116
rect 55752 1056 55816 1060
rect 55832 1116 55896 1120
rect 55832 1060 55836 1116
rect 55836 1060 55892 1116
rect 55892 1060 55896 1116
rect 55832 1056 55896 1060
rect 55912 1116 55976 1120
rect 55912 1060 55916 1116
rect 55916 1060 55972 1116
rect 55972 1060 55976 1116
rect 55912 1056 55976 1060
rect 55992 1116 56056 1120
rect 55992 1060 55996 1116
rect 55996 1060 56052 1116
rect 56052 1060 56056 1116
rect 55992 1056 56056 1060
rect 57352 1116 57416 1120
rect 57352 1060 57356 1116
rect 57356 1060 57412 1116
rect 57412 1060 57416 1116
rect 57352 1056 57416 1060
rect 57432 1116 57496 1120
rect 57432 1060 57436 1116
rect 57436 1060 57492 1116
rect 57492 1060 57496 1116
rect 57432 1056 57496 1060
rect 57512 1116 57576 1120
rect 57512 1060 57516 1116
rect 57516 1060 57572 1116
rect 57572 1060 57576 1116
rect 57512 1056 57576 1060
rect 57592 1116 57656 1120
rect 57592 1060 57596 1116
rect 57596 1060 57652 1116
rect 57652 1060 57656 1116
rect 57592 1056 57656 1060
rect 58952 1116 59016 1120
rect 58952 1060 58956 1116
rect 58956 1060 59012 1116
rect 59012 1060 59016 1116
rect 58952 1056 59016 1060
rect 59032 1116 59096 1120
rect 59032 1060 59036 1116
rect 59036 1060 59092 1116
rect 59092 1060 59096 1116
rect 59032 1056 59096 1060
rect 59112 1116 59176 1120
rect 59112 1060 59116 1116
rect 59116 1060 59172 1116
rect 59172 1060 59176 1116
rect 59112 1056 59176 1060
rect 59192 1116 59256 1120
rect 59192 1060 59196 1116
rect 59196 1060 59252 1116
rect 59252 1060 59256 1116
rect 59192 1056 59256 1060
rect 60552 1116 60616 1120
rect 60552 1060 60556 1116
rect 60556 1060 60612 1116
rect 60612 1060 60616 1116
rect 60552 1056 60616 1060
rect 60632 1116 60696 1120
rect 60632 1060 60636 1116
rect 60636 1060 60692 1116
rect 60692 1060 60696 1116
rect 60632 1056 60696 1060
rect 60712 1116 60776 1120
rect 60712 1060 60716 1116
rect 60716 1060 60772 1116
rect 60772 1060 60776 1116
rect 60712 1056 60776 1060
rect 60792 1116 60856 1120
rect 60792 1060 60796 1116
rect 60796 1060 60852 1116
rect 60852 1060 60856 1116
rect 60792 1056 60856 1060
rect 62152 1116 62216 1120
rect 62152 1060 62156 1116
rect 62156 1060 62212 1116
rect 62212 1060 62216 1116
rect 62152 1056 62216 1060
rect 62232 1116 62296 1120
rect 62232 1060 62236 1116
rect 62236 1060 62292 1116
rect 62292 1060 62296 1116
rect 62232 1056 62296 1060
rect 62312 1116 62376 1120
rect 62312 1060 62316 1116
rect 62316 1060 62372 1116
rect 62372 1060 62376 1116
rect 62312 1056 62376 1060
rect 62392 1116 62456 1120
rect 62392 1060 62396 1116
rect 62396 1060 62452 1116
rect 62452 1060 62456 1116
rect 62392 1056 62456 1060
rect 63752 1116 63816 1120
rect 63752 1060 63756 1116
rect 63756 1060 63812 1116
rect 63812 1060 63816 1116
rect 63752 1056 63816 1060
rect 63832 1116 63896 1120
rect 63832 1060 63836 1116
rect 63836 1060 63892 1116
rect 63892 1060 63896 1116
rect 63832 1056 63896 1060
rect 63912 1116 63976 1120
rect 63912 1060 63916 1116
rect 63916 1060 63972 1116
rect 63972 1060 63976 1116
rect 63912 1056 63976 1060
rect 63992 1116 64056 1120
rect 63992 1060 63996 1116
rect 63996 1060 64052 1116
rect 64052 1060 64056 1116
rect 63992 1056 64056 1060
rect 65352 1116 65416 1120
rect 65352 1060 65356 1116
rect 65356 1060 65412 1116
rect 65412 1060 65416 1116
rect 65352 1056 65416 1060
rect 65432 1116 65496 1120
rect 65432 1060 65436 1116
rect 65436 1060 65492 1116
rect 65492 1060 65496 1116
rect 65432 1056 65496 1060
rect 65512 1116 65576 1120
rect 65512 1060 65516 1116
rect 65516 1060 65572 1116
rect 65572 1060 65576 1116
rect 65512 1056 65576 1060
rect 65592 1116 65656 1120
rect 65592 1060 65596 1116
rect 65596 1060 65652 1116
rect 65652 1060 65656 1116
rect 65592 1056 65656 1060
rect 66952 1116 67016 1120
rect 66952 1060 66956 1116
rect 66956 1060 67012 1116
rect 67012 1060 67016 1116
rect 66952 1056 67016 1060
rect 67032 1116 67096 1120
rect 67032 1060 67036 1116
rect 67036 1060 67092 1116
rect 67092 1060 67096 1116
rect 67032 1056 67096 1060
rect 67112 1116 67176 1120
rect 67112 1060 67116 1116
rect 67116 1060 67172 1116
rect 67172 1060 67176 1116
rect 67112 1056 67176 1060
rect 67192 1116 67256 1120
rect 67192 1060 67196 1116
rect 67196 1060 67252 1116
rect 67252 1060 67256 1116
rect 67192 1056 67256 1060
rect 68552 1116 68616 1120
rect 68552 1060 68556 1116
rect 68556 1060 68612 1116
rect 68612 1060 68616 1116
rect 68552 1056 68616 1060
rect 68632 1116 68696 1120
rect 68632 1060 68636 1116
rect 68636 1060 68692 1116
rect 68692 1060 68696 1116
rect 68632 1056 68696 1060
rect 68712 1116 68776 1120
rect 68712 1060 68716 1116
rect 68716 1060 68772 1116
rect 68772 1060 68776 1116
rect 68712 1056 68776 1060
rect 68792 1116 68856 1120
rect 68792 1060 68796 1116
rect 68796 1060 68852 1116
rect 68852 1060 68856 1116
rect 68792 1056 68856 1060
rect 70152 1116 70216 1120
rect 70152 1060 70156 1116
rect 70156 1060 70212 1116
rect 70212 1060 70216 1116
rect 70152 1056 70216 1060
rect 70232 1116 70296 1120
rect 70232 1060 70236 1116
rect 70236 1060 70292 1116
rect 70292 1060 70296 1116
rect 70232 1056 70296 1060
rect 70312 1116 70376 1120
rect 70312 1060 70316 1116
rect 70316 1060 70372 1116
rect 70372 1060 70376 1116
rect 70312 1056 70376 1060
rect 70392 1116 70456 1120
rect 70392 1060 70396 1116
rect 70396 1060 70452 1116
rect 70452 1060 70456 1116
rect 70392 1056 70456 1060
rect 71752 1116 71816 1120
rect 71752 1060 71756 1116
rect 71756 1060 71812 1116
rect 71812 1060 71816 1116
rect 71752 1056 71816 1060
rect 71832 1116 71896 1120
rect 71832 1060 71836 1116
rect 71836 1060 71892 1116
rect 71892 1060 71896 1116
rect 71832 1056 71896 1060
rect 71912 1116 71976 1120
rect 71912 1060 71916 1116
rect 71916 1060 71972 1116
rect 71972 1060 71976 1116
rect 71912 1056 71976 1060
rect 71992 1116 72056 1120
rect 71992 1060 71996 1116
rect 71996 1060 72052 1116
rect 72052 1060 72056 1116
rect 71992 1056 72056 1060
rect 73352 1116 73416 1120
rect 73352 1060 73356 1116
rect 73356 1060 73412 1116
rect 73412 1060 73416 1116
rect 73352 1056 73416 1060
rect 73432 1116 73496 1120
rect 73432 1060 73436 1116
rect 73436 1060 73492 1116
rect 73492 1060 73496 1116
rect 73432 1056 73496 1060
rect 73512 1116 73576 1120
rect 73512 1060 73516 1116
rect 73516 1060 73572 1116
rect 73572 1060 73576 1116
rect 73512 1056 73576 1060
rect 73592 1116 73656 1120
rect 73592 1060 73596 1116
rect 73596 1060 73652 1116
rect 73652 1060 73656 1116
rect 73592 1056 73656 1060
rect 74952 1116 75016 1120
rect 74952 1060 74956 1116
rect 74956 1060 75012 1116
rect 75012 1060 75016 1116
rect 74952 1056 75016 1060
rect 75032 1116 75096 1120
rect 75032 1060 75036 1116
rect 75036 1060 75092 1116
rect 75092 1060 75096 1116
rect 75032 1056 75096 1060
rect 75112 1116 75176 1120
rect 75112 1060 75116 1116
rect 75116 1060 75172 1116
rect 75172 1060 75176 1116
rect 75112 1056 75176 1060
rect 75192 1116 75256 1120
rect 75192 1060 75196 1116
rect 75196 1060 75252 1116
rect 75252 1060 75256 1116
rect 75192 1056 75256 1060
rect 76552 1116 76616 1120
rect 76552 1060 76556 1116
rect 76556 1060 76612 1116
rect 76612 1060 76616 1116
rect 76552 1056 76616 1060
rect 76632 1116 76696 1120
rect 76632 1060 76636 1116
rect 76636 1060 76692 1116
rect 76692 1060 76696 1116
rect 76632 1056 76696 1060
rect 76712 1116 76776 1120
rect 76712 1060 76716 1116
rect 76716 1060 76772 1116
rect 76772 1060 76776 1116
rect 76712 1056 76776 1060
rect 76792 1116 76856 1120
rect 76792 1060 76796 1116
rect 76796 1060 76852 1116
rect 76852 1060 76856 1116
rect 76792 1056 76856 1060
rect 78152 1116 78216 1120
rect 78152 1060 78156 1116
rect 78156 1060 78212 1116
rect 78212 1060 78216 1116
rect 78152 1056 78216 1060
rect 78232 1116 78296 1120
rect 78232 1060 78236 1116
rect 78236 1060 78292 1116
rect 78292 1060 78296 1116
rect 78232 1056 78296 1060
rect 78312 1116 78376 1120
rect 78312 1060 78316 1116
rect 78316 1060 78372 1116
rect 78372 1060 78376 1116
rect 78312 1056 78376 1060
rect 78392 1116 78456 1120
rect 78392 1060 78396 1116
rect 78396 1060 78452 1116
rect 78452 1060 78456 1116
rect 78392 1056 78456 1060
rect 79752 1116 79816 1120
rect 79752 1060 79756 1116
rect 79756 1060 79812 1116
rect 79812 1060 79816 1116
rect 79752 1056 79816 1060
rect 79832 1116 79896 1120
rect 79832 1060 79836 1116
rect 79836 1060 79892 1116
rect 79892 1060 79896 1116
rect 79832 1056 79896 1060
rect 79912 1116 79976 1120
rect 79912 1060 79916 1116
rect 79916 1060 79972 1116
rect 79972 1060 79976 1116
rect 79912 1056 79976 1060
rect 79992 1116 80056 1120
rect 79992 1060 79996 1116
rect 79996 1060 80052 1116
rect 80052 1060 80056 1116
rect 79992 1056 80056 1060
rect 81352 1116 81416 1120
rect 81352 1060 81356 1116
rect 81356 1060 81412 1116
rect 81412 1060 81416 1116
rect 81352 1056 81416 1060
rect 81432 1116 81496 1120
rect 81432 1060 81436 1116
rect 81436 1060 81492 1116
rect 81492 1060 81496 1116
rect 81432 1056 81496 1060
rect 81512 1116 81576 1120
rect 81512 1060 81516 1116
rect 81516 1060 81572 1116
rect 81572 1060 81576 1116
rect 81512 1056 81576 1060
rect 81592 1116 81656 1120
rect 81592 1060 81596 1116
rect 81596 1060 81652 1116
rect 81652 1060 81656 1116
rect 81592 1056 81656 1060
rect 82952 1116 83016 1120
rect 82952 1060 82956 1116
rect 82956 1060 83012 1116
rect 83012 1060 83016 1116
rect 82952 1056 83016 1060
rect 83032 1116 83096 1120
rect 83032 1060 83036 1116
rect 83036 1060 83092 1116
rect 83092 1060 83096 1116
rect 83032 1056 83096 1060
rect 83112 1116 83176 1120
rect 83112 1060 83116 1116
rect 83116 1060 83172 1116
rect 83172 1060 83176 1116
rect 83112 1056 83176 1060
rect 83192 1116 83256 1120
rect 83192 1060 83196 1116
rect 83196 1060 83252 1116
rect 83252 1060 83256 1116
rect 83192 1056 83256 1060
rect 84552 1116 84616 1120
rect 84552 1060 84556 1116
rect 84556 1060 84612 1116
rect 84612 1060 84616 1116
rect 84552 1056 84616 1060
rect 84632 1116 84696 1120
rect 84632 1060 84636 1116
rect 84636 1060 84692 1116
rect 84692 1060 84696 1116
rect 84632 1056 84696 1060
rect 84712 1116 84776 1120
rect 84712 1060 84716 1116
rect 84716 1060 84772 1116
rect 84772 1060 84776 1116
rect 84712 1056 84776 1060
rect 84792 1116 84856 1120
rect 84792 1060 84796 1116
rect 84796 1060 84852 1116
rect 84852 1060 84856 1116
rect 84792 1056 84856 1060
rect 86152 1116 86216 1120
rect 86152 1060 86156 1116
rect 86156 1060 86212 1116
rect 86212 1060 86216 1116
rect 86152 1056 86216 1060
rect 86232 1116 86296 1120
rect 86232 1060 86236 1116
rect 86236 1060 86292 1116
rect 86292 1060 86296 1116
rect 86232 1056 86296 1060
rect 86312 1116 86376 1120
rect 86312 1060 86316 1116
rect 86316 1060 86372 1116
rect 86372 1060 86376 1116
rect 86312 1056 86376 1060
rect 86392 1116 86456 1120
rect 86392 1060 86396 1116
rect 86396 1060 86452 1116
rect 86452 1060 86456 1116
rect 86392 1056 86456 1060
rect 87752 1116 87816 1120
rect 87752 1060 87756 1116
rect 87756 1060 87812 1116
rect 87812 1060 87816 1116
rect 87752 1056 87816 1060
rect 87832 1116 87896 1120
rect 87832 1060 87836 1116
rect 87836 1060 87892 1116
rect 87892 1060 87896 1116
rect 87832 1056 87896 1060
rect 87912 1116 87976 1120
rect 87912 1060 87916 1116
rect 87916 1060 87972 1116
rect 87972 1060 87976 1116
rect 87912 1056 87976 1060
rect 87992 1116 88056 1120
rect 87992 1060 87996 1116
rect 87996 1060 88052 1116
rect 88052 1060 88056 1116
rect 87992 1056 88056 1060
rect 89352 1116 89416 1120
rect 89352 1060 89356 1116
rect 89356 1060 89412 1116
rect 89412 1060 89416 1116
rect 89352 1056 89416 1060
rect 89432 1116 89496 1120
rect 89432 1060 89436 1116
rect 89436 1060 89492 1116
rect 89492 1060 89496 1116
rect 89432 1056 89496 1060
rect 89512 1116 89576 1120
rect 89512 1060 89516 1116
rect 89516 1060 89572 1116
rect 89572 1060 89576 1116
rect 89512 1056 89576 1060
rect 89592 1116 89656 1120
rect 89592 1060 89596 1116
rect 89596 1060 89652 1116
rect 89652 1060 89656 1116
rect 89592 1056 89656 1060
rect 90952 1116 91016 1120
rect 90952 1060 90956 1116
rect 90956 1060 91012 1116
rect 91012 1060 91016 1116
rect 90952 1056 91016 1060
rect 91032 1116 91096 1120
rect 91032 1060 91036 1116
rect 91036 1060 91092 1116
rect 91092 1060 91096 1116
rect 91032 1056 91096 1060
rect 91112 1116 91176 1120
rect 91112 1060 91116 1116
rect 91116 1060 91172 1116
rect 91172 1060 91176 1116
rect 91112 1056 91176 1060
rect 91192 1116 91256 1120
rect 91192 1060 91196 1116
rect 91196 1060 91252 1116
rect 91252 1060 91256 1116
rect 91192 1056 91256 1060
rect 92552 1116 92616 1120
rect 92552 1060 92556 1116
rect 92556 1060 92612 1116
rect 92612 1060 92616 1116
rect 92552 1056 92616 1060
rect 92632 1116 92696 1120
rect 92632 1060 92636 1116
rect 92636 1060 92692 1116
rect 92692 1060 92696 1116
rect 92632 1056 92696 1060
rect 92712 1116 92776 1120
rect 92712 1060 92716 1116
rect 92716 1060 92772 1116
rect 92772 1060 92776 1116
rect 92712 1056 92776 1060
rect 92792 1116 92856 1120
rect 92792 1060 92796 1116
rect 92796 1060 92852 1116
rect 92852 1060 92856 1116
rect 92792 1056 92856 1060
rect 94152 1116 94216 1120
rect 94152 1060 94156 1116
rect 94156 1060 94212 1116
rect 94212 1060 94216 1116
rect 94152 1056 94216 1060
rect 94232 1116 94296 1120
rect 94232 1060 94236 1116
rect 94236 1060 94292 1116
rect 94292 1060 94296 1116
rect 94232 1056 94296 1060
rect 94312 1116 94376 1120
rect 94312 1060 94316 1116
rect 94316 1060 94372 1116
rect 94372 1060 94376 1116
rect 94312 1056 94376 1060
rect 94392 1116 94456 1120
rect 94392 1060 94396 1116
rect 94396 1060 94452 1116
rect 94452 1060 94456 1116
rect 94392 1056 94456 1060
rect 95752 1116 95816 1120
rect 95752 1060 95756 1116
rect 95756 1060 95812 1116
rect 95812 1060 95816 1116
rect 95752 1056 95816 1060
rect 95832 1116 95896 1120
rect 95832 1060 95836 1116
rect 95836 1060 95892 1116
rect 95892 1060 95896 1116
rect 95832 1056 95896 1060
rect 95912 1116 95976 1120
rect 95912 1060 95916 1116
rect 95916 1060 95972 1116
rect 95972 1060 95976 1116
rect 95912 1056 95976 1060
rect 95992 1116 96056 1120
rect 95992 1060 95996 1116
rect 95996 1060 96052 1116
rect 96052 1060 96056 1116
rect 95992 1056 96056 1060
rect 97352 1116 97416 1120
rect 97352 1060 97356 1116
rect 97356 1060 97412 1116
rect 97412 1060 97416 1116
rect 97352 1056 97416 1060
rect 97432 1116 97496 1120
rect 97432 1060 97436 1116
rect 97436 1060 97492 1116
rect 97492 1060 97496 1116
rect 97432 1056 97496 1060
rect 97512 1116 97576 1120
rect 97512 1060 97516 1116
rect 97516 1060 97572 1116
rect 97572 1060 97576 1116
rect 97512 1056 97576 1060
rect 97592 1116 97656 1120
rect 97592 1060 97596 1116
rect 97596 1060 97652 1116
rect 97652 1060 97656 1116
rect 97592 1056 97656 1060
rect 98952 1116 99016 1120
rect 98952 1060 98956 1116
rect 98956 1060 99012 1116
rect 99012 1060 99016 1116
rect 98952 1056 99016 1060
rect 99032 1116 99096 1120
rect 99032 1060 99036 1116
rect 99036 1060 99092 1116
rect 99092 1060 99096 1116
rect 99032 1056 99096 1060
rect 99112 1116 99176 1120
rect 99112 1060 99116 1116
rect 99116 1060 99172 1116
rect 99172 1060 99176 1116
rect 99112 1056 99176 1060
rect 99192 1116 99256 1120
rect 99192 1060 99196 1116
rect 99196 1060 99252 1116
rect 99252 1060 99256 1116
rect 99192 1056 99256 1060
rect 100552 1116 100616 1120
rect 100552 1060 100556 1116
rect 100556 1060 100612 1116
rect 100612 1060 100616 1116
rect 100552 1056 100616 1060
rect 100632 1116 100696 1120
rect 100632 1060 100636 1116
rect 100636 1060 100692 1116
rect 100692 1060 100696 1116
rect 100632 1056 100696 1060
rect 100712 1116 100776 1120
rect 100712 1060 100716 1116
rect 100716 1060 100772 1116
rect 100772 1060 100776 1116
rect 100712 1056 100776 1060
rect 100792 1116 100856 1120
rect 100792 1060 100796 1116
rect 100796 1060 100852 1116
rect 100852 1060 100856 1116
rect 100792 1056 100856 1060
rect 102152 1116 102216 1120
rect 102152 1060 102156 1116
rect 102156 1060 102212 1116
rect 102212 1060 102216 1116
rect 102152 1056 102216 1060
rect 102232 1116 102296 1120
rect 102232 1060 102236 1116
rect 102236 1060 102292 1116
rect 102292 1060 102296 1116
rect 102232 1056 102296 1060
rect 102312 1116 102376 1120
rect 102312 1060 102316 1116
rect 102316 1060 102372 1116
rect 102372 1060 102376 1116
rect 102312 1056 102376 1060
rect 102392 1116 102456 1120
rect 102392 1060 102396 1116
rect 102396 1060 102452 1116
rect 102452 1060 102456 1116
rect 102392 1056 102456 1060
rect 103752 1116 103816 1120
rect 103752 1060 103756 1116
rect 103756 1060 103812 1116
rect 103812 1060 103816 1116
rect 103752 1056 103816 1060
rect 103832 1116 103896 1120
rect 103832 1060 103836 1116
rect 103836 1060 103892 1116
rect 103892 1060 103896 1116
rect 103832 1056 103896 1060
rect 103912 1116 103976 1120
rect 103912 1060 103916 1116
rect 103916 1060 103972 1116
rect 103972 1060 103976 1116
rect 103912 1056 103976 1060
rect 103992 1116 104056 1120
rect 103992 1060 103996 1116
rect 103996 1060 104052 1116
rect 104052 1060 104056 1116
rect 103992 1056 104056 1060
rect 105352 1116 105416 1120
rect 105352 1060 105356 1116
rect 105356 1060 105412 1116
rect 105412 1060 105416 1116
rect 105352 1056 105416 1060
rect 105432 1116 105496 1120
rect 105432 1060 105436 1116
rect 105436 1060 105492 1116
rect 105492 1060 105496 1116
rect 105432 1056 105496 1060
rect 105512 1116 105576 1120
rect 105512 1060 105516 1116
rect 105516 1060 105572 1116
rect 105572 1060 105576 1116
rect 105512 1056 105576 1060
rect 105592 1116 105656 1120
rect 105592 1060 105596 1116
rect 105596 1060 105652 1116
rect 105652 1060 105656 1116
rect 105592 1056 105656 1060
rect 106952 1116 107016 1120
rect 106952 1060 106956 1116
rect 106956 1060 107012 1116
rect 107012 1060 107016 1116
rect 106952 1056 107016 1060
rect 107032 1116 107096 1120
rect 107032 1060 107036 1116
rect 107036 1060 107092 1116
rect 107092 1060 107096 1116
rect 107032 1056 107096 1060
rect 107112 1116 107176 1120
rect 107112 1060 107116 1116
rect 107116 1060 107172 1116
rect 107172 1060 107176 1116
rect 107112 1056 107176 1060
rect 107192 1116 107256 1120
rect 107192 1060 107196 1116
rect 107196 1060 107252 1116
rect 107252 1060 107256 1116
rect 107192 1056 107256 1060
rect 108552 1116 108616 1120
rect 108552 1060 108556 1116
rect 108556 1060 108612 1116
rect 108612 1060 108616 1116
rect 108552 1056 108616 1060
rect 108632 1116 108696 1120
rect 108632 1060 108636 1116
rect 108636 1060 108692 1116
rect 108692 1060 108696 1116
rect 108632 1056 108696 1060
rect 108712 1116 108776 1120
rect 108712 1060 108716 1116
rect 108716 1060 108772 1116
rect 108772 1060 108776 1116
rect 108712 1056 108776 1060
rect 108792 1116 108856 1120
rect 108792 1060 108796 1116
rect 108796 1060 108852 1116
rect 108852 1060 108856 1116
rect 108792 1056 108856 1060
rect 53052 852 53116 916
rect 93900 716 93964 780
rect 10732 580 10796 644
rect 27476 580 27540 644
rect 52316 580 52380 644
rect 41828 444 41892 508
<< metal4 >>
rect -1076 88634 -756 88676
rect -1076 88398 -1034 88634
rect -798 88398 -756 88634
rect -1076 82206 -756 88398
rect 2944 88634 3264 88676
rect 2944 88398 2986 88634
rect 3222 88398 3264 88634
rect -1076 81970 -1034 82206
rect -798 81970 -756 82206
rect -1076 6206 -756 81970
rect -1076 5970 -1034 6206
rect -798 5970 -756 6206
rect -1076 -814 -756 5970
rect -416 87974 -96 88016
rect -416 87738 -374 87974
rect -138 87738 -96 87974
rect -416 82866 -96 87738
rect -416 82630 -374 82866
rect -138 82630 -96 82866
rect -416 6866 -96 82630
rect 2944 85984 3264 88398
rect 2944 85920 2952 85984
rect 3016 85920 3032 85984
rect 3096 85920 3112 85984
rect 3176 85920 3192 85984
rect 3256 85920 3264 85984
rect 2944 84896 3264 85920
rect 2944 84832 2952 84896
rect 3016 84832 3032 84896
rect 3096 84832 3112 84896
rect 3176 84832 3192 84896
rect 3256 84832 3264 84896
rect 2944 83808 3264 84832
rect 2944 83744 2952 83808
rect 3016 83744 3032 83808
rect 3096 83744 3112 83808
rect 3176 83744 3192 83808
rect 3256 83744 3264 83808
rect 2944 82720 3264 83744
rect 2944 82656 2952 82720
rect 3016 82656 3032 82720
rect 3096 82656 3112 82720
rect 3176 82656 3192 82720
rect 3256 82656 3264 82720
rect 2944 82206 3264 82656
rect 2944 81970 2986 82206
rect 3222 81970 3264 82206
rect 2944 81632 3264 81970
rect 2944 81568 2952 81632
rect 3016 81568 3032 81632
rect 3096 81568 3112 81632
rect 3176 81568 3192 81632
rect 3256 81568 3264 81632
rect 2944 80544 3264 81568
rect 2944 80480 2952 80544
rect 3016 80480 3032 80544
rect 3096 80480 3112 80544
rect 3176 80480 3192 80544
rect 3256 80480 3264 80544
rect 2944 79456 3264 80480
rect 2944 79392 2952 79456
rect 3016 79392 3032 79456
rect 3096 79392 3112 79456
rect 3176 79392 3192 79456
rect 3256 79392 3264 79456
rect 2944 78368 3264 79392
rect 2944 78304 2952 78368
rect 3016 78304 3032 78368
rect 3096 78304 3112 78368
rect 3176 78304 3192 78368
rect 3256 78304 3264 78368
rect 2944 77280 3264 78304
rect 2944 77216 2952 77280
rect 3016 77216 3032 77280
rect 3096 77216 3112 77280
rect 3176 77216 3192 77280
rect 3256 77216 3264 77280
rect 2944 76192 3264 77216
rect 2944 76128 2952 76192
rect 3016 76128 3032 76192
rect 3096 76128 3112 76192
rect 3176 76128 3192 76192
rect 3256 76128 3264 76192
rect 2944 75104 3264 76128
rect 2944 75040 2952 75104
rect 3016 75040 3032 75104
rect 3096 75040 3112 75104
rect 3176 75040 3192 75104
rect 3256 75040 3264 75104
rect 2944 74016 3264 75040
rect 2944 73952 2952 74016
rect 3016 73952 3032 74016
rect 3096 73952 3112 74016
rect 3176 73952 3192 74016
rect 3256 73952 3264 74016
rect 2944 72928 3264 73952
rect 2944 72864 2952 72928
rect 3016 72864 3032 72928
rect 3096 72864 3112 72928
rect 3176 72864 3192 72928
rect 3256 72864 3264 72928
rect 795 71908 861 71909
rect 795 71844 796 71908
rect 860 71844 861 71908
rect 795 71843 861 71844
rect 798 37365 858 71843
rect 2944 71840 3264 72864
rect 2944 71776 2952 71840
rect 3016 71776 3032 71840
rect 3096 71776 3112 71840
rect 3176 71776 3192 71840
rect 3256 71776 3264 71840
rect 2944 70752 3264 71776
rect 2944 70688 2952 70752
rect 3016 70688 3032 70752
rect 3096 70688 3112 70752
rect 3176 70688 3192 70752
rect 3256 70688 3264 70752
rect 2944 69664 3264 70688
rect 2944 69600 2952 69664
rect 3016 69600 3032 69664
rect 3096 69600 3112 69664
rect 3176 69600 3192 69664
rect 3256 69600 3264 69664
rect 2944 68576 3264 69600
rect 2944 68512 2952 68576
rect 3016 68512 3032 68576
rect 3096 68512 3112 68576
rect 3176 68512 3192 68576
rect 3256 68512 3264 68576
rect 2944 67488 3264 68512
rect 2944 67424 2952 67488
rect 3016 67424 3032 67488
rect 3096 67424 3112 67488
rect 3176 67424 3192 67488
rect 3256 67424 3264 67488
rect 2944 66400 3264 67424
rect 2944 66336 2952 66400
rect 3016 66336 3032 66400
rect 3096 66336 3112 66400
rect 3176 66336 3192 66400
rect 3256 66336 3264 66400
rect 2944 65312 3264 66336
rect 2944 65248 2952 65312
rect 3016 65248 3032 65312
rect 3096 65248 3112 65312
rect 3176 65248 3192 65312
rect 3256 65248 3264 65312
rect 2944 64224 3264 65248
rect 2944 64160 2952 64224
rect 3016 64160 3032 64224
rect 3096 64160 3112 64224
rect 3176 64160 3192 64224
rect 3256 64160 3264 64224
rect 2944 63136 3264 64160
rect 2944 63072 2952 63136
rect 3016 63072 3032 63136
rect 3096 63072 3112 63136
rect 3176 63072 3192 63136
rect 3256 63072 3264 63136
rect 2944 62048 3264 63072
rect 2944 61984 2952 62048
rect 3016 61984 3032 62048
rect 3096 61984 3112 62048
rect 3176 61984 3192 62048
rect 3256 61984 3264 62048
rect 2944 60960 3264 61984
rect 2944 60896 2952 60960
rect 3016 60896 3032 60960
rect 3096 60896 3112 60960
rect 3176 60896 3192 60960
rect 3256 60896 3264 60960
rect 2944 59872 3264 60896
rect 2944 59808 2952 59872
rect 3016 59808 3032 59872
rect 3096 59808 3112 59872
rect 3176 59808 3192 59872
rect 3256 59808 3264 59872
rect 2944 58784 3264 59808
rect 2944 58720 2952 58784
rect 3016 58720 3032 58784
rect 3096 58720 3112 58784
rect 3176 58720 3192 58784
rect 3256 58720 3264 58784
rect 2944 57696 3264 58720
rect 2944 57632 2952 57696
rect 3016 57632 3032 57696
rect 3096 57632 3112 57696
rect 3176 57632 3192 57696
rect 3256 57632 3264 57696
rect 2944 56608 3264 57632
rect 2944 56544 2952 56608
rect 3016 56544 3032 56608
rect 3096 56544 3112 56608
rect 3176 56544 3192 56608
rect 3256 56544 3264 56608
rect 2944 55520 3264 56544
rect 2944 55456 2952 55520
rect 3016 55456 3032 55520
rect 3096 55456 3112 55520
rect 3176 55456 3192 55520
rect 3256 55456 3264 55520
rect 2944 54432 3264 55456
rect 2944 54368 2952 54432
rect 3016 54368 3032 54432
rect 3096 54368 3112 54432
rect 3176 54368 3192 54432
rect 3256 54368 3264 54432
rect 2944 53344 3264 54368
rect 2944 53280 2952 53344
rect 3016 53280 3032 53344
rect 3096 53280 3112 53344
rect 3176 53280 3192 53344
rect 3256 53280 3264 53344
rect 2944 52256 3264 53280
rect 2944 52192 2952 52256
rect 3016 52192 3032 52256
rect 3096 52192 3112 52256
rect 3176 52192 3192 52256
rect 3256 52192 3264 52256
rect 2944 51168 3264 52192
rect 2944 51104 2952 51168
rect 3016 51104 3032 51168
rect 3096 51104 3112 51168
rect 3176 51104 3192 51168
rect 3256 51104 3264 51168
rect 2944 50080 3264 51104
rect 2944 50016 2952 50080
rect 3016 50016 3032 50080
rect 3096 50016 3112 50080
rect 3176 50016 3192 50080
rect 3256 50016 3264 50080
rect 2944 48992 3264 50016
rect 2944 48928 2952 48992
rect 3016 48928 3032 48992
rect 3096 48928 3112 48992
rect 3176 48928 3192 48992
rect 3256 48928 3264 48992
rect 2944 47904 3264 48928
rect 2944 47840 2952 47904
rect 3016 47840 3032 47904
rect 3096 47840 3112 47904
rect 3176 47840 3192 47904
rect 3256 47840 3264 47904
rect 2944 46816 3264 47840
rect 2944 46752 2952 46816
rect 3016 46752 3032 46816
rect 3096 46752 3112 46816
rect 3176 46752 3192 46816
rect 3256 46752 3264 46816
rect 2944 45728 3264 46752
rect 2944 45664 2952 45728
rect 3016 45664 3032 45728
rect 3096 45664 3112 45728
rect 3176 45664 3192 45728
rect 3256 45664 3264 45728
rect 2944 44640 3264 45664
rect 2944 44576 2952 44640
rect 3016 44576 3032 44640
rect 3096 44576 3112 44640
rect 3176 44576 3192 44640
rect 3256 44576 3264 44640
rect 2944 43552 3264 44576
rect 2944 43488 2952 43552
rect 3016 43488 3032 43552
rect 3096 43488 3112 43552
rect 3176 43488 3192 43552
rect 3256 43488 3264 43552
rect 2944 42464 3264 43488
rect 2944 42400 2952 42464
rect 3016 42400 3032 42464
rect 3096 42400 3112 42464
rect 3176 42400 3192 42464
rect 3256 42400 3264 42464
rect 2944 41376 3264 42400
rect 2944 41312 2952 41376
rect 3016 41312 3032 41376
rect 3096 41312 3112 41376
rect 3176 41312 3192 41376
rect 3256 41312 3264 41376
rect 2944 40288 3264 41312
rect 2944 40224 2952 40288
rect 3016 40224 3032 40288
rect 3096 40224 3112 40288
rect 3176 40224 3192 40288
rect 3256 40224 3264 40288
rect 2944 39200 3264 40224
rect 2944 39136 2952 39200
rect 3016 39136 3032 39200
rect 3096 39136 3112 39200
rect 3176 39136 3192 39200
rect 3256 39136 3264 39200
rect 2944 38112 3264 39136
rect 2944 38048 2952 38112
rect 3016 38048 3032 38112
rect 3096 38048 3112 38112
rect 3176 38048 3192 38112
rect 3256 38048 3264 38112
rect 795 37364 861 37365
rect 795 37300 796 37364
rect 860 37300 861 37364
rect 795 37299 861 37300
rect -416 6630 -374 6866
rect -138 6630 -96 6866
rect -416 -154 -96 6630
rect -416 -390 -374 -154
rect -138 -390 -96 -154
rect -416 -432 -96 -390
rect 2944 37024 3264 38048
rect 2944 36960 2952 37024
rect 3016 36960 3032 37024
rect 3096 36960 3112 37024
rect 3176 36960 3192 37024
rect 3256 36960 3264 37024
rect 2944 35936 3264 36960
rect 2944 35872 2952 35936
rect 3016 35872 3032 35936
rect 3096 35872 3112 35936
rect 3176 35872 3192 35936
rect 3256 35872 3264 35936
rect 2944 34848 3264 35872
rect 2944 34784 2952 34848
rect 3016 34784 3032 34848
rect 3096 34784 3112 34848
rect 3176 34784 3192 34848
rect 3256 34784 3264 34848
rect 2944 33760 3264 34784
rect 2944 33696 2952 33760
rect 3016 33696 3032 33760
rect 3096 33696 3112 33760
rect 3176 33696 3192 33760
rect 3256 33696 3264 33760
rect 2944 32672 3264 33696
rect 2944 32608 2952 32672
rect 3016 32608 3032 32672
rect 3096 32608 3112 32672
rect 3176 32608 3192 32672
rect 3256 32608 3264 32672
rect 2944 31584 3264 32608
rect 2944 31520 2952 31584
rect 3016 31520 3032 31584
rect 3096 31520 3112 31584
rect 3176 31520 3192 31584
rect 3256 31520 3264 31584
rect 2944 30496 3264 31520
rect 2944 30432 2952 30496
rect 3016 30432 3032 30496
rect 3096 30432 3112 30496
rect 3176 30432 3192 30496
rect 3256 30432 3264 30496
rect 2944 29408 3264 30432
rect 2944 29344 2952 29408
rect 3016 29344 3032 29408
rect 3096 29344 3112 29408
rect 3176 29344 3192 29408
rect 3256 29344 3264 29408
rect 2944 28320 3264 29344
rect 2944 28256 2952 28320
rect 3016 28256 3032 28320
rect 3096 28256 3112 28320
rect 3176 28256 3192 28320
rect 3256 28256 3264 28320
rect 2944 27232 3264 28256
rect 2944 27168 2952 27232
rect 3016 27168 3032 27232
rect 3096 27168 3112 27232
rect 3176 27168 3192 27232
rect 3256 27168 3264 27232
rect 2944 26144 3264 27168
rect 2944 26080 2952 26144
rect 3016 26080 3032 26144
rect 3096 26080 3112 26144
rect 3176 26080 3192 26144
rect 3256 26080 3264 26144
rect 2944 25056 3264 26080
rect 2944 24992 2952 25056
rect 3016 24992 3032 25056
rect 3096 24992 3112 25056
rect 3176 24992 3192 25056
rect 3256 24992 3264 25056
rect 2944 23968 3264 24992
rect 2944 23904 2952 23968
rect 3016 23904 3032 23968
rect 3096 23904 3112 23968
rect 3176 23904 3192 23968
rect 3256 23904 3264 23968
rect 2944 22880 3264 23904
rect 2944 22816 2952 22880
rect 3016 22816 3032 22880
rect 3096 22816 3112 22880
rect 3176 22816 3192 22880
rect 3256 22816 3264 22880
rect 2944 21792 3264 22816
rect 2944 21728 2952 21792
rect 3016 21728 3032 21792
rect 3096 21728 3112 21792
rect 3176 21728 3192 21792
rect 3256 21728 3264 21792
rect 2944 20704 3264 21728
rect 2944 20640 2952 20704
rect 3016 20640 3032 20704
rect 3096 20640 3112 20704
rect 3176 20640 3192 20704
rect 3256 20640 3264 20704
rect 2944 19616 3264 20640
rect 2944 19552 2952 19616
rect 3016 19552 3032 19616
rect 3096 19552 3112 19616
rect 3176 19552 3192 19616
rect 3256 19552 3264 19616
rect 2944 18528 3264 19552
rect 2944 18464 2952 18528
rect 3016 18464 3032 18528
rect 3096 18464 3112 18528
rect 3176 18464 3192 18528
rect 3256 18464 3264 18528
rect 2944 17440 3264 18464
rect 2944 17376 2952 17440
rect 3016 17376 3032 17440
rect 3096 17376 3112 17440
rect 3176 17376 3192 17440
rect 3256 17376 3264 17440
rect 2944 16352 3264 17376
rect 2944 16288 2952 16352
rect 3016 16288 3032 16352
rect 3096 16288 3112 16352
rect 3176 16288 3192 16352
rect 3256 16288 3264 16352
rect 2944 15264 3264 16288
rect 2944 15200 2952 15264
rect 3016 15200 3032 15264
rect 3096 15200 3112 15264
rect 3176 15200 3192 15264
rect 3256 15200 3264 15264
rect 2944 14176 3264 15200
rect 2944 14112 2952 14176
rect 3016 14112 3032 14176
rect 3096 14112 3112 14176
rect 3176 14112 3192 14176
rect 3256 14112 3264 14176
rect 2944 13088 3264 14112
rect 2944 13024 2952 13088
rect 3016 13024 3032 13088
rect 3096 13024 3112 13088
rect 3176 13024 3192 13088
rect 3256 13024 3264 13088
rect 2944 12000 3264 13024
rect 2944 11936 2952 12000
rect 3016 11936 3032 12000
rect 3096 11936 3112 12000
rect 3176 11936 3192 12000
rect 3256 11936 3264 12000
rect 2944 10912 3264 11936
rect 2944 10848 2952 10912
rect 3016 10848 3032 10912
rect 3096 10848 3112 10912
rect 3176 10848 3192 10912
rect 3256 10848 3264 10912
rect 2944 9824 3264 10848
rect 2944 9760 2952 9824
rect 3016 9760 3032 9824
rect 3096 9760 3112 9824
rect 3176 9760 3192 9824
rect 3256 9760 3264 9824
rect 2944 8736 3264 9760
rect 2944 8672 2952 8736
rect 3016 8672 3032 8736
rect 3096 8672 3112 8736
rect 3176 8672 3192 8736
rect 3256 8672 3264 8736
rect 2944 7648 3264 8672
rect 2944 7584 2952 7648
rect 3016 7584 3032 7648
rect 3096 7584 3112 7648
rect 3176 7584 3192 7648
rect 3256 7584 3264 7648
rect 2944 6560 3264 7584
rect 2944 6496 2952 6560
rect 3016 6496 3032 6560
rect 3096 6496 3112 6560
rect 3176 6496 3192 6560
rect 3256 6496 3264 6560
rect 2944 6206 3264 6496
rect 2944 5970 2986 6206
rect 3222 5970 3264 6206
rect 2944 5472 3264 5970
rect 2944 5408 2952 5472
rect 3016 5408 3032 5472
rect 3096 5408 3112 5472
rect 3176 5408 3192 5472
rect 3256 5408 3264 5472
rect 2944 4384 3264 5408
rect 2944 4320 2952 4384
rect 3016 4320 3032 4384
rect 3096 4320 3112 4384
rect 3176 4320 3192 4384
rect 3256 4320 3264 4384
rect 2944 3296 3264 4320
rect 2944 3232 2952 3296
rect 3016 3232 3032 3296
rect 3096 3232 3112 3296
rect 3176 3232 3192 3296
rect 3256 3232 3264 3296
rect 2944 2208 3264 3232
rect 2944 2144 2952 2208
rect 3016 2144 3032 2208
rect 3096 2144 3112 2208
rect 3176 2144 3192 2208
rect 3256 2144 3264 2208
rect 2944 1120 3264 2144
rect 2944 1056 2952 1120
rect 3016 1056 3032 1120
rect 3096 1056 3112 1120
rect 3176 1056 3192 1120
rect 3256 1056 3264 1120
rect -1076 -1050 -1034 -814
rect -798 -1050 -756 -814
rect -1076 -1092 -756 -1050
rect 2944 -814 3264 1056
rect 2944 -1050 2986 -814
rect 3222 -1050 3264 -814
rect 2944 -1092 3264 -1050
rect 3604 87974 3924 88676
rect 3604 87738 3646 87974
rect 3882 87738 3924 87974
rect 3604 86528 3924 87738
rect 3604 86464 3612 86528
rect 3676 86464 3692 86528
rect 3756 86464 3772 86528
rect 3836 86464 3852 86528
rect 3916 86464 3924 86528
rect 3604 85440 3924 86464
rect 3604 85376 3612 85440
rect 3676 85376 3692 85440
rect 3756 85376 3772 85440
rect 3836 85376 3852 85440
rect 3916 85376 3924 85440
rect 3604 84352 3924 85376
rect 3604 84288 3612 84352
rect 3676 84288 3692 84352
rect 3756 84288 3772 84352
rect 3836 84288 3852 84352
rect 3916 84288 3924 84352
rect 3604 83264 3924 84288
rect 3604 83200 3612 83264
rect 3676 83200 3692 83264
rect 3756 83200 3772 83264
rect 3836 83200 3852 83264
rect 3916 83200 3924 83264
rect 3604 82866 3924 83200
rect 3604 82630 3646 82866
rect 3882 82630 3924 82866
rect 3604 82176 3924 82630
rect 3604 82112 3612 82176
rect 3676 82112 3692 82176
rect 3756 82112 3772 82176
rect 3836 82112 3852 82176
rect 3916 82112 3924 82176
rect 3604 81088 3924 82112
rect 3604 81024 3612 81088
rect 3676 81024 3692 81088
rect 3756 81024 3772 81088
rect 3836 81024 3852 81088
rect 3916 81024 3924 81088
rect 3604 80000 3924 81024
rect 3604 79936 3612 80000
rect 3676 79936 3692 80000
rect 3756 79936 3772 80000
rect 3836 79936 3852 80000
rect 3916 79936 3924 80000
rect 3604 78912 3924 79936
rect 3604 78848 3612 78912
rect 3676 78848 3692 78912
rect 3756 78848 3772 78912
rect 3836 78848 3852 78912
rect 3916 78848 3924 78912
rect 3604 77824 3924 78848
rect 3604 77760 3612 77824
rect 3676 77760 3692 77824
rect 3756 77760 3772 77824
rect 3836 77760 3852 77824
rect 3916 77760 3924 77824
rect 3604 76736 3924 77760
rect 3604 76672 3612 76736
rect 3676 76672 3692 76736
rect 3756 76672 3772 76736
rect 3836 76672 3852 76736
rect 3916 76672 3924 76736
rect 3604 75648 3924 76672
rect 3604 75584 3612 75648
rect 3676 75584 3692 75648
rect 3756 75584 3772 75648
rect 3836 75584 3852 75648
rect 3916 75584 3924 75648
rect 3604 74560 3924 75584
rect 3604 74496 3612 74560
rect 3676 74496 3692 74560
rect 3756 74496 3772 74560
rect 3836 74496 3852 74560
rect 3916 74496 3924 74560
rect 3604 73472 3924 74496
rect 3604 73408 3612 73472
rect 3676 73408 3692 73472
rect 3756 73408 3772 73472
rect 3836 73408 3852 73472
rect 3916 73408 3924 73472
rect 3604 72384 3924 73408
rect 3604 72320 3612 72384
rect 3676 72320 3692 72384
rect 3756 72320 3772 72384
rect 3836 72320 3852 72384
rect 3916 72320 3924 72384
rect 3604 71296 3924 72320
rect 3604 71232 3612 71296
rect 3676 71232 3692 71296
rect 3756 71232 3772 71296
rect 3836 71232 3852 71296
rect 3916 71232 3924 71296
rect 3604 70208 3924 71232
rect 3604 70144 3612 70208
rect 3676 70144 3692 70208
rect 3756 70144 3772 70208
rect 3836 70144 3852 70208
rect 3916 70144 3924 70208
rect 3604 69120 3924 70144
rect 3604 69056 3612 69120
rect 3676 69056 3692 69120
rect 3756 69056 3772 69120
rect 3836 69056 3852 69120
rect 3916 69056 3924 69120
rect 3604 68032 3924 69056
rect 3604 67968 3612 68032
rect 3676 67968 3692 68032
rect 3756 67968 3772 68032
rect 3836 67968 3852 68032
rect 3916 67968 3924 68032
rect 3604 66944 3924 67968
rect 3604 66880 3612 66944
rect 3676 66880 3692 66944
rect 3756 66880 3772 66944
rect 3836 66880 3852 66944
rect 3916 66880 3924 66944
rect 3604 65856 3924 66880
rect 3604 65792 3612 65856
rect 3676 65792 3692 65856
rect 3756 65792 3772 65856
rect 3836 65792 3852 65856
rect 3916 65792 3924 65856
rect 3604 64768 3924 65792
rect 3604 64704 3612 64768
rect 3676 64704 3692 64768
rect 3756 64704 3772 64768
rect 3836 64704 3852 64768
rect 3916 64704 3924 64768
rect 3604 63680 3924 64704
rect 3604 63616 3612 63680
rect 3676 63616 3692 63680
rect 3756 63616 3772 63680
rect 3836 63616 3852 63680
rect 3916 63616 3924 63680
rect 3604 62592 3924 63616
rect 3604 62528 3612 62592
rect 3676 62528 3692 62592
rect 3756 62528 3772 62592
rect 3836 62528 3852 62592
rect 3916 62528 3924 62592
rect 3604 61504 3924 62528
rect 3604 61440 3612 61504
rect 3676 61440 3692 61504
rect 3756 61440 3772 61504
rect 3836 61440 3852 61504
rect 3916 61440 3924 61504
rect 3604 60416 3924 61440
rect 3604 60352 3612 60416
rect 3676 60352 3692 60416
rect 3756 60352 3772 60416
rect 3836 60352 3852 60416
rect 3916 60352 3924 60416
rect 3604 59328 3924 60352
rect 3604 59264 3612 59328
rect 3676 59264 3692 59328
rect 3756 59264 3772 59328
rect 3836 59264 3852 59328
rect 3916 59264 3924 59328
rect 3604 58240 3924 59264
rect 3604 58176 3612 58240
rect 3676 58176 3692 58240
rect 3756 58176 3772 58240
rect 3836 58176 3852 58240
rect 3916 58176 3924 58240
rect 3604 57152 3924 58176
rect 3604 57088 3612 57152
rect 3676 57088 3692 57152
rect 3756 57088 3772 57152
rect 3836 57088 3852 57152
rect 3916 57088 3924 57152
rect 3604 56064 3924 57088
rect 3604 56000 3612 56064
rect 3676 56000 3692 56064
rect 3756 56000 3772 56064
rect 3836 56000 3852 56064
rect 3916 56000 3924 56064
rect 3604 54976 3924 56000
rect 3604 54912 3612 54976
rect 3676 54912 3692 54976
rect 3756 54912 3772 54976
rect 3836 54912 3852 54976
rect 3916 54912 3924 54976
rect 3604 53888 3924 54912
rect 3604 53824 3612 53888
rect 3676 53824 3692 53888
rect 3756 53824 3772 53888
rect 3836 53824 3852 53888
rect 3916 53824 3924 53888
rect 3604 52800 3924 53824
rect 3604 52736 3612 52800
rect 3676 52736 3692 52800
rect 3756 52736 3772 52800
rect 3836 52736 3852 52800
rect 3916 52736 3924 52800
rect 3604 51712 3924 52736
rect 3604 51648 3612 51712
rect 3676 51648 3692 51712
rect 3756 51648 3772 51712
rect 3836 51648 3852 51712
rect 3916 51648 3924 51712
rect 3604 50624 3924 51648
rect 3604 50560 3612 50624
rect 3676 50560 3692 50624
rect 3756 50560 3772 50624
rect 3836 50560 3852 50624
rect 3916 50560 3924 50624
rect 3604 49536 3924 50560
rect 3604 49472 3612 49536
rect 3676 49472 3692 49536
rect 3756 49472 3772 49536
rect 3836 49472 3852 49536
rect 3916 49472 3924 49536
rect 3604 48448 3924 49472
rect 3604 48384 3612 48448
rect 3676 48384 3692 48448
rect 3756 48384 3772 48448
rect 3836 48384 3852 48448
rect 3916 48384 3924 48448
rect 3604 47360 3924 48384
rect 3604 47296 3612 47360
rect 3676 47296 3692 47360
rect 3756 47296 3772 47360
rect 3836 47296 3852 47360
rect 3916 47296 3924 47360
rect 3604 46272 3924 47296
rect 3604 46208 3612 46272
rect 3676 46208 3692 46272
rect 3756 46208 3772 46272
rect 3836 46208 3852 46272
rect 3916 46208 3924 46272
rect 3604 45184 3924 46208
rect 3604 45120 3612 45184
rect 3676 45120 3692 45184
rect 3756 45120 3772 45184
rect 3836 45120 3852 45184
rect 3916 45120 3924 45184
rect 3604 44096 3924 45120
rect 3604 44032 3612 44096
rect 3676 44032 3692 44096
rect 3756 44032 3772 44096
rect 3836 44032 3852 44096
rect 3916 44032 3924 44096
rect 3604 43008 3924 44032
rect 3604 42944 3612 43008
rect 3676 42944 3692 43008
rect 3756 42944 3772 43008
rect 3836 42944 3852 43008
rect 3916 42944 3924 43008
rect 3604 41920 3924 42944
rect 3604 41856 3612 41920
rect 3676 41856 3692 41920
rect 3756 41856 3772 41920
rect 3836 41856 3852 41920
rect 3916 41856 3924 41920
rect 3604 40832 3924 41856
rect 3604 40768 3612 40832
rect 3676 40768 3692 40832
rect 3756 40768 3772 40832
rect 3836 40768 3852 40832
rect 3916 40768 3924 40832
rect 3604 39744 3924 40768
rect 3604 39680 3612 39744
rect 3676 39680 3692 39744
rect 3756 39680 3772 39744
rect 3836 39680 3852 39744
rect 3916 39680 3924 39744
rect 3604 38656 3924 39680
rect 3604 38592 3612 38656
rect 3676 38592 3692 38656
rect 3756 38592 3772 38656
rect 3836 38592 3852 38656
rect 3916 38592 3924 38656
rect 3604 37568 3924 38592
rect 3604 37504 3612 37568
rect 3676 37504 3692 37568
rect 3756 37504 3772 37568
rect 3836 37504 3852 37568
rect 3916 37504 3924 37568
rect 3604 36480 3924 37504
rect 3604 36416 3612 36480
rect 3676 36416 3692 36480
rect 3756 36416 3772 36480
rect 3836 36416 3852 36480
rect 3916 36416 3924 36480
rect 3604 35392 3924 36416
rect 3604 35328 3612 35392
rect 3676 35328 3692 35392
rect 3756 35328 3772 35392
rect 3836 35328 3852 35392
rect 3916 35328 3924 35392
rect 3604 34304 3924 35328
rect 3604 34240 3612 34304
rect 3676 34240 3692 34304
rect 3756 34240 3772 34304
rect 3836 34240 3852 34304
rect 3916 34240 3924 34304
rect 3604 33216 3924 34240
rect 3604 33152 3612 33216
rect 3676 33152 3692 33216
rect 3756 33152 3772 33216
rect 3836 33152 3852 33216
rect 3916 33152 3924 33216
rect 3604 32128 3924 33152
rect 3604 32064 3612 32128
rect 3676 32064 3692 32128
rect 3756 32064 3772 32128
rect 3836 32064 3852 32128
rect 3916 32064 3924 32128
rect 3604 31040 3924 32064
rect 3604 30976 3612 31040
rect 3676 30976 3692 31040
rect 3756 30976 3772 31040
rect 3836 30976 3852 31040
rect 3916 30976 3924 31040
rect 3604 29952 3924 30976
rect 3604 29888 3612 29952
rect 3676 29888 3692 29952
rect 3756 29888 3772 29952
rect 3836 29888 3852 29952
rect 3916 29888 3924 29952
rect 3604 28864 3924 29888
rect 3604 28800 3612 28864
rect 3676 28800 3692 28864
rect 3756 28800 3772 28864
rect 3836 28800 3852 28864
rect 3916 28800 3924 28864
rect 3604 27776 3924 28800
rect 3604 27712 3612 27776
rect 3676 27712 3692 27776
rect 3756 27712 3772 27776
rect 3836 27712 3852 27776
rect 3916 27712 3924 27776
rect 3604 26688 3924 27712
rect 3604 26624 3612 26688
rect 3676 26624 3692 26688
rect 3756 26624 3772 26688
rect 3836 26624 3852 26688
rect 3916 26624 3924 26688
rect 3604 25600 3924 26624
rect 3604 25536 3612 25600
rect 3676 25536 3692 25600
rect 3756 25536 3772 25600
rect 3836 25536 3852 25600
rect 3916 25536 3924 25600
rect 3604 24512 3924 25536
rect 3604 24448 3612 24512
rect 3676 24448 3692 24512
rect 3756 24448 3772 24512
rect 3836 24448 3852 24512
rect 3916 24448 3924 24512
rect 3604 23424 3924 24448
rect 3604 23360 3612 23424
rect 3676 23360 3692 23424
rect 3756 23360 3772 23424
rect 3836 23360 3852 23424
rect 3916 23360 3924 23424
rect 3604 22336 3924 23360
rect 3604 22272 3612 22336
rect 3676 22272 3692 22336
rect 3756 22272 3772 22336
rect 3836 22272 3852 22336
rect 3916 22272 3924 22336
rect 3604 21248 3924 22272
rect 3604 21184 3612 21248
rect 3676 21184 3692 21248
rect 3756 21184 3772 21248
rect 3836 21184 3852 21248
rect 3916 21184 3924 21248
rect 3604 20160 3924 21184
rect 3604 20096 3612 20160
rect 3676 20096 3692 20160
rect 3756 20096 3772 20160
rect 3836 20096 3852 20160
rect 3916 20096 3924 20160
rect 3604 19072 3924 20096
rect 3604 19008 3612 19072
rect 3676 19008 3692 19072
rect 3756 19008 3772 19072
rect 3836 19008 3852 19072
rect 3916 19008 3924 19072
rect 3604 17984 3924 19008
rect 3604 17920 3612 17984
rect 3676 17920 3692 17984
rect 3756 17920 3772 17984
rect 3836 17920 3852 17984
rect 3916 17920 3924 17984
rect 3604 16896 3924 17920
rect 3604 16832 3612 16896
rect 3676 16832 3692 16896
rect 3756 16832 3772 16896
rect 3836 16832 3852 16896
rect 3916 16832 3924 16896
rect 3604 15808 3924 16832
rect 3604 15744 3612 15808
rect 3676 15744 3692 15808
rect 3756 15744 3772 15808
rect 3836 15744 3852 15808
rect 3916 15744 3924 15808
rect 3604 14720 3924 15744
rect 3604 14656 3612 14720
rect 3676 14656 3692 14720
rect 3756 14656 3772 14720
rect 3836 14656 3852 14720
rect 3916 14656 3924 14720
rect 3604 13632 3924 14656
rect 3604 13568 3612 13632
rect 3676 13568 3692 13632
rect 3756 13568 3772 13632
rect 3836 13568 3852 13632
rect 3916 13568 3924 13632
rect 3604 12544 3924 13568
rect 3604 12480 3612 12544
rect 3676 12480 3692 12544
rect 3756 12480 3772 12544
rect 3836 12480 3852 12544
rect 3916 12480 3924 12544
rect 3604 11456 3924 12480
rect 3604 11392 3612 11456
rect 3676 11392 3692 11456
rect 3756 11392 3772 11456
rect 3836 11392 3852 11456
rect 3916 11392 3924 11456
rect 3604 10368 3924 11392
rect 3604 10304 3612 10368
rect 3676 10304 3692 10368
rect 3756 10304 3772 10368
rect 3836 10304 3852 10368
rect 3916 10304 3924 10368
rect 3604 9280 3924 10304
rect 3604 9216 3612 9280
rect 3676 9216 3692 9280
rect 3756 9216 3772 9280
rect 3836 9216 3852 9280
rect 3916 9216 3924 9280
rect 3604 8192 3924 9216
rect 3604 8128 3612 8192
rect 3676 8128 3692 8192
rect 3756 8128 3772 8192
rect 3836 8128 3852 8192
rect 3916 8128 3924 8192
rect 3604 7104 3924 8128
rect 3604 7040 3612 7104
rect 3676 7040 3692 7104
rect 3756 7040 3772 7104
rect 3836 7040 3852 7104
rect 3916 7040 3924 7104
rect 3604 6866 3924 7040
rect 3604 6630 3646 6866
rect 3882 6630 3924 6866
rect 3604 6016 3924 6630
rect 3604 5952 3612 6016
rect 3676 5952 3692 6016
rect 3756 5952 3772 6016
rect 3836 5952 3852 6016
rect 3916 5952 3924 6016
rect 3604 4928 3924 5952
rect 3604 4864 3612 4928
rect 3676 4864 3692 4928
rect 3756 4864 3772 4928
rect 3836 4864 3852 4928
rect 3916 4864 3924 4928
rect 3604 3840 3924 4864
rect 3604 3776 3612 3840
rect 3676 3776 3692 3840
rect 3756 3776 3772 3840
rect 3836 3776 3852 3840
rect 3916 3776 3924 3840
rect 3604 2752 3924 3776
rect 3604 2688 3612 2752
rect 3676 2688 3692 2752
rect 3756 2688 3772 2752
rect 3836 2688 3852 2752
rect 3916 2688 3924 2752
rect 3604 1664 3924 2688
rect 3604 1600 3612 1664
rect 3676 1600 3692 1664
rect 3756 1600 3772 1664
rect 3836 1600 3852 1664
rect 3916 1600 3924 1664
rect 3604 -154 3924 1600
rect 3604 -390 3646 -154
rect 3882 -390 3924 -154
rect 3604 -1092 3924 -390
rect 4544 88634 4864 88676
rect 4544 88398 4586 88634
rect 4822 88398 4864 88634
rect 4544 85984 4864 88398
rect 4544 85920 4552 85984
rect 4616 85920 4632 85984
rect 4696 85920 4712 85984
rect 4776 85920 4792 85984
rect 4856 85920 4864 85984
rect 4544 84896 4864 85920
rect 4544 84832 4552 84896
rect 4616 84832 4632 84896
rect 4696 84832 4712 84896
rect 4776 84832 4792 84896
rect 4856 84832 4864 84896
rect 4544 83808 4864 84832
rect 4544 83744 4552 83808
rect 4616 83744 4632 83808
rect 4696 83744 4712 83808
rect 4776 83744 4792 83808
rect 4856 83744 4864 83808
rect 4544 82720 4864 83744
rect 4544 82656 4552 82720
rect 4616 82656 4632 82720
rect 4696 82656 4712 82720
rect 4776 82656 4792 82720
rect 4856 82656 4864 82720
rect 4544 82206 4864 82656
rect 4544 81970 4586 82206
rect 4822 81970 4864 82206
rect 4544 81632 4864 81970
rect 4544 81568 4552 81632
rect 4616 81568 4632 81632
rect 4696 81568 4712 81632
rect 4776 81568 4792 81632
rect 4856 81568 4864 81632
rect 4544 80544 4864 81568
rect 4544 80480 4552 80544
rect 4616 80480 4632 80544
rect 4696 80480 4712 80544
rect 4776 80480 4792 80544
rect 4856 80480 4864 80544
rect 4544 79456 4864 80480
rect 4544 79392 4552 79456
rect 4616 79392 4632 79456
rect 4696 79392 4712 79456
rect 4776 79392 4792 79456
rect 4856 79392 4864 79456
rect 4544 78368 4864 79392
rect 4544 78304 4552 78368
rect 4616 78304 4632 78368
rect 4696 78304 4712 78368
rect 4776 78304 4792 78368
rect 4856 78304 4864 78368
rect 4544 77280 4864 78304
rect 4544 77216 4552 77280
rect 4616 77216 4632 77280
rect 4696 77216 4712 77280
rect 4776 77216 4792 77280
rect 4856 77216 4864 77280
rect 4544 76192 4864 77216
rect 4544 76128 4552 76192
rect 4616 76128 4632 76192
rect 4696 76128 4712 76192
rect 4776 76128 4792 76192
rect 4856 76128 4864 76192
rect 4544 75104 4864 76128
rect 4544 75040 4552 75104
rect 4616 75040 4632 75104
rect 4696 75040 4712 75104
rect 4776 75040 4792 75104
rect 4856 75040 4864 75104
rect 4544 74016 4864 75040
rect 4544 73952 4552 74016
rect 4616 73952 4632 74016
rect 4696 73952 4712 74016
rect 4776 73952 4792 74016
rect 4856 73952 4864 74016
rect 4544 72928 4864 73952
rect 4544 72864 4552 72928
rect 4616 72864 4632 72928
rect 4696 72864 4712 72928
rect 4776 72864 4792 72928
rect 4856 72864 4864 72928
rect 4544 71840 4864 72864
rect 4544 71776 4552 71840
rect 4616 71776 4632 71840
rect 4696 71776 4712 71840
rect 4776 71776 4792 71840
rect 4856 71776 4864 71840
rect 4544 70752 4864 71776
rect 4544 70688 4552 70752
rect 4616 70688 4632 70752
rect 4696 70688 4712 70752
rect 4776 70688 4792 70752
rect 4856 70688 4864 70752
rect 4544 69664 4864 70688
rect 4544 69600 4552 69664
rect 4616 69600 4632 69664
rect 4696 69600 4712 69664
rect 4776 69600 4792 69664
rect 4856 69600 4864 69664
rect 4544 68576 4864 69600
rect 4544 68512 4552 68576
rect 4616 68512 4632 68576
rect 4696 68512 4712 68576
rect 4776 68512 4792 68576
rect 4856 68512 4864 68576
rect 4544 67488 4864 68512
rect 4544 67424 4552 67488
rect 4616 67424 4632 67488
rect 4696 67424 4712 67488
rect 4776 67424 4792 67488
rect 4856 67424 4864 67488
rect 4544 66400 4864 67424
rect 4544 66336 4552 66400
rect 4616 66336 4632 66400
rect 4696 66336 4712 66400
rect 4776 66336 4792 66400
rect 4856 66336 4864 66400
rect 4544 65312 4864 66336
rect 4544 65248 4552 65312
rect 4616 65248 4632 65312
rect 4696 65248 4712 65312
rect 4776 65248 4792 65312
rect 4856 65248 4864 65312
rect 4544 64224 4864 65248
rect 4544 64160 4552 64224
rect 4616 64160 4632 64224
rect 4696 64160 4712 64224
rect 4776 64160 4792 64224
rect 4856 64160 4864 64224
rect 4544 63136 4864 64160
rect 4544 63072 4552 63136
rect 4616 63072 4632 63136
rect 4696 63072 4712 63136
rect 4776 63072 4792 63136
rect 4856 63072 4864 63136
rect 4544 62048 4864 63072
rect 4544 61984 4552 62048
rect 4616 61984 4632 62048
rect 4696 61984 4712 62048
rect 4776 61984 4792 62048
rect 4856 61984 4864 62048
rect 4544 60960 4864 61984
rect 4544 60896 4552 60960
rect 4616 60896 4632 60960
rect 4696 60896 4712 60960
rect 4776 60896 4792 60960
rect 4856 60896 4864 60960
rect 4544 59872 4864 60896
rect 4544 59808 4552 59872
rect 4616 59808 4632 59872
rect 4696 59808 4712 59872
rect 4776 59808 4792 59872
rect 4856 59808 4864 59872
rect 4544 58784 4864 59808
rect 4544 58720 4552 58784
rect 4616 58720 4632 58784
rect 4696 58720 4712 58784
rect 4776 58720 4792 58784
rect 4856 58720 4864 58784
rect 4544 57696 4864 58720
rect 4544 57632 4552 57696
rect 4616 57632 4632 57696
rect 4696 57632 4712 57696
rect 4776 57632 4792 57696
rect 4856 57632 4864 57696
rect 4544 56608 4864 57632
rect 4544 56544 4552 56608
rect 4616 56544 4632 56608
rect 4696 56544 4712 56608
rect 4776 56544 4792 56608
rect 4856 56544 4864 56608
rect 4544 55520 4864 56544
rect 4544 55456 4552 55520
rect 4616 55456 4632 55520
rect 4696 55456 4712 55520
rect 4776 55456 4792 55520
rect 4856 55456 4864 55520
rect 4544 54432 4864 55456
rect 4544 54368 4552 54432
rect 4616 54368 4632 54432
rect 4696 54368 4712 54432
rect 4776 54368 4792 54432
rect 4856 54368 4864 54432
rect 4544 53344 4864 54368
rect 4544 53280 4552 53344
rect 4616 53280 4632 53344
rect 4696 53280 4712 53344
rect 4776 53280 4792 53344
rect 4856 53280 4864 53344
rect 4544 52256 4864 53280
rect 4544 52192 4552 52256
rect 4616 52192 4632 52256
rect 4696 52192 4712 52256
rect 4776 52192 4792 52256
rect 4856 52192 4864 52256
rect 4544 51168 4864 52192
rect 4544 51104 4552 51168
rect 4616 51104 4632 51168
rect 4696 51104 4712 51168
rect 4776 51104 4792 51168
rect 4856 51104 4864 51168
rect 4544 50080 4864 51104
rect 4544 50016 4552 50080
rect 4616 50016 4632 50080
rect 4696 50016 4712 50080
rect 4776 50016 4792 50080
rect 4856 50016 4864 50080
rect 4544 48992 4864 50016
rect 4544 48928 4552 48992
rect 4616 48928 4632 48992
rect 4696 48928 4712 48992
rect 4776 48928 4792 48992
rect 4856 48928 4864 48992
rect 4544 47904 4864 48928
rect 4544 47840 4552 47904
rect 4616 47840 4632 47904
rect 4696 47840 4712 47904
rect 4776 47840 4792 47904
rect 4856 47840 4864 47904
rect 4544 46816 4864 47840
rect 4544 46752 4552 46816
rect 4616 46752 4632 46816
rect 4696 46752 4712 46816
rect 4776 46752 4792 46816
rect 4856 46752 4864 46816
rect 4544 45728 4864 46752
rect 4544 45664 4552 45728
rect 4616 45664 4632 45728
rect 4696 45664 4712 45728
rect 4776 45664 4792 45728
rect 4856 45664 4864 45728
rect 4544 44640 4864 45664
rect 4544 44576 4552 44640
rect 4616 44576 4632 44640
rect 4696 44576 4712 44640
rect 4776 44576 4792 44640
rect 4856 44576 4864 44640
rect 4544 43552 4864 44576
rect 4544 43488 4552 43552
rect 4616 43488 4632 43552
rect 4696 43488 4712 43552
rect 4776 43488 4792 43552
rect 4856 43488 4864 43552
rect 4544 42464 4864 43488
rect 4544 42400 4552 42464
rect 4616 42400 4632 42464
rect 4696 42400 4712 42464
rect 4776 42400 4792 42464
rect 4856 42400 4864 42464
rect 4544 41376 4864 42400
rect 4544 41312 4552 41376
rect 4616 41312 4632 41376
rect 4696 41312 4712 41376
rect 4776 41312 4792 41376
rect 4856 41312 4864 41376
rect 4544 40288 4864 41312
rect 4544 40224 4552 40288
rect 4616 40224 4632 40288
rect 4696 40224 4712 40288
rect 4776 40224 4792 40288
rect 4856 40224 4864 40288
rect 4544 39200 4864 40224
rect 4544 39136 4552 39200
rect 4616 39136 4632 39200
rect 4696 39136 4712 39200
rect 4776 39136 4792 39200
rect 4856 39136 4864 39200
rect 4544 38112 4864 39136
rect 4544 38048 4552 38112
rect 4616 38048 4632 38112
rect 4696 38048 4712 38112
rect 4776 38048 4792 38112
rect 4856 38048 4864 38112
rect 4544 37024 4864 38048
rect 4544 36960 4552 37024
rect 4616 36960 4632 37024
rect 4696 36960 4712 37024
rect 4776 36960 4792 37024
rect 4856 36960 4864 37024
rect 4544 35936 4864 36960
rect 4544 35872 4552 35936
rect 4616 35872 4632 35936
rect 4696 35872 4712 35936
rect 4776 35872 4792 35936
rect 4856 35872 4864 35936
rect 4544 34848 4864 35872
rect 4544 34784 4552 34848
rect 4616 34784 4632 34848
rect 4696 34784 4712 34848
rect 4776 34784 4792 34848
rect 4856 34784 4864 34848
rect 4544 33760 4864 34784
rect 4544 33696 4552 33760
rect 4616 33696 4632 33760
rect 4696 33696 4712 33760
rect 4776 33696 4792 33760
rect 4856 33696 4864 33760
rect 4544 32672 4864 33696
rect 4544 32608 4552 32672
rect 4616 32608 4632 32672
rect 4696 32608 4712 32672
rect 4776 32608 4792 32672
rect 4856 32608 4864 32672
rect 4544 31584 4864 32608
rect 4544 31520 4552 31584
rect 4616 31520 4632 31584
rect 4696 31520 4712 31584
rect 4776 31520 4792 31584
rect 4856 31520 4864 31584
rect 4544 30496 4864 31520
rect 4544 30432 4552 30496
rect 4616 30432 4632 30496
rect 4696 30432 4712 30496
rect 4776 30432 4792 30496
rect 4856 30432 4864 30496
rect 4544 29408 4864 30432
rect 4544 29344 4552 29408
rect 4616 29344 4632 29408
rect 4696 29344 4712 29408
rect 4776 29344 4792 29408
rect 4856 29344 4864 29408
rect 4544 28320 4864 29344
rect 4544 28256 4552 28320
rect 4616 28256 4632 28320
rect 4696 28256 4712 28320
rect 4776 28256 4792 28320
rect 4856 28256 4864 28320
rect 4544 27232 4864 28256
rect 4544 27168 4552 27232
rect 4616 27168 4632 27232
rect 4696 27168 4712 27232
rect 4776 27168 4792 27232
rect 4856 27168 4864 27232
rect 4544 26144 4864 27168
rect 4544 26080 4552 26144
rect 4616 26080 4632 26144
rect 4696 26080 4712 26144
rect 4776 26080 4792 26144
rect 4856 26080 4864 26144
rect 4544 25056 4864 26080
rect 4544 24992 4552 25056
rect 4616 24992 4632 25056
rect 4696 24992 4712 25056
rect 4776 24992 4792 25056
rect 4856 24992 4864 25056
rect 4544 23968 4864 24992
rect 4544 23904 4552 23968
rect 4616 23904 4632 23968
rect 4696 23904 4712 23968
rect 4776 23904 4792 23968
rect 4856 23904 4864 23968
rect 4544 22880 4864 23904
rect 4544 22816 4552 22880
rect 4616 22816 4632 22880
rect 4696 22816 4712 22880
rect 4776 22816 4792 22880
rect 4856 22816 4864 22880
rect 4544 21792 4864 22816
rect 4544 21728 4552 21792
rect 4616 21728 4632 21792
rect 4696 21728 4712 21792
rect 4776 21728 4792 21792
rect 4856 21728 4864 21792
rect 4544 20704 4864 21728
rect 4544 20640 4552 20704
rect 4616 20640 4632 20704
rect 4696 20640 4712 20704
rect 4776 20640 4792 20704
rect 4856 20640 4864 20704
rect 4544 19616 4864 20640
rect 4544 19552 4552 19616
rect 4616 19552 4632 19616
rect 4696 19552 4712 19616
rect 4776 19552 4792 19616
rect 4856 19552 4864 19616
rect 4544 18528 4864 19552
rect 4544 18464 4552 18528
rect 4616 18464 4632 18528
rect 4696 18464 4712 18528
rect 4776 18464 4792 18528
rect 4856 18464 4864 18528
rect 4544 17440 4864 18464
rect 4544 17376 4552 17440
rect 4616 17376 4632 17440
rect 4696 17376 4712 17440
rect 4776 17376 4792 17440
rect 4856 17376 4864 17440
rect 4544 16352 4864 17376
rect 4544 16288 4552 16352
rect 4616 16288 4632 16352
rect 4696 16288 4712 16352
rect 4776 16288 4792 16352
rect 4856 16288 4864 16352
rect 4544 15264 4864 16288
rect 4544 15200 4552 15264
rect 4616 15200 4632 15264
rect 4696 15200 4712 15264
rect 4776 15200 4792 15264
rect 4856 15200 4864 15264
rect 4544 14176 4864 15200
rect 4544 14112 4552 14176
rect 4616 14112 4632 14176
rect 4696 14112 4712 14176
rect 4776 14112 4792 14176
rect 4856 14112 4864 14176
rect 4544 13088 4864 14112
rect 4544 13024 4552 13088
rect 4616 13024 4632 13088
rect 4696 13024 4712 13088
rect 4776 13024 4792 13088
rect 4856 13024 4864 13088
rect 4544 12000 4864 13024
rect 4544 11936 4552 12000
rect 4616 11936 4632 12000
rect 4696 11936 4712 12000
rect 4776 11936 4792 12000
rect 4856 11936 4864 12000
rect 4544 10912 4864 11936
rect 4544 10848 4552 10912
rect 4616 10848 4632 10912
rect 4696 10848 4712 10912
rect 4776 10848 4792 10912
rect 4856 10848 4864 10912
rect 4544 9824 4864 10848
rect 4544 9760 4552 9824
rect 4616 9760 4632 9824
rect 4696 9760 4712 9824
rect 4776 9760 4792 9824
rect 4856 9760 4864 9824
rect 4544 8736 4864 9760
rect 4544 8672 4552 8736
rect 4616 8672 4632 8736
rect 4696 8672 4712 8736
rect 4776 8672 4792 8736
rect 4856 8672 4864 8736
rect 4544 7648 4864 8672
rect 4544 7584 4552 7648
rect 4616 7584 4632 7648
rect 4696 7584 4712 7648
rect 4776 7584 4792 7648
rect 4856 7584 4864 7648
rect 4544 6560 4864 7584
rect 4544 6496 4552 6560
rect 4616 6496 4632 6560
rect 4696 6496 4712 6560
rect 4776 6496 4792 6560
rect 4856 6496 4864 6560
rect 4544 6206 4864 6496
rect 4544 5970 4586 6206
rect 4822 5970 4864 6206
rect 4544 5472 4864 5970
rect 4544 5408 4552 5472
rect 4616 5408 4632 5472
rect 4696 5408 4712 5472
rect 4776 5408 4792 5472
rect 4856 5408 4864 5472
rect 4544 4384 4864 5408
rect 4544 4320 4552 4384
rect 4616 4320 4632 4384
rect 4696 4320 4712 4384
rect 4776 4320 4792 4384
rect 4856 4320 4864 4384
rect 4544 3296 4864 4320
rect 4544 3232 4552 3296
rect 4616 3232 4632 3296
rect 4696 3232 4712 3296
rect 4776 3232 4792 3296
rect 4856 3232 4864 3296
rect 4544 2208 4864 3232
rect 4544 2144 4552 2208
rect 4616 2144 4632 2208
rect 4696 2144 4712 2208
rect 4776 2144 4792 2208
rect 4856 2144 4864 2208
rect 4544 1120 4864 2144
rect 4544 1056 4552 1120
rect 4616 1056 4632 1120
rect 4696 1056 4712 1120
rect 4776 1056 4792 1120
rect 4856 1056 4864 1120
rect 4544 -814 4864 1056
rect 4544 -1050 4586 -814
rect 4822 -1050 4864 -814
rect 4544 -1092 4864 -1050
rect 5204 87974 5524 88676
rect 5204 87738 5246 87974
rect 5482 87738 5524 87974
rect 5204 86528 5524 87738
rect 5204 86464 5212 86528
rect 5276 86464 5292 86528
rect 5356 86464 5372 86528
rect 5436 86464 5452 86528
rect 5516 86464 5524 86528
rect 5204 85440 5524 86464
rect 5204 85376 5212 85440
rect 5276 85376 5292 85440
rect 5356 85376 5372 85440
rect 5436 85376 5452 85440
rect 5516 85376 5524 85440
rect 5204 84352 5524 85376
rect 5204 84288 5212 84352
rect 5276 84288 5292 84352
rect 5356 84288 5372 84352
rect 5436 84288 5452 84352
rect 5516 84288 5524 84352
rect 5204 83264 5524 84288
rect 5204 83200 5212 83264
rect 5276 83200 5292 83264
rect 5356 83200 5372 83264
rect 5436 83200 5452 83264
rect 5516 83200 5524 83264
rect 5204 82866 5524 83200
rect 5204 82630 5246 82866
rect 5482 82630 5524 82866
rect 5204 82176 5524 82630
rect 5204 82112 5212 82176
rect 5276 82112 5292 82176
rect 5356 82112 5372 82176
rect 5436 82112 5452 82176
rect 5516 82112 5524 82176
rect 5204 81088 5524 82112
rect 5204 81024 5212 81088
rect 5276 81024 5292 81088
rect 5356 81024 5372 81088
rect 5436 81024 5452 81088
rect 5516 81024 5524 81088
rect 5204 80000 5524 81024
rect 5204 79936 5212 80000
rect 5276 79936 5292 80000
rect 5356 79936 5372 80000
rect 5436 79936 5452 80000
rect 5516 79936 5524 80000
rect 5204 78912 5524 79936
rect 5204 78848 5212 78912
rect 5276 78848 5292 78912
rect 5356 78848 5372 78912
rect 5436 78848 5452 78912
rect 5516 78848 5524 78912
rect 5204 77824 5524 78848
rect 5204 77760 5212 77824
rect 5276 77760 5292 77824
rect 5356 77760 5372 77824
rect 5436 77760 5452 77824
rect 5516 77760 5524 77824
rect 5204 76736 5524 77760
rect 5204 76672 5212 76736
rect 5276 76672 5292 76736
rect 5356 76672 5372 76736
rect 5436 76672 5452 76736
rect 5516 76672 5524 76736
rect 5204 75648 5524 76672
rect 5204 75584 5212 75648
rect 5276 75584 5292 75648
rect 5356 75584 5372 75648
rect 5436 75584 5452 75648
rect 5516 75584 5524 75648
rect 5204 74560 5524 75584
rect 5204 74496 5212 74560
rect 5276 74496 5292 74560
rect 5356 74496 5372 74560
rect 5436 74496 5452 74560
rect 5516 74496 5524 74560
rect 5204 73472 5524 74496
rect 5204 73408 5212 73472
rect 5276 73408 5292 73472
rect 5356 73408 5372 73472
rect 5436 73408 5452 73472
rect 5516 73408 5524 73472
rect 5204 72384 5524 73408
rect 5204 72320 5212 72384
rect 5276 72320 5292 72384
rect 5356 72320 5372 72384
rect 5436 72320 5452 72384
rect 5516 72320 5524 72384
rect 5204 71296 5524 72320
rect 5204 71232 5212 71296
rect 5276 71232 5292 71296
rect 5356 71232 5372 71296
rect 5436 71232 5452 71296
rect 5516 71232 5524 71296
rect 5204 70208 5524 71232
rect 5204 70144 5212 70208
rect 5276 70144 5292 70208
rect 5356 70144 5372 70208
rect 5436 70144 5452 70208
rect 5516 70144 5524 70208
rect 5204 69120 5524 70144
rect 5204 69056 5212 69120
rect 5276 69056 5292 69120
rect 5356 69056 5372 69120
rect 5436 69056 5452 69120
rect 5516 69056 5524 69120
rect 5204 68032 5524 69056
rect 5204 67968 5212 68032
rect 5276 67968 5292 68032
rect 5356 67968 5372 68032
rect 5436 67968 5452 68032
rect 5516 67968 5524 68032
rect 5204 66944 5524 67968
rect 5204 66880 5212 66944
rect 5276 66880 5292 66944
rect 5356 66880 5372 66944
rect 5436 66880 5452 66944
rect 5516 66880 5524 66944
rect 5204 65856 5524 66880
rect 5204 65792 5212 65856
rect 5276 65792 5292 65856
rect 5356 65792 5372 65856
rect 5436 65792 5452 65856
rect 5516 65792 5524 65856
rect 5204 64768 5524 65792
rect 5204 64704 5212 64768
rect 5276 64704 5292 64768
rect 5356 64704 5372 64768
rect 5436 64704 5452 64768
rect 5516 64704 5524 64768
rect 5204 63680 5524 64704
rect 5204 63616 5212 63680
rect 5276 63616 5292 63680
rect 5356 63616 5372 63680
rect 5436 63616 5452 63680
rect 5516 63616 5524 63680
rect 5204 62592 5524 63616
rect 5204 62528 5212 62592
rect 5276 62528 5292 62592
rect 5356 62528 5372 62592
rect 5436 62528 5452 62592
rect 5516 62528 5524 62592
rect 5204 61504 5524 62528
rect 5204 61440 5212 61504
rect 5276 61440 5292 61504
rect 5356 61440 5372 61504
rect 5436 61440 5452 61504
rect 5516 61440 5524 61504
rect 5204 60416 5524 61440
rect 5204 60352 5212 60416
rect 5276 60352 5292 60416
rect 5356 60352 5372 60416
rect 5436 60352 5452 60416
rect 5516 60352 5524 60416
rect 5204 59328 5524 60352
rect 5204 59264 5212 59328
rect 5276 59264 5292 59328
rect 5356 59264 5372 59328
rect 5436 59264 5452 59328
rect 5516 59264 5524 59328
rect 5204 58240 5524 59264
rect 5204 58176 5212 58240
rect 5276 58176 5292 58240
rect 5356 58176 5372 58240
rect 5436 58176 5452 58240
rect 5516 58176 5524 58240
rect 5204 57152 5524 58176
rect 5204 57088 5212 57152
rect 5276 57088 5292 57152
rect 5356 57088 5372 57152
rect 5436 57088 5452 57152
rect 5516 57088 5524 57152
rect 5204 56064 5524 57088
rect 5204 56000 5212 56064
rect 5276 56000 5292 56064
rect 5356 56000 5372 56064
rect 5436 56000 5452 56064
rect 5516 56000 5524 56064
rect 5204 54976 5524 56000
rect 5204 54912 5212 54976
rect 5276 54912 5292 54976
rect 5356 54912 5372 54976
rect 5436 54912 5452 54976
rect 5516 54912 5524 54976
rect 5204 53888 5524 54912
rect 5204 53824 5212 53888
rect 5276 53824 5292 53888
rect 5356 53824 5372 53888
rect 5436 53824 5452 53888
rect 5516 53824 5524 53888
rect 5204 52800 5524 53824
rect 5204 52736 5212 52800
rect 5276 52736 5292 52800
rect 5356 52736 5372 52800
rect 5436 52736 5452 52800
rect 5516 52736 5524 52800
rect 5204 51712 5524 52736
rect 5204 51648 5212 51712
rect 5276 51648 5292 51712
rect 5356 51648 5372 51712
rect 5436 51648 5452 51712
rect 5516 51648 5524 51712
rect 5204 50624 5524 51648
rect 5204 50560 5212 50624
rect 5276 50560 5292 50624
rect 5356 50560 5372 50624
rect 5436 50560 5452 50624
rect 5516 50560 5524 50624
rect 5204 49536 5524 50560
rect 5204 49472 5212 49536
rect 5276 49472 5292 49536
rect 5356 49472 5372 49536
rect 5436 49472 5452 49536
rect 5516 49472 5524 49536
rect 5204 48448 5524 49472
rect 5204 48384 5212 48448
rect 5276 48384 5292 48448
rect 5356 48384 5372 48448
rect 5436 48384 5452 48448
rect 5516 48384 5524 48448
rect 5204 47360 5524 48384
rect 5204 47296 5212 47360
rect 5276 47296 5292 47360
rect 5356 47296 5372 47360
rect 5436 47296 5452 47360
rect 5516 47296 5524 47360
rect 5204 46272 5524 47296
rect 5204 46208 5212 46272
rect 5276 46208 5292 46272
rect 5356 46208 5372 46272
rect 5436 46208 5452 46272
rect 5516 46208 5524 46272
rect 5204 45184 5524 46208
rect 5204 45120 5212 45184
rect 5276 45120 5292 45184
rect 5356 45120 5372 45184
rect 5436 45120 5452 45184
rect 5516 45120 5524 45184
rect 5204 44096 5524 45120
rect 5204 44032 5212 44096
rect 5276 44032 5292 44096
rect 5356 44032 5372 44096
rect 5436 44032 5452 44096
rect 5516 44032 5524 44096
rect 5204 43008 5524 44032
rect 5204 42944 5212 43008
rect 5276 42944 5292 43008
rect 5356 42944 5372 43008
rect 5436 42944 5452 43008
rect 5516 42944 5524 43008
rect 5204 41920 5524 42944
rect 5204 41856 5212 41920
rect 5276 41856 5292 41920
rect 5356 41856 5372 41920
rect 5436 41856 5452 41920
rect 5516 41856 5524 41920
rect 5204 40832 5524 41856
rect 5204 40768 5212 40832
rect 5276 40768 5292 40832
rect 5356 40768 5372 40832
rect 5436 40768 5452 40832
rect 5516 40768 5524 40832
rect 5204 39744 5524 40768
rect 5204 39680 5212 39744
rect 5276 39680 5292 39744
rect 5356 39680 5372 39744
rect 5436 39680 5452 39744
rect 5516 39680 5524 39744
rect 5204 38656 5524 39680
rect 5204 38592 5212 38656
rect 5276 38592 5292 38656
rect 5356 38592 5372 38656
rect 5436 38592 5452 38656
rect 5516 38592 5524 38656
rect 5204 37568 5524 38592
rect 5204 37504 5212 37568
rect 5276 37504 5292 37568
rect 5356 37504 5372 37568
rect 5436 37504 5452 37568
rect 5516 37504 5524 37568
rect 5204 36480 5524 37504
rect 5204 36416 5212 36480
rect 5276 36416 5292 36480
rect 5356 36416 5372 36480
rect 5436 36416 5452 36480
rect 5516 36416 5524 36480
rect 5204 35392 5524 36416
rect 5204 35328 5212 35392
rect 5276 35328 5292 35392
rect 5356 35328 5372 35392
rect 5436 35328 5452 35392
rect 5516 35328 5524 35392
rect 5204 34304 5524 35328
rect 5204 34240 5212 34304
rect 5276 34240 5292 34304
rect 5356 34240 5372 34304
rect 5436 34240 5452 34304
rect 5516 34240 5524 34304
rect 5204 33216 5524 34240
rect 5204 33152 5212 33216
rect 5276 33152 5292 33216
rect 5356 33152 5372 33216
rect 5436 33152 5452 33216
rect 5516 33152 5524 33216
rect 5204 32128 5524 33152
rect 5204 32064 5212 32128
rect 5276 32064 5292 32128
rect 5356 32064 5372 32128
rect 5436 32064 5452 32128
rect 5516 32064 5524 32128
rect 5204 31040 5524 32064
rect 5204 30976 5212 31040
rect 5276 30976 5292 31040
rect 5356 30976 5372 31040
rect 5436 30976 5452 31040
rect 5516 30976 5524 31040
rect 5204 29952 5524 30976
rect 5204 29888 5212 29952
rect 5276 29888 5292 29952
rect 5356 29888 5372 29952
rect 5436 29888 5452 29952
rect 5516 29888 5524 29952
rect 5204 28864 5524 29888
rect 5204 28800 5212 28864
rect 5276 28800 5292 28864
rect 5356 28800 5372 28864
rect 5436 28800 5452 28864
rect 5516 28800 5524 28864
rect 5204 27776 5524 28800
rect 5204 27712 5212 27776
rect 5276 27712 5292 27776
rect 5356 27712 5372 27776
rect 5436 27712 5452 27776
rect 5516 27712 5524 27776
rect 5204 26688 5524 27712
rect 5204 26624 5212 26688
rect 5276 26624 5292 26688
rect 5356 26624 5372 26688
rect 5436 26624 5452 26688
rect 5516 26624 5524 26688
rect 5204 25600 5524 26624
rect 5204 25536 5212 25600
rect 5276 25536 5292 25600
rect 5356 25536 5372 25600
rect 5436 25536 5452 25600
rect 5516 25536 5524 25600
rect 5204 24512 5524 25536
rect 5204 24448 5212 24512
rect 5276 24448 5292 24512
rect 5356 24448 5372 24512
rect 5436 24448 5452 24512
rect 5516 24448 5524 24512
rect 5204 23424 5524 24448
rect 5204 23360 5212 23424
rect 5276 23360 5292 23424
rect 5356 23360 5372 23424
rect 5436 23360 5452 23424
rect 5516 23360 5524 23424
rect 5204 22336 5524 23360
rect 5204 22272 5212 22336
rect 5276 22272 5292 22336
rect 5356 22272 5372 22336
rect 5436 22272 5452 22336
rect 5516 22272 5524 22336
rect 5204 21248 5524 22272
rect 5204 21184 5212 21248
rect 5276 21184 5292 21248
rect 5356 21184 5372 21248
rect 5436 21184 5452 21248
rect 5516 21184 5524 21248
rect 5204 20160 5524 21184
rect 5204 20096 5212 20160
rect 5276 20096 5292 20160
rect 5356 20096 5372 20160
rect 5436 20096 5452 20160
rect 5516 20096 5524 20160
rect 5204 19072 5524 20096
rect 5204 19008 5212 19072
rect 5276 19008 5292 19072
rect 5356 19008 5372 19072
rect 5436 19008 5452 19072
rect 5516 19008 5524 19072
rect 5204 17984 5524 19008
rect 5204 17920 5212 17984
rect 5276 17920 5292 17984
rect 5356 17920 5372 17984
rect 5436 17920 5452 17984
rect 5516 17920 5524 17984
rect 5204 16896 5524 17920
rect 5204 16832 5212 16896
rect 5276 16832 5292 16896
rect 5356 16832 5372 16896
rect 5436 16832 5452 16896
rect 5516 16832 5524 16896
rect 5204 15808 5524 16832
rect 5204 15744 5212 15808
rect 5276 15744 5292 15808
rect 5356 15744 5372 15808
rect 5436 15744 5452 15808
rect 5516 15744 5524 15808
rect 5204 14720 5524 15744
rect 5204 14656 5212 14720
rect 5276 14656 5292 14720
rect 5356 14656 5372 14720
rect 5436 14656 5452 14720
rect 5516 14656 5524 14720
rect 5204 13632 5524 14656
rect 5204 13568 5212 13632
rect 5276 13568 5292 13632
rect 5356 13568 5372 13632
rect 5436 13568 5452 13632
rect 5516 13568 5524 13632
rect 5204 12544 5524 13568
rect 5204 12480 5212 12544
rect 5276 12480 5292 12544
rect 5356 12480 5372 12544
rect 5436 12480 5452 12544
rect 5516 12480 5524 12544
rect 5204 11456 5524 12480
rect 5204 11392 5212 11456
rect 5276 11392 5292 11456
rect 5356 11392 5372 11456
rect 5436 11392 5452 11456
rect 5516 11392 5524 11456
rect 5204 10368 5524 11392
rect 5204 10304 5212 10368
rect 5276 10304 5292 10368
rect 5356 10304 5372 10368
rect 5436 10304 5452 10368
rect 5516 10304 5524 10368
rect 5204 9280 5524 10304
rect 5204 9216 5212 9280
rect 5276 9216 5292 9280
rect 5356 9216 5372 9280
rect 5436 9216 5452 9280
rect 5516 9216 5524 9280
rect 5204 8192 5524 9216
rect 5204 8128 5212 8192
rect 5276 8128 5292 8192
rect 5356 8128 5372 8192
rect 5436 8128 5452 8192
rect 5516 8128 5524 8192
rect 5204 7104 5524 8128
rect 5204 7040 5212 7104
rect 5276 7040 5292 7104
rect 5356 7040 5372 7104
rect 5436 7040 5452 7104
rect 5516 7040 5524 7104
rect 5204 6866 5524 7040
rect 5204 6630 5246 6866
rect 5482 6630 5524 6866
rect 5204 6016 5524 6630
rect 5204 5952 5212 6016
rect 5276 5952 5292 6016
rect 5356 5952 5372 6016
rect 5436 5952 5452 6016
rect 5516 5952 5524 6016
rect 5204 4928 5524 5952
rect 5204 4864 5212 4928
rect 5276 4864 5292 4928
rect 5356 4864 5372 4928
rect 5436 4864 5452 4928
rect 5516 4864 5524 4928
rect 5204 3840 5524 4864
rect 5204 3776 5212 3840
rect 5276 3776 5292 3840
rect 5356 3776 5372 3840
rect 5436 3776 5452 3840
rect 5516 3776 5524 3840
rect 5204 2752 5524 3776
rect 5204 2688 5212 2752
rect 5276 2688 5292 2752
rect 5356 2688 5372 2752
rect 5436 2688 5452 2752
rect 5516 2688 5524 2752
rect 5204 1664 5524 2688
rect 5204 1600 5212 1664
rect 5276 1600 5292 1664
rect 5356 1600 5372 1664
rect 5436 1600 5452 1664
rect 5516 1600 5524 1664
rect 5204 -154 5524 1600
rect 5204 -390 5246 -154
rect 5482 -390 5524 -154
rect 5204 -1092 5524 -390
rect 6144 88634 6464 88676
rect 6144 88398 6186 88634
rect 6422 88398 6464 88634
rect 6144 85984 6464 88398
rect 6144 85920 6152 85984
rect 6216 85920 6232 85984
rect 6296 85920 6312 85984
rect 6376 85920 6392 85984
rect 6456 85920 6464 85984
rect 6144 84896 6464 85920
rect 6144 84832 6152 84896
rect 6216 84832 6232 84896
rect 6296 84832 6312 84896
rect 6376 84832 6392 84896
rect 6456 84832 6464 84896
rect 6144 83808 6464 84832
rect 6144 83744 6152 83808
rect 6216 83744 6232 83808
rect 6296 83744 6312 83808
rect 6376 83744 6392 83808
rect 6456 83744 6464 83808
rect 6144 82720 6464 83744
rect 6144 82656 6152 82720
rect 6216 82656 6232 82720
rect 6296 82656 6312 82720
rect 6376 82656 6392 82720
rect 6456 82656 6464 82720
rect 6144 82206 6464 82656
rect 6144 81970 6186 82206
rect 6422 81970 6464 82206
rect 6144 81632 6464 81970
rect 6144 81568 6152 81632
rect 6216 81568 6232 81632
rect 6296 81568 6312 81632
rect 6376 81568 6392 81632
rect 6456 81568 6464 81632
rect 6144 80544 6464 81568
rect 6144 80480 6152 80544
rect 6216 80480 6232 80544
rect 6296 80480 6312 80544
rect 6376 80480 6392 80544
rect 6456 80480 6464 80544
rect 6144 79456 6464 80480
rect 6144 79392 6152 79456
rect 6216 79392 6232 79456
rect 6296 79392 6312 79456
rect 6376 79392 6392 79456
rect 6456 79392 6464 79456
rect 6144 78368 6464 79392
rect 6144 78304 6152 78368
rect 6216 78304 6232 78368
rect 6296 78304 6312 78368
rect 6376 78304 6392 78368
rect 6456 78304 6464 78368
rect 6144 77280 6464 78304
rect 6144 77216 6152 77280
rect 6216 77216 6232 77280
rect 6296 77216 6312 77280
rect 6376 77216 6392 77280
rect 6456 77216 6464 77280
rect 6144 76192 6464 77216
rect 6144 76128 6152 76192
rect 6216 76128 6232 76192
rect 6296 76128 6312 76192
rect 6376 76128 6392 76192
rect 6456 76128 6464 76192
rect 6144 75104 6464 76128
rect 6144 75040 6152 75104
rect 6216 75040 6232 75104
rect 6296 75040 6312 75104
rect 6376 75040 6392 75104
rect 6456 75040 6464 75104
rect 6144 74016 6464 75040
rect 6144 73952 6152 74016
rect 6216 73952 6232 74016
rect 6296 73952 6312 74016
rect 6376 73952 6392 74016
rect 6456 73952 6464 74016
rect 6144 72928 6464 73952
rect 6144 72864 6152 72928
rect 6216 72864 6232 72928
rect 6296 72864 6312 72928
rect 6376 72864 6392 72928
rect 6456 72864 6464 72928
rect 6144 71840 6464 72864
rect 6144 71776 6152 71840
rect 6216 71776 6232 71840
rect 6296 71776 6312 71840
rect 6376 71776 6392 71840
rect 6456 71776 6464 71840
rect 6144 70752 6464 71776
rect 6144 70688 6152 70752
rect 6216 70688 6232 70752
rect 6296 70688 6312 70752
rect 6376 70688 6392 70752
rect 6456 70688 6464 70752
rect 6144 69664 6464 70688
rect 6144 69600 6152 69664
rect 6216 69600 6232 69664
rect 6296 69600 6312 69664
rect 6376 69600 6392 69664
rect 6456 69600 6464 69664
rect 6144 68576 6464 69600
rect 6144 68512 6152 68576
rect 6216 68512 6232 68576
rect 6296 68512 6312 68576
rect 6376 68512 6392 68576
rect 6456 68512 6464 68576
rect 6144 67488 6464 68512
rect 6144 67424 6152 67488
rect 6216 67424 6232 67488
rect 6296 67424 6312 67488
rect 6376 67424 6392 67488
rect 6456 67424 6464 67488
rect 6144 66400 6464 67424
rect 6144 66336 6152 66400
rect 6216 66336 6232 66400
rect 6296 66336 6312 66400
rect 6376 66336 6392 66400
rect 6456 66336 6464 66400
rect 6144 65312 6464 66336
rect 6144 65248 6152 65312
rect 6216 65248 6232 65312
rect 6296 65248 6312 65312
rect 6376 65248 6392 65312
rect 6456 65248 6464 65312
rect 6144 64224 6464 65248
rect 6144 64160 6152 64224
rect 6216 64160 6232 64224
rect 6296 64160 6312 64224
rect 6376 64160 6392 64224
rect 6456 64160 6464 64224
rect 6144 63136 6464 64160
rect 6144 63072 6152 63136
rect 6216 63072 6232 63136
rect 6296 63072 6312 63136
rect 6376 63072 6392 63136
rect 6456 63072 6464 63136
rect 6144 62048 6464 63072
rect 6144 61984 6152 62048
rect 6216 61984 6232 62048
rect 6296 61984 6312 62048
rect 6376 61984 6392 62048
rect 6456 61984 6464 62048
rect 6144 60960 6464 61984
rect 6144 60896 6152 60960
rect 6216 60896 6232 60960
rect 6296 60896 6312 60960
rect 6376 60896 6392 60960
rect 6456 60896 6464 60960
rect 6144 59872 6464 60896
rect 6144 59808 6152 59872
rect 6216 59808 6232 59872
rect 6296 59808 6312 59872
rect 6376 59808 6392 59872
rect 6456 59808 6464 59872
rect 6144 58784 6464 59808
rect 6144 58720 6152 58784
rect 6216 58720 6232 58784
rect 6296 58720 6312 58784
rect 6376 58720 6392 58784
rect 6456 58720 6464 58784
rect 6144 57696 6464 58720
rect 6144 57632 6152 57696
rect 6216 57632 6232 57696
rect 6296 57632 6312 57696
rect 6376 57632 6392 57696
rect 6456 57632 6464 57696
rect 6144 56608 6464 57632
rect 6144 56544 6152 56608
rect 6216 56544 6232 56608
rect 6296 56544 6312 56608
rect 6376 56544 6392 56608
rect 6456 56544 6464 56608
rect 6144 55520 6464 56544
rect 6144 55456 6152 55520
rect 6216 55456 6232 55520
rect 6296 55456 6312 55520
rect 6376 55456 6392 55520
rect 6456 55456 6464 55520
rect 6144 54432 6464 55456
rect 6144 54368 6152 54432
rect 6216 54368 6232 54432
rect 6296 54368 6312 54432
rect 6376 54368 6392 54432
rect 6456 54368 6464 54432
rect 6144 53344 6464 54368
rect 6144 53280 6152 53344
rect 6216 53280 6232 53344
rect 6296 53280 6312 53344
rect 6376 53280 6392 53344
rect 6456 53280 6464 53344
rect 6144 52256 6464 53280
rect 6144 52192 6152 52256
rect 6216 52192 6232 52256
rect 6296 52192 6312 52256
rect 6376 52192 6392 52256
rect 6456 52192 6464 52256
rect 6144 51168 6464 52192
rect 6144 51104 6152 51168
rect 6216 51104 6232 51168
rect 6296 51104 6312 51168
rect 6376 51104 6392 51168
rect 6456 51104 6464 51168
rect 6144 50080 6464 51104
rect 6144 50016 6152 50080
rect 6216 50016 6232 50080
rect 6296 50016 6312 50080
rect 6376 50016 6392 50080
rect 6456 50016 6464 50080
rect 6144 48992 6464 50016
rect 6144 48928 6152 48992
rect 6216 48928 6232 48992
rect 6296 48928 6312 48992
rect 6376 48928 6392 48992
rect 6456 48928 6464 48992
rect 6144 47904 6464 48928
rect 6144 47840 6152 47904
rect 6216 47840 6232 47904
rect 6296 47840 6312 47904
rect 6376 47840 6392 47904
rect 6456 47840 6464 47904
rect 6144 46816 6464 47840
rect 6144 46752 6152 46816
rect 6216 46752 6232 46816
rect 6296 46752 6312 46816
rect 6376 46752 6392 46816
rect 6456 46752 6464 46816
rect 6144 45728 6464 46752
rect 6144 45664 6152 45728
rect 6216 45664 6232 45728
rect 6296 45664 6312 45728
rect 6376 45664 6392 45728
rect 6456 45664 6464 45728
rect 6144 44640 6464 45664
rect 6144 44576 6152 44640
rect 6216 44576 6232 44640
rect 6296 44576 6312 44640
rect 6376 44576 6392 44640
rect 6456 44576 6464 44640
rect 6144 43552 6464 44576
rect 6144 43488 6152 43552
rect 6216 43488 6232 43552
rect 6296 43488 6312 43552
rect 6376 43488 6392 43552
rect 6456 43488 6464 43552
rect 6144 42464 6464 43488
rect 6144 42400 6152 42464
rect 6216 42400 6232 42464
rect 6296 42400 6312 42464
rect 6376 42400 6392 42464
rect 6456 42400 6464 42464
rect 6144 41376 6464 42400
rect 6144 41312 6152 41376
rect 6216 41312 6232 41376
rect 6296 41312 6312 41376
rect 6376 41312 6392 41376
rect 6456 41312 6464 41376
rect 6144 40288 6464 41312
rect 6144 40224 6152 40288
rect 6216 40224 6232 40288
rect 6296 40224 6312 40288
rect 6376 40224 6392 40288
rect 6456 40224 6464 40288
rect 6144 39200 6464 40224
rect 6144 39136 6152 39200
rect 6216 39136 6232 39200
rect 6296 39136 6312 39200
rect 6376 39136 6392 39200
rect 6456 39136 6464 39200
rect 6144 38112 6464 39136
rect 6144 38048 6152 38112
rect 6216 38048 6232 38112
rect 6296 38048 6312 38112
rect 6376 38048 6392 38112
rect 6456 38048 6464 38112
rect 6144 37024 6464 38048
rect 6144 36960 6152 37024
rect 6216 36960 6232 37024
rect 6296 36960 6312 37024
rect 6376 36960 6392 37024
rect 6456 36960 6464 37024
rect 6144 35936 6464 36960
rect 6144 35872 6152 35936
rect 6216 35872 6232 35936
rect 6296 35872 6312 35936
rect 6376 35872 6392 35936
rect 6456 35872 6464 35936
rect 6144 34848 6464 35872
rect 6144 34784 6152 34848
rect 6216 34784 6232 34848
rect 6296 34784 6312 34848
rect 6376 34784 6392 34848
rect 6456 34784 6464 34848
rect 6144 33760 6464 34784
rect 6144 33696 6152 33760
rect 6216 33696 6232 33760
rect 6296 33696 6312 33760
rect 6376 33696 6392 33760
rect 6456 33696 6464 33760
rect 6144 32672 6464 33696
rect 6144 32608 6152 32672
rect 6216 32608 6232 32672
rect 6296 32608 6312 32672
rect 6376 32608 6392 32672
rect 6456 32608 6464 32672
rect 6144 31584 6464 32608
rect 6144 31520 6152 31584
rect 6216 31520 6232 31584
rect 6296 31520 6312 31584
rect 6376 31520 6392 31584
rect 6456 31520 6464 31584
rect 6144 30496 6464 31520
rect 6144 30432 6152 30496
rect 6216 30432 6232 30496
rect 6296 30432 6312 30496
rect 6376 30432 6392 30496
rect 6456 30432 6464 30496
rect 6144 29408 6464 30432
rect 6144 29344 6152 29408
rect 6216 29344 6232 29408
rect 6296 29344 6312 29408
rect 6376 29344 6392 29408
rect 6456 29344 6464 29408
rect 6144 28320 6464 29344
rect 6144 28256 6152 28320
rect 6216 28256 6232 28320
rect 6296 28256 6312 28320
rect 6376 28256 6392 28320
rect 6456 28256 6464 28320
rect 6144 27232 6464 28256
rect 6144 27168 6152 27232
rect 6216 27168 6232 27232
rect 6296 27168 6312 27232
rect 6376 27168 6392 27232
rect 6456 27168 6464 27232
rect 6144 26144 6464 27168
rect 6144 26080 6152 26144
rect 6216 26080 6232 26144
rect 6296 26080 6312 26144
rect 6376 26080 6392 26144
rect 6456 26080 6464 26144
rect 6144 25056 6464 26080
rect 6144 24992 6152 25056
rect 6216 24992 6232 25056
rect 6296 24992 6312 25056
rect 6376 24992 6392 25056
rect 6456 24992 6464 25056
rect 6144 23968 6464 24992
rect 6144 23904 6152 23968
rect 6216 23904 6232 23968
rect 6296 23904 6312 23968
rect 6376 23904 6392 23968
rect 6456 23904 6464 23968
rect 6144 22880 6464 23904
rect 6144 22816 6152 22880
rect 6216 22816 6232 22880
rect 6296 22816 6312 22880
rect 6376 22816 6392 22880
rect 6456 22816 6464 22880
rect 6144 21792 6464 22816
rect 6144 21728 6152 21792
rect 6216 21728 6232 21792
rect 6296 21728 6312 21792
rect 6376 21728 6392 21792
rect 6456 21728 6464 21792
rect 6144 20704 6464 21728
rect 6144 20640 6152 20704
rect 6216 20640 6232 20704
rect 6296 20640 6312 20704
rect 6376 20640 6392 20704
rect 6456 20640 6464 20704
rect 6144 19616 6464 20640
rect 6144 19552 6152 19616
rect 6216 19552 6232 19616
rect 6296 19552 6312 19616
rect 6376 19552 6392 19616
rect 6456 19552 6464 19616
rect 6144 18528 6464 19552
rect 6144 18464 6152 18528
rect 6216 18464 6232 18528
rect 6296 18464 6312 18528
rect 6376 18464 6392 18528
rect 6456 18464 6464 18528
rect 6144 17440 6464 18464
rect 6144 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6392 17440
rect 6456 17376 6464 17440
rect 6144 16352 6464 17376
rect 6144 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6392 16352
rect 6456 16288 6464 16352
rect 6144 15264 6464 16288
rect 6144 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6392 15264
rect 6456 15200 6464 15264
rect 6144 14176 6464 15200
rect 6144 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6392 14176
rect 6456 14112 6464 14176
rect 6144 13088 6464 14112
rect 6144 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6392 13088
rect 6456 13024 6464 13088
rect 6144 12000 6464 13024
rect 6144 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6392 12000
rect 6456 11936 6464 12000
rect 6144 10912 6464 11936
rect 6144 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6392 10912
rect 6456 10848 6464 10912
rect 6144 9824 6464 10848
rect 6144 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6392 9824
rect 6456 9760 6464 9824
rect 6144 8736 6464 9760
rect 6144 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6392 8736
rect 6456 8672 6464 8736
rect 6144 7648 6464 8672
rect 6144 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6392 7648
rect 6456 7584 6464 7648
rect 6144 6560 6464 7584
rect 6144 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6392 6560
rect 6456 6496 6464 6560
rect 6144 6206 6464 6496
rect 6144 5970 6186 6206
rect 6422 5970 6464 6206
rect 6144 5472 6464 5970
rect 6144 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6392 5472
rect 6456 5408 6464 5472
rect 6144 4384 6464 5408
rect 6144 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6392 4384
rect 6456 4320 6464 4384
rect 6144 3296 6464 4320
rect 6144 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6392 3296
rect 6456 3232 6464 3296
rect 6144 2208 6464 3232
rect 6144 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6392 2208
rect 6456 2144 6464 2208
rect 6144 1120 6464 2144
rect 6144 1056 6152 1120
rect 6216 1056 6232 1120
rect 6296 1056 6312 1120
rect 6376 1056 6392 1120
rect 6456 1056 6464 1120
rect 6144 -814 6464 1056
rect 6144 -1050 6186 -814
rect 6422 -1050 6464 -814
rect 6144 -1092 6464 -1050
rect 6804 87974 7124 88676
rect 6804 87738 6846 87974
rect 7082 87738 7124 87974
rect 6804 86528 7124 87738
rect 6804 86464 6812 86528
rect 6876 86464 6892 86528
rect 6956 86464 6972 86528
rect 7036 86464 7052 86528
rect 7116 86464 7124 86528
rect 6804 85440 7124 86464
rect 6804 85376 6812 85440
rect 6876 85376 6892 85440
rect 6956 85376 6972 85440
rect 7036 85376 7052 85440
rect 7116 85376 7124 85440
rect 6804 84352 7124 85376
rect 6804 84288 6812 84352
rect 6876 84288 6892 84352
rect 6956 84288 6972 84352
rect 7036 84288 7052 84352
rect 7116 84288 7124 84352
rect 6804 83264 7124 84288
rect 6804 83200 6812 83264
rect 6876 83200 6892 83264
rect 6956 83200 6972 83264
rect 7036 83200 7052 83264
rect 7116 83200 7124 83264
rect 6804 82866 7124 83200
rect 6804 82630 6846 82866
rect 7082 82630 7124 82866
rect 6804 82176 7124 82630
rect 6804 82112 6812 82176
rect 6876 82112 6892 82176
rect 6956 82112 6972 82176
rect 7036 82112 7052 82176
rect 7116 82112 7124 82176
rect 6804 81088 7124 82112
rect 6804 81024 6812 81088
rect 6876 81024 6892 81088
rect 6956 81024 6972 81088
rect 7036 81024 7052 81088
rect 7116 81024 7124 81088
rect 6804 80000 7124 81024
rect 6804 79936 6812 80000
rect 6876 79936 6892 80000
rect 6956 79936 6972 80000
rect 7036 79936 7052 80000
rect 7116 79936 7124 80000
rect 6804 78912 7124 79936
rect 6804 78848 6812 78912
rect 6876 78848 6892 78912
rect 6956 78848 6972 78912
rect 7036 78848 7052 78912
rect 7116 78848 7124 78912
rect 6804 77824 7124 78848
rect 6804 77760 6812 77824
rect 6876 77760 6892 77824
rect 6956 77760 6972 77824
rect 7036 77760 7052 77824
rect 7116 77760 7124 77824
rect 6804 76736 7124 77760
rect 6804 76672 6812 76736
rect 6876 76672 6892 76736
rect 6956 76672 6972 76736
rect 7036 76672 7052 76736
rect 7116 76672 7124 76736
rect 6804 75648 7124 76672
rect 6804 75584 6812 75648
rect 6876 75584 6892 75648
rect 6956 75584 6972 75648
rect 7036 75584 7052 75648
rect 7116 75584 7124 75648
rect 6804 74560 7124 75584
rect 6804 74496 6812 74560
rect 6876 74496 6892 74560
rect 6956 74496 6972 74560
rect 7036 74496 7052 74560
rect 7116 74496 7124 74560
rect 6804 73472 7124 74496
rect 6804 73408 6812 73472
rect 6876 73408 6892 73472
rect 6956 73408 6972 73472
rect 7036 73408 7052 73472
rect 7116 73408 7124 73472
rect 6804 72384 7124 73408
rect 6804 72320 6812 72384
rect 6876 72320 6892 72384
rect 6956 72320 6972 72384
rect 7036 72320 7052 72384
rect 7116 72320 7124 72384
rect 6804 71296 7124 72320
rect 6804 71232 6812 71296
rect 6876 71232 6892 71296
rect 6956 71232 6972 71296
rect 7036 71232 7052 71296
rect 7116 71232 7124 71296
rect 6804 70208 7124 71232
rect 6804 70144 6812 70208
rect 6876 70144 6892 70208
rect 6956 70144 6972 70208
rect 7036 70144 7052 70208
rect 7116 70144 7124 70208
rect 6804 69120 7124 70144
rect 6804 69056 6812 69120
rect 6876 69056 6892 69120
rect 6956 69056 6972 69120
rect 7036 69056 7052 69120
rect 7116 69056 7124 69120
rect 6804 68032 7124 69056
rect 6804 67968 6812 68032
rect 6876 67968 6892 68032
rect 6956 67968 6972 68032
rect 7036 67968 7052 68032
rect 7116 67968 7124 68032
rect 6804 66944 7124 67968
rect 6804 66880 6812 66944
rect 6876 66880 6892 66944
rect 6956 66880 6972 66944
rect 7036 66880 7052 66944
rect 7116 66880 7124 66944
rect 6804 65856 7124 66880
rect 6804 65792 6812 65856
rect 6876 65792 6892 65856
rect 6956 65792 6972 65856
rect 7036 65792 7052 65856
rect 7116 65792 7124 65856
rect 6804 64768 7124 65792
rect 6804 64704 6812 64768
rect 6876 64704 6892 64768
rect 6956 64704 6972 64768
rect 7036 64704 7052 64768
rect 7116 64704 7124 64768
rect 6804 63680 7124 64704
rect 6804 63616 6812 63680
rect 6876 63616 6892 63680
rect 6956 63616 6972 63680
rect 7036 63616 7052 63680
rect 7116 63616 7124 63680
rect 6804 62592 7124 63616
rect 6804 62528 6812 62592
rect 6876 62528 6892 62592
rect 6956 62528 6972 62592
rect 7036 62528 7052 62592
rect 7116 62528 7124 62592
rect 6804 61504 7124 62528
rect 6804 61440 6812 61504
rect 6876 61440 6892 61504
rect 6956 61440 6972 61504
rect 7036 61440 7052 61504
rect 7116 61440 7124 61504
rect 6804 60416 7124 61440
rect 6804 60352 6812 60416
rect 6876 60352 6892 60416
rect 6956 60352 6972 60416
rect 7036 60352 7052 60416
rect 7116 60352 7124 60416
rect 6804 59328 7124 60352
rect 6804 59264 6812 59328
rect 6876 59264 6892 59328
rect 6956 59264 6972 59328
rect 7036 59264 7052 59328
rect 7116 59264 7124 59328
rect 6804 58240 7124 59264
rect 6804 58176 6812 58240
rect 6876 58176 6892 58240
rect 6956 58176 6972 58240
rect 7036 58176 7052 58240
rect 7116 58176 7124 58240
rect 6804 57152 7124 58176
rect 6804 57088 6812 57152
rect 6876 57088 6892 57152
rect 6956 57088 6972 57152
rect 7036 57088 7052 57152
rect 7116 57088 7124 57152
rect 6804 56064 7124 57088
rect 6804 56000 6812 56064
rect 6876 56000 6892 56064
rect 6956 56000 6972 56064
rect 7036 56000 7052 56064
rect 7116 56000 7124 56064
rect 6804 54976 7124 56000
rect 6804 54912 6812 54976
rect 6876 54912 6892 54976
rect 6956 54912 6972 54976
rect 7036 54912 7052 54976
rect 7116 54912 7124 54976
rect 6804 53888 7124 54912
rect 6804 53824 6812 53888
rect 6876 53824 6892 53888
rect 6956 53824 6972 53888
rect 7036 53824 7052 53888
rect 7116 53824 7124 53888
rect 6804 52800 7124 53824
rect 6804 52736 6812 52800
rect 6876 52736 6892 52800
rect 6956 52736 6972 52800
rect 7036 52736 7052 52800
rect 7116 52736 7124 52800
rect 6804 51712 7124 52736
rect 6804 51648 6812 51712
rect 6876 51648 6892 51712
rect 6956 51648 6972 51712
rect 7036 51648 7052 51712
rect 7116 51648 7124 51712
rect 6804 50624 7124 51648
rect 6804 50560 6812 50624
rect 6876 50560 6892 50624
rect 6956 50560 6972 50624
rect 7036 50560 7052 50624
rect 7116 50560 7124 50624
rect 6804 49536 7124 50560
rect 6804 49472 6812 49536
rect 6876 49472 6892 49536
rect 6956 49472 6972 49536
rect 7036 49472 7052 49536
rect 7116 49472 7124 49536
rect 6804 48448 7124 49472
rect 6804 48384 6812 48448
rect 6876 48384 6892 48448
rect 6956 48384 6972 48448
rect 7036 48384 7052 48448
rect 7116 48384 7124 48448
rect 6804 47360 7124 48384
rect 6804 47296 6812 47360
rect 6876 47296 6892 47360
rect 6956 47296 6972 47360
rect 7036 47296 7052 47360
rect 7116 47296 7124 47360
rect 6804 46272 7124 47296
rect 6804 46208 6812 46272
rect 6876 46208 6892 46272
rect 6956 46208 6972 46272
rect 7036 46208 7052 46272
rect 7116 46208 7124 46272
rect 6804 45184 7124 46208
rect 6804 45120 6812 45184
rect 6876 45120 6892 45184
rect 6956 45120 6972 45184
rect 7036 45120 7052 45184
rect 7116 45120 7124 45184
rect 6804 44096 7124 45120
rect 6804 44032 6812 44096
rect 6876 44032 6892 44096
rect 6956 44032 6972 44096
rect 7036 44032 7052 44096
rect 7116 44032 7124 44096
rect 6804 43008 7124 44032
rect 6804 42944 6812 43008
rect 6876 42944 6892 43008
rect 6956 42944 6972 43008
rect 7036 42944 7052 43008
rect 7116 42944 7124 43008
rect 6804 41920 7124 42944
rect 6804 41856 6812 41920
rect 6876 41856 6892 41920
rect 6956 41856 6972 41920
rect 7036 41856 7052 41920
rect 7116 41856 7124 41920
rect 6804 40832 7124 41856
rect 6804 40768 6812 40832
rect 6876 40768 6892 40832
rect 6956 40768 6972 40832
rect 7036 40768 7052 40832
rect 7116 40768 7124 40832
rect 6804 39744 7124 40768
rect 6804 39680 6812 39744
rect 6876 39680 6892 39744
rect 6956 39680 6972 39744
rect 7036 39680 7052 39744
rect 7116 39680 7124 39744
rect 6804 38656 7124 39680
rect 6804 38592 6812 38656
rect 6876 38592 6892 38656
rect 6956 38592 6972 38656
rect 7036 38592 7052 38656
rect 7116 38592 7124 38656
rect 6804 37568 7124 38592
rect 6804 37504 6812 37568
rect 6876 37504 6892 37568
rect 6956 37504 6972 37568
rect 7036 37504 7052 37568
rect 7116 37504 7124 37568
rect 6804 36480 7124 37504
rect 6804 36416 6812 36480
rect 6876 36416 6892 36480
rect 6956 36416 6972 36480
rect 7036 36416 7052 36480
rect 7116 36416 7124 36480
rect 6804 35392 7124 36416
rect 6804 35328 6812 35392
rect 6876 35328 6892 35392
rect 6956 35328 6972 35392
rect 7036 35328 7052 35392
rect 7116 35328 7124 35392
rect 6804 34304 7124 35328
rect 6804 34240 6812 34304
rect 6876 34240 6892 34304
rect 6956 34240 6972 34304
rect 7036 34240 7052 34304
rect 7116 34240 7124 34304
rect 6804 33216 7124 34240
rect 6804 33152 6812 33216
rect 6876 33152 6892 33216
rect 6956 33152 6972 33216
rect 7036 33152 7052 33216
rect 7116 33152 7124 33216
rect 6804 32128 7124 33152
rect 6804 32064 6812 32128
rect 6876 32064 6892 32128
rect 6956 32064 6972 32128
rect 7036 32064 7052 32128
rect 7116 32064 7124 32128
rect 6804 31040 7124 32064
rect 6804 30976 6812 31040
rect 6876 30976 6892 31040
rect 6956 30976 6972 31040
rect 7036 30976 7052 31040
rect 7116 30976 7124 31040
rect 6804 29952 7124 30976
rect 6804 29888 6812 29952
rect 6876 29888 6892 29952
rect 6956 29888 6972 29952
rect 7036 29888 7052 29952
rect 7116 29888 7124 29952
rect 6804 28864 7124 29888
rect 6804 28800 6812 28864
rect 6876 28800 6892 28864
rect 6956 28800 6972 28864
rect 7036 28800 7052 28864
rect 7116 28800 7124 28864
rect 6804 27776 7124 28800
rect 6804 27712 6812 27776
rect 6876 27712 6892 27776
rect 6956 27712 6972 27776
rect 7036 27712 7052 27776
rect 7116 27712 7124 27776
rect 6804 26688 7124 27712
rect 6804 26624 6812 26688
rect 6876 26624 6892 26688
rect 6956 26624 6972 26688
rect 7036 26624 7052 26688
rect 7116 26624 7124 26688
rect 6804 25600 7124 26624
rect 6804 25536 6812 25600
rect 6876 25536 6892 25600
rect 6956 25536 6972 25600
rect 7036 25536 7052 25600
rect 7116 25536 7124 25600
rect 6804 24512 7124 25536
rect 6804 24448 6812 24512
rect 6876 24448 6892 24512
rect 6956 24448 6972 24512
rect 7036 24448 7052 24512
rect 7116 24448 7124 24512
rect 6804 23424 7124 24448
rect 6804 23360 6812 23424
rect 6876 23360 6892 23424
rect 6956 23360 6972 23424
rect 7036 23360 7052 23424
rect 7116 23360 7124 23424
rect 6804 22336 7124 23360
rect 6804 22272 6812 22336
rect 6876 22272 6892 22336
rect 6956 22272 6972 22336
rect 7036 22272 7052 22336
rect 7116 22272 7124 22336
rect 6804 21248 7124 22272
rect 6804 21184 6812 21248
rect 6876 21184 6892 21248
rect 6956 21184 6972 21248
rect 7036 21184 7052 21248
rect 7116 21184 7124 21248
rect 6804 20160 7124 21184
rect 6804 20096 6812 20160
rect 6876 20096 6892 20160
rect 6956 20096 6972 20160
rect 7036 20096 7052 20160
rect 7116 20096 7124 20160
rect 6804 19072 7124 20096
rect 6804 19008 6812 19072
rect 6876 19008 6892 19072
rect 6956 19008 6972 19072
rect 7036 19008 7052 19072
rect 7116 19008 7124 19072
rect 6804 17984 7124 19008
rect 6804 17920 6812 17984
rect 6876 17920 6892 17984
rect 6956 17920 6972 17984
rect 7036 17920 7052 17984
rect 7116 17920 7124 17984
rect 6804 16896 7124 17920
rect 6804 16832 6812 16896
rect 6876 16832 6892 16896
rect 6956 16832 6972 16896
rect 7036 16832 7052 16896
rect 7116 16832 7124 16896
rect 6804 15808 7124 16832
rect 6804 15744 6812 15808
rect 6876 15744 6892 15808
rect 6956 15744 6972 15808
rect 7036 15744 7052 15808
rect 7116 15744 7124 15808
rect 6804 14720 7124 15744
rect 6804 14656 6812 14720
rect 6876 14656 6892 14720
rect 6956 14656 6972 14720
rect 7036 14656 7052 14720
rect 7116 14656 7124 14720
rect 6804 13632 7124 14656
rect 6804 13568 6812 13632
rect 6876 13568 6892 13632
rect 6956 13568 6972 13632
rect 7036 13568 7052 13632
rect 7116 13568 7124 13632
rect 6804 12544 7124 13568
rect 6804 12480 6812 12544
rect 6876 12480 6892 12544
rect 6956 12480 6972 12544
rect 7036 12480 7052 12544
rect 7116 12480 7124 12544
rect 6804 11456 7124 12480
rect 6804 11392 6812 11456
rect 6876 11392 6892 11456
rect 6956 11392 6972 11456
rect 7036 11392 7052 11456
rect 7116 11392 7124 11456
rect 6804 10368 7124 11392
rect 6804 10304 6812 10368
rect 6876 10304 6892 10368
rect 6956 10304 6972 10368
rect 7036 10304 7052 10368
rect 7116 10304 7124 10368
rect 6804 9280 7124 10304
rect 6804 9216 6812 9280
rect 6876 9216 6892 9280
rect 6956 9216 6972 9280
rect 7036 9216 7052 9280
rect 7116 9216 7124 9280
rect 6804 8192 7124 9216
rect 6804 8128 6812 8192
rect 6876 8128 6892 8192
rect 6956 8128 6972 8192
rect 7036 8128 7052 8192
rect 7116 8128 7124 8192
rect 6804 7104 7124 8128
rect 6804 7040 6812 7104
rect 6876 7040 6892 7104
rect 6956 7040 6972 7104
rect 7036 7040 7052 7104
rect 7116 7040 7124 7104
rect 6804 6866 7124 7040
rect 6804 6630 6846 6866
rect 7082 6630 7124 6866
rect 6804 6016 7124 6630
rect 6804 5952 6812 6016
rect 6876 5952 6892 6016
rect 6956 5952 6972 6016
rect 7036 5952 7052 6016
rect 7116 5952 7124 6016
rect 6804 4928 7124 5952
rect 6804 4864 6812 4928
rect 6876 4864 6892 4928
rect 6956 4864 6972 4928
rect 7036 4864 7052 4928
rect 7116 4864 7124 4928
rect 6804 3840 7124 4864
rect 6804 3776 6812 3840
rect 6876 3776 6892 3840
rect 6956 3776 6972 3840
rect 7036 3776 7052 3840
rect 7116 3776 7124 3840
rect 6804 2752 7124 3776
rect 6804 2688 6812 2752
rect 6876 2688 6892 2752
rect 6956 2688 6972 2752
rect 7036 2688 7052 2752
rect 7116 2688 7124 2752
rect 6804 1664 7124 2688
rect 6804 1600 6812 1664
rect 6876 1600 6892 1664
rect 6956 1600 6972 1664
rect 7036 1600 7052 1664
rect 7116 1600 7124 1664
rect 6804 -154 7124 1600
rect 6804 -390 6846 -154
rect 7082 -390 7124 -154
rect 6804 -1092 7124 -390
rect 7744 88634 8064 88676
rect 7744 88398 7786 88634
rect 8022 88398 8064 88634
rect 7744 85984 8064 88398
rect 7744 85920 7752 85984
rect 7816 85920 7832 85984
rect 7896 85920 7912 85984
rect 7976 85920 7992 85984
rect 8056 85920 8064 85984
rect 7744 84896 8064 85920
rect 7744 84832 7752 84896
rect 7816 84832 7832 84896
rect 7896 84832 7912 84896
rect 7976 84832 7992 84896
rect 8056 84832 8064 84896
rect 7744 83808 8064 84832
rect 7744 83744 7752 83808
rect 7816 83744 7832 83808
rect 7896 83744 7912 83808
rect 7976 83744 7992 83808
rect 8056 83744 8064 83808
rect 7744 82720 8064 83744
rect 7744 82656 7752 82720
rect 7816 82656 7832 82720
rect 7896 82656 7912 82720
rect 7976 82656 7992 82720
rect 8056 82656 8064 82720
rect 7744 82206 8064 82656
rect 7744 81970 7786 82206
rect 8022 81970 8064 82206
rect 7744 81632 8064 81970
rect 7744 81568 7752 81632
rect 7816 81568 7832 81632
rect 7896 81568 7912 81632
rect 7976 81568 7992 81632
rect 8056 81568 8064 81632
rect 7744 80544 8064 81568
rect 7744 80480 7752 80544
rect 7816 80480 7832 80544
rect 7896 80480 7912 80544
rect 7976 80480 7992 80544
rect 8056 80480 8064 80544
rect 7744 79456 8064 80480
rect 7744 79392 7752 79456
rect 7816 79392 7832 79456
rect 7896 79392 7912 79456
rect 7976 79392 7992 79456
rect 8056 79392 8064 79456
rect 7744 78368 8064 79392
rect 7744 78304 7752 78368
rect 7816 78304 7832 78368
rect 7896 78304 7912 78368
rect 7976 78304 7992 78368
rect 8056 78304 8064 78368
rect 7744 77280 8064 78304
rect 7744 77216 7752 77280
rect 7816 77216 7832 77280
rect 7896 77216 7912 77280
rect 7976 77216 7992 77280
rect 8056 77216 8064 77280
rect 7744 76192 8064 77216
rect 7744 76128 7752 76192
rect 7816 76128 7832 76192
rect 7896 76128 7912 76192
rect 7976 76128 7992 76192
rect 8056 76128 8064 76192
rect 7744 75104 8064 76128
rect 7744 75040 7752 75104
rect 7816 75040 7832 75104
rect 7896 75040 7912 75104
rect 7976 75040 7992 75104
rect 8056 75040 8064 75104
rect 7744 74016 8064 75040
rect 7744 73952 7752 74016
rect 7816 73952 7832 74016
rect 7896 73952 7912 74016
rect 7976 73952 7992 74016
rect 8056 73952 8064 74016
rect 7744 72928 8064 73952
rect 7744 72864 7752 72928
rect 7816 72864 7832 72928
rect 7896 72864 7912 72928
rect 7976 72864 7992 72928
rect 8056 72864 8064 72928
rect 7744 71840 8064 72864
rect 7744 71776 7752 71840
rect 7816 71776 7832 71840
rect 7896 71776 7912 71840
rect 7976 71776 7992 71840
rect 8056 71776 8064 71840
rect 7744 70752 8064 71776
rect 7744 70688 7752 70752
rect 7816 70688 7832 70752
rect 7896 70688 7912 70752
rect 7976 70688 7992 70752
rect 8056 70688 8064 70752
rect 7744 69664 8064 70688
rect 7744 69600 7752 69664
rect 7816 69600 7832 69664
rect 7896 69600 7912 69664
rect 7976 69600 7992 69664
rect 8056 69600 8064 69664
rect 7744 68576 8064 69600
rect 7744 68512 7752 68576
rect 7816 68512 7832 68576
rect 7896 68512 7912 68576
rect 7976 68512 7992 68576
rect 8056 68512 8064 68576
rect 7744 67488 8064 68512
rect 7744 67424 7752 67488
rect 7816 67424 7832 67488
rect 7896 67424 7912 67488
rect 7976 67424 7992 67488
rect 8056 67424 8064 67488
rect 7744 66400 8064 67424
rect 7744 66336 7752 66400
rect 7816 66336 7832 66400
rect 7896 66336 7912 66400
rect 7976 66336 7992 66400
rect 8056 66336 8064 66400
rect 7744 65312 8064 66336
rect 7744 65248 7752 65312
rect 7816 65248 7832 65312
rect 7896 65248 7912 65312
rect 7976 65248 7992 65312
rect 8056 65248 8064 65312
rect 7744 64224 8064 65248
rect 7744 64160 7752 64224
rect 7816 64160 7832 64224
rect 7896 64160 7912 64224
rect 7976 64160 7992 64224
rect 8056 64160 8064 64224
rect 7744 63136 8064 64160
rect 7744 63072 7752 63136
rect 7816 63072 7832 63136
rect 7896 63072 7912 63136
rect 7976 63072 7992 63136
rect 8056 63072 8064 63136
rect 7744 62048 8064 63072
rect 7744 61984 7752 62048
rect 7816 61984 7832 62048
rect 7896 61984 7912 62048
rect 7976 61984 7992 62048
rect 8056 61984 8064 62048
rect 7744 60960 8064 61984
rect 7744 60896 7752 60960
rect 7816 60896 7832 60960
rect 7896 60896 7912 60960
rect 7976 60896 7992 60960
rect 8056 60896 8064 60960
rect 7744 59872 8064 60896
rect 7744 59808 7752 59872
rect 7816 59808 7832 59872
rect 7896 59808 7912 59872
rect 7976 59808 7992 59872
rect 8056 59808 8064 59872
rect 7744 58784 8064 59808
rect 7744 58720 7752 58784
rect 7816 58720 7832 58784
rect 7896 58720 7912 58784
rect 7976 58720 7992 58784
rect 8056 58720 8064 58784
rect 7744 57696 8064 58720
rect 7744 57632 7752 57696
rect 7816 57632 7832 57696
rect 7896 57632 7912 57696
rect 7976 57632 7992 57696
rect 8056 57632 8064 57696
rect 7744 56608 8064 57632
rect 7744 56544 7752 56608
rect 7816 56544 7832 56608
rect 7896 56544 7912 56608
rect 7976 56544 7992 56608
rect 8056 56544 8064 56608
rect 7744 55520 8064 56544
rect 7744 55456 7752 55520
rect 7816 55456 7832 55520
rect 7896 55456 7912 55520
rect 7976 55456 7992 55520
rect 8056 55456 8064 55520
rect 7744 54432 8064 55456
rect 7744 54368 7752 54432
rect 7816 54368 7832 54432
rect 7896 54368 7912 54432
rect 7976 54368 7992 54432
rect 8056 54368 8064 54432
rect 7744 53344 8064 54368
rect 7744 53280 7752 53344
rect 7816 53280 7832 53344
rect 7896 53280 7912 53344
rect 7976 53280 7992 53344
rect 8056 53280 8064 53344
rect 7744 52256 8064 53280
rect 7744 52192 7752 52256
rect 7816 52192 7832 52256
rect 7896 52192 7912 52256
rect 7976 52192 7992 52256
rect 8056 52192 8064 52256
rect 7744 51168 8064 52192
rect 7744 51104 7752 51168
rect 7816 51104 7832 51168
rect 7896 51104 7912 51168
rect 7976 51104 7992 51168
rect 8056 51104 8064 51168
rect 7744 50080 8064 51104
rect 7744 50016 7752 50080
rect 7816 50016 7832 50080
rect 7896 50016 7912 50080
rect 7976 50016 7992 50080
rect 8056 50016 8064 50080
rect 7744 48992 8064 50016
rect 7744 48928 7752 48992
rect 7816 48928 7832 48992
rect 7896 48928 7912 48992
rect 7976 48928 7992 48992
rect 8056 48928 8064 48992
rect 7744 47904 8064 48928
rect 7744 47840 7752 47904
rect 7816 47840 7832 47904
rect 7896 47840 7912 47904
rect 7976 47840 7992 47904
rect 8056 47840 8064 47904
rect 7744 46816 8064 47840
rect 7744 46752 7752 46816
rect 7816 46752 7832 46816
rect 7896 46752 7912 46816
rect 7976 46752 7992 46816
rect 8056 46752 8064 46816
rect 7744 45728 8064 46752
rect 7744 45664 7752 45728
rect 7816 45664 7832 45728
rect 7896 45664 7912 45728
rect 7976 45664 7992 45728
rect 8056 45664 8064 45728
rect 7744 44640 8064 45664
rect 7744 44576 7752 44640
rect 7816 44576 7832 44640
rect 7896 44576 7912 44640
rect 7976 44576 7992 44640
rect 8056 44576 8064 44640
rect 7744 43552 8064 44576
rect 7744 43488 7752 43552
rect 7816 43488 7832 43552
rect 7896 43488 7912 43552
rect 7976 43488 7992 43552
rect 8056 43488 8064 43552
rect 7744 42464 8064 43488
rect 7744 42400 7752 42464
rect 7816 42400 7832 42464
rect 7896 42400 7912 42464
rect 7976 42400 7992 42464
rect 8056 42400 8064 42464
rect 7744 41376 8064 42400
rect 7744 41312 7752 41376
rect 7816 41312 7832 41376
rect 7896 41312 7912 41376
rect 7976 41312 7992 41376
rect 8056 41312 8064 41376
rect 7744 40288 8064 41312
rect 7744 40224 7752 40288
rect 7816 40224 7832 40288
rect 7896 40224 7912 40288
rect 7976 40224 7992 40288
rect 8056 40224 8064 40288
rect 7744 39200 8064 40224
rect 7744 39136 7752 39200
rect 7816 39136 7832 39200
rect 7896 39136 7912 39200
rect 7976 39136 7992 39200
rect 8056 39136 8064 39200
rect 7744 38112 8064 39136
rect 7744 38048 7752 38112
rect 7816 38048 7832 38112
rect 7896 38048 7912 38112
rect 7976 38048 7992 38112
rect 8056 38048 8064 38112
rect 7744 37024 8064 38048
rect 7744 36960 7752 37024
rect 7816 36960 7832 37024
rect 7896 36960 7912 37024
rect 7976 36960 7992 37024
rect 8056 36960 8064 37024
rect 7744 35936 8064 36960
rect 7744 35872 7752 35936
rect 7816 35872 7832 35936
rect 7896 35872 7912 35936
rect 7976 35872 7992 35936
rect 8056 35872 8064 35936
rect 7744 34848 8064 35872
rect 7744 34784 7752 34848
rect 7816 34784 7832 34848
rect 7896 34784 7912 34848
rect 7976 34784 7992 34848
rect 8056 34784 8064 34848
rect 7744 33760 8064 34784
rect 7744 33696 7752 33760
rect 7816 33696 7832 33760
rect 7896 33696 7912 33760
rect 7976 33696 7992 33760
rect 8056 33696 8064 33760
rect 7744 32672 8064 33696
rect 7744 32608 7752 32672
rect 7816 32608 7832 32672
rect 7896 32608 7912 32672
rect 7976 32608 7992 32672
rect 8056 32608 8064 32672
rect 7744 31584 8064 32608
rect 7744 31520 7752 31584
rect 7816 31520 7832 31584
rect 7896 31520 7912 31584
rect 7976 31520 7992 31584
rect 8056 31520 8064 31584
rect 7744 30496 8064 31520
rect 7744 30432 7752 30496
rect 7816 30432 7832 30496
rect 7896 30432 7912 30496
rect 7976 30432 7992 30496
rect 8056 30432 8064 30496
rect 7744 29408 8064 30432
rect 7744 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8064 29408
rect 7744 28320 8064 29344
rect 7744 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8064 28320
rect 7744 27232 8064 28256
rect 7744 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8064 27232
rect 7744 26144 8064 27168
rect 7744 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8064 26144
rect 7744 25056 8064 26080
rect 7744 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8064 25056
rect 7744 23968 8064 24992
rect 7744 23904 7752 23968
rect 7816 23904 7832 23968
rect 7896 23904 7912 23968
rect 7976 23904 7992 23968
rect 8056 23904 8064 23968
rect 7744 22880 8064 23904
rect 7744 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8064 22880
rect 7744 21792 8064 22816
rect 7744 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8064 21792
rect 7744 20704 8064 21728
rect 7744 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8064 20704
rect 7744 19616 8064 20640
rect 7744 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8064 19616
rect 7744 18528 8064 19552
rect 7744 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8064 18528
rect 7744 17440 8064 18464
rect 7744 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8064 17440
rect 7744 16352 8064 17376
rect 7744 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8064 16352
rect 7744 15264 8064 16288
rect 7744 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8064 15264
rect 7744 14176 8064 15200
rect 7744 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8064 14176
rect 7744 13088 8064 14112
rect 7744 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8064 13088
rect 7744 12000 8064 13024
rect 7744 11936 7752 12000
rect 7816 11936 7832 12000
rect 7896 11936 7912 12000
rect 7976 11936 7992 12000
rect 8056 11936 8064 12000
rect 7744 10912 8064 11936
rect 7744 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8064 10912
rect 7744 9824 8064 10848
rect 7744 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8064 9824
rect 7744 8736 8064 9760
rect 7744 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8064 8736
rect 7744 7648 8064 8672
rect 7744 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8064 7648
rect 7744 6560 8064 7584
rect 7744 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8064 6560
rect 7744 6206 8064 6496
rect 7744 5970 7786 6206
rect 8022 5970 8064 6206
rect 7744 5472 8064 5970
rect 7744 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8064 5472
rect 7744 4384 8064 5408
rect 7744 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8064 4384
rect 7744 3296 8064 4320
rect 7744 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8064 3296
rect 7744 2208 8064 3232
rect 7744 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8064 2208
rect 7744 1120 8064 2144
rect 7744 1056 7752 1120
rect 7816 1056 7832 1120
rect 7896 1056 7912 1120
rect 7976 1056 7992 1120
rect 8056 1056 8064 1120
rect 7744 -814 8064 1056
rect 7744 -1050 7786 -814
rect 8022 -1050 8064 -814
rect 7744 -1092 8064 -1050
rect 8404 87974 8724 88676
rect 8404 87738 8446 87974
rect 8682 87738 8724 87974
rect 8404 86528 8724 87738
rect 8404 86464 8412 86528
rect 8476 86464 8492 86528
rect 8556 86464 8572 86528
rect 8636 86464 8652 86528
rect 8716 86464 8724 86528
rect 8404 85440 8724 86464
rect 8404 85376 8412 85440
rect 8476 85376 8492 85440
rect 8556 85376 8572 85440
rect 8636 85376 8652 85440
rect 8716 85376 8724 85440
rect 8404 84352 8724 85376
rect 8404 84288 8412 84352
rect 8476 84288 8492 84352
rect 8556 84288 8572 84352
rect 8636 84288 8652 84352
rect 8716 84288 8724 84352
rect 8404 83264 8724 84288
rect 8404 83200 8412 83264
rect 8476 83200 8492 83264
rect 8556 83200 8572 83264
rect 8636 83200 8652 83264
rect 8716 83200 8724 83264
rect 8404 82866 8724 83200
rect 8404 82630 8446 82866
rect 8682 82630 8724 82866
rect 8404 82176 8724 82630
rect 8404 82112 8412 82176
rect 8476 82112 8492 82176
rect 8556 82112 8572 82176
rect 8636 82112 8652 82176
rect 8716 82112 8724 82176
rect 8404 81088 8724 82112
rect 8404 81024 8412 81088
rect 8476 81024 8492 81088
rect 8556 81024 8572 81088
rect 8636 81024 8652 81088
rect 8716 81024 8724 81088
rect 8404 80000 8724 81024
rect 8404 79936 8412 80000
rect 8476 79936 8492 80000
rect 8556 79936 8572 80000
rect 8636 79936 8652 80000
rect 8716 79936 8724 80000
rect 8404 78912 8724 79936
rect 8404 78848 8412 78912
rect 8476 78848 8492 78912
rect 8556 78848 8572 78912
rect 8636 78848 8652 78912
rect 8716 78848 8724 78912
rect 8404 77824 8724 78848
rect 8404 77760 8412 77824
rect 8476 77760 8492 77824
rect 8556 77760 8572 77824
rect 8636 77760 8652 77824
rect 8716 77760 8724 77824
rect 8404 76736 8724 77760
rect 8404 76672 8412 76736
rect 8476 76672 8492 76736
rect 8556 76672 8572 76736
rect 8636 76672 8652 76736
rect 8716 76672 8724 76736
rect 8404 75648 8724 76672
rect 8404 75584 8412 75648
rect 8476 75584 8492 75648
rect 8556 75584 8572 75648
rect 8636 75584 8652 75648
rect 8716 75584 8724 75648
rect 8404 74560 8724 75584
rect 8404 74496 8412 74560
rect 8476 74496 8492 74560
rect 8556 74496 8572 74560
rect 8636 74496 8652 74560
rect 8716 74496 8724 74560
rect 8404 73472 8724 74496
rect 8404 73408 8412 73472
rect 8476 73408 8492 73472
rect 8556 73408 8572 73472
rect 8636 73408 8652 73472
rect 8716 73408 8724 73472
rect 8404 72384 8724 73408
rect 8404 72320 8412 72384
rect 8476 72320 8492 72384
rect 8556 72320 8572 72384
rect 8636 72320 8652 72384
rect 8716 72320 8724 72384
rect 8404 71296 8724 72320
rect 8404 71232 8412 71296
rect 8476 71232 8492 71296
rect 8556 71232 8572 71296
rect 8636 71232 8652 71296
rect 8716 71232 8724 71296
rect 8404 70208 8724 71232
rect 8404 70144 8412 70208
rect 8476 70144 8492 70208
rect 8556 70144 8572 70208
rect 8636 70144 8652 70208
rect 8716 70144 8724 70208
rect 8404 69120 8724 70144
rect 8404 69056 8412 69120
rect 8476 69056 8492 69120
rect 8556 69056 8572 69120
rect 8636 69056 8652 69120
rect 8716 69056 8724 69120
rect 8404 68032 8724 69056
rect 8404 67968 8412 68032
rect 8476 67968 8492 68032
rect 8556 67968 8572 68032
rect 8636 67968 8652 68032
rect 8716 67968 8724 68032
rect 8404 66944 8724 67968
rect 8404 66880 8412 66944
rect 8476 66880 8492 66944
rect 8556 66880 8572 66944
rect 8636 66880 8652 66944
rect 8716 66880 8724 66944
rect 8404 65856 8724 66880
rect 8404 65792 8412 65856
rect 8476 65792 8492 65856
rect 8556 65792 8572 65856
rect 8636 65792 8652 65856
rect 8716 65792 8724 65856
rect 8404 64768 8724 65792
rect 8404 64704 8412 64768
rect 8476 64704 8492 64768
rect 8556 64704 8572 64768
rect 8636 64704 8652 64768
rect 8716 64704 8724 64768
rect 8404 63680 8724 64704
rect 8404 63616 8412 63680
rect 8476 63616 8492 63680
rect 8556 63616 8572 63680
rect 8636 63616 8652 63680
rect 8716 63616 8724 63680
rect 8404 62592 8724 63616
rect 8404 62528 8412 62592
rect 8476 62528 8492 62592
rect 8556 62528 8572 62592
rect 8636 62528 8652 62592
rect 8716 62528 8724 62592
rect 8404 61504 8724 62528
rect 8404 61440 8412 61504
rect 8476 61440 8492 61504
rect 8556 61440 8572 61504
rect 8636 61440 8652 61504
rect 8716 61440 8724 61504
rect 8404 60416 8724 61440
rect 8404 60352 8412 60416
rect 8476 60352 8492 60416
rect 8556 60352 8572 60416
rect 8636 60352 8652 60416
rect 8716 60352 8724 60416
rect 8404 59328 8724 60352
rect 8404 59264 8412 59328
rect 8476 59264 8492 59328
rect 8556 59264 8572 59328
rect 8636 59264 8652 59328
rect 8716 59264 8724 59328
rect 8404 58240 8724 59264
rect 8404 58176 8412 58240
rect 8476 58176 8492 58240
rect 8556 58176 8572 58240
rect 8636 58176 8652 58240
rect 8716 58176 8724 58240
rect 8404 57152 8724 58176
rect 8404 57088 8412 57152
rect 8476 57088 8492 57152
rect 8556 57088 8572 57152
rect 8636 57088 8652 57152
rect 8716 57088 8724 57152
rect 8404 56064 8724 57088
rect 8404 56000 8412 56064
rect 8476 56000 8492 56064
rect 8556 56000 8572 56064
rect 8636 56000 8652 56064
rect 8716 56000 8724 56064
rect 8404 54976 8724 56000
rect 8404 54912 8412 54976
rect 8476 54912 8492 54976
rect 8556 54912 8572 54976
rect 8636 54912 8652 54976
rect 8716 54912 8724 54976
rect 8404 53888 8724 54912
rect 8404 53824 8412 53888
rect 8476 53824 8492 53888
rect 8556 53824 8572 53888
rect 8636 53824 8652 53888
rect 8716 53824 8724 53888
rect 8404 52800 8724 53824
rect 8404 52736 8412 52800
rect 8476 52736 8492 52800
rect 8556 52736 8572 52800
rect 8636 52736 8652 52800
rect 8716 52736 8724 52800
rect 8404 51712 8724 52736
rect 8404 51648 8412 51712
rect 8476 51648 8492 51712
rect 8556 51648 8572 51712
rect 8636 51648 8652 51712
rect 8716 51648 8724 51712
rect 8404 50624 8724 51648
rect 8404 50560 8412 50624
rect 8476 50560 8492 50624
rect 8556 50560 8572 50624
rect 8636 50560 8652 50624
rect 8716 50560 8724 50624
rect 8404 49536 8724 50560
rect 8404 49472 8412 49536
rect 8476 49472 8492 49536
rect 8556 49472 8572 49536
rect 8636 49472 8652 49536
rect 8716 49472 8724 49536
rect 8404 48448 8724 49472
rect 8404 48384 8412 48448
rect 8476 48384 8492 48448
rect 8556 48384 8572 48448
rect 8636 48384 8652 48448
rect 8716 48384 8724 48448
rect 8404 47360 8724 48384
rect 8404 47296 8412 47360
rect 8476 47296 8492 47360
rect 8556 47296 8572 47360
rect 8636 47296 8652 47360
rect 8716 47296 8724 47360
rect 8404 46272 8724 47296
rect 8404 46208 8412 46272
rect 8476 46208 8492 46272
rect 8556 46208 8572 46272
rect 8636 46208 8652 46272
rect 8716 46208 8724 46272
rect 8404 45184 8724 46208
rect 8404 45120 8412 45184
rect 8476 45120 8492 45184
rect 8556 45120 8572 45184
rect 8636 45120 8652 45184
rect 8716 45120 8724 45184
rect 8404 44096 8724 45120
rect 8404 44032 8412 44096
rect 8476 44032 8492 44096
rect 8556 44032 8572 44096
rect 8636 44032 8652 44096
rect 8716 44032 8724 44096
rect 8404 43008 8724 44032
rect 8404 42944 8412 43008
rect 8476 42944 8492 43008
rect 8556 42944 8572 43008
rect 8636 42944 8652 43008
rect 8716 42944 8724 43008
rect 8404 41920 8724 42944
rect 8404 41856 8412 41920
rect 8476 41856 8492 41920
rect 8556 41856 8572 41920
rect 8636 41856 8652 41920
rect 8716 41856 8724 41920
rect 8404 40832 8724 41856
rect 8404 40768 8412 40832
rect 8476 40768 8492 40832
rect 8556 40768 8572 40832
rect 8636 40768 8652 40832
rect 8716 40768 8724 40832
rect 8404 39744 8724 40768
rect 8404 39680 8412 39744
rect 8476 39680 8492 39744
rect 8556 39680 8572 39744
rect 8636 39680 8652 39744
rect 8716 39680 8724 39744
rect 8404 38656 8724 39680
rect 8404 38592 8412 38656
rect 8476 38592 8492 38656
rect 8556 38592 8572 38656
rect 8636 38592 8652 38656
rect 8716 38592 8724 38656
rect 8404 37568 8724 38592
rect 8404 37504 8412 37568
rect 8476 37504 8492 37568
rect 8556 37504 8572 37568
rect 8636 37504 8652 37568
rect 8716 37504 8724 37568
rect 8404 36480 8724 37504
rect 8404 36416 8412 36480
rect 8476 36416 8492 36480
rect 8556 36416 8572 36480
rect 8636 36416 8652 36480
rect 8716 36416 8724 36480
rect 8404 35392 8724 36416
rect 8404 35328 8412 35392
rect 8476 35328 8492 35392
rect 8556 35328 8572 35392
rect 8636 35328 8652 35392
rect 8716 35328 8724 35392
rect 8404 34304 8724 35328
rect 8404 34240 8412 34304
rect 8476 34240 8492 34304
rect 8556 34240 8572 34304
rect 8636 34240 8652 34304
rect 8716 34240 8724 34304
rect 8404 33216 8724 34240
rect 8404 33152 8412 33216
rect 8476 33152 8492 33216
rect 8556 33152 8572 33216
rect 8636 33152 8652 33216
rect 8716 33152 8724 33216
rect 8404 32128 8724 33152
rect 8404 32064 8412 32128
rect 8476 32064 8492 32128
rect 8556 32064 8572 32128
rect 8636 32064 8652 32128
rect 8716 32064 8724 32128
rect 8404 31040 8724 32064
rect 8404 30976 8412 31040
rect 8476 30976 8492 31040
rect 8556 30976 8572 31040
rect 8636 30976 8652 31040
rect 8716 30976 8724 31040
rect 8404 29952 8724 30976
rect 8404 29888 8412 29952
rect 8476 29888 8492 29952
rect 8556 29888 8572 29952
rect 8636 29888 8652 29952
rect 8716 29888 8724 29952
rect 8404 28864 8724 29888
rect 8404 28800 8412 28864
rect 8476 28800 8492 28864
rect 8556 28800 8572 28864
rect 8636 28800 8652 28864
rect 8716 28800 8724 28864
rect 8404 27776 8724 28800
rect 8404 27712 8412 27776
rect 8476 27712 8492 27776
rect 8556 27712 8572 27776
rect 8636 27712 8652 27776
rect 8716 27712 8724 27776
rect 8404 26688 8724 27712
rect 8404 26624 8412 26688
rect 8476 26624 8492 26688
rect 8556 26624 8572 26688
rect 8636 26624 8652 26688
rect 8716 26624 8724 26688
rect 8404 25600 8724 26624
rect 8404 25536 8412 25600
rect 8476 25536 8492 25600
rect 8556 25536 8572 25600
rect 8636 25536 8652 25600
rect 8716 25536 8724 25600
rect 8404 24512 8724 25536
rect 8404 24448 8412 24512
rect 8476 24448 8492 24512
rect 8556 24448 8572 24512
rect 8636 24448 8652 24512
rect 8716 24448 8724 24512
rect 8404 23424 8724 24448
rect 8404 23360 8412 23424
rect 8476 23360 8492 23424
rect 8556 23360 8572 23424
rect 8636 23360 8652 23424
rect 8716 23360 8724 23424
rect 8404 22336 8724 23360
rect 8404 22272 8412 22336
rect 8476 22272 8492 22336
rect 8556 22272 8572 22336
rect 8636 22272 8652 22336
rect 8716 22272 8724 22336
rect 8404 21248 8724 22272
rect 8404 21184 8412 21248
rect 8476 21184 8492 21248
rect 8556 21184 8572 21248
rect 8636 21184 8652 21248
rect 8716 21184 8724 21248
rect 8404 20160 8724 21184
rect 8404 20096 8412 20160
rect 8476 20096 8492 20160
rect 8556 20096 8572 20160
rect 8636 20096 8652 20160
rect 8716 20096 8724 20160
rect 8404 19072 8724 20096
rect 8404 19008 8412 19072
rect 8476 19008 8492 19072
rect 8556 19008 8572 19072
rect 8636 19008 8652 19072
rect 8716 19008 8724 19072
rect 8404 17984 8724 19008
rect 8404 17920 8412 17984
rect 8476 17920 8492 17984
rect 8556 17920 8572 17984
rect 8636 17920 8652 17984
rect 8716 17920 8724 17984
rect 8404 16896 8724 17920
rect 8404 16832 8412 16896
rect 8476 16832 8492 16896
rect 8556 16832 8572 16896
rect 8636 16832 8652 16896
rect 8716 16832 8724 16896
rect 8404 15808 8724 16832
rect 8404 15744 8412 15808
rect 8476 15744 8492 15808
rect 8556 15744 8572 15808
rect 8636 15744 8652 15808
rect 8716 15744 8724 15808
rect 8404 14720 8724 15744
rect 8404 14656 8412 14720
rect 8476 14656 8492 14720
rect 8556 14656 8572 14720
rect 8636 14656 8652 14720
rect 8716 14656 8724 14720
rect 8404 13632 8724 14656
rect 8404 13568 8412 13632
rect 8476 13568 8492 13632
rect 8556 13568 8572 13632
rect 8636 13568 8652 13632
rect 8716 13568 8724 13632
rect 8404 12544 8724 13568
rect 8404 12480 8412 12544
rect 8476 12480 8492 12544
rect 8556 12480 8572 12544
rect 8636 12480 8652 12544
rect 8716 12480 8724 12544
rect 8404 11456 8724 12480
rect 8404 11392 8412 11456
rect 8476 11392 8492 11456
rect 8556 11392 8572 11456
rect 8636 11392 8652 11456
rect 8716 11392 8724 11456
rect 8404 10368 8724 11392
rect 8404 10304 8412 10368
rect 8476 10304 8492 10368
rect 8556 10304 8572 10368
rect 8636 10304 8652 10368
rect 8716 10304 8724 10368
rect 8404 9280 8724 10304
rect 8404 9216 8412 9280
rect 8476 9216 8492 9280
rect 8556 9216 8572 9280
rect 8636 9216 8652 9280
rect 8716 9216 8724 9280
rect 8404 8192 8724 9216
rect 8404 8128 8412 8192
rect 8476 8128 8492 8192
rect 8556 8128 8572 8192
rect 8636 8128 8652 8192
rect 8716 8128 8724 8192
rect 8404 7104 8724 8128
rect 8404 7040 8412 7104
rect 8476 7040 8492 7104
rect 8556 7040 8572 7104
rect 8636 7040 8652 7104
rect 8716 7040 8724 7104
rect 8404 6866 8724 7040
rect 8404 6630 8446 6866
rect 8682 6630 8724 6866
rect 8404 6016 8724 6630
rect 8404 5952 8412 6016
rect 8476 5952 8492 6016
rect 8556 5952 8572 6016
rect 8636 5952 8652 6016
rect 8716 5952 8724 6016
rect 8404 4928 8724 5952
rect 8404 4864 8412 4928
rect 8476 4864 8492 4928
rect 8556 4864 8572 4928
rect 8636 4864 8652 4928
rect 8716 4864 8724 4928
rect 8404 3840 8724 4864
rect 8404 3776 8412 3840
rect 8476 3776 8492 3840
rect 8556 3776 8572 3840
rect 8636 3776 8652 3840
rect 8716 3776 8724 3840
rect 8404 2752 8724 3776
rect 8404 2688 8412 2752
rect 8476 2688 8492 2752
rect 8556 2688 8572 2752
rect 8636 2688 8652 2752
rect 8716 2688 8724 2752
rect 8404 1664 8724 2688
rect 8404 1600 8412 1664
rect 8476 1600 8492 1664
rect 8556 1600 8572 1664
rect 8636 1600 8652 1664
rect 8716 1600 8724 1664
rect 8404 -154 8724 1600
rect 8404 -390 8446 -154
rect 8682 -390 8724 -154
rect 8404 -1092 8724 -390
rect 9344 88634 9664 88676
rect 9344 88398 9386 88634
rect 9622 88398 9664 88634
rect 9344 85984 9664 88398
rect 9344 85920 9352 85984
rect 9416 85920 9432 85984
rect 9496 85920 9512 85984
rect 9576 85920 9592 85984
rect 9656 85920 9664 85984
rect 9344 84896 9664 85920
rect 10004 87974 10324 88676
rect 10004 87738 10046 87974
rect 10282 87738 10324 87974
rect 10004 86528 10324 87738
rect 10004 86464 10012 86528
rect 10076 86464 10092 86528
rect 10156 86464 10172 86528
rect 10236 86464 10252 86528
rect 10316 86464 10324 86528
rect 10004 85496 10324 86464
rect 10944 88634 11264 88676
rect 10944 88398 10986 88634
rect 11222 88398 11264 88634
rect 10944 85984 11264 88398
rect 11604 87974 11924 88676
rect 11604 87738 11646 87974
rect 11882 87738 11924 87974
rect 11604 86528 11924 87738
rect 11604 86464 11612 86528
rect 11676 86464 11692 86528
rect 11756 86464 11772 86528
rect 11836 86464 11852 86528
rect 11916 86464 11924 86528
rect 11467 86188 11533 86189
rect 11467 86124 11468 86188
rect 11532 86124 11533 86188
rect 11467 86123 11533 86124
rect 10944 85920 10952 85984
rect 11016 85920 11032 85984
rect 11096 85920 11112 85984
rect 11176 85920 11192 85984
rect 11256 85920 11264 85984
rect 10944 85496 11264 85920
rect 9344 84832 9352 84896
rect 9416 84832 9432 84896
rect 9496 84832 9512 84896
rect 9576 84832 9592 84896
rect 9656 84832 9664 84896
rect 9344 83808 9664 84832
rect 10915 84284 10981 84285
rect 10915 84220 10916 84284
rect 10980 84220 10981 84284
rect 10915 84219 10981 84220
rect 9344 83744 9352 83808
rect 9416 83744 9432 83808
rect 9496 83744 9512 83808
rect 9576 83744 9592 83808
rect 9656 83744 9664 83808
rect 9344 82720 9664 83744
rect 9344 82656 9352 82720
rect 9416 82656 9432 82720
rect 9496 82656 9512 82720
rect 9576 82656 9592 82720
rect 9656 82656 9664 82720
rect 9344 82206 9664 82656
rect 9344 81970 9386 82206
rect 9622 81970 9664 82206
rect 9344 81632 9664 81970
rect 9344 81568 9352 81632
rect 9416 81568 9432 81632
rect 9496 81568 9512 81632
rect 9576 81568 9592 81632
rect 9656 81568 9664 81632
rect 9344 80544 9664 81568
rect 9344 80480 9352 80544
rect 9416 80480 9432 80544
rect 9496 80480 9512 80544
rect 9576 80480 9592 80544
rect 9656 80480 9664 80544
rect 9344 79456 9664 80480
rect 9344 79392 9352 79456
rect 9416 79392 9432 79456
rect 9496 79392 9512 79456
rect 9576 79392 9592 79456
rect 9656 79392 9664 79456
rect 9344 78368 9664 79392
rect 9344 78304 9352 78368
rect 9416 78304 9432 78368
rect 9496 78304 9512 78368
rect 9576 78304 9592 78368
rect 9656 78304 9664 78368
rect 9344 77280 9664 78304
rect 9344 77216 9352 77280
rect 9416 77216 9432 77280
rect 9496 77216 9512 77280
rect 9576 77216 9592 77280
rect 9656 77216 9664 77280
rect 9344 76192 9664 77216
rect 9344 76128 9352 76192
rect 9416 76128 9432 76192
rect 9496 76128 9512 76192
rect 9576 76128 9592 76192
rect 9656 76128 9664 76192
rect 9344 75104 9664 76128
rect 9344 75040 9352 75104
rect 9416 75040 9432 75104
rect 9496 75040 9512 75104
rect 9576 75040 9592 75104
rect 9656 75040 9664 75104
rect 9344 74016 9664 75040
rect 10918 74357 10978 84219
rect 10915 74356 10981 74357
rect 10915 74292 10916 74356
rect 10980 74292 10981 74356
rect 10915 74291 10981 74292
rect 9344 73952 9352 74016
rect 9416 73952 9432 74016
rect 9496 73952 9512 74016
rect 9576 73952 9592 74016
rect 9656 73952 9664 74016
rect 9344 72928 9664 73952
rect 9344 72864 9352 72928
rect 9416 72864 9432 72928
rect 9496 72864 9512 72928
rect 9576 72864 9592 72928
rect 9656 72864 9664 72928
rect 9344 71840 9664 72864
rect 9344 71776 9352 71840
rect 9416 71776 9432 71840
rect 9496 71776 9512 71840
rect 9576 71776 9592 71840
rect 9656 71776 9664 71840
rect 9344 70752 9664 71776
rect 9344 70688 9352 70752
rect 9416 70688 9432 70752
rect 9496 70688 9512 70752
rect 9576 70688 9592 70752
rect 9656 70688 9664 70752
rect 9344 69664 9664 70688
rect 10547 69868 10613 69869
rect 10547 69804 10548 69868
rect 10612 69804 10613 69868
rect 10547 69803 10613 69804
rect 9344 69600 9352 69664
rect 9416 69600 9432 69664
rect 9496 69600 9512 69664
rect 9576 69600 9592 69664
rect 9656 69600 9664 69664
rect 9344 68576 9664 69600
rect 9344 68512 9352 68576
rect 9416 68512 9432 68576
rect 9496 68512 9512 68576
rect 9576 68512 9592 68576
rect 9656 68512 9664 68576
rect 9344 67488 9664 68512
rect 9344 67424 9352 67488
rect 9416 67424 9432 67488
rect 9496 67424 9512 67488
rect 9576 67424 9592 67488
rect 9656 67424 9664 67488
rect 9344 66400 9664 67424
rect 9344 66336 9352 66400
rect 9416 66336 9432 66400
rect 9496 66336 9512 66400
rect 9576 66336 9592 66400
rect 9656 66336 9664 66400
rect 9344 65312 9664 66336
rect 9344 65248 9352 65312
rect 9416 65248 9432 65312
rect 9496 65248 9512 65312
rect 9576 65248 9592 65312
rect 9656 65248 9664 65312
rect 9344 64224 9664 65248
rect 9344 64160 9352 64224
rect 9416 64160 9432 64224
rect 9496 64160 9512 64224
rect 9576 64160 9592 64224
rect 9656 64160 9664 64224
rect 9344 63136 9664 64160
rect 9344 63072 9352 63136
rect 9416 63072 9432 63136
rect 9496 63072 9512 63136
rect 9576 63072 9592 63136
rect 9656 63072 9664 63136
rect 9344 62048 9664 63072
rect 9344 61984 9352 62048
rect 9416 61984 9432 62048
rect 9496 61984 9512 62048
rect 9576 61984 9592 62048
rect 9656 61984 9664 62048
rect 9344 60960 9664 61984
rect 9344 60896 9352 60960
rect 9416 60896 9432 60960
rect 9496 60896 9512 60960
rect 9576 60896 9592 60960
rect 9656 60896 9664 60960
rect 9344 59872 9664 60896
rect 9344 59808 9352 59872
rect 9416 59808 9432 59872
rect 9496 59808 9512 59872
rect 9576 59808 9592 59872
rect 9656 59808 9664 59872
rect 9344 58784 9664 59808
rect 9344 58720 9352 58784
rect 9416 58720 9432 58784
rect 9496 58720 9512 58784
rect 9576 58720 9592 58784
rect 9656 58720 9664 58784
rect 9344 57696 9664 58720
rect 9344 57632 9352 57696
rect 9416 57632 9432 57696
rect 9496 57632 9512 57696
rect 9576 57632 9592 57696
rect 9656 57632 9664 57696
rect 9344 56608 9664 57632
rect 9344 56544 9352 56608
rect 9416 56544 9432 56608
rect 9496 56544 9512 56608
rect 9576 56544 9592 56608
rect 9656 56544 9664 56608
rect 9344 55520 9664 56544
rect 9344 55456 9352 55520
rect 9416 55456 9432 55520
rect 9496 55456 9512 55520
rect 9576 55456 9592 55520
rect 9656 55456 9664 55520
rect 9344 54432 9664 55456
rect 9344 54368 9352 54432
rect 9416 54368 9432 54432
rect 9496 54368 9512 54432
rect 9576 54368 9592 54432
rect 9656 54368 9664 54432
rect 9344 53344 9664 54368
rect 9344 53280 9352 53344
rect 9416 53280 9432 53344
rect 9496 53280 9512 53344
rect 9576 53280 9592 53344
rect 9656 53280 9664 53344
rect 9344 52256 9664 53280
rect 9344 52192 9352 52256
rect 9416 52192 9432 52256
rect 9496 52192 9512 52256
rect 9576 52192 9592 52256
rect 9656 52192 9664 52256
rect 9344 51168 9664 52192
rect 9344 51104 9352 51168
rect 9416 51104 9432 51168
rect 9496 51104 9512 51168
rect 9576 51104 9592 51168
rect 9656 51104 9664 51168
rect 9344 50080 9664 51104
rect 9344 50016 9352 50080
rect 9416 50016 9432 50080
rect 9496 50016 9512 50080
rect 9576 50016 9592 50080
rect 9656 50016 9664 50080
rect 9344 48992 9664 50016
rect 9344 48928 9352 48992
rect 9416 48928 9432 48992
rect 9496 48928 9512 48992
rect 9576 48928 9592 48992
rect 9656 48928 9664 48992
rect 9344 47904 9664 48928
rect 9344 47840 9352 47904
rect 9416 47840 9432 47904
rect 9496 47840 9512 47904
rect 9576 47840 9592 47904
rect 9656 47840 9664 47904
rect 9344 46816 9664 47840
rect 9344 46752 9352 46816
rect 9416 46752 9432 46816
rect 9496 46752 9512 46816
rect 9576 46752 9592 46816
rect 9656 46752 9664 46816
rect 9344 45728 9664 46752
rect 9344 45664 9352 45728
rect 9416 45664 9432 45728
rect 9496 45664 9512 45728
rect 9576 45664 9592 45728
rect 9656 45664 9664 45728
rect 9344 44640 9664 45664
rect 9344 44576 9352 44640
rect 9416 44576 9432 44640
rect 9496 44576 9512 44640
rect 9576 44576 9592 44640
rect 9656 44576 9664 44640
rect 9344 43552 9664 44576
rect 9344 43488 9352 43552
rect 9416 43488 9432 43552
rect 9496 43488 9512 43552
rect 9576 43488 9592 43552
rect 9656 43488 9664 43552
rect 9344 42464 9664 43488
rect 9344 42400 9352 42464
rect 9416 42400 9432 42464
rect 9496 42400 9512 42464
rect 9576 42400 9592 42464
rect 9656 42400 9664 42464
rect 9344 41376 9664 42400
rect 9344 41312 9352 41376
rect 9416 41312 9432 41376
rect 9496 41312 9512 41376
rect 9576 41312 9592 41376
rect 9656 41312 9664 41376
rect 9344 40288 9664 41312
rect 9344 40224 9352 40288
rect 9416 40224 9432 40288
rect 9496 40224 9512 40288
rect 9576 40224 9592 40288
rect 9656 40224 9664 40288
rect 9344 39200 9664 40224
rect 9344 39136 9352 39200
rect 9416 39136 9432 39200
rect 9496 39136 9512 39200
rect 9576 39136 9592 39200
rect 9656 39136 9664 39200
rect 9344 38112 9664 39136
rect 10550 38453 10610 69803
rect 11099 69460 11165 69461
rect 11099 69396 11100 69460
rect 11164 69396 11165 69460
rect 11099 69395 11165 69396
rect 11102 39949 11162 69395
rect 11470 68917 11530 86123
rect 11604 85496 11924 86464
rect 12544 88634 12864 88676
rect 12544 88398 12586 88634
rect 12822 88398 12864 88634
rect 12544 85984 12864 88398
rect 12544 85920 12552 85984
rect 12616 85920 12632 85984
rect 12696 85920 12712 85984
rect 12776 85920 12792 85984
rect 12856 85920 12864 85984
rect 12544 85496 12864 85920
rect 13204 87974 13524 88676
rect 13204 87738 13246 87974
rect 13482 87738 13524 87974
rect 13204 86528 13524 87738
rect 13204 86464 13212 86528
rect 13276 86464 13292 86528
rect 13356 86464 13372 86528
rect 13436 86464 13452 86528
rect 13516 86464 13524 86528
rect 13204 85496 13524 86464
rect 14144 88634 14464 88676
rect 14144 88398 14186 88634
rect 14422 88398 14464 88634
rect 14144 85984 14464 88398
rect 14144 85920 14152 85984
rect 14216 85920 14232 85984
rect 14296 85920 14312 85984
rect 14376 85920 14392 85984
rect 14456 85920 14464 85984
rect 14144 85496 14464 85920
rect 14804 87974 15124 88676
rect 14804 87738 14846 87974
rect 15082 87738 15124 87974
rect 14804 86528 15124 87738
rect 14804 86464 14812 86528
rect 14876 86464 14892 86528
rect 14956 86464 14972 86528
rect 15036 86464 15052 86528
rect 15116 86464 15124 86528
rect 14804 85496 15124 86464
rect 15744 88634 16064 88676
rect 15744 88398 15786 88634
rect 16022 88398 16064 88634
rect 15744 85984 16064 88398
rect 15744 85920 15752 85984
rect 15816 85920 15832 85984
rect 15896 85920 15912 85984
rect 15976 85920 15992 85984
rect 16056 85920 16064 85984
rect 15744 85496 16064 85920
rect 16404 87974 16724 88676
rect 16404 87738 16446 87974
rect 16682 87738 16724 87974
rect 16404 86528 16724 87738
rect 16404 86464 16412 86528
rect 16476 86464 16492 86528
rect 16556 86464 16572 86528
rect 16636 86464 16652 86528
rect 16716 86464 16724 86528
rect 16404 85496 16724 86464
rect 17344 88634 17664 88676
rect 17344 88398 17386 88634
rect 17622 88398 17664 88634
rect 17344 85984 17664 88398
rect 17344 85920 17352 85984
rect 17416 85920 17432 85984
rect 17496 85920 17512 85984
rect 17576 85920 17592 85984
rect 17656 85920 17664 85984
rect 17344 85496 17664 85920
rect 18004 87974 18324 88676
rect 18004 87738 18046 87974
rect 18282 87738 18324 87974
rect 18004 86528 18324 87738
rect 18004 86464 18012 86528
rect 18076 86464 18092 86528
rect 18156 86464 18172 86528
rect 18236 86464 18252 86528
rect 18316 86464 18324 86528
rect 18004 85496 18324 86464
rect 18944 88634 19264 88676
rect 18944 88398 18986 88634
rect 19222 88398 19264 88634
rect 18944 85984 19264 88398
rect 18944 85920 18952 85984
rect 19016 85920 19032 85984
rect 19096 85920 19112 85984
rect 19176 85920 19192 85984
rect 19256 85920 19264 85984
rect 18944 85496 19264 85920
rect 19604 87974 19924 88676
rect 19604 87738 19646 87974
rect 19882 87738 19924 87974
rect 19604 86528 19924 87738
rect 19604 86464 19612 86528
rect 19676 86464 19692 86528
rect 19756 86464 19772 86528
rect 19836 86464 19852 86528
rect 19916 86464 19924 86528
rect 19604 85496 19924 86464
rect 20544 88634 20864 88676
rect 20544 88398 20586 88634
rect 20822 88398 20864 88634
rect 20544 85984 20864 88398
rect 20544 85920 20552 85984
rect 20616 85920 20632 85984
rect 20696 85920 20712 85984
rect 20776 85920 20792 85984
rect 20856 85920 20864 85984
rect 20544 85496 20864 85920
rect 21204 87974 21524 88676
rect 21204 87738 21246 87974
rect 21482 87738 21524 87974
rect 21204 86528 21524 87738
rect 21204 86464 21212 86528
rect 21276 86464 21292 86528
rect 21356 86464 21372 86528
rect 21436 86464 21452 86528
rect 21516 86464 21524 86528
rect 21204 85496 21524 86464
rect 22144 88634 22464 88676
rect 22144 88398 22186 88634
rect 22422 88398 22464 88634
rect 22144 85984 22464 88398
rect 22144 85920 22152 85984
rect 22216 85920 22232 85984
rect 22296 85920 22312 85984
rect 22376 85920 22392 85984
rect 22456 85920 22464 85984
rect 22144 85496 22464 85920
rect 22804 87974 23124 88676
rect 22804 87738 22846 87974
rect 23082 87738 23124 87974
rect 22804 86528 23124 87738
rect 22804 86464 22812 86528
rect 22876 86464 22892 86528
rect 22956 86464 22972 86528
rect 23036 86464 23052 86528
rect 23116 86464 23124 86528
rect 22804 85496 23124 86464
rect 23744 88634 24064 88676
rect 23744 88398 23786 88634
rect 24022 88398 24064 88634
rect 23744 85984 24064 88398
rect 23744 85920 23752 85984
rect 23816 85920 23832 85984
rect 23896 85920 23912 85984
rect 23976 85920 23992 85984
rect 24056 85920 24064 85984
rect 23744 85496 24064 85920
rect 24404 87974 24724 88676
rect 24404 87738 24446 87974
rect 24682 87738 24724 87974
rect 24404 86528 24724 87738
rect 24404 86464 24412 86528
rect 24476 86464 24492 86528
rect 24556 86464 24572 86528
rect 24636 86464 24652 86528
rect 24716 86464 24724 86528
rect 24404 85496 24724 86464
rect 25344 88634 25664 88676
rect 25344 88398 25386 88634
rect 25622 88398 25664 88634
rect 25344 85984 25664 88398
rect 25344 85920 25352 85984
rect 25416 85920 25432 85984
rect 25496 85920 25512 85984
rect 25576 85920 25592 85984
rect 25656 85920 25664 85984
rect 25344 85496 25664 85920
rect 26004 87974 26324 88676
rect 26004 87738 26046 87974
rect 26282 87738 26324 87974
rect 26004 86528 26324 87738
rect 26004 86464 26012 86528
rect 26076 86464 26092 86528
rect 26156 86464 26172 86528
rect 26236 86464 26252 86528
rect 26316 86464 26324 86528
rect 26004 85496 26324 86464
rect 26944 88634 27264 88676
rect 26944 88398 26986 88634
rect 27222 88398 27264 88634
rect 26944 85984 27264 88398
rect 26944 85920 26952 85984
rect 27016 85920 27032 85984
rect 27096 85920 27112 85984
rect 27176 85920 27192 85984
rect 27256 85920 27264 85984
rect 26944 85496 27264 85920
rect 27604 87974 27924 88676
rect 27604 87738 27646 87974
rect 27882 87738 27924 87974
rect 27604 86528 27924 87738
rect 27604 86464 27612 86528
rect 27676 86464 27692 86528
rect 27756 86464 27772 86528
rect 27836 86464 27852 86528
rect 27916 86464 27924 86528
rect 27604 85496 27924 86464
rect 28544 88634 28864 88676
rect 28544 88398 28586 88634
rect 28822 88398 28864 88634
rect 28544 85984 28864 88398
rect 28544 85920 28552 85984
rect 28616 85920 28632 85984
rect 28696 85920 28712 85984
rect 28776 85920 28792 85984
rect 28856 85920 28864 85984
rect 28544 85496 28864 85920
rect 29204 87974 29524 88676
rect 29204 87738 29246 87974
rect 29482 87738 29524 87974
rect 29204 86528 29524 87738
rect 29204 86464 29212 86528
rect 29276 86464 29292 86528
rect 29356 86464 29372 86528
rect 29436 86464 29452 86528
rect 29516 86464 29524 86528
rect 29204 85496 29524 86464
rect 30144 88634 30464 88676
rect 30144 88398 30186 88634
rect 30422 88398 30464 88634
rect 30144 85984 30464 88398
rect 30144 85920 30152 85984
rect 30216 85920 30232 85984
rect 30296 85920 30312 85984
rect 30376 85920 30392 85984
rect 30456 85920 30464 85984
rect 30144 85496 30464 85920
rect 30804 87974 31124 88676
rect 30804 87738 30846 87974
rect 31082 87738 31124 87974
rect 30804 86528 31124 87738
rect 30804 86464 30812 86528
rect 30876 86464 30892 86528
rect 30956 86464 30972 86528
rect 31036 86464 31052 86528
rect 31116 86464 31124 86528
rect 30804 85496 31124 86464
rect 31744 88634 32064 88676
rect 31744 88398 31786 88634
rect 32022 88398 32064 88634
rect 31744 85984 32064 88398
rect 31744 85920 31752 85984
rect 31816 85920 31832 85984
rect 31896 85920 31912 85984
rect 31976 85920 31992 85984
rect 32056 85920 32064 85984
rect 31744 85496 32064 85920
rect 32404 87974 32724 88676
rect 32404 87738 32446 87974
rect 32682 87738 32724 87974
rect 32404 86528 32724 87738
rect 32404 86464 32412 86528
rect 32476 86464 32492 86528
rect 32556 86464 32572 86528
rect 32636 86464 32652 86528
rect 32716 86464 32724 86528
rect 32404 85496 32724 86464
rect 33344 88634 33664 88676
rect 33344 88398 33386 88634
rect 33622 88398 33664 88634
rect 33344 85984 33664 88398
rect 33344 85920 33352 85984
rect 33416 85920 33432 85984
rect 33496 85920 33512 85984
rect 33576 85920 33592 85984
rect 33656 85920 33664 85984
rect 33344 85496 33664 85920
rect 34004 87974 34324 88676
rect 34004 87738 34046 87974
rect 34282 87738 34324 87974
rect 34004 86528 34324 87738
rect 34004 86464 34012 86528
rect 34076 86464 34092 86528
rect 34156 86464 34172 86528
rect 34236 86464 34252 86528
rect 34316 86464 34324 86528
rect 34004 85496 34324 86464
rect 34944 88634 35264 88676
rect 34944 88398 34986 88634
rect 35222 88398 35264 88634
rect 34944 85984 35264 88398
rect 34944 85920 34952 85984
rect 35016 85920 35032 85984
rect 35096 85920 35112 85984
rect 35176 85920 35192 85984
rect 35256 85920 35264 85984
rect 34944 85496 35264 85920
rect 35604 87974 35924 88676
rect 35604 87738 35646 87974
rect 35882 87738 35924 87974
rect 35604 86528 35924 87738
rect 35604 86464 35612 86528
rect 35676 86464 35692 86528
rect 35756 86464 35772 86528
rect 35836 86464 35852 86528
rect 35916 86464 35924 86528
rect 35604 85496 35924 86464
rect 36544 88634 36864 88676
rect 36544 88398 36586 88634
rect 36822 88398 36864 88634
rect 36544 85984 36864 88398
rect 36544 85920 36552 85984
rect 36616 85920 36632 85984
rect 36696 85920 36712 85984
rect 36776 85920 36792 85984
rect 36856 85920 36864 85984
rect 36544 85496 36864 85920
rect 37204 87974 37524 88676
rect 37204 87738 37246 87974
rect 37482 87738 37524 87974
rect 37204 86528 37524 87738
rect 37204 86464 37212 86528
rect 37276 86464 37292 86528
rect 37356 86464 37372 86528
rect 37436 86464 37452 86528
rect 37516 86464 37524 86528
rect 37204 85496 37524 86464
rect 38144 88634 38464 88676
rect 38144 88398 38186 88634
rect 38422 88398 38464 88634
rect 38144 85984 38464 88398
rect 38144 85920 38152 85984
rect 38216 85920 38232 85984
rect 38296 85920 38312 85984
rect 38376 85920 38392 85984
rect 38456 85920 38464 85984
rect 38144 85496 38464 85920
rect 38804 87974 39124 88676
rect 38804 87738 38846 87974
rect 39082 87738 39124 87974
rect 38804 86528 39124 87738
rect 38804 86464 38812 86528
rect 38876 86464 38892 86528
rect 38956 86464 38972 86528
rect 39036 86464 39052 86528
rect 39116 86464 39124 86528
rect 38804 85496 39124 86464
rect 39744 88634 40064 88676
rect 39744 88398 39786 88634
rect 40022 88398 40064 88634
rect 39744 85984 40064 88398
rect 39744 85920 39752 85984
rect 39816 85920 39832 85984
rect 39896 85920 39912 85984
rect 39976 85920 39992 85984
rect 40056 85920 40064 85984
rect 39744 85620 40064 85920
rect 40404 87974 40724 88676
rect 40404 87738 40446 87974
rect 40682 87738 40724 87974
rect 40404 86528 40724 87738
rect 40404 86464 40412 86528
rect 40476 86464 40492 86528
rect 40556 86464 40572 86528
rect 40636 86464 40652 86528
rect 40716 86464 40724 86528
rect 40171 85644 40237 85645
rect 40171 85580 40172 85644
rect 40236 85580 40237 85644
rect 40171 85579 40237 85580
rect 40174 84010 40234 85579
rect 40404 85496 40724 86464
rect 41344 88634 41664 88676
rect 41344 88398 41386 88634
rect 41622 88398 41664 88634
rect 41344 85984 41664 88398
rect 41344 85920 41352 85984
rect 41416 85920 41432 85984
rect 41496 85920 41512 85984
rect 41576 85920 41592 85984
rect 41656 85920 41664 85984
rect 41344 85620 41664 85920
rect 42004 87974 42324 88676
rect 42004 87738 42046 87974
rect 42282 87738 42324 87974
rect 42004 86528 42324 87738
rect 42004 86464 42012 86528
rect 42076 86464 42092 86528
rect 42156 86464 42172 86528
rect 42236 86464 42252 86528
rect 42316 86464 42324 86528
rect 41827 85644 41893 85645
rect 41827 85580 41828 85644
rect 41892 85580 41893 85644
rect 41827 85579 41893 85580
rect 41830 84010 41890 85579
rect 42004 85496 42324 86464
rect 42944 88634 43264 88676
rect 42944 88398 42986 88634
rect 43222 88398 43264 88634
rect 42944 85984 43264 88398
rect 42944 85920 42952 85984
rect 43016 85920 43032 85984
rect 43096 85920 43112 85984
rect 43176 85920 43192 85984
rect 43256 85920 43264 85984
rect 42944 85496 43264 85920
rect 43604 87974 43924 88676
rect 43604 87738 43646 87974
rect 43882 87738 43924 87974
rect 43604 86528 43924 87738
rect 43604 86464 43612 86528
rect 43676 86464 43692 86528
rect 43756 86464 43772 86528
rect 43836 86464 43852 86528
rect 43916 86464 43924 86528
rect 43604 85620 43924 86464
rect 44544 88634 44864 88676
rect 44544 88398 44586 88634
rect 44822 88398 44864 88634
rect 44544 85984 44864 88398
rect 44544 85920 44552 85984
rect 44616 85920 44632 85984
rect 44696 85920 44712 85984
rect 44776 85920 44792 85984
rect 44856 85920 44864 85984
rect 44035 85644 44101 85645
rect 44035 85580 44036 85644
rect 44100 85580 44101 85644
rect 44035 85579 44101 85580
rect 42563 84420 42629 84421
rect 42563 84356 42564 84420
rect 42628 84356 42629 84420
rect 42563 84355 42629 84356
rect 40160 83950 40234 84010
rect 41520 83950 41890 84010
rect 42566 84010 42626 84355
rect 44038 84010 44098 85579
rect 44544 85496 44864 85920
rect 45204 87974 45524 88676
rect 45204 87738 45246 87974
rect 45482 87738 45524 87974
rect 45204 86528 45524 87738
rect 45204 86464 45212 86528
rect 45276 86464 45292 86528
rect 45356 86464 45372 86528
rect 45436 86464 45452 86528
rect 45516 86464 45524 86528
rect 45204 85620 45524 86464
rect 46144 88634 46464 88676
rect 46144 88398 46186 88634
rect 46422 88398 46464 88634
rect 46144 85984 46464 88398
rect 46144 85920 46152 85984
rect 46216 85920 46232 85984
rect 46296 85920 46312 85984
rect 46376 85920 46392 85984
rect 46456 85920 46464 85984
rect 46144 85620 46464 85920
rect 46804 87974 47124 88676
rect 46804 87738 46846 87974
rect 47082 87738 47124 87974
rect 46804 86528 47124 87738
rect 46804 86464 46812 86528
rect 46876 86464 46892 86528
rect 46956 86464 46972 86528
rect 47036 86464 47052 86528
rect 47116 86464 47124 86528
rect 46611 85644 46677 85645
rect 46611 85580 46612 85644
rect 46676 85580 46677 85644
rect 46611 85579 46677 85580
rect 44771 84420 44837 84421
rect 44771 84356 44772 84420
rect 44836 84356 44837 84420
rect 44771 84355 44837 84356
rect 42566 83950 42668 84010
rect 40160 83394 40220 83950
rect 41520 83394 41580 83950
rect 42608 83394 42668 83950
rect 43968 83950 44098 84010
rect 44774 84010 44834 84355
rect 46614 84010 46674 85579
rect 46804 85496 47124 86464
rect 47744 88634 48064 88676
rect 47744 88398 47786 88634
rect 48022 88398 48064 88634
rect 47744 85984 48064 88398
rect 47744 85920 47752 85984
rect 47816 85920 47832 85984
rect 47896 85920 47912 85984
rect 47976 85920 47992 85984
rect 48056 85920 48064 85984
rect 47347 85644 47413 85645
rect 47347 85580 47348 85644
rect 47412 85580 47413 85644
rect 47744 85620 48064 85920
rect 48404 87974 48724 88676
rect 48404 87738 48446 87974
rect 48682 87738 48724 87974
rect 48404 86528 48724 87738
rect 48404 86464 48412 86528
rect 48476 86464 48492 86528
rect 48556 86464 48572 86528
rect 48636 86464 48652 86528
rect 48716 86464 48724 86528
rect 47347 85579 47413 85580
rect 44774 83950 45252 84010
rect 43968 83394 44028 83950
rect 45192 83394 45252 83950
rect 46552 83950 46674 84010
rect 47350 84010 47410 85579
rect 48404 85496 48724 86464
rect 49344 88634 49664 88676
rect 49344 88398 49386 88634
rect 49622 88398 49664 88634
rect 49344 85984 49664 88398
rect 49344 85920 49352 85984
rect 49416 85920 49432 85984
rect 49496 85920 49512 85984
rect 49576 85920 49592 85984
rect 49656 85920 49664 85984
rect 49003 85644 49069 85645
rect 49003 85580 49004 85644
rect 49068 85580 49069 85644
rect 49003 85579 49069 85580
rect 49006 84010 49066 85579
rect 49344 85496 49664 85920
rect 50004 87974 50324 88676
rect 50004 87738 50046 87974
rect 50282 87738 50324 87974
rect 50004 86528 50324 87738
rect 50004 86464 50012 86528
rect 50076 86464 50092 86528
rect 50156 86464 50172 86528
rect 50236 86464 50252 86528
rect 50316 86464 50324 86528
rect 50004 85620 50324 86464
rect 50944 88634 51264 88676
rect 50944 88398 50986 88634
rect 51222 88398 51264 88634
rect 50944 85984 51264 88398
rect 50944 85920 50952 85984
rect 51016 85920 51032 85984
rect 51096 85920 51112 85984
rect 51176 85920 51192 85984
rect 51256 85920 51264 85984
rect 50475 85644 50541 85645
rect 50475 85580 50476 85644
rect 50540 85580 50541 85644
rect 50944 85620 51264 85920
rect 51604 87974 51924 88676
rect 51604 87738 51646 87974
rect 51882 87738 51924 87974
rect 51604 86528 51924 87738
rect 51604 86464 51612 86528
rect 51676 86464 51692 86528
rect 51756 86464 51772 86528
rect 51836 86464 51852 86528
rect 51916 86464 51924 86528
rect 50475 85579 50541 85580
rect 50478 84010 50538 85579
rect 51604 85496 51924 86464
rect 52544 88634 52864 88676
rect 52544 88398 52586 88634
rect 52822 88398 52864 88634
rect 52544 85984 52864 88398
rect 52544 85920 52552 85984
rect 52616 85920 52632 85984
rect 52696 85920 52712 85984
rect 52776 85920 52792 85984
rect 52856 85920 52864 85984
rect 52544 85620 52864 85920
rect 53204 87974 53524 88676
rect 53204 87738 53246 87974
rect 53482 87738 53524 87974
rect 53204 86528 53524 87738
rect 53204 86464 53212 86528
rect 53276 86464 53292 86528
rect 53356 86464 53372 86528
rect 53436 86464 53452 86528
rect 53516 86464 53524 86528
rect 53204 85496 53524 86464
rect 54144 88634 54464 88676
rect 54144 88398 54186 88634
rect 54422 88398 54464 88634
rect 54144 85984 54464 88398
rect 54144 85920 54152 85984
rect 54216 85920 54232 85984
rect 54296 85920 54312 85984
rect 54376 85920 54392 85984
rect 54456 85920 54464 85984
rect 54144 85496 54464 85920
rect 54804 87974 55124 88676
rect 54804 87738 54846 87974
rect 55082 87738 55124 87974
rect 54804 86528 55124 87738
rect 54804 86464 54812 86528
rect 54876 86464 54892 86528
rect 54956 86464 54972 86528
rect 55036 86464 55052 86528
rect 55116 86464 55124 86528
rect 54804 85496 55124 86464
rect 55744 88634 56064 88676
rect 55744 88398 55786 88634
rect 56022 88398 56064 88634
rect 55744 85984 56064 88398
rect 55744 85920 55752 85984
rect 55816 85920 55832 85984
rect 55896 85920 55912 85984
rect 55976 85920 55992 85984
rect 56056 85920 56064 85984
rect 55259 85644 55325 85645
rect 55259 85580 55260 85644
rect 55324 85580 55325 85644
rect 55259 85579 55325 85580
rect 52499 84828 52565 84829
rect 52499 84764 52500 84828
rect 52564 84764 52565 84828
rect 52499 84763 52565 84764
rect 51211 84692 51277 84693
rect 51211 84628 51212 84692
rect 51276 84628 51277 84692
rect 51211 84627 51277 84628
rect 47350 83950 47836 84010
rect 46552 83394 46612 83950
rect 47776 83394 47836 83950
rect 48864 83950 49066 84010
rect 50224 83950 50538 84010
rect 51214 84010 51274 84627
rect 52502 84010 52562 84763
rect 53787 84692 53853 84693
rect 53787 84628 53788 84692
rect 53852 84628 53853 84692
rect 53787 84627 53853 84628
rect 53790 84010 53850 84627
rect 55262 84010 55322 85579
rect 55744 85496 56064 85920
rect 56404 87974 56724 88676
rect 56404 87738 56446 87974
rect 56682 87738 56724 87974
rect 56404 86528 56724 87738
rect 56404 86464 56412 86528
rect 56476 86464 56492 86528
rect 56556 86464 56572 86528
rect 56636 86464 56652 86528
rect 56716 86464 56724 86528
rect 56179 85644 56245 85645
rect 56179 85580 56180 85644
rect 56244 85580 56245 85644
rect 56404 85620 56724 86464
rect 57344 88634 57664 88676
rect 57344 88398 57386 88634
rect 57622 88398 57664 88634
rect 57344 85984 57664 88398
rect 57344 85920 57352 85984
rect 57416 85920 57432 85984
rect 57496 85920 57512 85984
rect 57576 85920 57592 85984
rect 57656 85920 57664 85984
rect 57344 85620 57664 85920
rect 58004 87974 58324 88676
rect 58004 87738 58046 87974
rect 58282 87738 58324 87974
rect 58004 86528 58324 87738
rect 58004 86464 58012 86528
rect 58076 86464 58092 86528
rect 58156 86464 58172 86528
rect 58236 86464 58252 86528
rect 58316 86464 58324 86528
rect 56179 85579 56245 85580
rect 51214 83950 51372 84010
rect 52502 83950 52732 84010
rect 53790 83950 53956 84010
rect 48864 83394 48924 83950
rect 50224 83394 50284 83950
rect 51312 83394 51372 83950
rect 52672 83394 52732 83950
rect 53896 83394 53956 83950
rect 55256 83950 55322 84010
rect 56182 84010 56242 85579
rect 58004 85496 58324 86464
rect 58944 88634 59264 88676
rect 58944 88398 58986 88634
rect 59222 88398 59264 88634
rect 58944 85984 59264 88398
rect 58944 85920 58952 85984
rect 59016 85920 59032 85984
rect 59096 85920 59112 85984
rect 59176 85920 59192 85984
rect 59256 85920 59264 85984
rect 58755 85644 58821 85645
rect 58755 85580 58756 85644
rect 58820 85580 58821 85644
rect 58944 85620 59264 85920
rect 59604 87974 59924 88676
rect 59604 87738 59646 87974
rect 59882 87738 59924 87974
rect 59604 86528 59924 87738
rect 59604 86464 59612 86528
rect 59676 86464 59692 86528
rect 59756 86464 59772 86528
rect 59836 86464 59852 86528
rect 59916 86464 59924 86528
rect 58755 85579 58821 85580
rect 57651 84556 57717 84557
rect 57651 84492 57652 84556
rect 57716 84492 57717 84556
rect 57651 84491 57717 84492
rect 57654 84010 57714 84491
rect 56182 83950 56404 84010
rect 55256 83394 55316 83950
rect 56344 83394 56404 83950
rect 57568 83950 57714 84010
rect 58758 84010 58818 85579
rect 59604 85496 59924 86464
rect 60544 88634 60864 88676
rect 60544 88398 60586 88634
rect 60822 88398 60864 88634
rect 60544 85984 60864 88398
rect 60544 85920 60552 85984
rect 60616 85920 60632 85984
rect 60696 85920 60712 85984
rect 60776 85920 60792 85984
rect 60856 85920 60864 85984
rect 60544 85496 60864 85920
rect 61204 87974 61524 88676
rect 61204 87738 61246 87974
rect 61482 87738 61524 87974
rect 61204 86528 61524 87738
rect 61204 86464 61212 86528
rect 61276 86464 61292 86528
rect 61356 86464 61372 86528
rect 61436 86464 61452 86528
rect 61516 86464 61524 86528
rect 60963 85916 61029 85917
rect 60963 85852 60964 85916
rect 61028 85852 61029 85916
rect 60963 85851 61029 85852
rect 60966 84210 61026 85851
rect 61204 85620 61524 86464
rect 62144 88634 62464 88676
rect 62144 88398 62186 88634
rect 62422 88398 62464 88634
rect 62144 85984 62464 88398
rect 62144 85920 62152 85984
rect 62216 85920 62232 85984
rect 62296 85920 62312 85984
rect 62376 85920 62392 85984
rect 62456 85920 62464 85984
rect 62144 85496 62464 85920
rect 62804 87974 63124 88676
rect 62804 87738 62846 87974
rect 63082 87738 63124 87974
rect 62804 86528 63124 87738
rect 62804 86464 62812 86528
rect 62876 86464 62892 86528
rect 62956 86464 62972 86528
rect 63036 86464 63052 86528
rect 63116 86464 63124 86528
rect 62619 85644 62685 85645
rect 62619 85580 62620 85644
rect 62684 85580 62685 85644
rect 62619 85579 62685 85580
rect 60966 84150 61394 84210
rect 61334 84010 61394 84150
rect 62622 84010 62682 85579
rect 62804 85496 63124 86464
rect 63744 88634 64064 88676
rect 63744 88398 63786 88634
rect 64022 88398 64064 88634
rect 63744 85984 64064 88398
rect 63744 85920 63752 85984
rect 63816 85920 63832 85984
rect 63896 85920 63912 85984
rect 63976 85920 63992 85984
rect 64056 85920 64064 85984
rect 63539 85916 63605 85917
rect 63539 85852 63540 85916
rect 63604 85852 63605 85916
rect 63539 85851 63605 85852
rect 63542 84210 63602 85851
rect 63744 85620 64064 85920
rect 64404 87974 64724 88676
rect 64404 87738 64446 87974
rect 64682 87738 64724 87974
rect 64404 86528 64724 87738
rect 64404 86464 64412 86528
rect 64476 86464 64492 86528
rect 64556 86464 64572 86528
rect 64636 86464 64652 86528
rect 64716 86464 64724 86528
rect 64404 85496 64724 86464
rect 65344 88634 65664 88676
rect 65344 88398 65386 88634
rect 65622 88398 65664 88634
rect 65344 85984 65664 88398
rect 65344 85920 65352 85984
rect 65416 85920 65432 85984
rect 65496 85920 65512 85984
rect 65576 85920 65592 85984
rect 65656 85920 65664 85984
rect 65344 85496 65664 85920
rect 66004 87974 66324 88676
rect 66004 87738 66046 87974
rect 66282 87738 66324 87974
rect 66004 86528 66324 87738
rect 66004 86464 66012 86528
rect 66076 86464 66092 86528
rect 66156 86464 66172 86528
rect 66236 86464 66252 86528
rect 66316 86464 66324 86528
rect 66004 85620 66324 86464
rect 66944 88634 67264 88676
rect 66944 88398 66986 88634
rect 67222 88398 67264 88634
rect 66944 85984 67264 88398
rect 66944 85920 66952 85984
rect 67016 85920 67032 85984
rect 67096 85920 67112 85984
rect 67176 85920 67192 85984
rect 67256 85920 67264 85984
rect 66944 85496 67264 85920
rect 67604 87974 67924 88676
rect 67604 87738 67646 87974
rect 67882 87738 67924 87974
rect 67604 86528 67924 87738
rect 67604 86464 67612 86528
rect 67676 86464 67692 86528
rect 67756 86464 67772 86528
rect 67836 86464 67852 86528
rect 67916 86464 67924 86528
rect 67604 85620 67924 86464
rect 68544 88634 68864 88676
rect 68544 88398 68586 88634
rect 68822 88398 68864 88634
rect 68544 85984 68864 88398
rect 68544 85920 68552 85984
rect 68616 85920 68632 85984
rect 68696 85920 68712 85984
rect 68776 85920 68792 85984
rect 68856 85920 68864 85984
rect 68139 85916 68205 85917
rect 68139 85852 68140 85916
rect 68204 85852 68205 85916
rect 68139 85851 68205 85852
rect 66299 84692 66365 84693
rect 66299 84628 66300 84692
rect 66364 84628 66365 84692
rect 66299 84627 66365 84628
rect 65011 84284 65077 84285
rect 65011 84220 65012 84284
rect 65076 84220 65077 84284
rect 65011 84219 65077 84220
rect 63542 84150 63970 84210
rect 58758 83950 58988 84010
rect 61334 83950 61572 84010
rect 57568 83394 57628 83950
rect 58928 83394 58988 83950
rect 60149 83740 60215 83741
rect 60149 83676 60150 83740
rect 60214 83676 60215 83740
rect 60149 83675 60215 83676
rect 60152 83394 60212 83675
rect 61512 83394 61572 83950
rect 62600 83950 62682 84010
rect 63910 84010 63970 84150
rect 65014 84010 65074 84219
rect 66302 84010 66362 84627
rect 68142 84210 68202 85851
rect 68323 85780 68389 85781
rect 68323 85716 68324 85780
rect 68388 85716 68389 85780
rect 68323 85715 68389 85716
rect 67774 84150 68202 84210
rect 68326 84210 68386 85715
rect 68544 85620 68864 85920
rect 69204 87974 69524 88676
rect 69204 87738 69246 87974
rect 69482 87738 69524 87974
rect 69204 86528 69524 87738
rect 69204 86464 69212 86528
rect 69276 86464 69292 86528
rect 69356 86464 69372 86528
rect 69436 86464 69452 86528
rect 69516 86464 69524 86528
rect 69204 85496 69524 86464
rect 70144 88634 70464 88676
rect 70144 88398 70186 88634
rect 70422 88398 70464 88634
rect 70144 85984 70464 88398
rect 70144 85920 70152 85984
rect 70216 85920 70232 85984
rect 70296 85920 70312 85984
rect 70376 85920 70392 85984
rect 70456 85920 70464 85984
rect 70144 85620 70464 85920
rect 70804 87974 71124 88676
rect 70804 87738 70846 87974
rect 71082 87738 71124 87974
rect 70804 86528 71124 87738
rect 70804 86464 70812 86528
rect 70876 86464 70892 86528
rect 70956 86464 70972 86528
rect 71036 86464 71052 86528
rect 71116 86464 71124 86528
rect 70804 85496 71124 86464
rect 71744 88634 72064 88676
rect 71744 88398 71786 88634
rect 72022 88398 72064 88634
rect 71744 85984 72064 88398
rect 71744 85920 71752 85984
rect 71816 85920 71832 85984
rect 71896 85920 71912 85984
rect 71976 85920 71992 85984
rect 72056 85920 72064 85984
rect 71744 85496 72064 85920
rect 72404 87974 72724 88676
rect 72404 87738 72446 87974
rect 72682 87738 72724 87974
rect 72404 86528 72724 87738
rect 72404 86464 72412 86528
rect 72476 86464 72492 86528
rect 72556 86464 72572 86528
rect 72636 86464 72652 86528
rect 72716 86464 72724 86528
rect 72187 85916 72253 85917
rect 72187 85852 72188 85916
rect 72252 85852 72253 85916
rect 72187 85851 72253 85852
rect 71267 84692 71333 84693
rect 71267 84628 71268 84692
rect 71332 84628 71333 84692
rect 71267 84627 71333 84628
rect 68326 84150 68754 84210
rect 67774 84010 67834 84150
rect 63910 83950 64020 84010
rect 65014 83950 65108 84010
rect 62600 83394 62660 83950
rect 63960 83394 64020 83950
rect 65048 83394 65108 83950
rect 66272 83950 66362 84010
rect 67632 83950 67834 84010
rect 68694 84010 68754 84150
rect 71270 84010 71330 84627
rect 72190 84210 72250 85851
rect 72404 85620 72724 86464
rect 73344 88634 73664 88676
rect 73344 88398 73386 88634
rect 73622 88398 73664 88634
rect 73344 85984 73664 88398
rect 73344 85920 73352 85984
rect 73416 85920 73432 85984
rect 73496 85920 73512 85984
rect 73576 85920 73592 85984
rect 73656 85920 73664 85984
rect 73344 85496 73664 85920
rect 74004 87974 74324 88676
rect 74004 87738 74046 87974
rect 74282 87738 74324 87974
rect 74004 86528 74324 87738
rect 74004 86464 74012 86528
rect 74076 86464 74092 86528
rect 74156 86464 74172 86528
rect 74236 86464 74252 86528
rect 74316 86464 74324 86528
rect 73843 85644 73909 85645
rect 73843 85580 73844 85644
rect 73908 85580 73909 85644
rect 74004 85620 74324 86464
rect 74944 88634 75264 88676
rect 74944 88398 74986 88634
rect 75222 88398 75264 88634
rect 74944 85984 75264 88398
rect 74944 85920 74952 85984
rect 75016 85920 75032 85984
rect 75096 85920 75112 85984
rect 75176 85920 75192 85984
rect 75256 85920 75264 85984
rect 74944 85620 75264 85920
rect 75604 87974 75924 88676
rect 75604 87738 75646 87974
rect 75882 87738 75924 87974
rect 75604 86528 75924 87738
rect 75604 86464 75612 86528
rect 75676 86464 75692 86528
rect 75756 86464 75772 86528
rect 75836 86464 75852 86528
rect 75916 86464 75924 86528
rect 73843 85579 73909 85580
rect 72190 84150 72618 84210
rect 72558 84010 72618 84150
rect 73846 84010 73906 85579
rect 75315 85508 75381 85509
rect 75315 85444 75316 85508
rect 75380 85444 75381 85508
rect 75604 85496 75924 86464
rect 76544 88634 76864 88676
rect 76544 88398 76586 88634
rect 76822 88398 76864 88634
rect 76544 85984 76864 88398
rect 76544 85920 76552 85984
rect 76616 85920 76632 85984
rect 76696 85920 76712 85984
rect 76776 85920 76792 85984
rect 76856 85920 76864 85984
rect 76235 85644 76301 85645
rect 76235 85580 76236 85644
rect 76300 85580 76301 85644
rect 76235 85579 76301 85580
rect 75315 85443 75381 85444
rect 75318 84010 75378 85443
rect 68694 83950 68916 84010
rect 71270 83950 71364 84010
rect 72558 83950 72724 84010
rect 73846 83950 73948 84010
rect 66272 83394 66332 83950
rect 67632 83394 67692 83950
rect 68856 83394 68916 83950
rect 70213 83740 70279 83741
rect 70213 83676 70214 83740
rect 70278 83676 70279 83740
rect 70213 83675 70279 83676
rect 70216 83394 70276 83675
rect 71304 83394 71364 83950
rect 72664 83394 72724 83950
rect 73888 83394 73948 83950
rect 75248 83950 75378 84010
rect 76238 84010 76298 85579
rect 76544 85496 76864 85920
rect 77204 87974 77524 88676
rect 77204 87738 77246 87974
rect 77482 87738 77524 87974
rect 77204 86528 77524 87738
rect 77204 86464 77212 86528
rect 77276 86464 77292 86528
rect 77356 86464 77372 86528
rect 77436 86464 77452 86528
rect 77516 86464 77524 86528
rect 77204 85620 77524 86464
rect 78144 88634 78464 88676
rect 78144 88398 78186 88634
rect 78422 88398 78464 88634
rect 78144 85984 78464 88398
rect 78144 85920 78152 85984
rect 78216 85920 78232 85984
rect 78296 85920 78312 85984
rect 78376 85920 78392 85984
rect 78456 85920 78464 85984
rect 77707 85644 77773 85645
rect 77707 85580 77708 85644
rect 77772 85580 77773 85644
rect 77707 85579 77773 85580
rect 77710 84010 77770 85579
rect 78144 85496 78464 85920
rect 78804 87974 79124 88676
rect 78804 87738 78846 87974
rect 79082 87738 79124 87974
rect 78804 86528 79124 87738
rect 78804 86464 78812 86528
rect 78876 86464 78892 86528
rect 78956 86464 78972 86528
rect 79036 86464 79052 86528
rect 79116 86464 79124 86528
rect 78804 85620 79124 86464
rect 79744 88634 80064 88676
rect 79744 88398 79786 88634
rect 80022 88398 80064 88634
rect 79744 85984 80064 88398
rect 79744 85920 79752 85984
rect 79816 85920 79832 85984
rect 79896 85920 79912 85984
rect 79976 85920 79992 85984
rect 80056 85920 80064 85984
rect 79744 85496 80064 85920
rect 80404 87974 80724 88676
rect 80404 87738 80446 87974
rect 80682 87738 80724 87974
rect 80404 86528 80724 87738
rect 80404 86464 80412 86528
rect 80476 86464 80492 86528
rect 80556 86464 80572 86528
rect 80636 86464 80652 86528
rect 80716 86464 80724 86528
rect 80404 85496 80724 86464
rect 81344 88634 81664 88676
rect 81344 88398 81386 88634
rect 81622 88398 81664 88634
rect 81344 85984 81664 88398
rect 81344 85920 81352 85984
rect 81416 85920 81432 85984
rect 81496 85920 81512 85984
rect 81576 85920 81592 85984
rect 81656 85920 81664 85984
rect 81344 85496 81664 85920
rect 82004 87974 82324 88676
rect 82004 87738 82046 87974
rect 82282 87738 82324 87974
rect 82004 86528 82324 87738
rect 82004 86464 82012 86528
rect 82076 86464 82092 86528
rect 82156 86464 82172 86528
rect 82236 86464 82252 86528
rect 82316 86464 82324 86528
rect 82004 85496 82324 86464
rect 82944 88634 83264 88676
rect 82944 88398 82986 88634
rect 83222 88398 83264 88634
rect 82944 85984 83264 88398
rect 82944 85920 82952 85984
rect 83016 85920 83032 85984
rect 83096 85920 83112 85984
rect 83176 85920 83192 85984
rect 83256 85920 83264 85984
rect 82944 85496 83264 85920
rect 83604 87974 83924 88676
rect 83604 87738 83646 87974
rect 83882 87738 83924 87974
rect 83604 86528 83924 87738
rect 83604 86464 83612 86528
rect 83676 86464 83692 86528
rect 83756 86464 83772 86528
rect 83836 86464 83852 86528
rect 83916 86464 83924 86528
rect 83604 85496 83924 86464
rect 84544 88634 84864 88676
rect 84544 88398 84586 88634
rect 84822 88398 84864 88634
rect 84544 85984 84864 88398
rect 84544 85920 84552 85984
rect 84616 85920 84632 85984
rect 84696 85920 84712 85984
rect 84776 85920 84792 85984
rect 84856 85920 84864 85984
rect 84544 85496 84864 85920
rect 85204 87974 85524 88676
rect 85204 87738 85246 87974
rect 85482 87738 85524 87974
rect 85204 86528 85524 87738
rect 85204 86464 85212 86528
rect 85276 86464 85292 86528
rect 85356 86464 85372 86528
rect 85436 86464 85452 86528
rect 85516 86464 85524 86528
rect 85204 85496 85524 86464
rect 86144 88634 86464 88676
rect 86144 88398 86186 88634
rect 86422 88398 86464 88634
rect 86144 85984 86464 88398
rect 86144 85920 86152 85984
rect 86216 85920 86232 85984
rect 86296 85920 86312 85984
rect 86376 85920 86392 85984
rect 86456 85920 86464 85984
rect 86144 85496 86464 85920
rect 86804 87974 87124 88676
rect 86804 87738 86846 87974
rect 87082 87738 87124 87974
rect 86804 86528 87124 87738
rect 86804 86464 86812 86528
rect 86876 86464 86892 86528
rect 86956 86464 86972 86528
rect 87036 86464 87052 86528
rect 87116 86464 87124 86528
rect 86804 85496 87124 86464
rect 87744 88634 88064 88676
rect 87744 88398 87786 88634
rect 88022 88398 88064 88634
rect 87744 85984 88064 88398
rect 87744 85920 87752 85984
rect 87816 85920 87832 85984
rect 87896 85920 87912 85984
rect 87976 85920 87992 85984
rect 88056 85920 88064 85984
rect 87744 85496 88064 85920
rect 88404 87974 88724 88676
rect 88404 87738 88446 87974
rect 88682 87738 88724 87974
rect 88404 86528 88724 87738
rect 88404 86464 88412 86528
rect 88476 86464 88492 86528
rect 88556 86464 88572 86528
rect 88636 86464 88652 86528
rect 88716 86464 88724 86528
rect 88404 85496 88724 86464
rect 89344 88634 89664 88676
rect 89344 88398 89386 88634
rect 89622 88398 89664 88634
rect 89344 85984 89664 88398
rect 89344 85920 89352 85984
rect 89416 85920 89432 85984
rect 89496 85920 89512 85984
rect 89576 85920 89592 85984
rect 89656 85920 89664 85984
rect 89344 85496 89664 85920
rect 90004 87974 90324 88676
rect 90004 87738 90046 87974
rect 90282 87738 90324 87974
rect 90004 86528 90324 87738
rect 90004 86464 90012 86528
rect 90076 86464 90092 86528
rect 90156 86464 90172 86528
rect 90236 86464 90252 86528
rect 90316 86464 90324 86528
rect 90004 85496 90324 86464
rect 90944 88634 91264 88676
rect 90944 88398 90986 88634
rect 91222 88398 91264 88634
rect 90944 85984 91264 88398
rect 90944 85920 90952 85984
rect 91016 85920 91032 85984
rect 91096 85920 91112 85984
rect 91176 85920 91192 85984
rect 91256 85920 91264 85984
rect 90944 85496 91264 85920
rect 91604 87974 91924 88676
rect 91604 87738 91646 87974
rect 91882 87738 91924 87974
rect 91604 86528 91924 87738
rect 91604 86464 91612 86528
rect 91676 86464 91692 86528
rect 91756 86464 91772 86528
rect 91836 86464 91852 86528
rect 91916 86464 91924 86528
rect 91604 85620 91924 86464
rect 92544 88634 92864 88676
rect 92544 88398 92586 88634
rect 92822 88398 92864 88634
rect 92544 85984 92864 88398
rect 92544 85920 92552 85984
rect 92616 85920 92632 85984
rect 92696 85920 92712 85984
rect 92776 85920 92792 85984
rect 92856 85920 92864 85984
rect 91507 85508 91573 85509
rect 91507 85444 91508 85508
rect 91572 85444 91573 85508
rect 92544 85496 92864 85920
rect 93204 87974 93524 88676
rect 93204 87738 93246 87974
rect 93482 87738 93524 87974
rect 93204 86528 93524 87738
rect 93204 86464 93212 86528
rect 93276 86464 93292 86528
rect 93356 86464 93372 86528
rect 93436 86464 93452 86528
rect 93516 86464 93524 86528
rect 93204 85496 93524 86464
rect 94144 88634 94464 88676
rect 94144 88398 94186 88634
rect 94422 88398 94464 88634
rect 94144 85984 94464 88398
rect 94144 85920 94152 85984
rect 94216 85920 94232 85984
rect 94296 85920 94312 85984
rect 94376 85920 94392 85984
rect 94456 85920 94464 85984
rect 94144 85496 94464 85920
rect 94804 87974 95124 88676
rect 94804 87738 94846 87974
rect 95082 87738 95124 87974
rect 94804 86528 95124 87738
rect 94804 86464 94812 86528
rect 94876 86464 94892 86528
rect 94956 86464 94972 86528
rect 95036 86464 95052 86528
rect 95116 86464 95124 86528
rect 94804 85496 95124 86464
rect 95744 88634 96064 88676
rect 95744 88398 95786 88634
rect 96022 88398 96064 88634
rect 95744 85984 96064 88398
rect 95744 85920 95752 85984
rect 95816 85920 95832 85984
rect 95896 85920 95912 85984
rect 95976 85920 95992 85984
rect 96056 85920 96064 85984
rect 95744 85496 96064 85920
rect 96404 87974 96724 88676
rect 96404 87738 96446 87974
rect 96682 87738 96724 87974
rect 96404 86528 96724 87738
rect 96404 86464 96412 86528
rect 96476 86464 96492 86528
rect 96556 86464 96572 86528
rect 96636 86464 96652 86528
rect 96716 86464 96724 86528
rect 96404 85496 96724 86464
rect 97344 88634 97664 88676
rect 97344 88398 97386 88634
rect 97622 88398 97664 88634
rect 97344 85984 97664 88398
rect 97344 85920 97352 85984
rect 97416 85920 97432 85984
rect 97496 85920 97512 85984
rect 97576 85920 97592 85984
rect 97656 85920 97664 85984
rect 97344 85496 97664 85920
rect 98004 87974 98324 88676
rect 98004 87738 98046 87974
rect 98282 87738 98324 87974
rect 98004 86528 98324 87738
rect 98004 86464 98012 86528
rect 98076 86464 98092 86528
rect 98156 86464 98172 86528
rect 98236 86464 98252 86528
rect 98316 86464 98324 86528
rect 98004 85496 98324 86464
rect 98944 88634 99264 88676
rect 98944 88398 98986 88634
rect 99222 88398 99264 88634
rect 98944 85984 99264 88398
rect 98944 85920 98952 85984
rect 99016 85920 99032 85984
rect 99096 85920 99112 85984
rect 99176 85920 99192 85984
rect 99256 85920 99264 85984
rect 98944 85496 99264 85920
rect 99604 87974 99924 88676
rect 99604 87738 99646 87974
rect 99882 87738 99924 87974
rect 99604 86528 99924 87738
rect 99604 86464 99612 86528
rect 99676 86464 99692 86528
rect 99756 86464 99772 86528
rect 99836 86464 99852 86528
rect 99916 86464 99924 86528
rect 99604 85496 99924 86464
rect 100544 88634 100864 88676
rect 100544 88398 100586 88634
rect 100822 88398 100864 88634
rect 100544 85984 100864 88398
rect 100544 85920 100552 85984
rect 100616 85920 100632 85984
rect 100696 85920 100712 85984
rect 100776 85920 100792 85984
rect 100856 85920 100864 85984
rect 100544 85496 100864 85920
rect 101204 87974 101524 88676
rect 101204 87738 101246 87974
rect 101482 87738 101524 87974
rect 101204 86528 101524 87738
rect 101204 86464 101212 86528
rect 101276 86464 101292 86528
rect 101356 86464 101372 86528
rect 101436 86464 101452 86528
rect 101516 86464 101524 86528
rect 101204 85496 101524 86464
rect 102144 88634 102464 88676
rect 102144 88398 102186 88634
rect 102422 88398 102464 88634
rect 102144 85984 102464 88398
rect 102144 85920 102152 85984
rect 102216 85920 102232 85984
rect 102296 85920 102312 85984
rect 102376 85920 102392 85984
rect 102456 85920 102464 85984
rect 101995 85644 102061 85645
rect 101995 85580 101996 85644
rect 102060 85580 102061 85644
rect 102144 85620 102464 85920
rect 102804 87974 103124 88676
rect 102804 87738 102846 87974
rect 103082 87738 103124 87974
rect 102804 86528 103124 87738
rect 102804 86464 102812 86528
rect 102876 86464 102892 86528
rect 102956 86464 102972 86528
rect 103036 86464 103052 86528
rect 103116 86464 103124 86528
rect 101995 85579 102061 85580
rect 91507 85443 91573 85444
rect 78627 84556 78693 84557
rect 78627 84492 78628 84556
rect 78692 84492 78693 84556
rect 78627 84491 78693 84492
rect 76238 83950 76396 84010
rect 75248 83394 75308 83950
rect 76336 83394 76396 83950
rect 77560 83950 77770 84010
rect 78630 84010 78690 84491
rect 91510 84010 91570 85443
rect 78630 83950 78980 84010
rect 77560 83394 77620 83950
rect 78920 83394 78980 83950
rect 91432 83950 91570 84010
rect 101998 84010 102058 85579
rect 102804 85496 103124 86464
rect 103744 88634 104064 88676
rect 103744 88398 103786 88634
rect 104022 88398 104064 88634
rect 103744 85984 104064 88398
rect 103744 85920 103752 85984
rect 103816 85920 103832 85984
rect 103896 85920 103912 85984
rect 103976 85920 103992 85984
rect 104056 85920 104064 85984
rect 103744 85496 104064 85920
rect 104404 87974 104724 88676
rect 104404 87738 104446 87974
rect 104682 87738 104724 87974
rect 104404 86528 104724 87738
rect 104404 86464 104412 86528
rect 104476 86464 104492 86528
rect 104556 86464 104572 86528
rect 104636 86464 104652 86528
rect 104716 86464 104724 86528
rect 104404 85496 104724 86464
rect 105344 88634 105664 88676
rect 105344 88398 105386 88634
rect 105622 88398 105664 88634
rect 105344 85984 105664 88398
rect 105344 85920 105352 85984
rect 105416 85920 105432 85984
rect 105496 85920 105512 85984
rect 105576 85920 105592 85984
rect 105656 85920 105664 85984
rect 105344 85496 105664 85920
rect 106004 87974 106324 88676
rect 106004 87738 106046 87974
rect 106282 87738 106324 87974
rect 106004 86528 106324 87738
rect 106004 86464 106012 86528
rect 106076 86464 106092 86528
rect 106156 86464 106172 86528
rect 106236 86464 106252 86528
rect 106316 86464 106324 86528
rect 106004 85496 106324 86464
rect 106944 88634 107264 88676
rect 106944 88398 106986 88634
rect 107222 88398 107264 88634
rect 106944 85984 107264 88398
rect 106944 85920 106952 85984
rect 107016 85920 107032 85984
rect 107096 85920 107112 85984
rect 107176 85920 107192 85984
rect 107256 85920 107264 85984
rect 106944 85496 107264 85920
rect 107604 87974 107924 88676
rect 107604 87738 107646 87974
rect 107882 87738 107924 87974
rect 107604 86528 107924 87738
rect 107604 86464 107612 86528
rect 107676 86464 107692 86528
rect 107756 86464 107772 86528
rect 107836 86464 107852 86528
rect 107916 86464 107924 86528
rect 107604 85496 107924 86464
rect 108544 88634 108864 88676
rect 108544 88398 108586 88634
rect 108822 88398 108864 88634
rect 108544 85984 108864 88398
rect 110696 88634 111016 88676
rect 110696 88398 110738 88634
rect 110974 88398 111016 88634
rect 108544 85920 108552 85984
rect 108616 85920 108632 85984
rect 108696 85920 108712 85984
rect 108776 85920 108792 85984
rect 108856 85920 108864 85984
rect 108544 85496 108864 85920
rect 110036 87974 110356 88016
rect 110036 87738 110078 87974
rect 110314 87738 110356 87974
rect 101998 83950 102100 84010
rect 91432 83394 91492 83950
rect 102040 83394 102100 83950
rect 110036 82866 110356 87738
rect 110036 82630 110078 82866
rect 110314 82630 110356 82866
rect 12272 82206 12620 82248
rect 12272 81970 12328 82206
rect 12564 81970 12620 82206
rect 12272 81928 12620 81970
rect 107336 82206 107684 82248
rect 107336 81970 107392 82206
rect 107628 81970 107684 82206
rect 107336 81928 107684 81970
rect 11467 68916 11533 68917
rect 11467 68852 11468 68916
rect 11532 68852 11533 68916
rect 11467 68851 11533 68852
rect 11835 66604 11901 66605
rect 11835 66540 11836 66604
rect 11900 66540 11901 66604
rect 11835 66539 11901 66540
rect 11099 39948 11165 39949
rect 11099 39884 11100 39948
rect 11164 39884 11165 39948
rect 11099 39883 11165 39884
rect 10547 38452 10613 38453
rect 10547 38388 10548 38452
rect 10612 38388 10613 38452
rect 10547 38387 10613 38388
rect 9344 38048 9352 38112
rect 9416 38048 9432 38112
rect 9496 38048 9512 38112
rect 9576 38048 9592 38112
rect 9656 38048 9664 38112
rect 9344 37024 9664 38048
rect 10731 37364 10797 37365
rect 10731 37300 10732 37364
rect 10796 37300 10797 37364
rect 10731 37299 10797 37300
rect 9344 36960 9352 37024
rect 9416 36960 9432 37024
rect 9496 36960 9512 37024
rect 9576 36960 9592 37024
rect 9656 36960 9664 37024
rect 9344 35936 9664 36960
rect 9344 35872 9352 35936
rect 9416 35872 9432 35936
rect 9496 35872 9512 35936
rect 9576 35872 9592 35936
rect 9656 35872 9664 35936
rect 9344 34848 9664 35872
rect 9344 34784 9352 34848
rect 9416 34784 9432 34848
rect 9496 34784 9512 34848
rect 9576 34784 9592 34848
rect 9656 34784 9664 34848
rect 9344 33760 9664 34784
rect 9344 33696 9352 33760
rect 9416 33696 9432 33760
rect 9496 33696 9512 33760
rect 9576 33696 9592 33760
rect 9656 33696 9664 33760
rect 9344 32672 9664 33696
rect 9344 32608 9352 32672
rect 9416 32608 9432 32672
rect 9496 32608 9512 32672
rect 9576 32608 9592 32672
rect 9656 32608 9664 32672
rect 9344 31584 9664 32608
rect 9344 31520 9352 31584
rect 9416 31520 9432 31584
rect 9496 31520 9512 31584
rect 9576 31520 9592 31584
rect 9656 31520 9664 31584
rect 9344 30496 9664 31520
rect 9344 30432 9352 30496
rect 9416 30432 9432 30496
rect 9496 30432 9512 30496
rect 9576 30432 9592 30496
rect 9656 30432 9664 30496
rect 9344 29408 9664 30432
rect 9344 29344 9352 29408
rect 9416 29344 9432 29408
rect 9496 29344 9512 29408
rect 9576 29344 9592 29408
rect 9656 29344 9664 29408
rect 9344 28320 9664 29344
rect 9344 28256 9352 28320
rect 9416 28256 9432 28320
rect 9496 28256 9512 28320
rect 9576 28256 9592 28320
rect 9656 28256 9664 28320
rect 9344 27232 9664 28256
rect 9344 27168 9352 27232
rect 9416 27168 9432 27232
rect 9496 27168 9512 27232
rect 9576 27168 9592 27232
rect 9656 27168 9664 27232
rect 9344 26144 9664 27168
rect 9344 26080 9352 26144
rect 9416 26080 9432 26144
rect 9496 26080 9512 26144
rect 9576 26080 9592 26144
rect 9656 26080 9664 26144
rect 9344 25056 9664 26080
rect 9344 24992 9352 25056
rect 9416 24992 9432 25056
rect 9496 24992 9512 25056
rect 9576 24992 9592 25056
rect 9656 24992 9664 25056
rect 9344 23968 9664 24992
rect 9344 23904 9352 23968
rect 9416 23904 9432 23968
rect 9496 23904 9512 23968
rect 9576 23904 9592 23968
rect 9656 23904 9664 23968
rect 9344 22880 9664 23904
rect 9344 22816 9352 22880
rect 9416 22816 9432 22880
rect 9496 22816 9512 22880
rect 9576 22816 9592 22880
rect 9656 22816 9664 22880
rect 9344 21792 9664 22816
rect 9344 21728 9352 21792
rect 9416 21728 9432 21792
rect 9496 21728 9512 21792
rect 9576 21728 9592 21792
rect 9656 21728 9664 21792
rect 9344 20704 9664 21728
rect 9344 20640 9352 20704
rect 9416 20640 9432 20704
rect 9496 20640 9512 20704
rect 9576 20640 9592 20704
rect 9656 20640 9664 20704
rect 9344 19616 9664 20640
rect 9344 19552 9352 19616
rect 9416 19552 9432 19616
rect 9496 19552 9512 19616
rect 9576 19552 9592 19616
rect 9656 19552 9664 19616
rect 9344 18528 9664 19552
rect 9344 18464 9352 18528
rect 9416 18464 9432 18528
rect 9496 18464 9512 18528
rect 9576 18464 9592 18528
rect 9656 18464 9664 18528
rect 9344 17440 9664 18464
rect 9344 17376 9352 17440
rect 9416 17376 9432 17440
rect 9496 17376 9512 17440
rect 9576 17376 9592 17440
rect 9656 17376 9664 17440
rect 9344 16352 9664 17376
rect 9344 16288 9352 16352
rect 9416 16288 9432 16352
rect 9496 16288 9512 16352
rect 9576 16288 9592 16352
rect 9656 16288 9664 16352
rect 9344 15264 9664 16288
rect 9344 15200 9352 15264
rect 9416 15200 9432 15264
rect 9496 15200 9512 15264
rect 9576 15200 9592 15264
rect 9656 15200 9664 15264
rect 9344 14176 9664 15200
rect 9344 14112 9352 14176
rect 9416 14112 9432 14176
rect 9496 14112 9512 14176
rect 9576 14112 9592 14176
rect 9656 14112 9664 14176
rect 9344 13088 9664 14112
rect 9344 13024 9352 13088
rect 9416 13024 9432 13088
rect 9496 13024 9512 13088
rect 9576 13024 9592 13088
rect 9656 13024 9664 13088
rect 9344 12000 9664 13024
rect 9344 11936 9352 12000
rect 9416 11936 9432 12000
rect 9496 11936 9512 12000
rect 9576 11936 9592 12000
rect 9656 11936 9664 12000
rect 9344 10912 9664 11936
rect 9344 10848 9352 10912
rect 9416 10848 9432 10912
rect 9496 10848 9512 10912
rect 9576 10848 9592 10912
rect 9656 10848 9664 10912
rect 9344 9824 9664 10848
rect 9344 9760 9352 9824
rect 9416 9760 9432 9824
rect 9496 9760 9512 9824
rect 9576 9760 9592 9824
rect 9656 9760 9664 9824
rect 9344 8736 9664 9760
rect 9344 8672 9352 8736
rect 9416 8672 9432 8736
rect 9496 8672 9512 8736
rect 9576 8672 9592 8736
rect 9656 8672 9664 8736
rect 9344 7648 9664 8672
rect 9344 7584 9352 7648
rect 9416 7584 9432 7648
rect 9496 7584 9512 7648
rect 9576 7584 9592 7648
rect 9656 7584 9664 7648
rect 9344 6560 9664 7584
rect 9344 6496 9352 6560
rect 9416 6496 9432 6560
rect 9496 6496 9512 6560
rect 9576 6496 9592 6560
rect 9656 6496 9664 6560
rect 9344 6206 9664 6496
rect 9344 5970 9386 6206
rect 9622 5970 9664 6206
rect 9344 5472 9664 5970
rect 9344 5408 9352 5472
rect 9416 5408 9432 5472
rect 9496 5408 9512 5472
rect 9576 5408 9592 5472
rect 9656 5408 9664 5472
rect 9344 4384 9664 5408
rect 9344 4320 9352 4384
rect 9416 4320 9432 4384
rect 9496 4320 9512 4384
rect 9576 4320 9592 4384
rect 9656 4320 9664 4384
rect 9344 3296 9664 4320
rect 9344 3232 9352 3296
rect 9416 3232 9432 3296
rect 9496 3232 9512 3296
rect 9576 3232 9592 3296
rect 9656 3232 9664 3296
rect 9344 2208 9664 3232
rect 9344 2144 9352 2208
rect 9416 2144 9432 2208
rect 9496 2144 9512 2208
rect 9576 2144 9592 2208
rect 9656 2144 9664 2208
rect 9344 1120 9664 2144
rect 9344 1056 9352 1120
rect 9416 1056 9432 1120
rect 9496 1056 9512 1120
rect 9576 1056 9592 1120
rect 9656 1056 9664 1120
rect 9344 -814 9664 1056
rect 9344 -1050 9386 -814
rect 9622 -1050 9664 -814
rect 9344 -1092 9664 -1050
rect 10004 1664 10324 2004
rect 10004 1600 10012 1664
rect 10076 1600 10092 1664
rect 10156 1600 10172 1664
rect 10236 1600 10252 1664
rect 10316 1600 10324 1664
rect 10004 -154 10324 1600
rect 10734 645 10794 37299
rect 11651 36412 11717 36413
rect 11651 36348 11652 36412
rect 11716 36348 11717 36412
rect 11651 36347 11717 36348
rect 11654 2141 11714 36347
rect 11838 34127 11898 66539
rect 11835 34126 11901 34127
rect 11835 34062 11836 34126
rect 11900 34062 11901 34126
rect 11835 34061 11901 34062
rect 11835 25804 11901 25805
rect 11835 25740 11836 25804
rect 11900 25740 11901 25804
rect 11835 25739 11901 25740
rect 11838 2685 11898 25739
rect 12952 6866 13300 6908
rect 12952 6630 13008 6866
rect 13244 6630 13300 6866
rect 12952 6588 13300 6630
rect 106656 6866 107004 6908
rect 106656 6630 106712 6866
rect 106948 6630 107004 6866
rect 106656 6588 107004 6630
rect 110036 6866 110356 82630
rect 110036 6630 110078 6866
rect 110314 6630 110356 6866
rect 12272 6206 12620 6248
rect 12272 5970 12328 6206
rect 12564 5970 12620 6206
rect 12272 5928 12620 5970
rect 107336 6206 107684 6248
rect 107336 5970 107392 6206
rect 107628 5970 107684 6206
rect 107336 5928 107684 5970
rect 17856 3909 17916 4080
rect 17853 3908 17919 3909
rect 17853 3844 17854 3908
rect 17918 3844 17919 3908
rect 17853 3843 17919 3844
rect 27512 3770 27572 4080
rect 28736 3773 28796 4080
rect 29824 3773 29884 4080
rect 27478 3710 27572 3770
rect 28733 3772 28799 3773
rect 11835 2684 11901 2685
rect 11835 2620 11836 2684
rect 11900 2620 11901 2684
rect 11835 2619 11901 2620
rect 11651 2140 11717 2141
rect 11651 2076 11652 2140
rect 11716 2076 11717 2140
rect 11651 2075 11717 2076
rect 10944 1120 11264 2004
rect 10944 1056 10952 1120
rect 11016 1056 11032 1120
rect 11096 1056 11112 1120
rect 11176 1056 11192 1120
rect 11256 1056 11264 1120
rect 10731 644 10797 645
rect 10731 580 10732 644
rect 10796 580 10797 644
rect 10731 579 10797 580
rect 10004 -390 10046 -154
rect 10282 -390 10324 -154
rect 10004 -1092 10324 -390
rect 10944 -814 11264 1056
rect 10944 -1050 10986 -814
rect 11222 -1050 11264 -814
rect 10944 -1092 11264 -1050
rect 11604 1664 11924 2004
rect 11604 1600 11612 1664
rect 11676 1600 11692 1664
rect 11756 1600 11772 1664
rect 11836 1600 11852 1664
rect 11916 1600 11924 1664
rect 11604 -154 11924 1600
rect 11604 -390 11646 -154
rect 11882 -390 11924 -154
rect 11604 -1092 11924 -390
rect 12544 1120 12864 2004
rect 12544 1056 12552 1120
rect 12616 1056 12632 1120
rect 12696 1056 12712 1120
rect 12776 1056 12792 1120
rect 12856 1056 12864 1120
rect 12544 -814 12864 1056
rect 12544 -1050 12586 -814
rect 12822 -1050 12864 -814
rect 12544 -1092 12864 -1050
rect 13204 1664 13524 2004
rect 13204 1600 13212 1664
rect 13276 1600 13292 1664
rect 13356 1600 13372 1664
rect 13436 1600 13452 1664
rect 13516 1600 13524 1664
rect 13204 -154 13524 1600
rect 13204 -390 13246 -154
rect 13482 -390 13524 -154
rect 13204 -1092 13524 -390
rect 14144 1120 14464 2004
rect 14144 1056 14152 1120
rect 14216 1056 14232 1120
rect 14296 1056 14312 1120
rect 14376 1056 14392 1120
rect 14456 1056 14464 1120
rect 14144 -814 14464 1056
rect 14144 -1050 14186 -814
rect 14422 -1050 14464 -814
rect 14144 -1092 14464 -1050
rect 14804 1664 15124 2004
rect 14804 1600 14812 1664
rect 14876 1600 14892 1664
rect 14956 1600 14972 1664
rect 15036 1600 15052 1664
rect 15116 1600 15124 1664
rect 14804 -154 15124 1600
rect 14804 -390 14846 -154
rect 15082 -390 15124 -154
rect 14804 -1092 15124 -390
rect 15744 1120 16064 2004
rect 15744 1056 15752 1120
rect 15816 1056 15832 1120
rect 15896 1056 15912 1120
rect 15976 1056 15992 1120
rect 16056 1056 16064 1120
rect 15744 -814 16064 1056
rect 15744 -1050 15786 -814
rect 16022 -1050 16064 -814
rect 15744 -1092 16064 -1050
rect 16404 1664 16724 2004
rect 16404 1600 16412 1664
rect 16476 1600 16492 1664
rect 16556 1600 16572 1664
rect 16636 1600 16652 1664
rect 16716 1600 16724 1664
rect 16404 -154 16724 1600
rect 16404 -390 16446 -154
rect 16682 -390 16724 -154
rect 16404 -1092 16724 -390
rect 17344 1120 17664 2004
rect 17344 1056 17352 1120
rect 17416 1056 17432 1120
rect 17496 1056 17512 1120
rect 17576 1056 17592 1120
rect 17656 1056 17664 1120
rect 17344 -814 17664 1056
rect 17344 -1050 17386 -814
rect 17622 -1050 17664 -814
rect 17344 -1092 17664 -1050
rect 18004 1664 18324 1880
rect 18004 1600 18012 1664
rect 18076 1600 18092 1664
rect 18156 1600 18172 1664
rect 18236 1600 18252 1664
rect 18316 1600 18324 1664
rect 18004 -154 18324 1600
rect 18004 -390 18046 -154
rect 18282 -390 18324 -154
rect 18004 -1092 18324 -390
rect 18944 1120 19264 2004
rect 18944 1056 18952 1120
rect 19016 1056 19032 1120
rect 19096 1056 19112 1120
rect 19176 1056 19192 1120
rect 19256 1056 19264 1120
rect 18944 -814 19264 1056
rect 18944 -1050 18986 -814
rect 19222 -1050 19264 -814
rect 18944 -1092 19264 -1050
rect 19604 1664 19924 2004
rect 19604 1600 19612 1664
rect 19676 1600 19692 1664
rect 19756 1600 19772 1664
rect 19836 1600 19852 1664
rect 19916 1600 19924 1664
rect 19604 -154 19924 1600
rect 19604 -390 19646 -154
rect 19882 -390 19924 -154
rect 19604 -1092 19924 -390
rect 20544 1120 20864 2004
rect 20544 1056 20552 1120
rect 20616 1056 20632 1120
rect 20696 1056 20712 1120
rect 20776 1056 20792 1120
rect 20856 1056 20864 1120
rect 20544 -814 20864 1056
rect 20544 -1050 20586 -814
rect 20822 -1050 20864 -814
rect 20544 -1092 20864 -1050
rect 21204 1664 21524 2004
rect 21204 1600 21212 1664
rect 21276 1600 21292 1664
rect 21356 1600 21372 1664
rect 21436 1600 21452 1664
rect 21516 1600 21524 1664
rect 21204 -154 21524 1600
rect 21204 -390 21246 -154
rect 21482 -390 21524 -154
rect 21204 -1092 21524 -390
rect 22144 1120 22464 2004
rect 22144 1056 22152 1120
rect 22216 1056 22232 1120
rect 22296 1056 22312 1120
rect 22376 1056 22392 1120
rect 22456 1056 22464 1120
rect 22144 -814 22464 1056
rect 22144 -1050 22186 -814
rect 22422 -1050 22464 -814
rect 22144 -1092 22464 -1050
rect 22804 1664 23124 2004
rect 22804 1600 22812 1664
rect 22876 1600 22892 1664
rect 22956 1600 22972 1664
rect 23036 1600 23052 1664
rect 23116 1600 23124 1664
rect 22804 -154 23124 1600
rect 22804 -390 22846 -154
rect 23082 -390 23124 -154
rect 22804 -1092 23124 -390
rect 23744 1120 24064 2004
rect 23744 1056 23752 1120
rect 23816 1056 23832 1120
rect 23896 1056 23912 1120
rect 23976 1056 23992 1120
rect 24056 1056 24064 1120
rect 23744 -814 24064 1056
rect 23744 -1050 23786 -814
rect 24022 -1050 24064 -814
rect 23744 -1092 24064 -1050
rect 24404 1664 24724 2004
rect 24404 1600 24412 1664
rect 24476 1600 24492 1664
rect 24556 1600 24572 1664
rect 24636 1600 24652 1664
rect 24716 1600 24724 1664
rect 24404 -154 24724 1600
rect 24404 -390 24446 -154
rect 24682 -390 24724 -154
rect 24404 -1092 24724 -390
rect 25344 1120 25664 2004
rect 25344 1056 25352 1120
rect 25416 1056 25432 1120
rect 25496 1056 25512 1120
rect 25576 1056 25592 1120
rect 25656 1056 25664 1120
rect 25344 -814 25664 1056
rect 25344 -1050 25386 -814
rect 25622 -1050 25664 -814
rect 25344 -1092 25664 -1050
rect 26004 1664 26324 2004
rect 26004 1600 26012 1664
rect 26076 1600 26092 1664
rect 26156 1600 26172 1664
rect 26236 1600 26252 1664
rect 26316 1600 26324 1664
rect 26004 -154 26324 1600
rect 26004 -390 26046 -154
rect 26282 -390 26324 -154
rect 26004 -1092 26324 -390
rect 26944 1120 27264 2004
rect 26944 1056 26952 1120
rect 27016 1056 27032 1120
rect 27096 1056 27112 1120
rect 27176 1056 27192 1120
rect 27256 1056 27264 1120
rect 26944 -814 27264 1056
rect 27478 645 27538 3710
rect 28733 3708 28734 3772
rect 28798 3708 28799 3772
rect 28733 3707 28799 3708
rect 29821 3772 29887 3773
rect 29821 3708 29822 3772
rect 29886 3708 29887 3772
rect 31184 3770 31244 4080
rect 32136 3770 32196 4080
rect 33360 3770 33420 4080
rect 34584 3770 34644 4080
rect 35672 3770 35732 4080
rect 31184 3710 31402 3770
rect 29821 3707 29887 3708
rect 27604 1664 27924 1880
rect 27604 1600 27612 1664
rect 27676 1600 27692 1664
rect 27756 1600 27772 1664
rect 27836 1600 27852 1664
rect 27916 1600 27924 1664
rect 27475 644 27541 645
rect 27475 580 27476 644
rect 27540 580 27541 644
rect 27475 579 27541 580
rect 26944 -1050 26986 -814
rect 27222 -1050 27264 -814
rect 26944 -1092 27264 -1050
rect 27604 -154 27924 1600
rect 27604 -390 27646 -154
rect 27882 -390 27924 -154
rect 27604 -1092 27924 -390
rect 28544 1120 28864 1880
rect 28544 1056 28552 1120
rect 28616 1056 28632 1120
rect 28696 1056 28712 1120
rect 28776 1056 28792 1120
rect 28856 1056 28864 1120
rect 28544 -814 28864 1056
rect 28544 -1050 28586 -814
rect 28822 -1050 28864 -814
rect 28544 -1092 28864 -1050
rect 29204 1664 29524 2004
rect 29204 1600 29212 1664
rect 29276 1600 29292 1664
rect 29356 1600 29372 1664
rect 29436 1600 29452 1664
rect 29516 1600 29524 1664
rect 29204 -154 29524 1600
rect 29204 -390 29246 -154
rect 29482 -390 29524 -154
rect 29204 -1092 29524 -390
rect 30144 1120 30464 2004
rect 30144 1056 30152 1120
rect 30216 1056 30232 1120
rect 30296 1056 30312 1120
rect 30376 1056 30392 1120
rect 30456 1056 30464 1120
rect 30144 -814 30464 1056
rect 30144 -1050 30186 -814
rect 30422 -1050 30464 -814
rect 30144 -1092 30464 -1050
rect 30804 1664 31124 1880
rect 30804 1600 30812 1664
rect 30876 1600 30892 1664
rect 30956 1600 30972 1664
rect 31036 1600 31052 1664
rect 31116 1600 31124 1664
rect 30804 -154 31124 1600
rect 31342 1325 31402 3710
rect 32078 3710 32196 3770
rect 33182 3710 33420 3770
rect 34470 3710 34644 3770
rect 35574 3710 35732 3770
rect 37032 3770 37092 4080
rect 38120 3770 38180 4080
rect 39208 3909 39268 4080
rect 40296 3909 40356 4080
rect 39205 3908 39271 3909
rect 39205 3844 39206 3908
rect 39270 3844 39271 3908
rect 39205 3843 39271 3844
rect 40293 3908 40359 3909
rect 40293 3844 40294 3908
rect 40358 3844 40359 3908
rect 40293 3843 40359 3844
rect 37032 3710 37106 3770
rect 32078 2413 32138 3710
rect 32075 2412 32141 2413
rect 32075 2348 32076 2412
rect 32140 2348 32141 2412
rect 32075 2347 32141 2348
rect 31339 1324 31405 1325
rect 31339 1260 31340 1324
rect 31404 1260 31405 1324
rect 31339 1259 31405 1260
rect 30804 -390 30846 -154
rect 31082 -390 31124 -154
rect 30804 -1092 31124 -390
rect 31744 1120 32064 1880
rect 31744 1056 31752 1120
rect 31816 1056 31832 1120
rect 31896 1056 31912 1120
rect 31976 1056 31992 1120
rect 32056 1056 32064 1120
rect 31744 -814 32064 1056
rect 31744 -1050 31786 -814
rect 32022 -1050 32064 -814
rect 31744 -1092 32064 -1050
rect 32404 1664 32724 2004
rect 32404 1600 32412 1664
rect 32476 1600 32492 1664
rect 32556 1600 32572 1664
rect 32636 1600 32652 1664
rect 32716 1600 32724 1664
rect 32404 -154 32724 1600
rect 33182 1325 33242 3710
rect 33179 1324 33245 1325
rect 33179 1260 33180 1324
rect 33244 1260 33245 1324
rect 33179 1259 33245 1260
rect 32404 -390 32446 -154
rect 32682 -390 32724 -154
rect 32404 -1092 32724 -390
rect 33344 1120 33664 1880
rect 33344 1056 33352 1120
rect 33416 1056 33432 1120
rect 33496 1056 33512 1120
rect 33576 1056 33592 1120
rect 33656 1056 33664 1120
rect 33344 -814 33664 1056
rect 33344 -1050 33386 -814
rect 33622 -1050 33664 -814
rect 33344 -1092 33664 -1050
rect 34004 1664 34324 2004
rect 34004 1600 34012 1664
rect 34076 1600 34092 1664
rect 34156 1600 34172 1664
rect 34236 1600 34252 1664
rect 34316 1600 34324 1664
rect 34004 -154 34324 1600
rect 34470 1325 34530 3710
rect 35574 2685 35634 3710
rect 37046 2685 37106 3710
rect 37966 3710 38180 3770
rect 41656 3770 41716 4080
rect 42744 3770 42804 4080
rect 43832 3770 43892 4080
rect 45056 3909 45116 4080
rect 46144 3909 46204 4080
rect 45053 3908 45119 3909
rect 45053 3844 45054 3908
rect 45118 3844 45119 3908
rect 45053 3843 45119 3844
rect 46141 3908 46207 3909
rect 46141 3844 46142 3908
rect 46206 3844 46207 3908
rect 46141 3843 46207 3844
rect 47504 3773 47564 4080
rect 47501 3772 47567 3773
rect 41656 3710 41890 3770
rect 42744 3710 42810 3770
rect 43832 3710 43914 3770
rect 35571 2684 35637 2685
rect 35571 2620 35572 2684
rect 35636 2620 35637 2684
rect 35571 2619 35637 2620
rect 37043 2684 37109 2685
rect 37043 2620 37044 2684
rect 37108 2620 37109 2684
rect 37043 2619 37109 2620
rect 34467 1324 34533 1325
rect 34467 1260 34468 1324
rect 34532 1260 34533 1324
rect 34467 1259 34533 1260
rect 34004 -390 34046 -154
rect 34282 -390 34324 -154
rect 34004 -1092 34324 -390
rect 34944 1120 35264 2004
rect 34944 1056 34952 1120
rect 35016 1056 35032 1120
rect 35096 1056 35112 1120
rect 35176 1056 35192 1120
rect 35256 1056 35264 1120
rect 34944 -814 35264 1056
rect 34944 -1050 34986 -814
rect 35222 -1050 35264 -814
rect 34944 -1092 35264 -1050
rect 35604 1664 35924 1880
rect 35604 1600 35612 1664
rect 35676 1600 35692 1664
rect 35756 1600 35772 1664
rect 35836 1600 35852 1664
rect 35916 1600 35924 1664
rect 35604 -154 35924 1600
rect 35604 -390 35646 -154
rect 35882 -390 35924 -154
rect 35604 -1092 35924 -390
rect 36544 1120 36864 2004
rect 36544 1056 36552 1120
rect 36616 1056 36632 1120
rect 36696 1056 36712 1120
rect 36776 1056 36792 1120
rect 36856 1056 36864 1120
rect 36544 -814 36864 1056
rect 36544 -1050 36586 -814
rect 36822 -1050 36864 -814
rect 36544 -1092 36864 -1050
rect 37204 1664 37524 1880
rect 37204 1600 37212 1664
rect 37276 1600 37292 1664
rect 37356 1600 37372 1664
rect 37436 1600 37452 1664
rect 37516 1600 37524 1664
rect 37204 -154 37524 1600
rect 37966 1325 38026 3710
rect 37963 1324 38029 1325
rect 37963 1260 37964 1324
rect 38028 1260 38029 1324
rect 37963 1259 38029 1260
rect 37204 -390 37246 -154
rect 37482 -390 37524 -154
rect 37204 -1092 37524 -390
rect 38144 1120 38464 1880
rect 38144 1056 38152 1120
rect 38216 1056 38232 1120
rect 38296 1056 38312 1120
rect 38376 1056 38392 1120
rect 38456 1056 38464 1120
rect 38144 -814 38464 1056
rect 38144 -1050 38186 -814
rect 38422 -1050 38464 -814
rect 38144 -1092 38464 -1050
rect 38804 1664 39124 1880
rect 38804 1600 38812 1664
rect 38876 1600 38892 1664
rect 38956 1600 38972 1664
rect 39036 1600 39052 1664
rect 39116 1600 39124 1664
rect 38804 -154 39124 1600
rect 38804 -390 38846 -154
rect 39082 -390 39124 -154
rect 38804 -1092 39124 -390
rect 39744 1120 40064 1880
rect 39744 1056 39752 1120
rect 39816 1056 39832 1120
rect 39896 1056 39912 1120
rect 39976 1056 39992 1120
rect 40056 1056 40064 1120
rect 39744 -814 40064 1056
rect 39744 -1050 39786 -814
rect 40022 -1050 40064 -814
rect 39744 -1092 40064 -1050
rect 40404 1664 40724 1880
rect 40404 1600 40412 1664
rect 40476 1600 40492 1664
rect 40556 1600 40572 1664
rect 40636 1600 40652 1664
rect 40716 1600 40724 1664
rect 40404 -154 40724 1600
rect 40404 -390 40446 -154
rect 40682 -390 40724 -154
rect 40404 -1092 40724 -390
rect 41344 1120 41664 1880
rect 41344 1056 41352 1120
rect 41416 1056 41432 1120
rect 41496 1056 41512 1120
rect 41576 1056 41592 1120
rect 41656 1056 41664 1120
rect 41344 -814 41664 1056
rect 41830 509 41890 3710
rect 42750 2413 42810 3710
rect 43854 2413 43914 3710
rect 47501 3708 47502 3772
rect 47566 3708 47567 3772
rect 48592 3770 48652 4080
rect 49680 3770 49740 4080
rect 50904 3909 50964 4080
rect 50901 3908 50967 3909
rect 50901 3844 50902 3908
rect 50966 3844 50967 3908
rect 50901 3843 50967 3844
rect 52264 3770 52324 4080
rect 53352 3770 53412 4080
rect 54440 3909 54500 4080
rect 54437 3908 54503 3909
rect 54437 3844 54438 3908
rect 54502 3844 54503 3908
rect 54437 3843 54503 3844
rect 55528 3770 55588 4080
rect 48592 3710 48698 3770
rect 49680 3710 49802 3770
rect 52264 3710 52378 3770
rect 47501 3707 47567 3708
rect 48638 2413 48698 3710
rect 49742 2685 49802 3710
rect 49739 2684 49805 2685
rect 49739 2620 49740 2684
rect 49804 2620 49805 2684
rect 49739 2619 49805 2620
rect 42747 2412 42813 2413
rect 42747 2348 42748 2412
rect 42812 2348 42813 2412
rect 42747 2347 42813 2348
rect 43851 2412 43917 2413
rect 43851 2348 43852 2412
rect 43916 2348 43917 2412
rect 43851 2347 43917 2348
rect 48635 2412 48701 2413
rect 48635 2348 48636 2412
rect 48700 2348 48701 2412
rect 48635 2347 48701 2348
rect 42004 1664 42324 1880
rect 42004 1600 42012 1664
rect 42076 1600 42092 1664
rect 42156 1600 42172 1664
rect 42236 1600 42252 1664
rect 42316 1600 42324 1664
rect 41827 508 41893 509
rect 41827 444 41828 508
rect 41892 444 41893 508
rect 41827 443 41893 444
rect 41344 -1050 41386 -814
rect 41622 -1050 41664 -814
rect 41344 -1092 41664 -1050
rect 42004 -154 42324 1600
rect 42004 -390 42046 -154
rect 42282 -390 42324 -154
rect 42004 -1092 42324 -390
rect 42944 1120 43264 2004
rect 42944 1056 42952 1120
rect 43016 1056 43032 1120
rect 43096 1056 43112 1120
rect 43176 1056 43192 1120
rect 43256 1056 43264 1120
rect 42944 -814 43264 1056
rect 42944 -1050 42986 -814
rect 43222 -1050 43264 -814
rect 42944 -1092 43264 -1050
rect 43604 1664 43924 1880
rect 43604 1600 43612 1664
rect 43676 1600 43692 1664
rect 43756 1600 43772 1664
rect 43836 1600 43852 1664
rect 43916 1600 43924 1664
rect 43604 -154 43924 1600
rect 43604 -390 43646 -154
rect 43882 -390 43924 -154
rect 43604 -1092 43924 -390
rect 44544 1120 44864 2004
rect 44544 1056 44552 1120
rect 44616 1056 44632 1120
rect 44696 1056 44712 1120
rect 44776 1056 44792 1120
rect 44856 1056 44864 1120
rect 44544 -814 44864 1056
rect 44544 -1050 44586 -814
rect 44822 -1050 44864 -814
rect 44544 -1092 44864 -1050
rect 45204 1664 45524 1880
rect 45204 1600 45212 1664
rect 45276 1600 45292 1664
rect 45356 1600 45372 1664
rect 45436 1600 45452 1664
rect 45516 1600 45524 1664
rect 45204 -154 45524 1600
rect 45204 -390 45246 -154
rect 45482 -390 45524 -154
rect 45204 -1092 45524 -390
rect 46144 1120 46464 1880
rect 46144 1056 46152 1120
rect 46216 1056 46232 1120
rect 46296 1056 46312 1120
rect 46376 1056 46392 1120
rect 46456 1056 46464 1120
rect 46144 -814 46464 1056
rect 46144 -1050 46186 -814
rect 46422 -1050 46464 -814
rect 46144 -1092 46464 -1050
rect 46804 1664 47124 2004
rect 46804 1600 46812 1664
rect 46876 1600 46892 1664
rect 46956 1600 46972 1664
rect 47036 1600 47052 1664
rect 47116 1600 47124 1664
rect 46804 -154 47124 1600
rect 46804 -390 46846 -154
rect 47082 -390 47124 -154
rect 46804 -1092 47124 -390
rect 47744 1120 48064 1880
rect 47744 1056 47752 1120
rect 47816 1056 47832 1120
rect 47896 1056 47912 1120
rect 47976 1056 47992 1120
rect 48056 1056 48064 1120
rect 47744 -814 48064 1056
rect 47744 -1050 47786 -814
rect 48022 -1050 48064 -814
rect 47744 -1092 48064 -1050
rect 48404 1664 48724 1880
rect 48404 1600 48412 1664
rect 48476 1600 48492 1664
rect 48556 1600 48572 1664
rect 48636 1600 48652 1664
rect 48716 1600 48724 1664
rect 48404 -154 48724 1600
rect 48404 -390 48446 -154
rect 48682 -390 48724 -154
rect 48404 -1092 48724 -390
rect 49344 1120 49664 1880
rect 49344 1056 49352 1120
rect 49416 1056 49432 1120
rect 49496 1056 49512 1120
rect 49576 1056 49592 1120
rect 49656 1056 49664 1120
rect 49344 -814 49664 1056
rect 49344 -1050 49386 -814
rect 49622 -1050 49664 -814
rect 49344 -1092 49664 -1050
rect 50004 1664 50324 1880
rect 50004 1600 50012 1664
rect 50076 1600 50092 1664
rect 50156 1600 50172 1664
rect 50236 1600 50252 1664
rect 50316 1600 50324 1664
rect 50004 -154 50324 1600
rect 50004 -390 50046 -154
rect 50282 -390 50324 -154
rect 50004 -1092 50324 -390
rect 50944 1120 51264 1880
rect 50944 1056 50952 1120
rect 51016 1056 51032 1120
rect 51096 1056 51112 1120
rect 51176 1056 51192 1120
rect 51256 1056 51264 1120
rect 50944 -814 51264 1056
rect 50944 -1050 50986 -814
rect 51222 -1050 51264 -814
rect 50944 -1092 51264 -1050
rect 51604 1664 51924 2004
rect 51604 1600 51612 1664
rect 51676 1600 51692 1664
rect 51756 1600 51772 1664
rect 51836 1600 51852 1664
rect 51916 1600 51924 1664
rect 51604 -154 51924 1600
rect 52318 645 52378 3710
rect 53054 3710 53412 3770
rect 55446 3710 55588 3770
rect 56888 3770 56948 4080
rect 57976 3770 58036 4080
rect 59064 3770 59124 4080
rect 60288 3770 60348 4080
rect 61376 3770 61436 4080
rect 62736 3770 62796 4080
rect 63824 3770 63884 4080
rect 64912 3770 64972 4080
rect 66000 3770 66060 4080
rect 56888 3710 56978 3770
rect 57976 3710 58082 3770
rect 52544 1120 52864 1880
rect 52544 1056 52552 1120
rect 52616 1056 52632 1120
rect 52696 1056 52712 1120
rect 52776 1056 52792 1120
rect 52856 1056 52864 1120
rect 52315 644 52381 645
rect 52315 580 52316 644
rect 52380 580 52381 644
rect 52315 579 52381 580
rect 51604 -390 51646 -154
rect 51882 -390 51924 -154
rect 51604 -1092 51924 -390
rect 52544 -814 52864 1056
rect 53054 917 53114 3710
rect 55446 2685 55506 3710
rect 55443 2684 55509 2685
rect 55443 2620 55444 2684
rect 55508 2620 55509 2684
rect 55443 2619 55509 2620
rect 53204 1664 53524 1880
rect 53204 1600 53212 1664
rect 53276 1600 53292 1664
rect 53356 1600 53372 1664
rect 53436 1600 53452 1664
rect 53516 1600 53524 1664
rect 53051 916 53117 917
rect 53051 852 53052 916
rect 53116 852 53117 916
rect 53051 851 53117 852
rect 52544 -1050 52586 -814
rect 52822 -1050 52864 -814
rect 52544 -1092 52864 -1050
rect 53204 -154 53524 1600
rect 53204 -390 53246 -154
rect 53482 -390 53524 -154
rect 53204 -1092 53524 -390
rect 54144 1120 54464 1880
rect 54144 1056 54152 1120
rect 54216 1056 54232 1120
rect 54296 1056 54312 1120
rect 54376 1056 54392 1120
rect 54456 1056 54464 1120
rect 54144 -814 54464 1056
rect 54144 -1050 54186 -814
rect 54422 -1050 54464 -814
rect 54144 -1092 54464 -1050
rect 54804 1664 55124 1880
rect 54804 1600 54812 1664
rect 54876 1600 54892 1664
rect 54956 1600 54972 1664
rect 55036 1600 55052 1664
rect 55116 1600 55124 1664
rect 54804 -154 55124 1600
rect 54804 -390 54846 -154
rect 55082 -390 55124 -154
rect 54804 -1092 55124 -390
rect 55744 1120 56064 2004
rect 55744 1056 55752 1120
rect 55816 1056 55832 1120
rect 55896 1056 55912 1120
rect 55976 1056 55992 1120
rect 56056 1056 56064 1120
rect 55744 -814 56064 1056
rect 55744 -1050 55786 -814
rect 56022 -1050 56064 -814
rect 55744 -1092 56064 -1050
rect 56404 1664 56724 1880
rect 56404 1600 56412 1664
rect 56476 1600 56492 1664
rect 56556 1600 56572 1664
rect 56636 1600 56652 1664
rect 56716 1600 56724 1664
rect 56404 -154 56724 1600
rect 56918 1325 56978 3710
rect 58022 2685 58082 3710
rect 58758 3710 59124 3770
rect 60230 3710 60348 3770
rect 60966 3710 61436 3770
rect 62622 3710 62796 3770
rect 63542 3710 63884 3770
rect 64646 3710 64972 3770
rect 65750 3710 66060 3770
rect 67224 3770 67284 4080
rect 68584 3770 68644 4080
rect 69672 3770 69732 4080
rect 93899 3908 93965 3909
rect 93899 3844 93900 3908
rect 93964 3844 93965 3908
rect 93899 3843 93965 3844
rect 67224 3710 67466 3770
rect 58019 2684 58085 2685
rect 58019 2620 58020 2684
rect 58084 2620 58085 2684
rect 58019 2619 58085 2620
rect 56915 1324 56981 1325
rect 56915 1260 56916 1324
rect 56980 1260 56981 1324
rect 56915 1259 56981 1260
rect 56404 -390 56446 -154
rect 56682 -390 56724 -154
rect 56404 -1092 56724 -390
rect 57344 1120 57664 1880
rect 57344 1056 57352 1120
rect 57416 1056 57432 1120
rect 57496 1056 57512 1120
rect 57576 1056 57592 1120
rect 57656 1056 57664 1120
rect 57344 -814 57664 1056
rect 57344 -1050 57386 -814
rect 57622 -1050 57664 -814
rect 57344 -1092 57664 -1050
rect 58004 1664 58324 1880
rect 58004 1600 58012 1664
rect 58076 1600 58092 1664
rect 58156 1600 58172 1664
rect 58236 1600 58252 1664
rect 58316 1600 58324 1664
rect 58004 -154 58324 1600
rect 58758 1325 58818 3710
rect 58755 1324 58821 1325
rect 58755 1260 58756 1324
rect 58820 1260 58821 1324
rect 58755 1259 58821 1260
rect 58004 -390 58046 -154
rect 58282 -390 58324 -154
rect 58004 -1092 58324 -390
rect 58944 1120 59264 1880
rect 58944 1056 58952 1120
rect 59016 1056 59032 1120
rect 59096 1056 59112 1120
rect 59176 1056 59192 1120
rect 59256 1056 59264 1120
rect 58944 -814 59264 1056
rect 58944 -1050 58986 -814
rect 59222 -1050 59264 -814
rect 58944 -1092 59264 -1050
rect 59604 1664 59924 1880
rect 59604 1600 59612 1664
rect 59676 1600 59692 1664
rect 59756 1600 59772 1664
rect 59836 1600 59852 1664
rect 59916 1600 59924 1664
rect 59604 -154 59924 1600
rect 60230 1325 60290 3710
rect 60227 1324 60293 1325
rect 60227 1260 60228 1324
rect 60292 1260 60293 1324
rect 60227 1259 60293 1260
rect 59604 -390 59646 -154
rect 59882 -390 59924 -154
rect 59604 -1092 59924 -390
rect 60544 1120 60864 2004
rect 60966 1325 61026 3710
rect 61204 1664 61524 1880
rect 61204 1600 61212 1664
rect 61276 1600 61292 1664
rect 61356 1600 61372 1664
rect 61436 1600 61452 1664
rect 61516 1600 61524 1664
rect 60963 1324 61029 1325
rect 60963 1260 60964 1324
rect 61028 1260 61029 1324
rect 60963 1259 61029 1260
rect 60544 1056 60552 1120
rect 60616 1056 60632 1120
rect 60696 1056 60712 1120
rect 60776 1056 60792 1120
rect 60856 1056 60864 1120
rect 60544 -814 60864 1056
rect 60544 -1050 60586 -814
rect 60822 -1050 60864 -814
rect 60544 -1092 60864 -1050
rect 61204 -154 61524 1600
rect 61204 -390 61246 -154
rect 61482 -390 61524 -154
rect 61204 -1092 61524 -390
rect 62144 1120 62464 2004
rect 62622 1325 62682 3710
rect 62804 1664 63124 1880
rect 62804 1600 62812 1664
rect 62876 1600 62892 1664
rect 62956 1600 62972 1664
rect 63036 1600 63052 1664
rect 63116 1600 63124 1664
rect 62619 1324 62685 1325
rect 62619 1260 62620 1324
rect 62684 1260 62685 1324
rect 62619 1259 62685 1260
rect 62144 1056 62152 1120
rect 62216 1056 62232 1120
rect 62296 1056 62312 1120
rect 62376 1056 62392 1120
rect 62456 1056 62464 1120
rect 62144 -814 62464 1056
rect 62144 -1050 62186 -814
rect 62422 -1050 62464 -814
rect 62144 -1092 62464 -1050
rect 62804 -154 63124 1600
rect 63542 1325 63602 3710
rect 64646 2410 64706 3710
rect 64646 2350 65074 2410
rect 63539 1324 63605 1325
rect 63539 1260 63540 1324
rect 63604 1260 63605 1324
rect 63539 1259 63605 1260
rect 62804 -390 62846 -154
rect 63082 -390 63124 -154
rect 62804 -1092 63124 -390
rect 63744 1120 64064 1880
rect 63744 1056 63752 1120
rect 63816 1056 63832 1120
rect 63896 1056 63912 1120
rect 63976 1056 63992 1120
rect 64056 1056 64064 1120
rect 63744 -814 64064 1056
rect 63744 -1050 63786 -814
rect 64022 -1050 64064 -814
rect 63744 -1092 64064 -1050
rect 64404 1664 64724 2004
rect 64404 1600 64412 1664
rect 64476 1600 64492 1664
rect 64556 1600 64572 1664
rect 64636 1600 64652 1664
rect 64716 1600 64724 1664
rect 64404 -154 64724 1600
rect 65014 1325 65074 2350
rect 65011 1324 65077 1325
rect 65011 1260 65012 1324
rect 65076 1260 65077 1324
rect 65011 1259 65077 1260
rect 64404 -390 64446 -154
rect 64682 -390 64724 -154
rect 64404 -1092 64724 -390
rect 65344 1120 65664 1880
rect 65750 1325 65810 3710
rect 66004 1664 66324 1880
rect 66004 1600 66012 1664
rect 66076 1600 66092 1664
rect 66156 1600 66172 1664
rect 66236 1600 66252 1664
rect 66316 1600 66324 1664
rect 65747 1324 65813 1325
rect 65747 1260 65748 1324
rect 65812 1260 65813 1324
rect 65747 1259 65813 1260
rect 65344 1056 65352 1120
rect 65416 1056 65432 1120
rect 65496 1056 65512 1120
rect 65576 1056 65592 1120
rect 65656 1056 65664 1120
rect 65344 -814 65664 1056
rect 65344 -1050 65386 -814
rect 65622 -1050 65664 -814
rect 65344 -1092 65664 -1050
rect 66004 -154 66324 1600
rect 66004 -390 66046 -154
rect 66282 -390 66324 -154
rect 66004 -1092 66324 -390
rect 66944 1120 67264 1880
rect 67406 1325 67466 3710
rect 68326 3710 68644 3770
rect 69614 3710 69732 3770
rect 67604 1664 67924 1880
rect 67604 1600 67612 1664
rect 67676 1600 67692 1664
rect 67756 1600 67772 1664
rect 67836 1600 67852 1664
rect 67916 1600 67924 1664
rect 67403 1324 67469 1325
rect 67403 1260 67404 1324
rect 67468 1260 67469 1324
rect 67403 1259 67469 1260
rect 66944 1056 66952 1120
rect 67016 1056 67032 1120
rect 67096 1056 67112 1120
rect 67176 1056 67192 1120
rect 67256 1056 67264 1120
rect 66944 -814 67264 1056
rect 66944 -1050 66986 -814
rect 67222 -1050 67264 -814
rect 66944 -1092 67264 -1050
rect 67604 -154 67924 1600
rect 68326 1325 68386 3710
rect 68323 1324 68389 1325
rect 68323 1260 68324 1324
rect 68388 1260 68389 1324
rect 68323 1259 68389 1260
rect 67604 -390 67646 -154
rect 67882 -390 67924 -154
rect 67604 -1092 67924 -390
rect 68544 1120 68864 1880
rect 68544 1056 68552 1120
rect 68616 1056 68632 1120
rect 68696 1056 68712 1120
rect 68776 1056 68792 1120
rect 68856 1056 68864 1120
rect 68544 -814 68864 1056
rect 68544 -1050 68586 -814
rect 68822 -1050 68864 -814
rect 68544 -1092 68864 -1050
rect 69204 1664 69524 2004
rect 69204 1600 69212 1664
rect 69276 1600 69292 1664
rect 69356 1600 69372 1664
rect 69436 1600 69452 1664
rect 69516 1600 69524 1664
rect 69204 -154 69524 1600
rect 69614 1325 69674 3710
rect 69611 1324 69677 1325
rect 69611 1260 69612 1324
rect 69676 1260 69677 1324
rect 69611 1259 69677 1260
rect 69204 -390 69246 -154
rect 69482 -390 69524 -154
rect 69204 -1092 69524 -390
rect 70144 1120 70464 2004
rect 70144 1056 70152 1120
rect 70216 1056 70232 1120
rect 70296 1056 70312 1120
rect 70376 1056 70392 1120
rect 70456 1056 70464 1120
rect 70144 -814 70464 1056
rect 70144 -1050 70186 -814
rect 70422 -1050 70464 -814
rect 70144 -1092 70464 -1050
rect 70804 1664 71124 2004
rect 70804 1600 70812 1664
rect 70876 1600 70892 1664
rect 70956 1600 70972 1664
rect 71036 1600 71052 1664
rect 71116 1600 71124 1664
rect 70804 -154 71124 1600
rect 70804 -390 70846 -154
rect 71082 -390 71124 -154
rect 70804 -1092 71124 -390
rect 71744 1120 72064 2004
rect 71744 1056 71752 1120
rect 71816 1056 71832 1120
rect 71896 1056 71912 1120
rect 71976 1056 71992 1120
rect 72056 1056 72064 1120
rect 71744 -814 72064 1056
rect 71744 -1050 71786 -814
rect 72022 -1050 72064 -814
rect 71744 -1092 72064 -1050
rect 72404 1664 72724 1880
rect 72404 1600 72412 1664
rect 72476 1600 72492 1664
rect 72556 1600 72572 1664
rect 72636 1600 72652 1664
rect 72716 1600 72724 1664
rect 72404 -154 72724 1600
rect 72404 -390 72446 -154
rect 72682 -390 72724 -154
rect 72404 -1092 72724 -390
rect 73344 1120 73664 2004
rect 73344 1056 73352 1120
rect 73416 1056 73432 1120
rect 73496 1056 73512 1120
rect 73576 1056 73592 1120
rect 73656 1056 73664 1120
rect 73344 -814 73664 1056
rect 73344 -1050 73386 -814
rect 73622 -1050 73664 -814
rect 73344 -1092 73664 -1050
rect 74004 1664 74324 1880
rect 74004 1600 74012 1664
rect 74076 1600 74092 1664
rect 74156 1600 74172 1664
rect 74236 1600 74252 1664
rect 74316 1600 74324 1664
rect 74004 -154 74324 1600
rect 74004 -390 74046 -154
rect 74282 -390 74324 -154
rect 74004 -1092 74324 -390
rect 74944 1120 75264 1880
rect 74944 1056 74952 1120
rect 75016 1056 75032 1120
rect 75096 1056 75112 1120
rect 75176 1056 75192 1120
rect 75256 1056 75264 1120
rect 74944 -814 75264 1056
rect 74944 -1050 74986 -814
rect 75222 -1050 75264 -814
rect 74944 -1092 75264 -1050
rect 75604 1664 75924 2004
rect 75604 1600 75612 1664
rect 75676 1600 75692 1664
rect 75756 1600 75772 1664
rect 75836 1600 75852 1664
rect 75916 1600 75924 1664
rect 75604 -154 75924 1600
rect 75604 -390 75646 -154
rect 75882 -390 75924 -154
rect 75604 -1092 75924 -390
rect 76544 1120 76864 2004
rect 76544 1056 76552 1120
rect 76616 1056 76632 1120
rect 76696 1056 76712 1120
rect 76776 1056 76792 1120
rect 76856 1056 76864 1120
rect 76544 -814 76864 1056
rect 76544 -1050 76586 -814
rect 76822 -1050 76864 -814
rect 76544 -1092 76864 -1050
rect 77204 1664 77524 1880
rect 77204 1600 77212 1664
rect 77276 1600 77292 1664
rect 77356 1600 77372 1664
rect 77436 1600 77452 1664
rect 77516 1600 77524 1664
rect 77204 -154 77524 1600
rect 77204 -390 77246 -154
rect 77482 -390 77524 -154
rect 77204 -1092 77524 -390
rect 78144 1120 78464 2004
rect 78144 1056 78152 1120
rect 78216 1056 78232 1120
rect 78296 1056 78312 1120
rect 78376 1056 78392 1120
rect 78456 1056 78464 1120
rect 78144 -814 78464 1056
rect 78144 -1050 78186 -814
rect 78422 -1050 78464 -814
rect 78144 -1092 78464 -1050
rect 78804 1664 79124 1880
rect 78804 1600 78812 1664
rect 78876 1600 78892 1664
rect 78956 1600 78972 1664
rect 79036 1600 79052 1664
rect 79116 1600 79124 1664
rect 78804 -154 79124 1600
rect 78804 -390 78846 -154
rect 79082 -390 79124 -154
rect 78804 -1092 79124 -390
rect 79744 1120 80064 2004
rect 79744 1056 79752 1120
rect 79816 1056 79832 1120
rect 79896 1056 79912 1120
rect 79976 1056 79992 1120
rect 80056 1056 80064 1120
rect 79744 -814 80064 1056
rect 79744 -1050 79786 -814
rect 80022 -1050 80064 -814
rect 79744 -1092 80064 -1050
rect 80404 1664 80724 2004
rect 80404 1600 80412 1664
rect 80476 1600 80492 1664
rect 80556 1600 80572 1664
rect 80636 1600 80652 1664
rect 80716 1600 80724 1664
rect 80404 -154 80724 1600
rect 80404 -390 80446 -154
rect 80682 -390 80724 -154
rect 80404 -1092 80724 -390
rect 81344 1120 81664 2004
rect 81344 1056 81352 1120
rect 81416 1056 81432 1120
rect 81496 1056 81512 1120
rect 81576 1056 81592 1120
rect 81656 1056 81664 1120
rect 81344 -814 81664 1056
rect 81344 -1050 81386 -814
rect 81622 -1050 81664 -814
rect 81344 -1092 81664 -1050
rect 82004 1664 82324 2004
rect 82004 1600 82012 1664
rect 82076 1600 82092 1664
rect 82156 1600 82172 1664
rect 82236 1600 82252 1664
rect 82316 1600 82324 1664
rect 82004 -154 82324 1600
rect 82004 -390 82046 -154
rect 82282 -390 82324 -154
rect 82004 -1092 82324 -390
rect 82944 1120 83264 2004
rect 82944 1056 82952 1120
rect 83016 1056 83032 1120
rect 83096 1056 83112 1120
rect 83176 1056 83192 1120
rect 83256 1056 83264 1120
rect 82944 -814 83264 1056
rect 82944 -1050 82986 -814
rect 83222 -1050 83264 -814
rect 82944 -1092 83264 -1050
rect 83604 1664 83924 2004
rect 83604 1600 83612 1664
rect 83676 1600 83692 1664
rect 83756 1600 83772 1664
rect 83836 1600 83852 1664
rect 83916 1600 83924 1664
rect 83604 -154 83924 1600
rect 83604 -390 83646 -154
rect 83882 -390 83924 -154
rect 83604 -1092 83924 -390
rect 84544 1120 84864 2004
rect 84544 1056 84552 1120
rect 84616 1056 84632 1120
rect 84696 1056 84712 1120
rect 84776 1056 84792 1120
rect 84856 1056 84864 1120
rect 84544 -814 84864 1056
rect 84544 -1050 84586 -814
rect 84822 -1050 84864 -814
rect 84544 -1092 84864 -1050
rect 85204 1664 85524 2004
rect 85204 1600 85212 1664
rect 85276 1600 85292 1664
rect 85356 1600 85372 1664
rect 85436 1600 85452 1664
rect 85516 1600 85524 1664
rect 85204 -154 85524 1600
rect 85204 -390 85246 -154
rect 85482 -390 85524 -154
rect 85204 -1092 85524 -390
rect 86144 1120 86464 2004
rect 86144 1056 86152 1120
rect 86216 1056 86232 1120
rect 86296 1056 86312 1120
rect 86376 1056 86392 1120
rect 86456 1056 86464 1120
rect 86144 -814 86464 1056
rect 86144 -1050 86186 -814
rect 86422 -1050 86464 -814
rect 86144 -1092 86464 -1050
rect 86804 1664 87124 2004
rect 86804 1600 86812 1664
rect 86876 1600 86892 1664
rect 86956 1600 86972 1664
rect 87036 1600 87052 1664
rect 87116 1600 87124 1664
rect 86804 -154 87124 1600
rect 86804 -390 86846 -154
rect 87082 -390 87124 -154
rect 86804 -1092 87124 -390
rect 87744 1120 88064 2004
rect 87744 1056 87752 1120
rect 87816 1056 87832 1120
rect 87896 1056 87912 1120
rect 87976 1056 87992 1120
rect 88056 1056 88064 1120
rect 87744 -814 88064 1056
rect 87744 -1050 87786 -814
rect 88022 -1050 88064 -814
rect 87744 -1092 88064 -1050
rect 88404 1664 88724 2004
rect 88404 1600 88412 1664
rect 88476 1600 88492 1664
rect 88556 1600 88572 1664
rect 88636 1600 88652 1664
rect 88716 1600 88724 1664
rect 88404 -154 88724 1600
rect 88404 -390 88446 -154
rect 88682 -390 88724 -154
rect 88404 -1092 88724 -390
rect 89344 1120 89664 2004
rect 89344 1056 89352 1120
rect 89416 1056 89432 1120
rect 89496 1056 89512 1120
rect 89576 1056 89592 1120
rect 89656 1056 89664 1120
rect 89344 -814 89664 1056
rect 89344 -1050 89386 -814
rect 89622 -1050 89664 -814
rect 89344 -1092 89664 -1050
rect 90004 1664 90324 2004
rect 90004 1600 90012 1664
rect 90076 1600 90092 1664
rect 90156 1600 90172 1664
rect 90236 1600 90252 1664
rect 90316 1600 90324 1664
rect 90004 -154 90324 1600
rect 90004 -390 90046 -154
rect 90282 -390 90324 -154
rect 90004 -1092 90324 -390
rect 90944 1120 91264 2004
rect 90944 1056 90952 1120
rect 91016 1056 91032 1120
rect 91096 1056 91112 1120
rect 91176 1056 91192 1120
rect 91256 1056 91264 1120
rect 90944 -814 91264 1056
rect 90944 -1050 90986 -814
rect 91222 -1050 91264 -814
rect 90944 -1092 91264 -1050
rect 91604 1664 91924 2004
rect 91604 1600 91612 1664
rect 91676 1600 91692 1664
rect 91756 1600 91772 1664
rect 91836 1600 91852 1664
rect 91916 1600 91924 1664
rect 91604 -154 91924 1600
rect 91604 -390 91646 -154
rect 91882 -390 91924 -154
rect 91604 -1092 91924 -390
rect 92544 1120 92864 2004
rect 92544 1056 92552 1120
rect 92616 1056 92632 1120
rect 92696 1056 92712 1120
rect 92776 1056 92792 1120
rect 92856 1056 92864 1120
rect 92544 -814 92864 1056
rect 92544 -1050 92586 -814
rect 92822 -1050 92864 -814
rect 92544 -1092 92864 -1050
rect 93204 1664 93524 2004
rect 93204 1600 93212 1664
rect 93276 1600 93292 1664
rect 93356 1600 93372 1664
rect 93436 1600 93452 1664
rect 93516 1600 93524 1664
rect 93204 -154 93524 1600
rect 93902 781 93962 3843
rect 94696 3770 94756 4080
rect 94832 3770 94892 4080
rect 94968 3909 95028 4080
rect 94965 3908 95031 3909
rect 94965 3844 94966 3908
rect 95030 3844 95031 3908
rect 94965 3843 95031 3844
rect 95104 3770 95164 4080
rect 94638 3710 94756 3770
rect 94822 3710 94892 3770
rect 95006 3710 95164 3770
rect 94638 2005 94698 3710
rect 94822 2549 94882 3710
rect 95006 2549 95066 3710
rect 94819 2548 94885 2549
rect 94819 2484 94820 2548
rect 94884 2484 94885 2548
rect 94819 2483 94885 2484
rect 95003 2548 95069 2549
rect 95003 2484 95004 2548
rect 95068 2484 95069 2548
rect 95003 2483 95069 2484
rect 94635 2004 94701 2005
rect 94144 1120 94464 2004
rect 94635 1940 94636 2004
rect 94700 1940 94701 2004
rect 94635 1939 94701 1940
rect 94144 1056 94152 1120
rect 94216 1056 94232 1120
rect 94296 1056 94312 1120
rect 94376 1056 94392 1120
rect 94456 1056 94464 1120
rect 93899 780 93965 781
rect 93899 716 93900 780
rect 93964 716 93965 780
rect 93899 715 93965 716
rect 93204 -390 93246 -154
rect 93482 -390 93524 -154
rect 93204 -1092 93524 -390
rect 94144 -814 94464 1056
rect 94144 -1050 94186 -814
rect 94422 -1050 94464 -814
rect 94144 -1092 94464 -1050
rect 94804 1664 95124 1880
rect 94804 1600 94812 1664
rect 94876 1600 94892 1664
rect 94956 1600 94972 1664
rect 95036 1600 95052 1664
rect 95116 1600 95124 1664
rect 94804 -154 95124 1600
rect 94804 -390 94846 -154
rect 95082 -390 95124 -154
rect 94804 -1092 95124 -390
rect 95744 1120 96064 2004
rect 95744 1056 95752 1120
rect 95816 1056 95832 1120
rect 95896 1056 95912 1120
rect 95976 1056 95992 1120
rect 96056 1056 96064 1120
rect 95744 -814 96064 1056
rect 95744 -1050 95786 -814
rect 96022 -1050 96064 -814
rect 95744 -1092 96064 -1050
rect 96404 1664 96724 2004
rect 96404 1600 96412 1664
rect 96476 1600 96492 1664
rect 96556 1600 96572 1664
rect 96636 1600 96652 1664
rect 96716 1600 96724 1664
rect 96404 -154 96724 1600
rect 96404 -390 96446 -154
rect 96682 -390 96724 -154
rect 96404 -1092 96724 -390
rect 97344 1120 97664 2004
rect 97344 1056 97352 1120
rect 97416 1056 97432 1120
rect 97496 1056 97512 1120
rect 97576 1056 97592 1120
rect 97656 1056 97664 1120
rect 97344 -814 97664 1056
rect 97344 -1050 97386 -814
rect 97622 -1050 97664 -814
rect 97344 -1092 97664 -1050
rect 98004 1664 98324 2004
rect 98004 1600 98012 1664
rect 98076 1600 98092 1664
rect 98156 1600 98172 1664
rect 98236 1600 98252 1664
rect 98316 1600 98324 1664
rect 98004 -154 98324 1600
rect 98004 -390 98046 -154
rect 98282 -390 98324 -154
rect 98004 -1092 98324 -390
rect 98944 1120 99264 2004
rect 98944 1056 98952 1120
rect 99016 1056 99032 1120
rect 99096 1056 99112 1120
rect 99176 1056 99192 1120
rect 99256 1056 99264 1120
rect 98944 -814 99264 1056
rect 98944 -1050 98986 -814
rect 99222 -1050 99264 -814
rect 98944 -1092 99264 -1050
rect 99604 1664 99924 2004
rect 99604 1600 99612 1664
rect 99676 1600 99692 1664
rect 99756 1600 99772 1664
rect 99836 1600 99852 1664
rect 99916 1600 99924 1664
rect 99604 -154 99924 1600
rect 99604 -390 99646 -154
rect 99882 -390 99924 -154
rect 99604 -1092 99924 -390
rect 100544 1120 100864 2004
rect 100544 1056 100552 1120
rect 100616 1056 100632 1120
rect 100696 1056 100712 1120
rect 100776 1056 100792 1120
rect 100856 1056 100864 1120
rect 100544 -814 100864 1056
rect 100544 -1050 100586 -814
rect 100822 -1050 100864 -814
rect 100544 -1092 100864 -1050
rect 101204 1664 101524 2004
rect 101204 1600 101212 1664
rect 101276 1600 101292 1664
rect 101356 1600 101372 1664
rect 101436 1600 101452 1664
rect 101516 1600 101524 1664
rect 101204 -154 101524 1600
rect 101204 -390 101246 -154
rect 101482 -390 101524 -154
rect 101204 -1092 101524 -390
rect 102144 1120 102464 2004
rect 102144 1056 102152 1120
rect 102216 1056 102232 1120
rect 102296 1056 102312 1120
rect 102376 1056 102392 1120
rect 102456 1056 102464 1120
rect 102144 -814 102464 1056
rect 102144 -1050 102186 -814
rect 102422 -1050 102464 -814
rect 102144 -1092 102464 -1050
rect 102804 1664 103124 2004
rect 102804 1600 102812 1664
rect 102876 1600 102892 1664
rect 102956 1600 102972 1664
rect 103036 1600 103052 1664
rect 103116 1600 103124 1664
rect 102804 -154 103124 1600
rect 102804 -390 102846 -154
rect 103082 -390 103124 -154
rect 102804 -1092 103124 -390
rect 103744 1120 104064 2004
rect 103744 1056 103752 1120
rect 103816 1056 103832 1120
rect 103896 1056 103912 1120
rect 103976 1056 103992 1120
rect 104056 1056 104064 1120
rect 103744 -814 104064 1056
rect 103744 -1050 103786 -814
rect 104022 -1050 104064 -814
rect 103744 -1092 104064 -1050
rect 104404 1664 104724 2004
rect 104404 1600 104412 1664
rect 104476 1600 104492 1664
rect 104556 1600 104572 1664
rect 104636 1600 104652 1664
rect 104716 1600 104724 1664
rect 104404 -154 104724 1600
rect 104404 -390 104446 -154
rect 104682 -390 104724 -154
rect 104404 -1092 104724 -390
rect 105344 1120 105664 2004
rect 105344 1056 105352 1120
rect 105416 1056 105432 1120
rect 105496 1056 105512 1120
rect 105576 1056 105592 1120
rect 105656 1056 105664 1120
rect 105344 -814 105664 1056
rect 105344 -1050 105386 -814
rect 105622 -1050 105664 -814
rect 105344 -1092 105664 -1050
rect 106004 1664 106324 2004
rect 106004 1600 106012 1664
rect 106076 1600 106092 1664
rect 106156 1600 106172 1664
rect 106236 1600 106252 1664
rect 106316 1600 106324 1664
rect 106004 -154 106324 1600
rect 106004 -390 106046 -154
rect 106282 -390 106324 -154
rect 106004 -1092 106324 -390
rect 106944 1120 107264 2004
rect 106944 1056 106952 1120
rect 107016 1056 107032 1120
rect 107096 1056 107112 1120
rect 107176 1056 107192 1120
rect 107256 1056 107264 1120
rect 106944 -814 107264 1056
rect 106944 -1050 106986 -814
rect 107222 -1050 107264 -814
rect 106944 -1092 107264 -1050
rect 107604 1664 107924 2004
rect 107604 1600 107612 1664
rect 107676 1600 107692 1664
rect 107756 1600 107772 1664
rect 107836 1600 107852 1664
rect 107916 1600 107924 1664
rect 107604 -154 107924 1600
rect 107604 -390 107646 -154
rect 107882 -390 107924 -154
rect 107604 -1092 107924 -390
rect 108544 1120 108864 2004
rect 108544 1056 108552 1120
rect 108616 1056 108632 1120
rect 108696 1056 108712 1120
rect 108776 1056 108792 1120
rect 108856 1056 108864 1120
rect 108544 -814 108864 1056
rect 110036 -154 110356 6630
rect 110036 -390 110078 -154
rect 110314 -390 110356 -154
rect 110036 -432 110356 -390
rect 110696 82206 111016 88398
rect 110696 81970 110738 82206
rect 110974 81970 111016 82206
rect 110696 6206 111016 81970
rect 110696 5970 110738 6206
rect 110974 5970 111016 6206
rect 108544 -1050 108586 -814
rect 108822 -1050 108864 -814
rect 108544 -1092 108864 -1050
rect 110696 -814 111016 5970
rect 110696 -1050 110738 -814
rect 110974 -1050 111016 -814
rect 110696 -1092 111016 -1050
<< via4 >>
rect -1034 88398 -798 88634
rect 2986 88398 3222 88634
rect -1034 81970 -798 82206
rect -1034 5970 -798 6206
rect -374 87738 -138 87974
rect -374 82630 -138 82866
rect 2986 81970 3222 82206
rect -374 6630 -138 6866
rect -374 -390 -138 -154
rect 2986 5970 3222 6206
rect -1034 -1050 -798 -814
rect 2986 -1050 3222 -814
rect 3646 87738 3882 87974
rect 3646 82630 3882 82866
rect 3646 6630 3882 6866
rect 3646 -390 3882 -154
rect 4586 88398 4822 88634
rect 4586 81970 4822 82206
rect 4586 5970 4822 6206
rect 4586 -1050 4822 -814
rect 5246 87738 5482 87974
rect 5246 82630 5482 82866
rect 5246 6630 5482 6866
rect 5246 -390 5482 -154
rect 6186 88398 6422 88634
rect 6186 81970 6422 82206
rect 6186 5970 6422 6206
rect 6186 -1050 6422 -814
rect 6846 87738 7082 87974
rect 6846 82630 7082 82866
rect 6846 6630 7082 6866
rect 6846 -390 7082 -154
rect 7786 88398 8022 88634
rect 7786 81970 8022 82206
rect 7786 5970 8022 6206
rect 7786 -1050 8022 -814
rect 8446 87738 8682 87974
rect 8446 82630 8682 82866
rect 8446 6630 8682 6866
rect 8446 -390 8682 -154
rect 9386 88398 9622 88634
rect 10046 87738 10282 87974
rect 10986 88398 11222 88634
rect 11646 87738 11882 87974
rect 9386 81970 9622 82206
rect 12586 88398 12822 88634
rect 13246 87738 13482 87974
rect 14186 88398 14422 88634
rect 14846 87738 15082 87974
rect 15786 88398 16022 88634
rect 16446 87738 16682 87974
rect 17386 88398 17622 88634
rect 18046 87738 18282 87974
rect 18986 88398 19222 88634
rect 19646 87738 19882 87974
rect 20586 88398 20822 88634
rect 21246 87738 21482 87974
rect 22186 88398 22422 88634
rect 22846 87738 23082 87974
rect 23786 88398 24022 88634
rect 24446 87738 24682 87974
rect 25386 88398 25622 88634
rect 26046 87738 26282 87974
rect 26986 88398 27222 88634
rect 27646 87738 27882 87974
rect 28586 88398 28822 88634
rect 29246 87738 29482 87974
rect 30186 88398 30422 88634
rect 30846 87738 31082 87974
rect 31786 88398 32022 88634
rect 32446 87738 32682 87974
rect 33386 88398 33622 88634
rect 34046 87738 34282 87974
rect 34986 88398 35222 88634
rect 35646 87738 35882 87974
rect 36586 88398 36822 88634
rect 37246 87738 37482 87974
rect 38186 88398 38422 88634
rect 38846 87738 39082 87974
rect 39786 88398 40022 88634
rect 40446 87738 40682 87974
rect 41386 88398 41622 88634
rect 42046 87738 42282 87974
rect 42986 88398 43222 88634
rect 43646 87738 43882 87974
rect 44586 88398 44822 88634
rect 45246 87738 45482 87974
rect 46186 88398 46422 88634
rect 46846 87738 47082 87974
rect 47786 88398 48022 88634
rect 48446 87738 48682 87974
rect 49386 88398 49622 88634
rect 50046 87738 50282 87974
rect 50986 88398 51222 88634
rect 51646 87738 51882 87974
rect 52586 88398 52822 88634
rect 53246 87738 53482 87974
rect 54186 88398 54422 88634
rect 54846 87738 55082 87974
rect 55786 88398 56022 88634
rect 56446 87738 56682 87974
rect 57386 88398 57622 88634
rect 58046 87738 58282 87974
rect 58986 88398 59222 88634
rect 59646 87738 59882 87974
rect 60586 88398 60822 88634
rect 61246 87738 61482 87974
rect 62186 88398 62422 88634
rect 62846 87738 63082 87974
rect 63786 88398 64022 88634
rect 64446 87738 64682 87974
rect 65386 88398 65622 88634
rect 66046 87738 66282 87974
rect 66986 88398 67222 88634
rect 67646 87738 67882 87974
rect 68586 88398 68822 88634
rect 69246 87738 69482 87974
rect 70186 88398 70422 88634
rect 70846 87738 71082 87974
rect 71786 88398 72022 88634
rect 72446 87738 72682 87974
rect 73386 88398 73622 88634
rect 74046 87738 74282 87974
rect 74986 88398 75222 88634
rect 75646 87738 75882 87974
rect 76586 88398 76822 88634
rect 77246 87738 77482 87974
rect 78186 88398 78422 88634
rect 78846 87738 79082 87974
rect 79786 88398 80022 88634
rect 80446 87738 80682 87974
rect 81386 88398 81622 88634
rect 82046 87738 82282 87974
rect 82986 88398 83222 88634
rect 83646 87738 83882 87974
rect 84586 88398 84822 88634
rect 85246 87738 85482 87974
rect 86186 88398 86422 88634
rect 86846 87738 87082 87974
rect 87786 88398 88022 88634
rect 88446 87738 88682 87974
rect 89386 88398 89622 88634
rect 90046 87738 90282 87974
rect 90986 88398 91222 88634
rect 91646 87738 91882 87974
rect 92586 88398 92822 88634
rect 93246 87738 93482 87974
rect 94186 88398 94422 88634
rect 94846 87738 95082 87974
rect 95786 88398 96022 88634
rect 96446 87738 96682 87974
rect 97386 88398 97622 88634
rect 98046 87738 98282 87974
rect 98986 88398 99222 88634
rect 99646 87738 99882 87974
rect 100586 88398 100822 88634
rect 101246 87738 101482 87974
rect 102186 88398 102422 88634
rect 102846 87738 103082 87974
rect 103786 88398 104022 88634
rect 104446 87738 104682 87974
rect 105386 88398 105622 88634
rect 106046 87738 106282 87974
rect 106986 88398 107222 88634
rect 107646 87738 107882 87974
rect 108586 88398 108822 88634
rect 110738 88398 110974 88634
rect 110078 87738 110314 87974
rect 110078 82630 110314 82866
rect 12328 81970 12564 82206
rect 107392 81970 107628 82206
rect 9386 5970 9622 6206
rect 9386 -1050 9622 -814
rect 13008 6630 13244 6866
rect 106712 6630 106948 6866
rect 110078 6630 110314 6866
rect 12328 5970 12564 6206
rect 107392 5970 107628 6206
rect 10046 -390 10282 -154
rect 10986 -1050 11222 -814
rect 11646 -390 11882 -154
rect 12586 -1050 12822 -814
rect 13246 -390 13482 -154
rect 14186 -1050 14422 -814
rect 14846 -390 15082 -154
rect 15786 -1050 16022 -814
rect 16446 -390 16682 -154
rect 17386 -1050 17622 -814
rect 18046 -390 18282 -154
rect 18986 -1050 19222 -814
rect 19646 -390 19882 -154
rect 20586 -1050 20822 -814
rect 21246 -390 21482 -154
rect 22186 -1050 22422 -814
rect 22846 -390 23082 -154
rect 23786 -1050 24022 -814
rect 24446 -390 24682 -154
rect 25386 -1050 25622 -814
rect 26046 -390 26282 -154
rect 26986 -1050 27222 -814
rect 27646 -390 27882 -154
rect 28586 -1050 28822 -814
rect 29246 -390 29482 -154
rect 30186 -1050 30422 -814
rect 30846 -390 31082 -154
rect 31786 -1050 32022 -814
rect 32446 -390 32682 -154
rect 33386 -1050 33622 -814
rect 34046 -390 34282 -154
rect 34986 -1050 35222 -814
rect 35646 -390 35882 -154
rect 36586 -1050 36822 -814
rect 37246 -390 37482 -154
rect 38186 -1050 38422 -814
rect 38846 -390 39082 -154
rect 39786 -1050 40022 -814
rect 40446 -390 40682 -154
rect 41386 -1050 41622 -814
rect 42046 -390 42282 -154
rect 42986 -1050 43222 -814
rect 43646 -390 43882 -154
rect 44586 -1050 44822 -814
rect 45246 -390 45482 -154
rect 46186 -1050 46422 -814
rect 46846 -390 47082 -154
rect 47786 -1050 48022 -814
rect 48446 -390 48682 -154
rect 49386 -1050 49622 -814
rect 50046 -390 50282 -154
rect 50986 -1050 51222 -814
rect 51646 -390 51882 -154
rect 52586 -1050 52822 -814
rect 53246 -390 53482 -154
rect 54186 -1050 54422 -814
rect 54846 -390 55082 -154
rect 55786 -1050 56022 -814
rect 56446 -390 56682 -154
rect 57386 -1050 57622 -814
rect 58046 -390 58282 -154
rect 58986 -1050 59222 -814
rect 59646 -390 59882 -154
rect 60586 -1050 60822 -814
rect 61246 -390 61482 -154
rect 62186 -1050 62422 -814
rect 62846 -390 63082 -154
rect 63786 -1050 64022 -814
rect 64446 -390 64682 -154
rect 65386 -1050 65622 -814
rect 66046 -390 66282 -154
rect 66986 -1050 67222 -814
rect 67646 -390 67882 -154
rect 68586 -1050 68822 -814
rect 69246 -390 69482 -154
rect 70186 -1050 70422 -814
rect 70846 -390 71082 -154
rect 71786 -1050 72022 -814
rect 72446 -390 72682 -154
rect 73386 -1050 73622 -814
rect 74046 -390 74282 -154
rect 74986 -1050 75222 -814
rect 75646 -390 75882 -154
rect 76586 -1050 76822 -814
rect 77246 -390 77482 -154
rect 78186 -1050 78422 -814
rect 78846 -390 79082 -154
rect 79786 -1050 80022 -814
rect 80446 -390 80682 -154
rect 81386 -1050 81622 -814
rect 82046 -390 82282 -154
rect 82986 -1050 83222 -814
rect 83646 -390 83882 -154
rect 84586 -1050 84822 -814
rect 85246 -390 85482 -154
rect 86186 -1050 86422 -814
rect 86846 -390 87082 -154
rect 87786 -1050 88022 -814
rect 88446 -390 88682 -154
rect 89386 -1050 89622 -814
rect 90046 -390 90282 -154
rect 90986 -1050 91222 -814
rect 91646 -390 91882 -154
rect 92586 -1050 92822 -814
rect 93246 -390 93482 -154
rect 94186 -1050 94422 -814
rect 94846 -390 95082 -154
rect 95786 -1050 96022 -814
rect 96446 -390 96682 -154
rect 97386 -1050 97622 -814
rect 98046 -390 98282 -154
rect 98986 -1050 99222 -814
rect 99646 -390 99882 -154
rect 100586 -1050 100822 -814
rect 101246 -390 101482 -154
rect 102186 -1050 102422 -814
rect 102846 -390 103082 -154
rect 103786 -1050 104022 -814
rect 104446 -390 104682 -154
rect 105386 -1050 105622 -814
rect 106046 -390 106282 -154
rect 106986 -1050 107222 -814
rect 107646 -390 107882 -154
rect 110078 -390 110314 -154
rect 110738 81970 110974 82206
rect 110738 5970 110974 6206
rect 108586 -1050 108822 -814
rect 110738 -1050 110974 -814
<< metal5 >>
rect -1076 88634 111016 88676
rect -1076 88398 -1034 88634
rect -798 88398 2986 88634
rect 3222 88398 4586 88634
rect 4822 88398 6186 88634
rect 6422 88398 7786 88634
rect 8022 88398 9386 88634
rect 9622 88398 10986 88634
rect 11222 88398 12586 88634
rect 12822 88398 14186 88634
rect 14422 88398 15786 88634
rect 16022 88398 17386 88634
rect 17622 88398 18986 88634
rect 19222 88398 20586 88634
rect 20822 88398 22186 88634
rect 22422 88398 23786 88634
rect 24022 88398 25386 88634
rect 25622 88398 26986 88634
rect 27222 88398 28586 88634
rect 28822 88398 30186 88634
rect 30422 88398 31786 88634
rect 32022 88398 33386 88634
rect 33622 88398 34986 88634
rect 35222 88398 36586 88634
rect 36822 88398 38186 88634
rect 38422 88398 39786 88634
rect 40022 88398 41386 88634
rect 41622 88398 42986 88634
rect 43222 88398 44586 88634
rect 44822 88398 46186 88634
rect 46422 88398 47786 88634
rect 48022 88398 49386 88634
rect 49622 88398 50986 88634
rect 51222 88398 52586 88634
rect 52822 88398 54186 88634
rect 54422 88398 55786 88634
rect 56022 88398 57386 88634
rect 57622 88398 58986 88634
rect 59222 88398 60586 88634
rect 60822 88398 62186 88634
rect 62422 88398 63786 88634
rect 64022 88398 65386 88634
rect 65622 88398 66986 88634
rect 67222 88398 68586 88634
rect 68822 88398 70186 88634
rect 70422 88398 71786 88634
rect 72022 88398 73386 88634
rect 73622 88398 74986 88634
rect 75222 88398 76586 88634
rect 76822 88398 78186 88634
rect 78422 88398 79786 88634
rect 80022 88398 81386 88634
rect 81622 88398 82986 88634
rect 83222 88398 84586 88634
rect 84822 88398 86186 88634
rect 86422 88398 87786 88634
rect 88022 88398 89386 88634
rect 89622 88398 90986 88634
rect 91222 88398 92586 88634
rect 92822 88398 94186 88634
rect 94422 88398 95786 88634
rect 96022 88398 97386 88634
rect 97622 88398 98986 88634
rect 99222 88398 100586 88634
rect 100822 88398 102186 88634
rect 102422 88398 103786 88634
rect 104022 88398 105386 88634
rect 105622 88398 106986 88634
rect 107222 88398 108586 88634
rect 108822 88398 110738 88634
rect 110974 88398 111016 88634
rect -1076 88356 111016 88398
rect -416 87974 110356 88016
rect -416 87738 -374 87974
rect -138 87738 3646 87974
rect 3882 87738 5246 87974
rect 5482 87738 6846 87974
rect 7082 87738 8446 87974
rect 8682 87738 10046 87974
rect 10282 87738 11646 87974
rect 11882 87738 13246 87974
rect 13482 87738 14846 87974
rect 15082 87738 16446 87974
rect 16682 87738 18046 87974
rect 18282 87738 19646 87974
rect 19882 87738 21246 87974
rect 21482 87738 22846 87974
rect 23082 87738 24446 87974
rect 24682 87738 26046 87974
rect 26282 87738 27646 87974
rect 27882 87738 29246 87974
rect 29482 87738 30846 87974
rect 31082 87738 32446 87974
rect 32682 87738 34046 87974
rect 34282 87738 35646 87974
rect 35882 87738 37246 87974
rect 37482 87738 38846 87974
rect 39082 87738 40446 87974
rect 40682 87738 42046 87974
rect 42282 87738 43646 87974
rect 43882 87738 45246 87974
rect 45482 87738 46846 87974
rect 47082 87738 48446 87974
rect 48682 87738 50046 87974
rect 50282 87738 51646 87974
rect 51882 87738 53246 87974
rect 53482 87738 54846 87974
rect 55082 87738 56446 87974
rect 56682 87738 58046 87974
rect 58282 87738 59646 87974
rect 59882 87738 61246 87974
rect 61482 87738 62846 87974
rect 63082 87738 64446 87974
rect 64682 87738 66046 87974
rect 66282 87738 67646 87974
rect 67882 87738 69246 87974
rect 69482 87738 70846 87974
rect 71082 87738 72446 87974
rect 72682 87738 74046 87974
rect 74282 87738 75646 87974
rect 75882 87738 77246 87974
rect 77482 87738 78846 87974
rect 79082 87738 80446 87974
rect 80682 87738 82046 87974
rect 82282 87738 83646 87974
rect 83882 87738 85246 87974
rect 85482 87738 86846 87974
rect 87082 87738 88446 87974
rect 88682 87738 90046 87974
rect 90282 87738 91646 87974
rect 91882 87738 93246 87974
rect 93482 87738 94846 87974
rect 95082 87738 96446 87974
rect 96682 87738 98046 87974
rect 98282 87738 99646 87974
rect 99882 87738 101246 87974
rect 101482 87738 102846 87974
rect 103082 87738 104446 87974
rect 104682 87738 106046 87974
rect 106282 87738 107646 87974
rect 107882 87738 110078 87974
rect 110314 87738 110356 87974
rect -416 87696 110356 87738
rect -1076 82866 111016 82908
rect -1076 82630 -374 82866
rect -138 82630 3646 82866
rect 3882 82630 5246 82866
rect 5482 82630 6846 82866
rect 7082 82630 8446 82866
rect 8682 82630 110078 82866
rect 110314 82630 111016 82866
rect -1076 82588 111016 82630
rect -1076 82206 111016 82248
rect -1076 81970 -1034 82206
rect -798 81970 2986 82206
rect 3222 81970 4586 82206
rect 4822 81970 6186 82206
rect 6422 81970 7786 82206
rect 8022 81970 9386 82206
rect 9622 81970 12328 82206
rect 12564 81970 107392 82206
rect 107628 81970 110738 82206
rect 110974 81970 111016 82206
rect -1076 81928 111016 81970
rect -1076 6866 111016 6908
rect -1076 6630 -374 6866
rect -138 6630 3646 6866
rect 3882 6630 5246 6866
rect 5482 6630 6846 6866
rect 7082 6630 8446 6866
rect 8682 6630 13008 6866
rect 13244 6630 106712 6866
rect 106948 6630 110078 6866
rect 110314 6630 111016 6866
rect -1076 6588 111016 6630
rect -1076 6206 111016 6248
rect -1076 5970 -1034 6206
rect -798 5970 2986 6206
rect 3222 5970 4586 6206
rect 4822 5970 6186 6206
rect 6422 5970 7786 6206
rect 8022 5970 9386 6206
rect 9622 5970 12328 6206
rect 12564 5970 107392 6206
rect 107628 5970 110738 6206
rect 110974 5970 111016 6206
rect -1076 5928 111016 5970
rect -416 -154 110356 -112
rect -416 -390 -374 -154
rect -138 -390 3646 -154
rect 3882 -390 5246 -154
rect 5482 -390 6846 -154
rect 7082 -390 8446 -154
rect 8682 -390 10046 -154
rect 10282 -390 11646 -154
rect 11882 -390 13246 -154
rect 13482 -390 14846 -154
rect 15082 -390 16446 -154
rect 16682 -390 18046 -154
rect 18282 -390 19646 -154
rect 19882 -390 21246 -154
rect 21482 -390 22846 -154
rect 23082 -390 24446 -154
rect 24682 -390 26046 -154
rect 26282 -390 27646 -154
rect 27882 -390 29246 -154
rect 29482 -390 30846 -154
rect 31082 -390 32446 -154
rect 32682 -390 34046 -154
rect 34282 -390 35646 -154
rect 35882 -390 37246 -154
rect 37482 -390 38846 -154
rect 39082 -390 40446 -154
rect 40682 -390 42046 -154
rect 42282 -390 43646 -154
rect 43882 -390 45246 -154
rect 45482 -390 46846 -154
rect 47082 -390 48446 -154
rect 48682 -390 50046 -154
rect 50282 -390 51646 -154
rect 51882 -390 53246 -154
rect 53482 -390 54846 -154
rect 55082 -390 56446 -154
rect 56682 -390 58046 -154
rect 58282 -390 59646 -154
rect 59882 -390 61246 -154
rect 61482 -390 62846 -154
rect 63082 -390 64446 -154
rect 64682 -390 66046 -154
rect 66282 -390 67646 -154
rect 67882 -390 69246 -154
rect 69482 -390 70846 -154
rect 71082 -390 72446 -154
rect 72682 -390 74046 -154
rect 74282 -390 75646 -154
rect 75882 -390 77246 -154
rect 77482 -390 78846 -154
rect 79082 -390 80446 -154
rect 80682 -390 82046 -154
rect 82282 -390 83646 -154
rect 83882 -390 85246 -154
rect 85482 -390 86846 -154
rect 87082 -390 88446 -154
rect 88682 -390 90046 -154
rect 90282 -390 91646 -154
rect 91882 -390 93246 -154
rect 93482 -390 94846 -154
rect 95082 -390 96446 -154
rect 96682 -390 98046 -154
rect 98282 -390 99646 -154
rect 99882 -390 101246 -154
rect 101482 -390 102846 -154
rect 103082 -390 104446 -154
rect 104682 -390 106046 -154
rect 106282 -390 107646 -154
rect 107882 -390 110078 -154
rect 110314 -390 110356 -154
rect -416 -432 110356 -390
rect -1076 -814 111016 -772
rect -1076 -1050 -1034 -814
rect -798 -1050 2986 -814
rect 3222 -1050 4586 -814
rect 4822 -1050 6186 -814
rect 6422 -1050 7786 -814
rect 8022 -1050 9386 -814
rect 9622 -1050 10986 -814
rect 11222 -1050 12586 -814
rect 12822 -1050 14186 -814
rect 14422 -1050 15786 -814
rect 16022 -1050 17386 -814
rect 17622 -1050 18986 -814
rect 19222 -1050 20586 -814
rect 20822 -1050 22186 -814
rect 22422 -1050 23786 -814
rect 24022 -1050 25386 -814
rect 25622 -1050 26986 -814
rect 27222 -1050 28586 -814
rect 28822 -1050 30186 -814
rect 30422 -1050 31786 -814
rect 32022 -1050 33386 -814
rect 33622 -1050 34986 -814
rect 35222 -1050 36586 -814
rect 36822 -1050 38186 -814
rect 38422 -1050 39786 -814
rect 40022 -1050 41386 -814
rect 41622 -1050 42986 -814
rect 43222 -1050 44586 -814
rect 44822 -1050 46186 -814
rect 46422 -1050 47786 -814
rect 48022 -1050 49386 -814
rect 49622 -1050 50986 -814
rect 51222 -1050 52586 -814
rect 52822 -1050 54186 -814
rect 54422 -1050 55786 -814
rect 56022 -1050 57386 -814
rect 57622 -1050 58986 -814
rect 59222 -1050 60586 -814
rect 60822 -1050 62186 -814
rect 62422 -1050 63786 -814
rect 64022 -1050 65386 -814
rect 65622 -1050 66986 -814
rect 67222 -1050 68586 -814
rect 68822 -1050 70186 -814
rect 70422 -1050 71786 -814
rect 72022 -1050 73386 -814
rect 73622 -1050 74986 -814
rect 75222 -1050 76586 -814
rect 76822 -1050 78186 -814
rect 78422 -1050 79786 -814
rect 80022 -1050 81386 -814
rect 81622 -1050 82986 -814
rect 83222 -1050 84586 -814
rect 84822 -1050 86186 -814
rect 86422 -1050 87786 -814
rect 88022 -1050 89386 -814
rect 89622 -1050 90986 -814
rect 91222 -1050 92586 -814
rect 92822 -1050 94186 -814
rect 94422 -1050 95786 -814
rect 96022 -1050 97386 -814
rect 97622 -1050 98986 -814
rect 99222 -1050 100586 -814
rect 100822 -1050 102186 -814
rect 102422 -1050 103786 -814
rect 104022 -1050 105386 -814
rect 105622 -1050 106986 -814
rect 107222 -1050 108586 -814
rect 108822 -1050 110738 -814
rect 110974 -1050 111016 -814
rect -1076 -1092 111016 -1050
use sky130_fd_sc_hd__or2_1  _173_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _174_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _175_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _176_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _177_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _178_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _179_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _180_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _181_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _182_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _183_
timestamp 1688980957
transform 1 0 6992 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1688980957
transform 1 0 8188 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _185_
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _186_
timestamp 1688980957
transform 1 0 4508 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _187_
timestamp 1688980957
transform 1 0 8004 0 1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1688980957
transform 1 0 7452 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _189_
timestamp 1688980957
transform 1 0 6624 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _190_
timestamp 1688980957
transform 1 0 7636 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _191_
timestamp 1688980957
transform 1 0 8832 0 -1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _192_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _193_
timestamp 1688980957
transform 1 0 6256 0 1 51136
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1688980957
transform 1 0 8096 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _195_
timestamp 1688980957
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _196_
timestamp 1688980957
transform 1 0 5152 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _197_
timestamp 1688980957
transform 1 0 8464 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 1688980957
transform 1 0 6992 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _199_
timestamp 1688980957
transform 1 0 6624 0 -1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _200_
timestamp 1688980957
transform 1 0 8924 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _201_
timestamp 1688980957
transform 1 0 7912 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _202_
timestamp 1688980957
transform 1 0 8004 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _203_
timestamp 1688980957
transform 1 0 4784 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform 1 0 4508 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _205_
timestamp 1688980957
transform 1 0 4232 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _206_
timestamp 1688980957
transform 1 0 4140 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1688980957
transform 1 0 8004 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _210_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1688980957
transform 1 0 7728 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _212_
timestamp 1688980957
transform 1 0 4140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1688980957
transform 1 0 8832 0 -1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _214_
timestamp 1688980957
transform 1 0 5980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1688980957
transform 1 0 6440 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _216_
timestamp 1688980957
transform 1 0 3956 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _217_
timestamp 1688980957
transform 1 0 8832 0 -1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _218_
timestamp 1688980957
transform 1 0 8280 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _219_
timestamp 1688980957
transform 1 0 6716 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _220_
timestamp 1688980957
transform 1 0 4140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1688980957
transform 1 0 8004 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _222_
timestamp 1688980957
transform 1 0 8924 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _223_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1688980957
transform 1 0 6992 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _225_
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _226_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _227_
timestamp 1688980957
transform 1 0 8832 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1688980957
transform 1 0 6900 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _229_
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1688980957
transform 1 0 8832 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _231_
timestamp 1688980957
transform 1 0 8556 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1688980957
transform 1 0 4324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1688980957
transform 1 0 8832 0 -1 71808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _235_
timestamp 1688980957
transform 1 0 8924 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1688980957
transform 1 0 6532 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _237_
timestamp 1688980957
transform 1 0 4048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1688980957
transform 1 0 8832 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _239_
timestamp 1688980957
transform 1 0 7728 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1688980957
transform 1 0 6624 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _241_
timestamp 1688980957
transform 1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _242_
timestamp 1688980957
transform 1 0 7360 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1688980957
transform 1 0 7728 0 -1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _244_
timestamp 1688980957
transform 1 0 4324 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1688980957
transform 1 0 6624 0 1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _246_
timestamp 1688980957
transform 1 0 4508 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _247_
timestamp 1688980957
transform 1 0 7176 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1688980957
transform 1 0 4232 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1688980957
transform 1 0 7452 0 1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1688980957
transform 1 0 4232 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1688980957
transform 1 0 6440 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _252_
timestamp 1688980957
transform 1 0 4232 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp 1688980957
transform 1 0 4784 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1688980957
transform 1 0 8004 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _255_
timestamp 1688980957
transform 1 0 4140 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _256_
timestamp 1688980957
transform 1 0 8004 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1688980957
transform 1 0 4508 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1688980957
transform 1 0 8096 0 -1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1688980957
transform 1 0 4508 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1688980957
transform 1 0 5428 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1688980957
transform 1 0 3772 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1688980957
transform 1 0 6348 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1688980957
transform 1 0 2116 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _264_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _265_
timestamp 1688980957
transform 1 0 24380 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _266_
timestamp 1688980957
transform 1 0 8924 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _267_
timestamp 1688980957
transform 1 0 33488 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _268_
timestamp 1688980957
transform 1 0 8556 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _269_
timestamp 1688980957
transform 1 0 37260 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _270_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 73984
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _271_
timestamp 1688980957
transform 1 0 26956 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _272_
timestamp 1688980957
transform 1 0 9200 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _273_
timestamp 1688980957
transform 1 0 29808 0 1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 1688980957
transform 1 0 8096 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1688980957
transform 1 0 7636 0 1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1688980957
transform 1 0 4140 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _277_
timestamp 1688980957
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1688980957
transform 1 0 7268 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _279_
timestamp 1688980957
transform 1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _280_
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1688980957
transform 1 0 8004 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _282_
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _283_
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _285_
timestamp 1688980957
transform 1 0 7268 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _286_
timestamp 1688980957
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _288_
timestamp 1688980957
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _290_
timestamp 1688980957
transform 1 0 9108 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _291_
timestamp 1688980957
transform 1 0 6992 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _292_
timestamp 1688980957
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1688980957
transform 1 0 6808 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _294_
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _295_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _297_
timestamp 1688980957
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _298_
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _299_
timestamp 1688980957
transform 1 0 28428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _300_
timestamp 1688980957
transform 1 0 4416 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _301_
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _302_
timestamp 1688980957
transform 1 0 26128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp 1688980957
transform 1 0 7360 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _304_
timestamp 1688980957
transform 1 0 7268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp 1688980957
transform 1 0 7176 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _306_
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _307_
timestamp 1688980957
transform 1 0 6992 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _308_
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _309_
timestamp 1688980957
transform 1 0 7912 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _310_
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _313_
timestamp 1688980957
transform 1 0 7452 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1688980957
transform 1 0 22724 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _315_
timestamp 1688980957
transform 1 0 7176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _316_
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _317_
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _318_
timestamp 1688980957
transform 1 0 8188 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _319_
timestamp 1688980957
transform 1 0 27508 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _320_
timestamp 1688980957
transform 1 0 8004 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _321_
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _322_
timestamp 1688980957
transform 1 0 7912 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _323_
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _324_
timestamp 1688980957
transform 1 0 8004 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _325_
timestamp 1688980957
transform 1 0 30452 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _326_
timestamp 1688980957
transform 1 0 8004 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _327_
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _328_
timestamp 1688980957
transform 1 0 8004 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _329_
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_2  _330_
timestamp 1688980957
transform 1 0 8004 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _331_
timestamp 1688980957
transform 1 0 33580 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_4  _332_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _333_
timestamp 1688980957
transform 1 0 37444 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__o21bai_1  _334_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _335_
timestamp 1688980957
transform 1 0 4324 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _336_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _337_
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _338_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _339_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _340_
timestamp 1688980957
transform 1 0 7820 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _341_
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _342_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1688980957
transform 1 0 7176 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _344_
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _345_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _346_
timestamp 1688980957
transform 1 0 6900 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _347_
timestamp 1688980957
transform 1 0 5336 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _348_
timestamp 1688980957
transform 1 0 6532 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1688980957
transform 1 0 8096 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _350_
timestamp 1688980957
transform 1 0 7176 0 1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _351_
timestamp 1688980957
transform 1 0 4784 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _352_
timestamp 1688980957
transform 1 0 4968 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _353_
timestamp 1688980957
transform 1 0 4692 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _354_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 60928
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _355_
timestamp 1688980957
transform 1 0 5152 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _356_
timestamp 1688980957
transform 1 0 6072 0 1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _357_
timestamp 1688980957
transform 1 0 4232 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _358_
timestamp 1688980957
transform 1 0 7268 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _359_
timestamp 1688980957
transform 1 0 4508 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _360_
timestamp 1688980957
transform 1 0 6532 0 1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  _361_
timestamp 1688980957
transform 1 0 4048 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _362_
timestamp 1688980957
transform 1 0 5336 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _363_
timestamp 1688980957
transform 1 0 4140 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _364_
timestamp 1688980957
transform 1 0 6348 0 1 71808
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _365_
timestamp 1688980957
transform 1 0 6808 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_2  _366_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _367_
timestamp 1688980957
transform 1 0 5244 0 -1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_2  _368_
timestamp 1688980957
transform 1 0 7176 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _369_
timestamp 1688980957
transform 1 0 6992 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1688980957
transform 1 0 7728 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _371_
timestamp 1688980957
transform 1 0 6624 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _372_
timestamp 1688980957
transform 1 0 4140 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _373_
timestamp 1688980957
transform 1 0 8464 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _374_
timestamp 1688980957
transform 1 0 5336 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _375_
timestamp 1688980957
transform 1 0 5704 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _376_
timestamp 1688980957
transform 1 0 5060 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1688980957
transform 1 0 8004 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _378_
timestamp 1688980957
transform 1 0 4876 0 -1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _379_
timestamp 1688980957
transform 1 0 4784 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _380_
timestamp 1688980957
transform 1 0 7268 0 1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _381_
timestamp 1688980957
transform 1 0 7084 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _382_
timestamp 1688980957
transform 1 0 5520 0 1 72896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _383_
timestamp 1688980957
transform 1 0 5336 0 1 71808
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _384_
timestamp 1688980957
transform 1 0 3956 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _385_
timestamp 1688980957
transform 1 0 7636 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _386_
timestamp 1688980957
transform 1 0 7544 0 1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1688980957
transform 1 0 7636 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _388_
timestamp 1688980957
transform 1 0 7452 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _389_
timestamp 1688980957
transform 1 0 6900 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _390_
timestamp 1688980957
transform 1 0 4416 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1688980957
transform 1 0 8004 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _392_
timestamp 1688980957
transform 1 0 6992 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _393_
timestamp 1688980957
transform 1 0 6440 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _394_
timestamp 1688980957
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _395_
timestamp 1688980957
transform 1 0 7912 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _396_
timestamp 1688980957
transform 1 0 7728 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _397_
timestamp 1688980957
transform 1 0 7176 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1688980957
transform 1 0 8004 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _399_
timestamp 1688980957
transform 1 0 8464 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _400_
timestamp 1688980957
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _401_
timestamp 1688980957
transform 1 0 4416 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1688980957
transform 1 0 7176 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _403_
timestamp 1688980957
transform 1 0 4968 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _404_
timestamp 1688980957
transform 1 0 6992 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _405_
timestamp 1688980957
transform 1 0 8096 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _406_
timestamp 1688980957
transform 1 0 8924 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _407_
timestamp 1688980957
transform 1 0 6348 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _408_
timestamp 1688980957
transform 1 0 4324 0 -1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1688980957
transform 1 0 6348 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _410_
timestamp 1688980957
transform 1 0 7176 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _411_
timestamp 1688980957
transform 1 0 4784 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1688980957
transform 1 0 8648 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _413_
timestamp 1688980957
transform 1 0 6532 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _414_
timestamp 1688980957
transform 1 0 6624 0 -1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _415_
timestamp 1688980957
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _416_
timestamp 1688980957
transform 1 0 7912 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _417_
timestamp 1688980957
transform 1 0 6624 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__dlxtn_1  _418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _419_
timestamp 1688980957
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _420_
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _421_
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _422_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp 1688980957
transform 1 0 6624 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp 1688980957
transform 1 0 6716 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _425_
timestamp 1688980957
transform 1 0 6624 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp 1688980957
transform 1 0 6716 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _427_
timestamp 1688980957
transform 1 0 6624 0 -1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp 1688980957
transform 1 0 6624 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp 1688980957
transform 1 0 3772 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp 1688980957
transform 1 0 6716 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp 1688980957
transform 1 0 6624 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _432_
timestamp 1688980957
transform 1 0 6716 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1688980957
transform 1 0 6716 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1688980957
transform 1 0 6348 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _435_
timestamp 1688980957
transform 1 0 6716 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1688980957
transform 1 0 6716 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1688980957
transform 1 0 6716 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _438_
timestamp 1688980957
transform 1 0 7268 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _439_
timestamp 1688980957
transform 1 0 5888 0 1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _440_
timestamp 1688980957
transform 1 0 6532 0 -1 63104
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _441_
timestamp 1688980957
transform 1 0 5704 0 1 64192
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1688980957
transform 1 0 4784 0 -1 67456
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1688980957
transform 1 0 6440 0 -1 64192
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1688980957
transform 1 0 6624 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _445_
timestamp 1688980957
transform 1 0 6716 0 -1 60928
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1688980957
transform 1 0 4324 0 1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1688980957
transform 1 0 6348 0 -1 71808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1688980957
transform 1 0 35052 0 1 85952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1688980957
transform -1 0 49312 0 1 85952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1688980957
transform 1 0 55292 0 1 85952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1688980957
transform 1 0 40572 0 1 85952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1688980957
transform 1 0 43424 0 1 85952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1688980957
transform 1 0 7084 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1688980957
transform 1 0 6348 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1688980957
transform 1 0 5428 0 1 58752
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35788 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 38548 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 52992 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 7544 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 8464 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 61180 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 7452 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 50324 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 7452 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 6900 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 49864 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 7636 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 9108 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 52440 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 6808 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 6624 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 6900 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1688980957
transform 1 0 50692 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1688980957
transform 1 0 8188 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1688980957
transform 1 0 5980 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1688980957
transform 1 0 38824 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1688980957
transform 1 0 8096 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1688980957
transform 1 0 7636 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1688980957
transform 1 0 51152 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1688980957
transform 1 0 51520 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1688980957
transform 1 0 6808 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1688980957
transform 1 0 51888 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1688980957
transform 1 0 39192 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1688980957
transform 1 0 39560 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1688980957
transform 1 0 40020 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1688980957
transform 1 0 40388 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1688980957
transform 1 0 42872 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1688980957
transform 1 0 43240 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1688980957
transform 1 0 47288 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1688980957
transform -1 0 49680 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 53360 0 1 85952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 44988 0 1 85952
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_233 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_243
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_257
timestamp 1688980957
transform 1 0 24748 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_275 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26404 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_285
timestamp 1688980957
transform 1 0 27324 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_313
timestamp 1688980957
transform 1 0 29900 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_317
timestamp 1688980957
transform 1 0 30268 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_323
timestamp 1688980957
transform 1 0 30820 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_347 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33028 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_375
timestamp 1688980957
transform 1 0 35604 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_379
timestamp 1688980957
transform 1 0 35972 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_409
timestamp 1688980957
transform 1 0 38732 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1688980957
transform 1 0 46092 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 1688980957
transform 1 0 47196 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 1688980957
transform 1 0 47564 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 1688980957
transform 1 0 48668 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1688980957
transform 1 0 49772 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 1688980957
transform 1 0 50140 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1688980957
transform 1 0 51244 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1688980957
transform 1 0 52348 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 1688980957
transform 1 0 52716 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 1688980957
transform 1 0 53820 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1688980957
transform 1 0 54924 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 1688980957
transform 1 0 56396 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 1688980957
transform 1 0 57500 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_617
timestamp 1688980957
transform 1 0 57868 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_629
timestamp 1688980957
transform 1 0 58972 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_641
timestamp 1688980957
transform 1 0 60076 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_645
timestamp 1688980957
transform 1 0 60444 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_657
timestamp 1688980957
transform 1 0 61548 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_669
timestamp 1688980957
transform 1 0 62652 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_673
timestamp 1688980957
transform 1 0 63020 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_685
timestamp 1688980957
transform 1 0 64124 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_697
timestamp 1688980957
transform 1 0 65228 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_701
timestamp 1688980957
transform 1 0 65596 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_713
timestamp 1688980957
transform 1 0 66700 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_725
timestamp 1688980957
transform 1 0 67804 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_729
timestamp 1688980957
transform 1 0 68172 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_741
timestamp 1688980957
transform 1 0 69276 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_753
timestamp 1688980957
transform 1 0 70380 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_757
timestamp 1688980957
transform 1 0 70748 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_769
timestamp 1688980957
transform 1 0 71852 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_781
timestamp 1688980957
transform 1 0 72956 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_785
timestamp 1688980957
transform 1 0 73324 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_797
timestamp 1688980957
transform 1 0 74428 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_809
timestamp 1688980957
transform 1 0 75532 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_813
timestamp 1688980957
transform 1 0 75900 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_825
timestamp 1688980957
transform 1 0 77004 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_837
timestamp 1688980957
transform 1 0 78108 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_841
timestamp 1688980957
transform 1 0 78476 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_853
timestamp 1688980957
transform 1 0 79580 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_865
timestamp 1688980957
transform 1 0 80684 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_869
timestamp 1688980957
transform 1 0 81052 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_881
timestamp 1688980957
transform 1 0 82156 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_893
timestamp 1688980957
transform 1 0 83260 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_897
timestamp 1688980957
transform 1 0 83628 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_909
timestamp 1688980957
transform 1 0 84732 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_921
timestamp 1688980957
transform 1 0 85836 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_925
timestamp 1688980957
transform 1 0 86204 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_937
timestamp 1688980957
transform 1 0 87308 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_949
timestamp 1688980957
transform 1 0 88412 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_953
timestamp 1688980957
transform 1 0 88780 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_965
timestamp 1688980957
transform 1 0 89884 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_977
timestamp 1688980957
transform 1 0 90988 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_981
timestamp 1688980957
transform 1 0 91356 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_993
timestamp 1688980957
transform 1 0 92460 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1005
timestamp 1688980957
transform 1 0 93564 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1009
timestamp 1688980957
transform 1 0 93932 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1021
timestamp 1688980957
transform 1 0 95036 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1033
timestamp 1688980957
transform 1 0 96140 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1037
timestamp 1688980957
transform 1 0 96508 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1049
timestamp 1688980957
transform 1 0 97612 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1061
timestamp 1688980957
transform 1 0 98716 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1065
timestamp 1688980957
transform 1 0 99084 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1077
timestamp 1688980957
transform 1 0 100188 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1089
timestamp 1688980957
transform 1 0 101292 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1093
timestamp 1688980957
transform 1 0 101660 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1105
timestamp 1688980957
transform 1 0 102764 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1117
timestamp 1688980957
transform 1 0 103868 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1121
timestamp 1688980957
transform 1 0 104236 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1133
timestamp 1688980957
transform 1 0 105340 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1145
timestamp 1688980957
transform 1 0 106444 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1149
timestamp 1688980957
transform 1 0 106812 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1161
timestamp 1688980957
transform 1 0 107916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1167
timestamp 1688980957
transform 1 0 108468 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_21
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1688980957
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_33
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_21
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_71
timestamp 1688980957
transform 1 0 7636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_21
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_71
timestamp 1688980957
transform 1 0 7636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_73
timestamp 1688980957
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_21
timestamp 1688980957
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_45
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_21
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_45
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_21
timestamp 1688980957
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_33
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_45
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_72
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_84
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_92
timestamp 1688980957
transform 1 0 9568 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_74
timestamp 1688980957
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_82
timestamp 1688980957
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_21
timestamp 1688980957
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_14
timestamp 1688980957
transform 1 0 2392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_73
timestamp 1688980957
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_21
timestamp 1688980957
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_65
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_71
timestamp 1688980957
transform 1 0 7636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_83
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_91
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_21
timestamp 1688980957
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_35
timestamp 1688980957
transform 1 0 4324 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_47
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_59
timestamp 1688980957
transform 1 0 6532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_71
timestamp 1688980957
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_7
timestamp 1688980957
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_19
timestamp 1688980957
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_31
timestamp 1688980957
transform 1 0 3956 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_38
timestamp 1688980957
transform 1 0 4600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_50
timestamp 1688980957
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_75
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_87
timestamp 1688980957
transform 1 0 9108 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_36
timestamp 1688980957
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_48
timestamp 1688980957
transform 1 0 5520 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_60
timestamp 1688980957
transform 1 0 6624 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_72
timestamp 1688980957
transform 1 0 7728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_6
timestamp 1688980957
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_18
timestamp 1688980957
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_30
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_34
timestamp 1688980957
transform 1 0 4232 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_38
timestamp 1688980957
transform 1 0 4600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_50
timestamp 1688980957
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_36
timestamp 1688980957
transform 1 0 4416 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_48
timestamp 1688980957
transform 1 0 5520 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_60
timestamp 1688980957
transform 1 0 6624 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_66
timestamp 1688980957
transform 1 0 7176 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_72
timestamp 1688980957
transform 1 0 7728 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_7
timestamp 1688980957
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_19
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_31
timestamp 1688980957
transform 1 0 3956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_36
timestamp 1688980957
transform 1 0 4416 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_48
timestamp 1688980957
transform 1 0 5520 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_61
timestamp 1688980957
transform 1 0 6716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_64
timestamp 1688980957
transform 1 0 6992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_84
timestamp 1688980957
transform 1 0 8832 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_91
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_21
timestamp 1688980957
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_34
timestamp 1688980957
transform 1 0 4232 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_46
timestamp 1688980957
transform 1 0 5336 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_58
timestamp 1688980957
transform 1 0 6440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_65
timestamp 1688980957
transform 1 0 7084 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_76
timestamp 1688980957
transform 1 0 8096 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_88
timestamp 1688980957
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_92
timestamp 1688980957
transform 1 0 9568 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_9
timestamp 1688980957
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_21
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_70
timestamp 1688980957
transform 1 0 7544 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_82
timestamp 1688980957
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_6
timestamp 1688980957
transform 1 0 1656 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_18
timestamp 1688980957
transform 1 0 2760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_74
timestamp 1688980957
transform 1 0 7912 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_70
timestamp 1688980957
transform 1 0 7544 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_76
timestamp 1688980957
transform 1 0 8096 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_86
timestamp 1688980957
transform 1 0 9016 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_92
timestamp 1688980957
transform 1 0 9568 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_6
timestamp 1688980957
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_18
timestamp 1688980957
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_6
timestamp 1688980957
transform 1 0 1656 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_18
timestamp 1688980957
transform 1 0 2760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_30
timestamp 1688980957
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_42
timestamp 1688980957
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_54
timestamp 1688980957
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_72
timestamp 1688980957
transform 1 0 7728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_84
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_92
timestamp 1688980957
transform 1 0 9568 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_6
timestamp 1688980957
transform 1 0 1656 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_18
timestamp 1688980957
transform 1 0 2760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_30
timestamp 1688980957
transform 1 0 3864 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_42
timestamp 1688980957
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_54
timestamp 1688980957
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_61
timestamp 1688980957
transform 1 0 6716 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_73
timestamp 1688980957
transform 1 0 7820 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_9
timestamp 1688980957
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_21
timestamp 1688980957
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_33
timestamp 1688980957
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_45
timestamp 1688980957
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_53
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_61
timestamp 1688980957
transform 1 0 6716 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_71
timestamp 1688980957
transform 1 0 7636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_83
timestamp 1688980957
transform 1 0 8740 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_91
timestamp 1688980957
transform 1 0 9476 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_73
timestamp 1688980957
transform 1 0 7820 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_9
timestamp 1688980957
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_21
timestamp 1688980957
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_33
timestamp 1688980957
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_45
timestamp 1688980957
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_53
timestamp 1688980957
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_84
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_92
timestamp 1688980957
transform 1 0 9568 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_73
timestamp 1688980957
transform 1 0 7820 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_84
timestamp 1688980957
transform 1 0 8832 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_92
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_21
timestamp 1688980957
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_71
timestamp 1688980957
transform 1 0 7636 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_92
timestamp 1688980957
transform 1 0 9568 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_9
timestamp 1688980957
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_21
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_61
timestamp 1688980957
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_64
timestamp 1688980957
transform 1 0 6992 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_75
timestamp 1688980957
transform 1 0 8004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_9
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_21
timestamp 1688980957
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_33
timestamp 1688980957
transform 1 0 4140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_45
timestamp 1688980957
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_53
timestamp 1688980957
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_78
timestamp 1688980957
transform 1 0 8280 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_90
timestamp 1688980957
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_78
timestamp 1688980957
transform 1 0 8280 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_9
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_21
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_33
timestamp 1688980957
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_45
timestamp 1688980957
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_53
timestamp 1688980957
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_62
timestamp 1688980957
transform 1 0 6808 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_9
timestamp 1688980957
transform 1 0 1932 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_21
timestamp 1688980957
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_33
timestamp 1688980957
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_45
timestamp 1688980957
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_53
timestamp 1688980957
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_90
timestamp 1688980957
transform 1 0 9384 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_35
timestamp 1688980957
transform 1 0 4324 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_40
timestamp 1688980957
transform 1 0 4784 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_52
timestamp 1688980957
transform 1 0 5888 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_73
timestamp 1688980957
transform 1 0 7820 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_81
timestamp 1688980957
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_9
timestamp 1688980957
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_21
timestamp 1688980957
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_33
timestamp 1688980957
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_45
timestamp 1688980957
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_53
timestamp 1688980957
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_9
timestamp 1688980957
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_21
timestamp 1688980957
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_40
timestamp 1688980957
transform 1 0 4784 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_52
timestamp 1688980957
transform 1 0 5888 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_64
timestamp 1688980957
transform 1 0 6992 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_76
timestamp 1688980957
transform 1 0 8096 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_77
timestamp 1688980957
transform 1 0 8188 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_89
timestamp 1688980957
transform 1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_9
timestamp 1688980957
transform 1 0 1932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_21
timestamp 1688980957
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_51
timestamp 1688980957
transform 1 0 5796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_57
timestamp 1688980957
transform 1 0 6348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_67
timestamp 1688980957
transform 1 0 7268 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_79
timestamp 1688980957
transform 1 0 8372 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_77
timestamp 1688980957
transform 1 0 8188 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_89
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_6
timestamp 1688980957
transform 1 0 1656 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_18
timestamp 1688980957
transform 1 0 2760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78_26
timestamp 1688980957
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_33
timestamp 1688980957
transform 1 0 4140 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_40
timestamp 1688980957
transform 1 0 4784 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_52
timestamp 1688980957
transform 1 0 5888 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_60
timestamp 1688980957
transform 1 0 6624 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_47
timestamp 1688980957
transform 1 0 5428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_77
timestamp 1688980957
transform 1 0 8188 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_89
timestamp 1688980957
transform 1 0 9292 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_6
timestamp 1688980957
transform 1 0 1656 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_18
timestamp 1688980957
transform 1 0 2760 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_26
timestamp 1688980957
transform 1 0 3496 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_50
timestamp 1688980957
transform 1 0 5704 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80_58
timestamp 1688980957
transform 1 0 6440 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_70
timestamp 1688980957
transform 1 0 7544 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80_82
timestamp 1688980957
transform 1 0 8648 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_9
timestamp 1688980957
transform 1 0 1932 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_21
timestamp 1688980957
transform 1 0 3036 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81_33
timestamp 1688980957
transform 1 0 4140 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_43
timestamp 1688980957
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_65
timestamp 1688980957
transform 1 0 7084 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_72
timestamp 1688980957
transform 1 0 7728 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_80
timestamp 1688980957
transform 1 0 8464 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_92
timestamp 1688980957
transform 1 0 9568 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1688980957
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1688980957
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1688980957
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_59
timestamp 1688980957
transform 1 0 6532 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_76
timestamp 1688980957
transform 1 0 8096 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82_91
timestamp 1688980957
transform 1 0 9476 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_9
timestamp 1688980957
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_21
timestamp 1688980957
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_33
timestamp 1688980957
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_45
timestamp 1688980957
transform 1 0 5244 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_49
timestamp 1688980957
transform 1 0 5612 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1688980957
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1688980957
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1688980957
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_45
timestamp 1688980957
transform 1 0 5244 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_84_57
timestamp 1688980957
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1688980957
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1688980957
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_85
timestamp 1688980957
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_9
timestamp 1688980957
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_21
timestamp 1688980957
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_33
timestamp 1688980957
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_45
timestamp 1688980957
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85_53
timestamp 1688980957
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_57
timestamp 1688980957
transform 1 0 6348 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1688980957
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1688980957
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 1688980957
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 1688980957
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1688980957
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1688980957
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1688980957
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_53
timestamp 1688980957
transform 1 0 5980 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_59
timestamp 1688980957
transform 1 0 6532 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_76
timestamp 1688980957
transform 1 0 8096 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_85
timestamp 1688980957
transform 1 0 8924 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_9
timestamp 1688980957
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_21
timestamp 1688980957
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_33
timestamp 1688980957
transform 1 0 4140 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_40
timestamp 1688980957
transform 1 0 4784 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_87_57
timestamp 1688980957
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_76
timestamp 1688980957
transform 1 0 8096 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_88
timestamp 1688980957
transform 1 0 9200 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_92
timestamp 1688980957
transform 1 0 9568 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_9
timestamp 1688980957
transform 1 0 1932 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_21
timestamp 1688980957
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1688980957
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1688980957
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1688980957
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88_53
timestamp 1688980957
transform 1 0 5980 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1688980957
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_85
timestamp 1688980957
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 1688980957
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 1688980957
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_27
timestamp 1688980957
transform 1 0 3588 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_33
timestamp 1688980957
transform 1 0 4140 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_45
timestamp 1688980957
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_89_53
timestamp 1688980957
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_89_57
timestamp 1688980957
transform 1 0 6348 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_79
timestamp 1688980957
transform 1 0 8372 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89_91
timestamp 1688980957
transform 1 0 9476 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_9
timestamp 1688980957
transform 1 0 1932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_21
timestamp 1688980957
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1688980957
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1688980957
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1688980957
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1688980957
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1688980957
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1688980957
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1688980957
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90_85
timestamp 1688980957
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1688980957
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1688980957
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 1688980957
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 1688980957
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 1688980957
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 1688980957
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_76
timestamp 1688980957
transform 1 0 8096 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_88
timestamp 1688980957
transform 1 0 9200 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_92
timestamp 1688980957
transform 1 0 9568 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_9
timestamp 1688980957
transform 1 0 1932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_21
timestamp 1688980957
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1688980957
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1688980957
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 1688980957
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_92_53
timestamp 1688980957
transform 1 0 5980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 1688980957
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_85
timestamp 1688980957
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1688980957
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1688980957
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_27
timestamp 1688980957
transform 1 0 3588 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_38
timestamp 1688980957
transform 1 0 4600 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_50
timestamp 1688980957
transform 1 0 5704 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_57
timestamp 1688980957
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_77
timestamp 1688980957
transform 1 0 8188 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_89
timestamp 1688980957
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_9
timestamp 1688980957
transform 1 0 1932 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_21
timestamp 1688980957
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1688980957
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1688980957
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1688980957
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_56
timestamp 1688980957
transform 1 0 6256 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_60
timestamp 1688980957
transform 1 0 6624 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 1688980957
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 1688980957
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_85
timestamp 1688980957
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_9
timestamp 1688980957
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_21
timestamp 1688980957
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_33
timestamp 1688980957
transform 1 0 4140 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_45
timestamp 1688980957
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_95_53
timestamp 1688980957
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_57
timestamp 1688980957
transform 1 0 6348 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_63
timestamp 1688980957
transform 1 0 6900 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_78
timestamp 1688980957
transform 1 0 8280 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_95_90
timestamp 1688980957
transform 1 0 9384 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1688980957
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1688980957
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1688980957
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_29
timestamp 1688980957
transform 1 0 3772 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_37
timestamp 1688980957
transform 1 0 4508 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_44
timestamp 1688980957
transform 1 0 5152 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_56
timestamp 1688980957
transform 1 0 6256 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_69
timestamp 1688980957
transform 1 0 7452 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_75
timestamp 1688980957
transform 1 0 8004 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1688980957
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_85
timestamp 1688980957
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_9
timestamp 1688980957
transform 1 0 1932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_21
timestamp 1688980957
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_33
timestamp 1688980957
transform 1 0 4140 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_40
timestamp 1688980957
transform 1 0 4784 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_52
timestamp 1688980957
transform 1 0 5888 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_57
timestamp 1688980957
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_65
timestamp 1688980957
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_76
timestamp 1688980957
transform 1 0 8096 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_88
timestamp 1688980957
transform 1 0 9200 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_92
timestamp 1688980957
transform 1 0 9568 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 1688980957
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 1688980957
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1688980957
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_29
timestamp 1688980957
transform 1 0 3772 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_33
timestamp 1688980957
transform 1 0 4140 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_37
timestamp 1688980957
transform 1 0 4508 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_49
timestamp 1688980957
transform 1 0 5612 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98_57
timestamp 1688980957
transform 1 0 6348 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_64
timestamp 1688980957
transform 1 0 6992 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_76
timestamp 1688980957
transform 1 0 8096 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_85
timestamp 1688980957
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_9
timestamp 1688980957
transform 1 0 1932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_21
timestamp 1688980957
transform 1 0 3036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_33
timestamp 1688980957
transform 1 0 4140 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_45
timestamp 1688980957
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_53
timestamp 1688980957
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1688980957
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1688980957
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1688980957
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1688980957
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1688980957
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1688980957
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_29
timestamp 1688980957
transform 1 0 3772 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_35
timestamp 1688980957
transform 1 0 4324 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_47
timestamp 1688980957
transform 1 0 5428 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_59
timestamp 1688980957
transform 1 0 6532 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_63
timestamp 1688980957
transform 1 0 6900 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_74
timestamp 1688980957
transform 1 0 7912 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_82
timestamp 1688980957
transform 1 0 8648 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_85
timestamp 1688980957
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_9
timestamp 1688980957
transform 1 0 1932 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_21
timestamp 1688980957
transform 1 0 3036 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_33
timestamp 1688980957
transform 1 0 4140 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_40
timestamp 1688980957
transform 1 0 4784 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_52
timestamp 1688980957
transform 1 0 5888 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_57
timestamp 1688980957
transform 1 0 6348 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_65
timestamp 1688980957
transform 1 0 7084 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_72
timestamp 1688980957
transform 1 0 7728 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_84
timestamp 1688980957
transform 1 0 8832 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_92
timestamp 1688980957
transform 1 0 9568 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_9
timestamp 1688980957
transform 1 0 1932 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_102_21
timestamp 1688980957
transform 1 0 3036 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102_27
timestamp 1688980957
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102_29
timestamp 1688980957
transform 1 0 3772 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_36
timestamp 1688980957
transform 1 0 4416 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_102_48
timestamp 1688980957
transform 1 0 5520 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_60
timestamp 1688980957
transform 1 0 6624 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102_68
timestamp 1688980957
transform 1 0 7360 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_73
timestamp 1688980957
transform 1 0 7820 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_102_81
timestamp 1688980957
transform 1 0 8556 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102_85
timestamp 1688980957
transform 1 0 8924 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_3
timestamp 1688980957
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_15
timestamp 1688980957
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103_27
timestamp 1688980957
transform 1 0 3588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_40
timestamp 1688980957
transform 1 0 4784 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103_52
timestamp 1688980957
transform 1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_103_78
timestamp 1688980957
transform 1 0 8280 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103_90
timestamp 1688980957
transform 1 0 9384 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_9
timestamp 1688980957
transform 1 0 1932 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104_21
timestamp 1688980957
transform 1 0 3036 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_27
timestamp 1688980957
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_29
timestamp 1688980957
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_104_41
timestamp 1688980957
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104_53
timestamp 1688980957
transform 1 0 5980 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104_61
timestamp 1688980957
transform 1 0 6716 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104_88
timestamp 1688980957
transform 1 0 9200 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_104_92
timestamp 1688980957
transform 1 0 9568 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_3
timestamp 1688980957
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_15
timestamp 1688980957
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_27
timestamp 1688980957
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_105_39
timestamp 1688980957
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105_51
timestamp 1688980957
transform 1 0 5796 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105_57
timestamp 1688980957
transform 1 0 6348 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105_69
timestamp 1688980957
transform 1 0 7452 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105_84
timestamp 1688980957
transform 1 0 8832 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_105_92
timestamp 1688980957
transform 1 0 9568 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_9
timestamp 1688980957
transform 1 0 1932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106_21
timestamp 1688980957
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_27
timestamp 1688980957
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_106_29
timestamp 1688980957
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106_41
timestamp 1688980957
transform 1 0 4876 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106_63
timestamp 1688980957
transform 1 0 6900 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_106_81
timestamp 1688980957
transform 1 0 8556 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106_85
timestamp 1688980957
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_3
timestamp 1688980957
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_15
timestamp 1688980957
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107_27
timestamp 1688980957
transform 1 0 3588 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_32
timestamp 1688980957
transform 1 0 4048 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_36
timestamp 1688980957
transform 1 0 4416 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_107_40
timestamp 1688980957
transform 1 0 4784 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107_46
timestamp 1688980957
transform 1 0 5336 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107_54
timestamp 1688980957
transform 1 0 6072 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_107_57
timestamp 1688980957
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107_69
timestamp 1688980957
transform 1 0 7452 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_9
timestamp 1688980957
transform 1 0 1932 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_108_21
timestamp 1688980957
transform 1 0 3036 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_27
timestamp 1688980957
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_29
timestamp 1688980957
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_41
timestamp 1688980957
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_108_53
timestamp 1688980957
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108_65
timestamp 1688980957
transform 1 0 7084 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108_83
timestamp 1688980957
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108_85
timestamp 1688980957
transform 1 0 8924 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_6
timestamp 1688980957
transform 1 0 1656 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_18
timestamp 1688980957
transform 1 0 2760 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109_30
timestamp 1688980957
transform 1 0 3864 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_109_45
timestamp 1688980957
transform 1 0 5244 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109_53
timestamp 1688980957
transform 1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_57
timestamp 1688980957
transform 1 0 6348 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_109_77
timestamp 1688980957
transform 1 0 8188 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_109_89
timestamp 1688980957
transform 1 0 9292 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_3
timestamp 1688980957
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_15
timestamp 1688980957
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_27
timestamp 1688980957
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_29
timestamp 1688980957
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_41
timestamp 1688980957
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_110_53
timestamp 1688980957
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_65
timestamp 1688980957
transform 1 0 7084 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_110_88
timestamp 1688980957
transform 1 0 9200 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110_92
timestamp 1688980957
transform 1 0 9568 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_7
timestamp 1688980957
transform 1 0 1748 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_19
timestamp 1688980957
transform 1 0 2852 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_31
timestamp 1688980957
transform 1 0 3956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_111_43
timestamp 1688980957
transform 1 0 5060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111_55
timestamp 1688980957
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_111_57
timestamp 1688980957
transform 1 0 6348 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_111_85
timestamp 1688980957
transform 1 0 8924 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_3
timestamp 1688980957
transform 1 0 1380 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_14
timestamp 1688980957
transform 1 0 2392 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_112_26
timestamp 1688980957
transform 1 0 3496 0 1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_29
timestamp 1688980957
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_112_41
timestamp 1688980957
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_112_53
timestamp 1688980957
transform 1 0 5980 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112_59
timestamp 1688980957
transform 1 0 6532 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_112_81
timestamp 1688980957
transform 1 0 8556 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_112_85
timestamp 1688980957
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_9
timestamp 1688980957
transform 1 0 1932 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_21
timestamp 1688980957
transform 1 0 3036 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_33
timestamp 1688980957
transform 1 0 4140 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113_39
timestamp 1688980957
transform 1 0 4692 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113_44
timestamp 1688980957
transform 1 0 5152 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113_57
timestamp 1688980957
transform 1 0 6348 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113_87
timestamp 1688980957
transform 1 0 9108 0 -1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_3
timestamp 1688980957
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_15
timestamp 1688980957
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_27
timestamp 1688980957
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_29
timestamp 1688980957
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_114_41
timestamp 1688980957
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_53
timestamp 1688980957
transform 1 0 5980 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114_57
timestamp 1688980957
transform 1 0 6348 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_114_67
timestamp 1688980957
transform 1 0 7268 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114_73
timestamp 1688980957
transform 1 0 7820 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_114_85
timestamp 1688980957
transform 1 0 8924 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_7
timestamp 1688980957
transform 1 0 1748 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_19
timestamp 1688980957
transform 1 0 2852 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_31
timestamp 1688980957
transform 1 0 3956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_115_43
timestamp 1688980957
transform 1 0 5060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_55
timestamp 1688980957
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115_57
timestamp 1688980957
transform 1 0 6348 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_74
timestamp 1688980957
transform 1 0 7912 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115_78
timestamp 1688980957
transform 1 0 8280 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115_89
timestamp 1688980957
transform 1 0 9292 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_7
timestamp 1688980957
transform 1 0 1748 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_19
timestamp 1688980957
transform 1 0 2852 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_27
timestamp 1688980957
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116_29
timestamp 1688980957
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_41
timestamp 1688980957
transform 1 0 4876 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_49
timestamp 1688980957
transform 1 0 5612 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_66
timestamp 1688980957
transform 1 0 7176 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116_74
timestamp 1688980957
transform 1 0 7912 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116_85
timestamp 1688980957
transform 1 0 8924 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_3
timestamp 1688980957
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_15
timestamp 1688980957
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_117_27
timestamp 1688980957
transform 1 0 3588 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_33
timestamp 1688980957
transform 1 0 4140 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117_40
timestamp 1688980957
transform 1 0 4784 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_44
timestamp 1688980957
transform 1 0 5152 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117_55
timestamp 1688980957
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_117_57
timestamp 1688980957
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117_78
timestamp 1688980957
transform 1 0 8280 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117_82
timestamp 1688980957
transform 1 0 8648 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_7
timestamp 1688980957
transform 1 0 1748 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_19
timestamp 1688980957
transform 1 0 2852 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_27
timestamp 1688980957
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_29
timestamp 1688980957
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_118_41
timestamp 1688980957
transform 1 0 4876 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118_50
timestamp 1688980957
transform 1 0 5704 0 1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118_68
timestamp 1688980957
transform 1 0 7360 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118_80
timestamp 1688980957
transform 1 0 8464 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118_85
timestamp 1688980957
transform 1 0 8924 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_3
timestamp 1688980957
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_15
timestamp 1688980957
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119_27
timestamp 1688980957
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119_39
timestamp 1688980957
transform 1 0 4692 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119_43
timestamp 1688980957
transform 1 0 5060 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_119_57
timestamp 1688980957
transform 1 0 6348 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_119_65
timestamp 1688980957
transform 1 0 7084 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119_85
timestamp 1688980957
transform 1 0 8924 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120_7
timestamp 1688980957
transform 1 0 1748 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_19
timestamp 1688980957
transform 1 0 2852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120_27
timestamp 1688980957
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_29
timestamp 1688980957
transform 1 0 3772 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_37
timestamp 1688980957
transform 1 0 4508 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_120_43
timestamp 1688980957
transform 1 0 5060 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_120_51
timestamp 1688980957
transform 1 0 5796 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120_64
timestamp 1688980957
transform 1 0 6992 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_3
timestamp 1688980957
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_121_15
timestamp 1688980957
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_121_27
timestamp 1688980957
transform 1 0 3588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121_33
timestamp 1688980957
transform 1 0 4140 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121_57
timestamp 1688980957
transform 1 0 6348 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121_67
timestamp 1688980957
transform 1 0 7268 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121_71
timestamp 1688980957
transform 1 0 7636 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121_91
timestamp 1688980957
transform 1 0 9476 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_7
timestamp 1688980957
transform 1 0 1748 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_19
timestamp 1688980957
transform 1 0 2852 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_27
timestamp 1688980957
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_29
timestamp 1688980957
transform 1 0 3772 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122_43
timestamp 1688980957
transform 1 0 5060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_55
timestamp 1688980957
transform 1 0 6164 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_122_63
timestamp 1688980957
transform 1 0 6900 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_69
timestamp 1688980957
transform 1 0 7452 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122_79
timestamp 1688980957
transform 1 0 8372 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122_83
timestamp 1688980957
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_122_85
timestamp 1688980957
transform 1 0 8924 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_7
timestamp 1688980957
transform 1 0 1748 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_19
timestamp 1688980957
transform 1 0 2852 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123_31
timestamp 1688980957
transform 1 0 3956 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_39
timestamp 1688980957
transform 1 0 4692 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_43
timestamp 1688980957
transform 1 0 5060 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123_55
timestamp 1688980957
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_57
timestamp 1688980957
transform 1 0 6348 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123_69
timestamp 1688980957
transform 1 0 7452 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_123_81
timestamp 1688980957
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_3
timestamp 1688980957
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_124_15
timestamp 1688980957
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_27
timestamp 1688980957
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_124_29
timestamp 1688980957
transform 1 0 3772 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124_51
timestamp 1688980957
transform 1 0 5796 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124_55
timestamp 1688980957
transform 1 0 6164 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_124_75
timestamp 1688980957
transform 1 0 8004 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124_79
timestamp 1688980957
transform 1 0 8372 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_83
timestamp 1688980957
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124_88
timestamp 1688980957
transform 1 0 9200 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124_92
timestamp 1688980957
transform 1 0 9568 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_7
timestamp 1688980957
transform 1 0 1748 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_19
timestamp 1688980957
transform 1 0 2852 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_31
timestamp 1688980957
transform 1 0 3956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125_43
timestamp 1688980957
transform 1 0 5060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125_55
timestamp 1688980957
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125_66
timestamp 1688980957
transform 1 0 7176 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125_72
timestamp 1688980957
transform 1 0 7728 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125_91
timestamp 1688980957
transform 1 0 9476 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_3
timestamp 1688980957
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_15
timestamp 1688980957
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_27
timestamp 1688980957
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_126_29
timestamp 1688980957
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126_41
timestamp 1688980957
transform 1 0 4876 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126_45
timestamp 1688980957
transform 1 0 5244 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_126_81
timestamp 1688980957
transform 1 0 8556 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126_85
timestamp 1688980957
transform 1 0 8924 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_126_89
timestamp 1688980957
transform 1 0 9292 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_7
timestamp 1688980957
transform 1 0 1748 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_19
timestamp 1688980957
transform 1 0 2852 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_31
timestamp 1688980957
transform 1 0 3956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_127_43
timestamp 1688980957
transform 1 0 5060 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_55
timestamp 1688980957
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127_57
timestamp 1688980957
transform 1 0 6348 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_61
timestamp 1688980957
transform 1 0 6716 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127_70
timestamp 1688980957
transform 1 0 7544 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127_79
timestamp 1688980957
transform 1 0 8372 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_3
timestamp 1688980957
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_15
timestamp 1688980957
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128_27
timestamp 1688980957
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_29
timestamp 1688980957
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128_41
timestamp 1688980957
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_128_53
timestamp 1688980957
transform 1 0 5980 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_128_69
timestamp 1688980957
transform 1 0 7452 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_128_73
timestamp 1688980957
transform 1 0 7820 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_128_91
timestamp 1688980957
transform 1 0 9476 0 1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_7
timestamp 1688980957
transform 1 0 1748 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_19
timestamp 1688980957
transform 1 0 2852 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_31
timestamp 1688980957
transform 1 0 3956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_129_43
timestamp 1688980957
transform 1 0 5060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129_55
timestamp 1688980957
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_129_81
timestamp 1688980957
transform 1 0 8556 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_7
timestamp 1688980957
transform 1 0 1748 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_19
timestamp 1688980957
transform 1 0 2852 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_27
timestamp 1688980957
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_130_29
timestamp 1688980957
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130_41
timestamp 1688980957
transform 1 0 4876 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_45
timestamp 1688980957
transform 1 0 5244 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_56
timestamp 1688980957
transform 1 0 6256 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_130_74
timestamp 1688980957
transform 1 0 7912 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130_79
timestamp 1688980957
transform 1 0 8372 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_130_83
timestamp 1688980957
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130_85
timestamp 1688980957
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_3
timestamp 1688980957
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_15
timestamp 1688980957
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_27
timestamp 1688980957
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_131_39
timestamp 1688980957
transform 1 0 4692 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131_51
timestamp 1688980957
transform 1 0 5796 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_55
timestamp 1688980957
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_57
timestamp 1688980957
transform 1 0 6348 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131_73
timestamp 1688980957
transform 1 0 7820 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131_91
timestamp 1688980957
transform 1 0 9476 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_7
timestamp 1688980957
transform 1 0 1748 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132_19
timestamp 1688980957
transform 1 0 2852 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_27
timestamp 1688980957
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_132_29
timestamp 1688980957
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_132_41
timestamp 1688980957
transform 1 0 4876 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_47
timestamp 1688980957
transform 1 0 5428 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_132_58
timestamp 1688980957
transform 1 0 6440 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_132_71
timestamp 1688980957
transform 1 0 7636 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_132_81
timestamp 1688980957
transform 1 0 8556 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132_92
timestamp 1688980957
transform 1 0 9568 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_3
timestamp 1688980957
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_15
timestamp 1688980957
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_27
timestamp 1688980957
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_133_39
timestamp 1688980957
transform 1 0 4692 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_51
timestamp 1688980957
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_55
timestamp 1688980957
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133_57
timestamp 1688980957
transform 1 0 6348 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133_67
timestamp 1688980957
transform 1 0 7268 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133_78
timestamp 1688980957
transform 1 0 8280 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133_82
timestamp 1688980957
transform 1 0 8648 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_7
timestamp 1688980957
transform 1 0 1748 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134_19
timestamp 1688980957
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134_27
timestamp 1688980957
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_29
timestamp 1688980957
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_41
timestamp 1688980957
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_53
timestamp 1688980957
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_134_65
timestamp 1688980957
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134_77
timestamp 1688980957
transform 1 0 8188 0 1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_3
timestamp 1688980957
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_15
timestamp 1688980957
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_27
timestamp 1688980957
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_39
timestamp 1688980957
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135_51
timestamp 1688980957
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_55
timestamp 1688980957
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_135_57
timestamp 1688980957
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_135_69
timestamp 1688980957
transform 1 0 7452 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135_75
timestamp 1688980957
transform 1 0 8004 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_7
timestamp 1688980957
transform 1 0 1748 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_136_19
timestamp 1688980957
transform 1 0 2852 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_27
timestamp 1688980957
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_29
timestamp 1688980957
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_41
timestamp 1688980957
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_53
timestamp 1688980957
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_136_65
timestamp 1688980957
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_136_77
timestamp 1688980957
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136_83
timestamp 1688980957
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_7
timestamp 1688980957
transform 1 0 1748 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_19
timestamp 1688980957
transform 1 0 2852 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_31
timestamp 1688980957
transform 1 0 3956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_43
timestamp 1688980957
transform 1 0 5060 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137_55
timestamp 1688980957
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_57
timestamp 1688980957
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_69
timestamp 1688980957
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_137_81
timestamp 1688980957
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_3
timestamp 1688980957
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_15
timestamp 1688980957
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_138_27
timestamp 1688980957
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_29
timestamp 1688980957
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_41
timestamp 1688980957
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_138_53
timestamp 1688980957
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_65
timestamp 1688980957
transform 1 0 7084 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138_73
timestamp 1688980957
transform 1 0 7820 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_138_85
timestamp 1688980957
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_7
timestamp 1688980957
transform 1 0 1748 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_19
timestamp 1688980957
transform 1 0 2852 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_31
timestamp 1688980957
transform 1 0 3956 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_43
timestamp 1688980957
transform 1 0 5060 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139_55
timestamp 1688980957
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_57
timestamp 1688980957
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_139_69
timestamp 1688980957
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_139_81
timestamp 1688980957
transform 1 0 8556 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_3
timestamp 1688980957
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_15
timestamp 1688980957
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_27
timestamp 1688980957
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_29
timestamp 1688980957
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_41
timestamp 1688980957
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_53
timestamp 1688980957
transform 1 0 5980 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_140_65
timestamp 1688980957
transform 1 0 7084 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_140_77
timestamp 1688980957
transform 1 0 8188 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_140_83
timestamp 1688980957
transform 1 0 8740 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_140_85
timestamp 1688980957
transform 1 0 8924 0 1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_7
timestamp 1688980957
transform 1 0 1748 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_19
timestamp 1688980957
transform 1 0 2852 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_31
timestamp 1688980957
transform 1 0 3956 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_43
timestamp 1688980957
transform 1 0 5060 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141_55
timestamp 1688980957
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_57
timestamp 1688980957
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_69
timestamp 1688980957
transform 1 0 7452 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141_81
timestamp 1688980957
transform 1 0 8556 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_3
timestamp 1688980957
transform 1 0 1380 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_15
timestamp 1688980957
transform 1 0 2484 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_27
timestamp 1688980957
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_29
timestamp 1688980957
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_41
timestamp 1688980957
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_53
timestamp 1688980957
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_142_65
timestamp 1688980957
transform 1 0 7084 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_142_77
timestamp 1688980957
transform 1 0 8188 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_142_83
timestamp 1688980957
transform 1 0 8740 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_142_85
timestamp 1688980957
transform 1 0 8924 0 1 78336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_7
timestamp 1688980957
transform 1 0 1748 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_19
timestamp 1688980957
transform 1 0 2852 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_31
timestamp 1688980957
transform 1 0 3956 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_43
timestamp 1688980957
transform 1 0 5060 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143_55
timestamp 1688980957
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_57
timestamp 1688980957
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_69
timestamp 1688980957
transform 1 0 7452 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_143_81
timestamp 1688980957
transform 1 0 8556 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_7
timestamp 1688980957
transform 1 0 1748 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144_19
timestamp 1688980957
transform 1 0 2852 0 1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_27
timestamp 1688980957
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_29
timestamp 1688980957
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_41
timestamp 1688980957
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_53
timestamp 1688980957
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_144_65
timestamp 1688980957
transform 1 0 7084 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_144_77
timestamp 1688980957
transform 1 0 8188 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144_83
timestamp 1688980957
transform 1 0 8740 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144_85
timestamp 1688980957
transform 1 0 8924 0 1 79424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_3
timestamp 1688980957
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_15
timestamp 1688980957
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_27
timestamp 1688980957
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_39
timestamp 1688980957
transform 1 0 4692 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145_51
timestamp 1688980957
transform 1 0 5796 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145_55
timestamp 1688980957
transform 1 0 6164 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_57
timestamp 1688980957
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_69
timestamp 1688980957
transform 1 0 7452 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_145_81
timestamp 1688980957
transform 1 0 8556 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_7
timestamp 1688980957
transform 1 0 1748 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146_19
timestamp 1688980957
transform 1 0 2852 0 1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_27
timestamp 1688980957
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_29
timestamp 1688980957
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_41
timestamp 1688980957
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_53
timestamp 1688980957
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_146_65
timestamp 1688980957
transform 1 0 7084 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146_77
timestamp 1688980957
transform 1 0 8188 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146_83
timestamp 1688980957
transform 1 0 8740 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146_85
timestamp 1688980957
transform 1 0 8924 0 1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_3
timestamp 1688980957
transform 1 0 1380 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_15
timestamp 1688980957
transform 1 0 2484 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_27
timestamp 1688980957
transform 1 0 3588 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_39
timestamp 1688980957
transform 1 0 4692 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147_51
timestamp 1688980957
transform 1 0 5796 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147_55
timestamp 1688980957
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_57
timestamp 1688980957
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_69
timestamp 1688980957
transform 1 0 7452 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147_81
timestamp 1688980957
transform 1 0 8556 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_7
timestamp 1688980957
transform 1 0 1748 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_148_19
timestamp 1688980957
transform 1 0 2852 0 1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_27
timestamp 1688980957
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_29
timestamp 1688980957
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_41
timestamp 1688980957
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_53
timestamp 1688980957
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_148_65
timestamp 1688980957
transform 1 0 7084 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_148_77
timestamp 1688980957
transform 1 0 8188 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148_83
timestamp 1688980957
transform 1 0 8740 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_148_85
timestamp 1688980957
transform 1 0 8924 0 1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_3
timestamp 1688980957
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_15
timestamp 1688980957
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_27
timestamp 1688980957
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_39
timestamp 1688980957
transform 1 0 4692 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149_51
timestamp 1688980957
transform 1 0 5796 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149_55
timestamp 1688980957
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_57
timestamp 1688980957
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_69
timestamp 1688980957
transform 1 0 7452 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_149_81
timestamp 1688980957
transform 1 0 8556 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_7
timestamp 1688980957
transform 1 0 1748 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_150_19
timestamp 1688980957
transform 1 0 2852 0 1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_27
timestamp 1688980957
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_29
timestamp 1688980957
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_41
timestamp 1688980957
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_53
timestamp 1688980957
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_150_65
timestamp 1688980957
transform 1 0 7084 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_150_77
timestamp 1688980957
transform 1 0 8188 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_150_83
timestamp 1688980957
transform 1 0 8740 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_150_85
timestamp 1688980957
transform 1 0 8924 0 1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_7
timestamp 1688980957
transform 1 0 1748 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_19
timestamp 1688980957
transform 1 0 2852 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_31
timestamp 1688980957
transform 1 0 3956 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_43
timestamp 1688980957
transform 1 0 5060 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151_55
timestamp 1688980957
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_57
timestamp 1688980957
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_69
timestamp 1688980957
transform 1 0 7452 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_151_81
timestamp 1688980957
transform 1 0 8556 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_3
timestamp 1688980957
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_15
timestamp 1688980957
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_27
timestamp 1688980957
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_29
timestamp 1688980957
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_41
timestamp 1688980957
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_53
timestamp 1688980957
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_152_65
timestamp 1688980957
transform 1 0 7084 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_152_77
timestamp 1688980957
transform 1 0 8188 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152_83
timestamp 1688980957
transform 1 0 8740 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_152_85
timestamp 1688980957
transform 1 0 8924 0 1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_7
timestamp 1688980957
transform 1 0 1748 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_19
timestamp 1688980957
transform 1 0 2852 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_31
timestamp 1688980957
transform 1 0 3956 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_43
timestamp 1688980957
transform 1 0 5060 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153_55
timestamp 1688980957
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_57
timestamp 1688980957
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_69
timestamp 1688980957
transform 1 0 7452 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153_81
timestamp 1688980957
transform 1 0 8556 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_3
timestamp 1688980957
transform 1 0 1380 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_15
timestamp 1688980957
transform 1 0 2484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_27
timestamp 1688980957
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_29
timestamp 1688980957
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_41
timestamp 1688980957
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_53
timestamp 1688980957
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154_65
timestamp 1688980957
transform 1 0 7084 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154_77
timestamp 1688980957
transform 1 0 8188 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154_83
timestamp 1688980957
transform 1 0 8740 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_154_85
timestamp 1688980957
transform 1 0 8924 0 1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_3
timestamp 1688980957
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_15
timestamp 1688980957
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_27
timestamp 1688980957
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_39
timestamp 1688980957
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_155_51
timestamp 1688980957
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155_55
timestamp 1688980957
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_57
timestamp 1688980957
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_69
timestamp 1688980957
transform 1 0 7452 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_155_81
timestamp 1688980957
transform 1 0 8556 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_3
timestamp 1688980957
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_15
timestamp 1688980957
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_27
timestamp 1688980957
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_29
timestamp 1688980957
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_41
timestamp 1688980957
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_53
timestamp 1688980957
transform 1 0 5980 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_57
timestamp 1688980957
transform 1 0 6348 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_69
timestamp 1688980957
transform 1 0 7452 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_81
timestamp 1688980957
transform 1 0 8556 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_85
timestamp 1688980957
transform 1 0 8924 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_97
timestamp 1688980957
transform 1 0 10028 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_109
timestamp 1688980957
transform 1 0 11132 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_113
timestamp 1688980957
transform 1 0 11500 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_125
timestamp 1688980957
transform 1 0 12604 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_137
timestamp 1688980957
transform 1 0 13708 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_141
timestamp 1688980957
transform 1 0 14076 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_153
timestamp 1688980957
transform 1 0 15180 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_165
timestamp 1688980957
transform 1 0 16284 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_169
timestamp 1688980957
transform 1 0 16652 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_181
timestamp 1688980957
transform 1 0 17756 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_193
timestamp 1688980957
transform 1 0 18860 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_197
timestamp 1688980957
transform 1 0 19228 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_207
timestamp 1688980957
transform 1 0 20148 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_219
timestamp 1688980957
transform 1 0 21252 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_223
timestamp 1688980957
transform 1 0 21620 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_225
timestamp 1688980957
transform 1 0 21804 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_237
timestamp 1688980957
transform 1 0 22908 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_249
timestamp 1688980957
transform 1 0 24012 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_262
timestamp 1688980957
transform 1 0 25208 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156_274
timestamp 1688980957
transform 1 0 26312 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_290
timestamp 1688980957
transform 1 0 27784 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156_302
timestamp 1688980957
transform 1 0 28888 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_309
timestamp 1688980957
transform 1 0 29532 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_321
timestamp 1688980957
transform 1 0 30636 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_333
timestamp 1688980957
transform 1 0 31740 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_337
timestamp 1688980957
transform 1 0 32108 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_349
timestamp 1688980957
transform 1 0 33212 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_361
timestamp 1688980957
transform 1 0 34316 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_365
timestamp 1688980957
transform 1 0 34684 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156_385
timestamp 1688980957
transform 1 0 36524 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_391
timestamp 1688980957
transform 1 0 37076 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156_402
timestamp 1688980957
transform 1 0 38088 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_412
timestamp 1688980957
transform 1 0 39008 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_416
timestamp 1688980957
transform 1 0 39376 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_421
timestamp 1688980957
transform 1 0 39836 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_425
timestamp 1688980957
transform 1 0 40204 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_445
timestamp 1688980957
transform 1 0 42044 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_449
timestamp 1688980957
transform 1 0 42412 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_453
timestamp 1688980957
transform 1 0 42780 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_456
timestamp 1688980957
transform 1 0 43056 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_497
timestamp 1688980957
transform 1 0 46828 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_501
timestamp 1688980957
transform 1 0 47196 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_505
timestamp 1688980957
transform 1 0 47564 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_524
timestamp 1688980957
transform 1 0 49312 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_528
timestamp 1688980957
transform 1 0 49680 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_533
timestamp 1688980957
transform 1 0 50140 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_537
timestamp 1688980957
transform 1 0 50508 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_541
timestamp 1688980957
transform 1 0 50876 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_546
timestamp 1688980957
transform 1 0 51336 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_550
timestamp 1688980957
transform 1 0 51704 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_554
timestamp 1688980957
transform 1 0 52072 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_561
timestamp 1688980957
transform 1 0 52716 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156_566
timestamp 1688980957
transform 1 0 53176 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156_605
timestamp 1688980957
transform 1 0 56764 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_613
timestamp 1688980957
transform 1 0 57500 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_617
timestamp 1688980957
transform 1 0 57868 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_629
timestamp 1688980957
transform 1 0 58972 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_641
timestamp 1688980957
transform 1 0 60076 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156_645
timestamp 1688980957
transform 1 0 60444 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_655
timestamp 1688980957
transform 1 0 61364 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_667
timestamp 1688980957
transform 1 0 62468 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_671
timestamp 1688980957
transform 1 0 62836 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_673
timestamp 1688980957
transform 1 0 63020 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_685
timestamp 1688980957
transform 1 0 64124 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_697
timestamp 1688980957
transform 1 0 65228 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_701
timestamp 1688980957
transform 1 0 65596 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_713
timestamp 1688980957
transform 1 0 66700 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_725
timestamp 1688980957
transform 1 0 67804 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_729
timestamp 1688980957
transform 1 0 68172 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_741
timestamp 1688980957
transform 1 0 69276 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_753
timestamp 1688980957
transform 1 0 70380 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_757
timestamp 1688980957
transform 1 0 70748 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_769
timestamp 1688980957
transform 1 0 71852 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_781
timestamp 1688980957
transform 1 0 72956 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_785
timestamp 1688980957
transform 1 0 73324 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_797
timestamp 1688980957
transform 1 0 74428 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_809
timestamp 1688980957
transform 1 0 75532 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_813
timestamp 1688980957
transform 1 0 75900 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_825
timestamp 1688980957
transform 1 0 77004 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_837
timestamp 1688980957
transform 1 0 78108 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_841
timestamp 1688980957
transform 1 0 78476 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_853
timestamp 1688980957
transform 1 0 79580 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_865
timestamp 1688980957
transform 1 0 80684 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_869
timestamp 1688980957
transform 1 0 81052 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_881
timestamp 1688980957
transform 1 0 82156 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_893
timestamp 1688980957
transform 1 0 83260 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_897
timestamp 1688980957
transform 1 0 83628 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_909
timestamp 1688980957
transform 1 0 84732 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_921
timestamp 1688980957
transform 1 0 85836 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_925
timestamp 1688980957
transform 1 0 86204 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_937
timestamp 1688980957
transform 1 0 87308 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_949
timestamp 1688980957
transform 1 0 88412 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_953
timestamp 1688980957
transform 1 0 88780 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_965
timestamp 1688980957
transform 1 0 89884 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_977
timestamp 1688980957
transform 1 0 90988 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_981
timestamp 1688980957
transform 1 0 91356 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_993
timestamp 1688980957
transform 1 0 92460 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1005
timestamp 1688980957
transform 1 0 93564 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1009
timestamp 1688980957
transform 1 0 93932 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1021
timestamp 1688980957
transform 1 0 95036 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1033
timestamp 1688980957
transform 1 0 96140 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1037
timestamp 1688980957
transform 1 0 96508 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1049
timestamp 1688980957
transform 1 0 97612 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1061
timestamp 1688980957
transform 1 0 98716 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1065
timestamp 1688980957
transform 1 0 99084 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1077
timestamp 1688980957
transform 1 0 100188 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1089
timestamp 1688980957
transform 1 0 101292 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1093
timestamp 1688980957
transform 1 0 101660 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1105
timestamp 1688980957
transform 1 0 102764 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1117
timestamp 1688980957
transform 1 0 103868 0 1 85952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1121
timestamp 1688980957
transform 1 0 104236 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156_1133
timestamp 1688980957
transform 1 0 105340 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1145
timestamp 1688980957
transform 1 0 106444 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156_1149
timestamp 1688980957
transform 1 0 106812 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156_1157
timestamp 1688980957
transform 1 0 107548 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156_1163
timestamp 1688980957
transform 1 0 108100 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156_1167
timestamp 1688980957
transform 1 0 108468 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1380 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1688980957
transform 1 0 1380 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1688980957
transform 1 0 1380 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1688980957
transform 1 0 1380 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1688980957
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1688980957
transform 1 0 1380 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1688980957
transform 1 0 1380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1688980957
transform 1 0 1380 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1688980957
transform 1 0 1380 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 1380 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1688980957
transform 1 0 1380 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1688980957
transform 1 0 1380 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1688980957
transform 1 0 1380 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1688980957
transform 1 0 1380 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1688980957
transform 1 0 1380 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1688980957
transform 1 0 1380 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1688980957
transform 1 0 1380 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 1688980957
transform 1 0 1380 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1688980957
transform 1 0 1380 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1688980957
transform 1 0 1380 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1688980957
transform 1 0 1380 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1688980957
transform 1 0 1380 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input45
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1688980957
transform 1 0 1380 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1688980957
transform 1 0 1380 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input48
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input49
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input50
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_sram_1kbyte_1rw1r_32x256_8  memory_cell
timestamp 0
transform 1 0 12000 0 1 4000
box 0 0 95956 79500
use sky130_fd_sc_hd__conb_1  memory_cell_87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 107824 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output56
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output57
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 1380 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform 1 0 1380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1688980957
transform 1 0 1380 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 1380 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 1380 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 1380 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 1380 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 1380 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 1380 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 1380 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 1380 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 108836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 9936 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 9936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 9936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 9936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 9936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 9936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 9936 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 9936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 9936 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 9936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 9936 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 9936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 9936 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 9936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 9936 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 9936 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 9936 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 9936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 9936 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 9936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 9936 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 9936 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 9936 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 9936 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 9936 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 9936 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 9936 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 9936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 9936 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 9936 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 9936 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 9936 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 9936 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 9936 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 9936 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 9936 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 9936 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 9936 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 9936 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 9936 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 9936 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 9936 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1688980957
transform -1 0 9936 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1688980957
transform -1 0 9936 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1688980957
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1688980957
transform -1 0 9936 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1688980957
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1688980957
transform -1 0 9936 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1688980957
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1688980957
transform -1 0 9936 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1688980957
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1688980957
transform -1 0 9936 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1688980957
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1688980957
transform -1 0 9936 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1688980957
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1688980957
transform -1 0 9936 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1688980957
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1688980957
transform -1 0 9936 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1688980957
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1688980957
transform -1 0 9936 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1688980957
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1688980957
transform -1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1688980957
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1688980957
transform -1 0 9936 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1688980957
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1688980957
transform -1 0 9936 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1688980957
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1688980957
transform -1 0 9936 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1688980957
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1688980957
transform -1 0 9936 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1688980957
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1688980957
transform -1 0 9936 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1688980957
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1688980957
transform -1 0 9936 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1688980957
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1688980957
transform -1 0 9936 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1688980957
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1688980957
transform -1 0 9936 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1688980957
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1688980957
transform -1 0 9936 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1688980957
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1688980957
transform -1 0 9936 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1688980957
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1688980957
transform -1 0 9936 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1688980957
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1688980957
transform -1 0 9936 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1688980957
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1688980957
transform -1 0 9936 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1688980957
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1688980957
transform -1 0 9936 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1688980957
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1688980957
transform -1 0 9936 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1688980957
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1688980957
transform -1 0 9936 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1688980957
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1688980957
transform -1 0 9936 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1688980957
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1688980957
transform -1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1688980957
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1688980957
transform -1 0 9936 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1688980957
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1688980957
transform -1 0 9936 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1688980957
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1688980957
transform -1 0 9936 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1688980957
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1688980957
transform -1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1688980957
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1688980957
transform -1 0 9936 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1688980957
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1688980957
transform -1 0 9936 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1688980957
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1688980957
transform -1 0 9936 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1688980957
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1688980957
transform -1 0 9936 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1688980957
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1688980957
transform -1 0 9936 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1688980957
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1688980957
transform -1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1688980957
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1688980957
transform -1 0 9936 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1688980957
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1688980957
transform -1 0 9936 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1688980957
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1688980957
transform -1 0 9936 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1688980957
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1688980957
transform -1 0 9936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1688980957
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1688980957
transform -1 0 9936 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1688980957
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1688980957
transform -1 0 9936 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1688980957
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1688980957
transform -1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1688980957
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1688980957
transform -1 0 9936 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1688980957
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1688980957
transform -1 0 9936 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1688980957
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1688980957
transform -1 0 9936 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1688980957
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1688980957
transform -1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1688980957
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1688980957
transform -1 0 9936 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1688980957
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1688980957
transform -1 0 9936 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1688980957
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1688980957
transform -1 0 9936 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1688980957
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1688980957
transform -1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1688980957
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1688980957
transform -1 0 9936 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1688980957
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1688980957
transform -1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1688980957
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1688980957
transform -1 0 9936 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1688980957
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1688980957
transform -1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1688980957
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1688980957
transform -1 0 9936 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1688980957
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1688980957
transform -1 0 9936 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1688980957
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1688980957
transform -1 0 9936 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1688980957
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1688980957
transform -1 0 9936 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1688980957
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1688980957
transform -1 0 9936 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1688980957
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1688980957
transform -1 0 9936 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1688980957
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1688980957
transform -1 0 9936 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1688980957
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1688980957
transform -1 0 9936 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1688980957
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1688980957
transform -1 0 9936 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1688980957
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1688980957
transform -1 0 9936 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1688980957
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1688980957
transform -1 0 9936 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1688980957
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1688980957
transform -1 0 9936 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1688980957
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1688980957
transform -1 0 9936 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1688980957
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1688980957
transform -1 0 9936 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1688980957
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1688980957
transform -1 0 9936 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1688980957
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1688980957
transform -1 0 9936 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1688980957
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1688980957
transform -1 0 9936 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1688980957
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1688980957
transform -1 0 108836 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 47472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 50048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 52624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 55200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 57776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 60352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 62928 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 65504 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 68080 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 70656 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 73232 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 75808 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 78384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 80960 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 83536 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 86112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 88688 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 91264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 93840 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 96416 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 98992 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 101568 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 104144 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 106720 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 8832 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 8832 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 8832 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 8832 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 8832 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 8832 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 8832 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 6256 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 8832 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 11408 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 13984 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 16560 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 19136 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 21712 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 26864 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 29440 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 32016 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 34592 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 37168 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 39744 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 42320 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 44896 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 47472 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 50048 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 52624 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 55200 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 57776 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 60352 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 62928 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 65504 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 68080 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 70656 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 73232 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 75808 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 78384 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 80960 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 83536 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 86112 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 88688 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 91264 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 93840 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 96416 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 98992 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 101568 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 104144 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 106720 0 1 85952
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 22478 800 22538 0 FreeSans 480 0 0 0 C0
port 0 nsew signal input
flabel metal3 s 0 23430 800 23490 0 FreeSans 480 0 0 0 C1
port 1 nsew signal input
flabel metal3 s 0 24382 800 24442 0 FreeSans 480 0 0 0 C2
port 2 nsew signal input
flabel metal3 s 0 25334 800 25394 0 FreeSans 480 0 0 0 C3
port 3 nsew signal input
flabel metal3 s 0 60558 800 60618 0 FreeSans 480 0 0 0 C4
port 4 nsew signal input
flabel metal3 s 0 61510 800 61570 0 FreeSans 480 0 0 0 C5
port 5 nsew signal input
flabel metal2 s 54956 0 54984 800 0 FreeSans 224 90 0 0 clk
port 6 nsew signal input
flabel metal3 s 0 18670 800 18730 0 FreeSans 480 0 0 0 rd_addr[0]
port 7 nsew signal input
flabel metal3 s 0 19622 800 19682 0 FreeSans 480 0 0 0 rd_addr[1]
port 8 nsew signal input
flabel metal3 s 0 20574 800 20634 0 FreeSans 480 0 0 0 rd_addr[2]
port 9 nsew signal input
flabel metal3 s 0 21526 800 21586 0 FreeSans 480 0 0 0 rd_addr[3]
port 10 nsew signal input
flabel metal3 s 0 26286 800 26346 0 FreeSans 480 0 0 0 rd_addr[4]
port 11 nsew signal input
flabel metal3 s 0 27238 800 27298 0 FreeSans 480 0 0 0 rd_addr[5]
port 12 nsew signal input
flabel metal3 s 0 35806 800 35866 0 FreeSans 480 0 0 0 rd_addr[6]
port 13 nsew signal input
flabel metal3 s 0 36758 800 36818 0 FreeSans 480 0 0 0 rd_addr[7]
port 14 nsew signal input
flabel metal3 s 0 17718 800 17778 0 FreeSans 480 0 0 0 rd_data[0]
port 15 nsew signal tristate
flabel metal3 s 0 8198 800 8258 0 FreeSans 480 0 0 0 rd_data[10]
port 16 nsew signal tristate
flabel metal3 s 0 7246 800 7306 0 FreeSans 480 0 0 0 rd_data[11]
port 17 nsew signal tristate
flabel metal3 s 0 3438 800 3498 0 FreeSans 480 0 0 0 rd_data[12]
port 18 nsew signal tristate
flabel metal3 s 0 4390 800 4450 0 FreeSans 480 0 0 0 rd_data[13]
port 19 nsew signal tristate
flabel metal3 s 0 5342 800 5402 0 FreeSans 480 0 0 0 rd_data[14]
port 20 nsew signal tristate
flabel metal3 s 0 6294 800 6354 0 FreeSans 480 0 0 0 rd_data[15]
port 21 nsew signal tristate
flabel metal3 s 0 45326 800 45386 0 FreeSans 480 0 0 0 rd_data[16]
port 22 nsew signal tristate
flabel metal3 s 0 46278 800 46338 0 FreeSans 480 0 0 0 rd_data[17]
port 23 nsew signal tristate
flabel metal3 s 0 47230 800 47290 0 FreeSans 480 0 0 0 rd_data[18]
port 24 nsew signal tristate
flabel metal3 s 0 48182 800 48242 0 FreeSans 480 0 0 0 rd_data[19]
port 25 nsew signal tristate
flabel metal3 s 0 16766 800 16826 0 FreeSans 480 0 0 0 rd_data[1]
port 26 nsew signal tristate
flabel metal3 s 0 49134 800 49194 0 FreeSans 480 0 0 0 rd_data[20]
port 27 nsew signal tristate
flabel metal3 s 0 50086 800 50146 0 FreeSans 480 0 0 0 rd_data[21]
port 28 nsew signal tristate
flabel metal3 s 0 51038 800 51098 0 FreeSans 480 0 0 0 rd_data[22]
port 29 nsew signal tristate
flabel metal3 s 0 51990 800 52050 0 FreeSans 480 0 0 0 rd_data[23]
port 30 nsew signal tristate
flabel metal3 s 0 52942 800 53002 0 FreeSans 480 0 0 0 rd_data[24]
port 31 nsew signal tristate
flabel metal3 s 0 53894 800 53954 0 FreeSans 480 0 0 0 rd_data[25]
port 32 nsew signal tristate
flabel metal3 s 0 54846 800 54906 0 FreeSans 480 0 0 0 rd_data[26]
port 33 nsew signal tristate
flabel metal3 s 0 55798 800 55858 0 FreeSans 480 0 0 0 rd_data[27]
port 34 nsew signal tristate
flabel metal3 s 0 56750 800 56810 0 FreeSans 480 0 0 0 rd_data[28]
port 35 nsew signal tristate
flabel metal3 s 0 57702 800 57762 0 FreeSans 480 0 0 0 rd_data[29]
port 36 nsew signal tristate
flabel metal3 s 0 15814 800 15874 0 FreeSans 480 0 0 0 rd_data[2]
port 37 nsew signal tristate
flabel metal3 s 0 58654 800 58714 0 FreeSans 480 0 0 0 rd_data[30]
port 38 nsew signal tristate
flabel metal3 s 0 59606 800 59666 0 FreeSans 480 0 0 0 rd_data[31]
port 39 nsew signal tristate
flabel metal3 s 0 14862 800 14922 0 FreeSans 480 0 0 0 rd_data[3]
port 40 nsew signal tristate
flabel metal3 s 0 13910 800 13970 0 FreeSans 480 0 0 0 rd_data[4]
port 41 nsew signal tristate
flabel metal3 s 0 12958 800 13018 0 FreeSans 480 0 0 0 rd_data[5]
port 42 nsew signal tristate
flabel metal3 s 0 12006 800 12066 0 FreeSans 480 0 0 0 rd_data[6]
port 43 nsew signal tristate
flabel metal3 s 0 11054 800 11114 0 FreeSans 480 0 0 0 rd_data[7]
port 44 nsew signal tristate
flabel metal3 s 0 10102 800 10162 0 FreeSans 480 0 0 0 rd_data[8]
port 45 nsew signal tristate
flabel metal3 s 0 9150 800 9210 0 FreeSans 480 0 0 0 rd_data[9]
port 46 nsew signal tristate
flabel metal4 s -416 -432 -96 88016 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal5 s -416 -432 110356 -112 0 FreeSans 2560 0 0 0 vccd1
port 47 nsew power bidirectional
flabel metal5 s -416 87696 110356 88016 0 FreeSans 2560 0 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 110036 -432 110356 88016 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 3604 -1092 3924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 5204 -1092 5524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 6804 -1092 7124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 8404 -1092 8724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 10004 -1092 10324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 10004 85496 10324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 11604 -1092 11924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 11604 85496 11924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 13204 -1092 13524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 13204 85496 13524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 14804 -1092 15124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 14804 85496 15124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 16404 -1092 16724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 16404 85496 16724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 18004 -1092 18324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 18004 85496 18324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 19604 -1092 19924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 19604 85496 19924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 21204 -1092 21524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 21204 85496 21524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 22804 -1092 23124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 22804 85496 23124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 24404 -1092 24724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 24404 85496 24724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 26004 -1092 26324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 26004 85496 26324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 27604 -1092 27924 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 27604 85496 27924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 29204 -1092 29524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 29204 85496 29524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 30804 -1092 31124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 30804 85496 31124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 32404 -1092 32724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 32404 85496 32724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 34004 -1092 34324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 34004 85496 34324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 35604 -1092 35924 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 35604 85496 35924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 37204 -1092 37524 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 37204 85496 37524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 38804 -1092 39124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 38804 85496 39124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 40404 -1092 40724 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 40404 85496 40724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 42004 -1092 42324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 42004 85496 42324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 43604 -1092 43924 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 43604 85620 43924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 45204 -1092 45524 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 45204 85620 45524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 46804 -1092 47124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 46804 85496 47124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 48404 -1092 48724 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 48404 85496 48724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 50004 -1092 50324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 50004 85620 50324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 51604 -1092 51924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 51604 85496 51924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 53204 -1092 53524 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 53204 85496 53524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 54804 -1092 55124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 54804 85496 55124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 56404 -1092 56724 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 56404 85620 56724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 58004 -1092 58324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 58004 85496 58324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 59604 -1092 59924 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 59604 85496 59924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 61204 -1092 61524 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 61204 85620 61524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 62804 -1092 63124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 62804 85496 63124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 64404 -1092 64724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 64404 85496 64724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 66004 -1092 66324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 66004 85620 66324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 67604 -1092 67924 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 67604 85620 67924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 69204 -1092 69524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 69204 85496 69524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 70804 -1092 71124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 70804 85496 71124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 72404 -1092 72724 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 72404 85620 72724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 74004 -1092 74324 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 74004 85620 74324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 75604 -1092 75924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 75604 85496 75924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 77204 -1092 77524 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 77204 85620 77524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 78804 -1092 79124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 78804 85620 79124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 80404 -1092 80724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 80404 85496 80724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 82004 -1092 82324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 82004 85496 82324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 83604 -1092 83924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 83604 85496 83924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 85204 -1092 85524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 85204 85496 85524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 86804 -1092 87124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 86804 85496 87124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 88404 -1092 88724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 88404 85496 88724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 90004 -1092 90324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 90004 85496 90324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 91604 -1092 91924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 91604 85620 91924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 93204 -1092 93524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 93204 85496 93524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 94804 -1092 95124 1880 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 94804 85496 95124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 96404 -1092 96724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 96404 85496 96724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 98004 -1092 98324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 98004 85496 98324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 99604 -1092 99924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 99604 85496 99924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 101204 -1092 101524 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 101204 85496 101524 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 102804 -1092 103124 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 102804 85496 103124 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 104404 -1092 104724 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 104404 85496 104724 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 106004 -1092 106324 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 106004 85496 106324 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 107604 -1092 107924 2004 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s 107604 85496 107924 88676 0 FreeSans 1920 90 0 0 vccd1
port 47 nsew power bidirectional
flabel metal5 s -1076 6588 111016 6908 0 FreeSans 2560 0 0 0 vccd1
port 47 nsew power bidirectional
flabel metal5 s -1076 82588 111016 82908 0 FreeSans 2560 0 0 0 vccd1
port 47 nsew power bidirectional
flabel metal4 s -1076 -1092 -756 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal5 s -1076 -1092 111016 -772 0 FreeSans 2560 0 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal5 s -1076 88356 111016 88676 0 FreeSans 2560 0 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 110696 -1092 111016 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 2944 -1092 3264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 4544 -1092 4864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 6144 -1092 6464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 7744 -1092 8064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 9344 -1092 9664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 10944 -1092 11264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 10944 85496 11264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 12544 -1092 12864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 12544 85496 12864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 14144 -1092 14464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 14144 85496 14464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 15744 -1092 16064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 15744 85496 16064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 17344 -1092 17664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 17344 85496 17664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 18944 -1092 19264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 18944 85496 19264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 20544 -1092 20864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 20544 85496 20864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 22144 -1092 22464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 22144 85496 22464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 23744 -1092 24064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 23744 85496 24064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 25344 -1092 25664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 25344 85496 25664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 26944 -1092 27264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 26944 85496 27264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 28544 -1092 28864 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 28544 85496 28864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 30144 -1092 30464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 30144 85496 30464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 31744 -1092 32064 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 31744 85496 32064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 33344 -1092 33664 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 33344 85496 33664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 34944 -1092 35264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 34944 85496 35264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 36544 -1092 36864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 36544 85496 36864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 38144 -1092 38464 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 38144 85496 38464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 39744 -1092 40064 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 39744 85620 40064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 41344 -1092 41664 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 41344 85620 41664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 42944 -1092 43264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 42944 85496 43264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 44544 -1092 44864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 44544 85496 44864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 46144 -1092 46464 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 46144 85620 46464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 47744 -1092 48064 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 47744 85620 48064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 49344 -1092 49664 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 49344 85496 49664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 50944 -1092 51264 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 50944 85620 51264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 52544 -1092 52864 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 52544 85620 52864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 54144 -1092 54464 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 54144 85496 54464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 55744 -1092 56064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 55744 85496 56064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 57344 -1092 57664 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 57344 85620 57664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 58944 -1092 59264 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 58944 85620 59264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 60544 -1092 60864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 60544 85496 60864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 62144 -1092 62464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 62144 85496 62464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 63744 -1092 64064 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 63744 85620 64064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 65344 -1092 65664 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 65344 85496 65664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 66944 -1092 67264 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 66944 85496 67264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 68544 -1092 68864 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 68544 85620 68864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 70144 -1092 70464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 70144 85620 70464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 71744 -1092 72064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 71744 85496 72064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 73344 -1092 73664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 73344 85496 73664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 74944 -1092 75264 1880 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 74944 85620 75264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 76544 -1092 76864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 76544 85496 76864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 78144 -1092 78464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 78144 85496 78464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 79744 -1092 80064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 79744 85496 80064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 81344 -1092 81664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 81344 85496 81664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 82944 -1092 83264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 82944 85496 83264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 84544 -1092 84864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 84544 85496 84864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 86144 -1092 86464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 86144 85496 86464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 87744 -1092 88064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 87744 85496 88064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 89344 -1092 89664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 89344 85496 89664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 90944 -1092 91264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 90944 85496 91264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 92544 -1092 92864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 92544 85496 92864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 94144 -1092 94464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 94144 85496 94464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 95744 -1092 96064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 95744 85496 96064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 97344 -1092 97664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 97344 85496 97664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 98944 -1092 99264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 98944 85496 99264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 100544 -1092 100864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 100544 85496 100864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 102144 -1092 102464 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 102144 85620 102464 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 103744 -1092 104064 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 103744 85496 104064 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 105344 -1092 105664 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 105344 85496 105664 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 106944 -1092 107264 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 106944 85496 107264 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 108544 -1092 108864 2004 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal4 s 108544 85496 108864 88676 0 FreeSans 1920 90 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal5 s -1076 5928 111016 6248 0 FreeSans 2560 0 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal5 s -1076 81928 111016 82248 0 FreeSans 2560 0 0 0 vssd1
port 48 nsew ground bidirectional
flabel metal3 s 0 62462 800 62522 0 FreeSans 480 0 0 0 wr_addr[0]
port 49 nsew signal input
flabel metal3 s 0 63414 800 63474 0 FreeSans 480 0 0 0 wr_addr[1]
port 50 nsew signal input
flabel metal3 s 0 64366 800 64426 0 FreeSans 480 0 0 0 wr_addr[2]
port 51 nsew signal input
flabel metal3 s 0 65318 800 65378 0 FreeSans 480 0 0 0 wr_addr[3]
port 52 nsew signal input
flabel metal3 s 0 66270 800 66330 0 FreeSans 480 0 0 0 wr_addr[4]
port 53 nsew signal input
flabel metal3 s 0 67222 800 67282 0 FreeSans 480 0 0 0 wr_addr[5]
port 54 nsew signal input
flabel metal3 s 0 68174 800 68234 0 FreeSans 480 0 0 0 wr_addr[6]
port 55 nsew signal input
flabel metal3 s 0 69126 800 69186 0 FreeSans 480 0 0 0 wr_addr[7]
port 56 nsew signal input
flabel metal3 s 0 37710 800 37770 0 FreeSans 480 0 0 0 wr_data[0]
port 57 nsew signal input
flabel metal3 s 0 28190 800 28250 0 FreeSans 480 0 0 0 wr_data[10]
port 58 nsew signal input
flabel metal3 s 0 29142 800 29202 0 FreeSans 480 0 0 0 wr_data[11]
port 59 nsew signal input
flabel metal3 s 0 30094 800 30154 0 FreeSans 480 0 0 0 wr_data[12]
port 60 nsew signal input
flabel metal3 s 0 31046 800 31106 0 FreeSans 480 0 0 0 wr_data[13]
port 61 nsew signal input
flabel metal3 s 0 43422 800 43482 0 FreeSans 480 0 0 0 wr_data[14]
port 62 nsew signal input
flabel metal3 s 0 44374 800 44434 0 FreeSans 480 0 0 0 wr_data[15]
port 63 nsew signal input
flabel metal3 s 0 70078 800 70138 0 FreeSans 480 0 0 0 wr_data[16]
port 64 nsew signal input
flabel metal3 s 0 71030 800 71090 0 FreeSans 480 0 0 0 wr_data[17]
port 65 nsew signal input
flabel metal3 s 0 71982 800 72042 0 FreeSans 480 0 0 0 wr_data[18]
port 66 nsew signal input
flabel metal3 s 0 72934 800 72994 0 FreeSans 480 0 0 0 wr_data[19]
port 67 nsew signal input
flabel metal3 s 0 38662 800 38722 0 FreeSans 480 0 0 0 wr_data[1]
port 68 nsew signal input
flabel metal3 s 0 73886 800 73946 0 FreeSans 480 0 0 0 wr_data[20]
port 69 nsew signal input
flabel metal3 s 0 74838 800 74898 0 FreeSans 480 0 0 0 wr_data[21]
port 70 nsew signal input
flabel metal3 s 0 75790 800 75850 0 FreeSans 480 0 0 0 wr_data[22]
port 71 nsew signal input
flabel metal3 s 0 76742 800 76802 0 FreeSans 480 0 0 0 wr_data[23]
port 72 nsew signal input
flabel metal3 s 0 77694 800 77754 0 FreeSans 480 0 0 0 wr_data[24]
port 73 nsew signal input
flabel metal3 s 0 78646 800 78706 0 FreeSans 480 0 0 0 wr_data[25]
port 74 nsew signal input
flabel metal3 s 0 79598 800 79658 0 FreeSans 480 0 0 0 wr_data[26]
port 75 nsew signal input
flabel metal3 s 0 80550 800 80610 0 FreeSans 480 0 0 0 wr_data[27]
port 76 nsew signal input
flabel metal3 s 0 81502 800 81562 0 FreeSans 480 0 0 0 wr_data[28]
port 77 nsew signal input
flabel metal3 s 0 82454 800 82514 0 FreeSans 480 0 0 0 wr_data[29]
port 78 nsew signal input
flabel metal3 s 0 39614 800 39674 0 FreeSans 480 0 0 0 wr_data[2]
port 79 nsew signal input
flabel metal3 s 0 83406 800 83466 0 FreeSans 480 0 0 0 wr_data[30]
port 80 nsew signal input
flabel metal3 s 0 84358 800 84418 0 FreeSans 480 0 0 0 wr_data[31]
port 81 nsew signal input
flabel metal3 s 0 40566 800 40626 0 FreeSans 480 0 0 0 wr_data[3]
port 82 nsew signal input
flabel metal3 s 0 41518 800 41578 0 FreeSans 480 0 0 0 wr_data[4]
port 83 nsew signal input
flabel metal3 s 0 42470 800 42530 0 FreeSans 480 0 0 0 wr_data[5]
port 84 nsew signal input
flabel metal3 s 0 31998 800 32058 0 FreeSans 480 0 0 0 wr_data[6]
port 85 nsew signal input
flabel metal3 s 0 32950 800 33010 0 FreeSans 480 0 0 0 wr_data[7]
port 86 nsew signal input
flabel metal3 s 0 33902 800 33962 0 FreeSans 480 0 0 0 wr_data[8]
port 87 nsew signal input
flabel metal3 s 0 34854 800 34914 0 FreeSans 480 0 0 0 wr_data[9]
port 88 nsew signal input
rlabel via4 106830 6748 106830 6748 0 vccd1
rlabel via4 107510 82088 107510 82088 0 vssd1
rlabel metal3 820 22508 820 22508 0 C0
rlabel metal3 820 23460 820 23460 0 C1
rlabel metal3 820 24412 820 24412 0 C2
rlabel metal3 820 25364 820 25364 0 C3
rlabel metal3 820 60588 820 60588 0 C4
rlabel metal3 820 61540 820 61540 0 C5
rlabel metal1 7774 11050 7774 11050 0 _000_
rlabel metal2 8096 13940 8096 13940 0 _001_
rlabel metal1 8372 16490 8372 16490 0 _002_
rlabel metal1 8878 11764 8878 11764 0 _003_
rlabel metal1 7590 11186 7590 11186 0 _004_
rlabel metal2 7590 55556 7590 55556 0 _005_
rlabel metal1 4968 58990 4968 58990 0 _006_
rlabel metal1 6670 67660 6670 67660 0 _007_
rlabel metal1 9246 67116 9246 67116 0 _008_
rlabel metal1 7498 57902 7498 57902 0 _009_
rlabel metal1 5520 44982 5520 44982 0 _010_
rlabel metal1 4186 57426 4186 57426 0 _011_
rlabel metal1 3772 64974 3772 64974 0 _012_
rlabel metal1 4692 66470 4692 66470 0 _013_
rlabel metal1 5106 66130 5106 66130 0 _014_
rlabel metal2 8786 64192 8786 64192 0 _015_
rlabel metal1 7590 66708 7590 66708 0 _016_
rlabel metal1 7452 69870 7452 69870 0 _017_
rlabel via1 7405 66606 7405 66606 0 _018_
rlabel metal2 8602 67405 8602 67405 0 _019_
rlabel metal1 7222 70516 7222 70516 0 _020_
rlabel metal1 4830 69870 4830 69870 0 _021_
rlabel metal1 6072 70006 6072 70006 0 _022_
rlabel metal2 9292 67558 9292 67558 0 _023_
rlabel metal2 9798 73134 9798 73134 0 _024_
rlabel metal1 6992 66674 6992 66674 0 _025_
rlabel metal1 4278 57562 4278 57562 0 _026_
rlabel metal1 6072 65042 6072 65042 0 _027_
rlabel metal1 11454 53720 11454 53720 0 _028_
rlabel metal1 7958 53108 7958 53108 0 _029_
rlabel metal2 9706 51187 9706 51187 0 _030_
rlabel metal2 4646 45152 4646 45152 0 _031_
rlabel metal1 8556 51374 8556 51374 0 _032_
rlabel metal1 5888 48722 5888 48722 0 _033_
rlabel metal1 5750 44846 5750 44846 0 _034_
rlabel metal2 1150 63172 1150 63172 0 _035_
rlabel metal1 4922 59398 4922 59398 0 _036_
rlabel metal1 6256 69938 6256 69938 0 _037_
rlabel metal1 7774 72250 7774 72250 0 _038_
rlabel metal1 7738 67728 7738 67728 0 _039_
rlabel metal1 8142 73202 8142 73202 0 _040_
rlabel via2 8418 72675 8418 72675 0 _041_
rlabel metal2 1288 59500 1288 59500 0 _042_
rlabel metal2 8326 70652 8326 70652 0 _043_
rlabel metal1 7498 54162 7498 54162 0 _044_
rlabel metal2 7682 53516 7682 53516 0 _045_
rlabel metal1 4882 44846 4882 44846 0 _046_
rlabel metal2 7222 59772 7222 59772 0 _047_
rlabel metal1 8188 54230 8188 54230 0 _048_
rlabel metal2 7038 72845 7038 72845 0 _049_
rlabel metal2 8970 71264 8970 71264 0 _050_
rlabel metal2 8050 73100 8050 73100 0 _051_
rlabel metal1 4922 45390 4922 45390 0 _052_
rlabel metal1 8234 53142 8234 53142 0 _053_
rlabel metal1 8970 51238 8970 51238 0 _054_
rlabel metal1 4922 45492 4922 45492 0 _055_
rlabel metal1 4554 64838 4554 64838 0 _056_
rlabel metal1 5244 58854 5244 58854 0 _057_
rlabel metal1 7590 73066 7590 73066 0 _058_
rlabel viali 6577 68782 6577 68782 0 _059_
rlabel metal2 8510 73219 8510 73219 0 _060_
rlabel metal1 4278 53074 4278 53074 0 _061_
rlabel metal1 5198 53006 5198 53006 0 _062_
rlabel metal1 5290 44404 5290 44404 0 _063_
rlabel metal1 6808 58514 6808 58514 0 _064_
rlabel metal1 2392 50966 2392 50966 0 _065_
rlabel metal1 7084 73542 7084 73542 0 _066_
rlabel metal2 5658 71774 5658 71774 0 _067_
rlabel metal1 6946 68340 6946 68340 0 _068_
rlabel metal2 1012 63036 1012 63036 0 _069_
rlabel metal2 6210 52666 6210 52666 0 _070_
rlabel metal2 6716 46342 6716 46342 0 _071_
rlabel metal1 8510 57426 8510 57426 0 _072_
rlabel metal1 7176 53074 7176 53074 0 _073_
rlabel metal1 8326 71536 8326 71536 0 _074_
rlabel metal1 6394 71638 6394 71638 0 _075_
rlabel metal1 8786 66130 8786 66130 0 _076_
rlabel metal1 7038 53142 7038 53142 0 _077_
rlabel metal1 8372 51374 8372 51374 0 _078_
rlabel metal1 5152 42670 5152 42670 0 _079_
rlabel metal1 7912 55726 7912 55726 0 _080_
rlabel metal1 2530 42296 2530 42296 0 _081_
rlabel metal1 7498 69734 7498 69734 0 _082_
rlabel metal2 7585 66198 7585 66198 0 _083_
rlabel metal1 7774 65076 7774 65076 0 _084_
rlabel metal1 6348 51374 6348 51374 0 _085_
rlabel metal1 8326 51272 8326 51272 0 _086_
rlabel metal1 6992 42670 6992 42670 0 _087_
rlabel metal1 9062 60214 9062 60214 0 _088_
rlabel metal1 3634 41718 3634 41718 0 _089_
rlabel metal1 9430 66674 9430 66674 0 _090_
rlabel metal1 8234 63308 8234 63308 0 _091_
rlabel metal1 8234 63444 8234 63444 0 _092_
rlabel metal2 2346 56338 2346 56338 0 _093_
rlabel metal1 4830 48722 4830 48722 0 _094_
rlabel metal1 4784 41582 4784 41582 0 _095_
rlabel metal1 10350 71502 10350 71502 0 _096_
rlabel metal2 20010 85918 20010 85918 0 _097_
rlabel metal2 9430 60044 9430 60044 0 _098_
rlabel metal1 8326 39814 8326 39814 0 _099_
rlabel metal1 6006 58547 6006 58547 0 _100_
rlabel metal1 4646 42330 4646 42330 0 _101_
rlabel metal2 2576 68204 2576 68204 0 _102_
rlabel metal2 9108 39100 9108 39100 0 _103_
rlabel metal2 598 71638 598 71638 0 _104_
rlabel metal1 7406 37774 7406 37774 0 _105_
rlabel metal1 6348 40358 6348 40358 0 _106_
rlabel metal2 17342 86666 17342 86666 0 _107_
rlabel metal1 6394 40154 6394 40154 0 _108_
rlabel metal1 9752 58514 9752 58514 0 _109_
rlabel metal1 9292 40086 9292 40086 0 _110_
rlabel metal1 10120 57902 10120 57902 0 _111_
rlabel metal1 6302 39270 6302 39270 0 _112_
rlabel metal1 5060 58106 5060 58106 0 _113_
rlabel metal1 4324 21998 4324 21998 0 _114_
rlabel metal1 7912 58446 7912 58446 0 _115_
rlabel metal1 6900 58310 6900 58310 0 _116_
rlabel metal1 5290 54162 5290 54162 0 _117_
rlabel metal1 5152 54230 5152 54230 0 _118_
rlabel metal1 9200 58650 9200 58650 0 _119_
rlabel metal1 6026 63206 6026 63206 0 _120_
rlabel metal1 6072 66062 6072 66062 0 _121_
rlabel metal1 5474 56814 5474 56814 0 _122_
rlabel metal2 5152 60588 5152 60588 0 _123_
rlabel metal1 7958 60282 7958 60282 0 _124_
rlabel metal2 4002 62798 4002 62798 0 _125_
rlabel metal2 5612 66266 5612 66266 0 _126_
rlabel metal2 25070 86054 25070 86054 0 _127_
rlabel metal1 17158 86258 17158 86258 0 _128_
rlabel metal1 13846 86360 13846 86360 0 _129_
rlabel metal2 37398 85102 37398 85102 0 _130_
rlabel metal2 4186 82333 4186 82333 0 _131_
rlabel via1 16974 86275 16974 86275 0 _132_
rlabel metal1 7498 58106 7498 58106 0 _133_
rlabel metal1 7682 17714 7682 17714 0 _134_
rlabel metal1 8832 19822 8832 19822 0 _135_
rlabel metal1 7544 27642 7544 27642 0 _136_
rlabel metal1 9062 20434 9062 20434 0 _137_
rlabel metal1 8510 22066 8510 22066 0 _138_
rlabel metal1 8372 23086 8372 23086 0 _139_
rlabel metal1 9108 23086 9108 23086 0 _140_
rlabel metal1 9246 24242 9246 24242 0 _141_
rlabel metal1 7268 31926 7268 31926 0 _142_
rlabel metal1 8602 25942 8602 25942 0 _143_
rlabel metal1 7498 18700 7498 18700 0 _144_
rlabel metal1 6578 25738 6578 25738 0 _145_
rlabel metal2 7728 21964 7728 21964 0 _146_
rlabel metal1 7912 14518 7912 14518 0 _147_
rlabel metal1 7360 18734 7360 18734 0 _148_
rlabel metal1 9039 986 9039 986 0 _149_
rlabel metal2 8694 33762 8694 33762 0 _150_
rlabel metal1 7590 36006 7590 36006 0 _151_
rlabel metal1 9568 14382 9568 14382 0 _152_
rlabel metal1 9614 16558 9614 16558 0 _153_
rlabel metal2 1058 16626 1058 16626 0 _154_
rlabel metal1 6440 15470 6440 15470 0 _155_
rlabel metal1 17250 1360 17250 1360 0 _156_
rlabel metal1 8694 33524 8694 33524 0 _157_
rlabel metal1 9798 37638 9798 37638 0 _158_
rlabel metal2 27554 2074 27554 2074 0 _159_
rlabel metal2 32154 2312 32154 2312 0 _160_
rlabel metal1 9292 33014 9292 33014 0 _161_
rlabel metal2 1150 17272 1150 17272 0 _162_
rlabel metal3 20194 3332 20194 3332 0 _163_
rlabel metal2 34730 2040 34730 2040 0 _164_
rlabel metal1 1104 35258 1104 35258 0 _165_
rlabel metal1 37536 1326 37536 1326 0 _166_
rlabel metal1 4508 39270 4508 39270 0 _167_
rlabel metal1 7406 25466 7406 25466 0 _168_
rlabel metal1 8004 18734 8004 18734 0 _169_
rlabel metal2 8326 17034 8326 17034 0 _170_
rlabel metal1 7544 17170 7544 17170 0 _171_
rlabel metal2 54970 823 54970 823 0 clk
rlabel metal1 17250 86156 17250 86156 0 clknet_0_clk
rlabel metal2 17894 3927 17894 3927 0 clknet_2_0__leaf_clk
rlabel metal2 6762 51646 6762 51646 0 clknet_2_1__leaf_clk
rlabel metal2 6394 57494 6394 57494 0 clknet_2_2__leaf_clk
rlabel metal4 102070 83702 102070 83702 0 clknet_2_3__leaf_clk
rlabel metal3 11761 11246 11761 11246 0 memWriteEnable
rlabel metal4 40190 83702 40190 83702 0 mem_dout\[0\]
rlabel metal4 52702 83702 52702 83702 0 mem_dout\[10\]
rlabel metal4 53926 83702 53926 83702 0 mem_dout\[11\]
rlabel metal4 55286 83702 55286 83702 0 mem_dout\[12\]
rlabel metal4 56374 83702 56374 83702 0 mem_dout\[13\]
rlabel metal4 57598 83702 57598 83702 0 mem_dout\[14\]
rlabel metal4 58958 83702 58958 83702 0 mem_dout\[15\]
rlabel metal4 60182 83566 60182 83566 0 mem_dout\[16\]
rlabel metal4 61542 83702 61542 83702 0 mem_dout\[17\]
rlabel metal4 62630 83702 62630 83702 0 mem_dout\[18\]
rlabel metal4 63990 83702 63990 83702 0 mem_dout\[19\]
rlabel metal1 9614 69530 9614 69530 0 mem_dout\[1\]
rlabel metal4 65078 83702 65078 83702 0 mem_dout\[20\]
rlabel metal4 66302 83702 66302 83702 0 mem_dout\[21\]
rlabel metal4 67662 83702 67662 83702 0 mem_dout\[22\]
rlabel metal4 68886 83702 68886 83702 0 mem_dout\[23\]
rlabel metal4 70246 83566 70246 83566 0 mem_dout\[24\]
rlabel metal4 71334 83702 71334 83702 0 mem_dout\[25\]
rlabel metal4 72694 83702 72694 83702 0 mem_dout\[26\]
rlabel metal4 73918 83702 73918 83702 0 mem_dout\[27\]
rlabel metal4 75278 83702 75278 83702 0 mem_dout\[28\]
rlabel metal4 76366 83702 76366 83702 0 mem_dout\[29\]
rlabel metal1 10120 68306 10120 68306 0 mem_dout\[2\]
rlabel metal4 77590 83702 77590 83702 0 mem_dout\[30\]
rlabel metal4 78950 83702 78950 83702 0 mem_dout\[31\]
rlabel via2 38870 86139 38870 86139 0 mem_dout\[3\]
rlabel metal2 11822 76500 11822 76500 0 mem_dout\[4\]
rlabel metal1 10350 67320 10350 67320 0 mem_dout\[5\]
rlabel metal2 36570 87312 36570 87312 0 mem_dout\[6\]
rlabel metal2 11730 74732 11730 74732 0 mem_dout\[7\]
rlabel metal2 11454 78744 11454 78744 0 mem_dout\[8\]
rlabel metal4 51342 83702 51342 83702 0 mem_dout\[9\]
rlabel metal2 28750 3553 28750 3553 0 mem_wr_mask\[0\]
rlabel metal2 29854 3621 29854 3621 0 mem_wr_mask\[1\]
rlabel metal4 31293 3740 31293 3740 0 mem_wr_mask\[2\]
rlabel metal2 32062 2465 32062 2465 0 mem_wr_mask\[3\]
rlabel metal2 45034 3757 45034 3757 0 muxedDataIn\[10\]
rlabel via2 46138 3859 46138 3859 0 muxedDataIn\[11\]
rlabel metal2 47518 3451 47518 3451 0 muxedDataIn\[12\]
rlabel metal2 48622 2261 48622 2261 0 muxedDataIn\[13\]
rlabel metal2 828 16560 828 16560 0 muxedDataIn\[14\]
rlabel metal2 50922 3791 50922 3791 0 muxedDataIn\[15\]
rlabel metal2 32246 663 32246 663 0 muxedDataIn\[16\]
rlabel metal4 53084 2312 53084 2312 0 muxedDataIn\[17\]
rlabel via2 54418 3893 54418 3893 0 muxedDataIn\[18\]
rlabel metal2 55430 2533 55430 2533 0 muxedDataIn\[19\]
rlabel metal2 56626 1071 56626 1071 0 muxedDataIn\[20\]
rlabel metal2 58006 2499 58006 2499 0 muxedDataIn\[21\]
rlabel metal2 58006 765 58006 765 0 muxedDataIn\[22\]
rlabel via2 59386 1275 59386 1275 0 muxedDataIn\[23\]
rlabel metal2 60950 1003 60950 1003 0 muxedDataIn\[24\]
rlabel metal2 62514 901 62514 901 0 muxedDataIn\[25\]
rlabel metal2 63526 833 63526 833 0 muxedDataIn\[26\]
rlabel metal4 64676 3060 64676 3060 0 muxedDataIn\[27\]
rlabel metal2 65182 1139 65182 1139 0 muxedDataIn\[28\]
rlabel metal2 37398 952 37398 952 0 muxedDataIn\[29\]
rlabel metal2 33902 1122 33902 1122 0 muxedDataIn\[30\]
rlabel metal2 37766 986 37766 986 0 muxedDataIn\[31\]
rlabel metal2 42826 2193 42826 2193 0 muxedDataIn\[8\]
rlabel metal2 43838 2431 43838 2431 0 muxedDataIn\[9\]
rlabel metal1 4922 24106 4922 24106 0 net1
rlabel metal3 57040 3604 57040 3604 0 net10
rlabel metal2 94990 2295 94990 2295 0 net11
rlabel metal4 94668 2856 94668 2856 0 net12
rlabel metal1 1472 36074 1472 36074 0 net13
rlabel metal1 2070 37162 2070 37162 0 net14
rlabel metal4 27525 3740 27525 3740 0 net15
rlabel metal2 1610 63648 1610 63648 0 net16
rlabel metal2 1610 64192 1610 64192 0 net17
rlabel metal2 2162 65263 2162 65263 0 net18
rlabel metal3 11945 34094 11945 34094 0 net19
rlabel viali 6023 25874 6023 25874 0 net2
rlabel metal2 1104 51060 1104 51060 0 net20
rlabel metal2 506 48907 506 48907 0 net21
rlabel via2 2162 69275 2162 69275 0 net22
rlabel metal1 2070 37638 2070 37638 0 net23
rlabel metal2 1426 28288 1426 28288 0 net24
rlabel metal1 6624 27098 6624 27098 0 net25
rlabel metal1 6348 26282 6348 26282 0 net26
rlabel metal2 7498 29818 7498 29818 0 net27
rlabel metal1 8556 32334 8556 32334 0 net28
rlabel metal2 2622 40947 2622 40947 0 net29
rlabel metal1 1242 24582 1242 24582 0 net3
rlabel metal1 1150 70618 1150 70618 0 net30
rlabel metal1 598 40460 598 40460 0 net31
rlabel metal3 1219 71876 1219 71876 0 net32
rlabel metal2 1380 57960 1380 57960 0 net33
rlabel metal2 2714 26044 2714 26044 0 net34
rlabel metal1 1794 74086 1794 74086 0 net35
rlabel metal1 2208 75242 2208 75242 0 net36
rlabel metal1 8096 38182 8096 38182 0 net37
rlabel metal1 2162 76874 2162 76874 0 net38
rlabel metal2 6670 36380 6670 36380 0 net39
rlabel metal1 2162 31178 2162 31178 0 net4
rlabel metal1 1426 78982 1426 78982 0 net40
rlabel metal1 1886 79594 1886 79594 0 net41
rlabel metal1 1794 80682 1794 80682 0 net42
rlabel metal1 1748 81770 1748 81770 0 net43
rlabel metal1 1978 82858 1978 82858 0 net44
rlabel metal1 2254 39814 2254 39814 0 net45
rlabel metal1 2852 83402 2852 83402 0 net46
rlabel metal1 1702 36176 1702 36176 0 net47
rlabel metal2 37030 2431 37030 2431 0 net48
rlabel metal2 37306 1241 37306 1241 0 net49
rlabel metal2 2806 60316 2806 60316 0 net5
rlabel metal2 39238 3723 39238 3723 0 net50
rlabel metal2 40342 3825 40342 3825 0 net51
rlabel metal4 41860 2108 41860 2108 0 net52
rlabel metal1 2484 33830 2484 33830 0 net53
rlabel metal1 2254 34918 2254 34918 0 net54
rlabel metal2 2622 20145 2622 20145 0 net55
rlabel metal1 1656 8534 1656 8534 0 net56
rlabel metal1 2438 7446 2438 7446 0 net57
rlabel metal1 1932 3502 1932 3502 0 net58
rlabel metal1 2898 4590 2898 4590 0 net59
rlabel metal1 8602 57834 8602 57834 0 net6
rlabel metal1 2760 5678 2760 5678 0 net60
rlabel metal1 1840 6766 1840 6766 0 net61
rlabel metal2 1610 51421 1610 51421 0 net62
rlabel metal1 2622 50898 2622 50898 0 net63
rlabel metal1 2116 47702 2116 47702 0 net64
rlabel metal1 3588 54502 3588 54502 0 net65
rlabel metal1 1794 17238 1794 17238 0 net66
rlabel metal2 2714 55667 2714 55667 0 net67
rlabel metal1 2438 50286 2438 50286 0 net68
rlabel metal2 1518 53788 1518 53788 0 net69
rlabel metal4 91462 83702 91462 83702 0 net7
rlabel metal2 4278 54808 4278 54808 0 net70
rlabel metal2 2806 56270 2806 56270 0 net71
rlabel metal2 1518 57868 1518 57868 0 net72
rlabel metal1 1978 55318 1978 55318 0 net73
rlabel metal1 2438 56406 2438 56406 0 net74
rlabel metal2 2438 68238 2438 68238 0 net75
rlabel metal1 2116 57902 2116 57902 0 net76
rlabel metal1 2944 16150 2944 16150 0 net77
rlabel metal3 5658 71468 5658 71468 0 net78
rlabel metal2 1518 59874 1518 59874 0 net79
rlabel metal3 56902 3468 56902 3468 0 net8
rlabel metal1 2990 15062 2990 15062 0 net80
rlabel metal1 2806 14382 2806 14382 0 net81
rlabel metal1 1702 13294 1702 13294 0 net82
rlabel metal1 1748 12206 1748 12206 0 net83
rlabel metal1 2024 11118 2024 11118 0 net84
rlabel metal1 1886 10710 1886 10710 0 net85
rlabel metal1 2852 9622 2852 9622 0 net86
rlabel metal3 108004 80470 108004 80470 0 net87
rlabel via2 107943 18428 107943 18428 0 net9
rlabel metal3 820 18700 820 18700 0 rd_addr[0]
rlabel metal3 820 19652 820 19652 0 rd_addr[1]
rlabel metal3 1050 20604 1050 20604 0 rd_addr[2]
rlabel metal3 820 21556 820 21556 0 rd_addr[3]
rlabel metal3 820 26316 820 26316 0 rd_addr[4]
rlabel metal3 820 27268 820 27268 0 rd_addr[5]
rlabel metal3 1050 35836 1050 35836 0 rd_addr[6]
rlabel metal3 866 36788 866 36788 0 rd_addr[7]
rlabel metal3 1142 17748 1142 17748 0 rd_data[0]
rlabel metal3 1050 8228 1050 8228 0 rd_data[10]
rlabel metal3 820 7276 820 7276 0 rd_data[11]
rlabel metal3 820 3468 820 3468 0 rd_data[12]
rlabel metal3 820 4420 820 4420 0 rd_data[13]
rlabel metal3 751 5372 751 5372 0 rd_data[14]
rlabel metal3 820 6324 820 6324 0 rd_data[15]
rlabel metal3 820 45356 820 45356 0 rd_data[16]
rlabel metal3 820 46308 820 46308 0 rd_data[17]
rlabel metal3 820 47260 820 47260 0 rd_data[18]
rlabel metal3 1142 48212 1142 48212 0 rd_data[19]
rlabel metal3 820 16796 820 16796 0 rd_data[1]
rlabel metal3 820 49164 820 49164 0 rd_data[20]
rlabel metal3 820 50116 820 50116 0 rd_data[21]
rlabel metal3 820 51068 820 51068 0 rd_data[22]
rlabel metal3 751 52020 751 52020 0 rd_data[23]
rlabel metal3 820 52972 820 52972 0 rd_data[24]
rlabel metal3 820 53924 820 53924 0 rd_data[25]
rlabel metal3 820 54876 820 54876 0 rd_data[26]
rlabel metal3 820 55828 820 55828 0 rd_data[27]
rlabel metal3 820 56780 820 56780 0 rd_data[28]
rlabel metal3 1142 57732 1142 57732 0 rd_data[29]
rlabel metal3 820 15844 820 15844 0 rd_data[2]
rlabel metal3 820 58684 820 58684 0 rd_data[30]
rlabel metal3 820 59636 820 59636 0 rd_data[31]
rlabel metal3 820 14892 820 14892 0 rd_data[3]
rlabel metal3 820 13940 820 13940 0 rd_data[4]
rlabel metal3 820 12988 820 12988 0 rd_data[5]
rlabel metal3 820 12036 820 12036 0 rd_data[6]
rlabel metal3 820 11084 820 11084 0 rd_data[7]
rlabel metal3 820 10132 820 10132 0 rd_data[8]
rlabel metal3 820 9180 820 9180 0 rd_data[9]
rlabel metal1 5842 46376 5842 46376 0 rd_dout_additional_register\[0\]
rlabel metal1 7682 44846 7682 44846 0 rd_dout_additional_register\[10\]
rlabel metal1 8188 40426 8188 40426 0 rd_dout_additional_register\[11\]
rlabel metal1 7268 40154 7268 40154 0 rd_dout_additional_register\[12\]
rlabel metal1 8602 43622 8602 43622 0 rd_dout_additional_register\[13\]
rlabel metal1 7314 39338 7314 39338 0 rd_dout_additional_register\[14\]
rlabel metal1 7268 37910 7268 37910 0 rd_dout_additional_register\[15\]
rlabel metal1 8280 58650 8280 58650 0 rd_dout_additional_register\[16\]
rlabel metal1 7222 62254 7222 62254 0 rd_dout_additional_register\[17\]
rlabel metal2 7682 61948 7682 61948 0 rd_dout_additional_register\[18\]
rlabel metal1 7774 62322 7774 62322 0 rd_dout_additional_register\[19\]
rlabel metal1 7268 47430 7268 47430 0 rd_dout_additional_register\[1\]
rlabel metal1 6854 63410 6854 63410 0 rd_dout_additional_register\[20\]
rlabel metal1 8418 63002 8418 63002 0 rd_dout_additional_register\[21\]
rlabel metal1 8280 61234 8280 61234 0 rd_dout_additional_register\[22\]
rlabel metal1 8234 60554 8234 60554 0 rd_dout_additional_register\[23\]
rlabel metal1 5842 66198 5842 66198 0 rd_dout_additional_register\[24\]
rlabel metal2 6854 69734 6854 69734 0 rd_dout_additional_register\[25\]
rlabel metal2 36478 85884 36478 85884 0 rd_dout_additional_register\[26\]
rlabel metal1 34040 86122 34040 86122 0 rd_dout_additional_register\[27\]
rlabel metal2 56718 85918 56718 85918 0 rd_dout_additional_register\[28\]
rlabel metal2 27554 86802 27554 86802 0 rd_dout_additional_register\[29\]
rlabel metal1 8234 49402 8234 49402 0 rd_dout_additional_register\[2\]
rlabel metal2 30406 86666 30406 86666 0 rd_dout_additional_register\[30\]
rlabel metal1 8234 57902 8234 57902 0 rd_dout_additional_register\[31\]
rlabel metal2 7498 46614 7498 46614 0 rd_dout_additional_register\[3\]
rlabel metal1 7406 52666 7406 52666 0 rd_dout_additional_register\[4\]
rlabel metal1 9062 46104 9062 46104 0 rd_dout_additional_register\[5\]
rlabel metal2 8326 47872 8326 47872 0 rd_dout_additional_register\[6\]
rlabel metal1 4232 43962 4232 43962 0 rd_dout_additional_register\[7\]
rlabel metal1 8188 39950 8188 39950 0 rd_dout_additional_register\[8\]
rlabel metal1 7176 42534 7176 42534 0 rd_dout_additional_register\[9\]
rlabel metal1 7171 51306 7171 51306 0 rd_dout_muxed\[0\]
rlabel metal1 9195 49130 9195 49130 0 rd_dout_muxed\[10\]
rlabel metal2 9108 57868 9108 57868 0 rd_dout_muxed\[11\]
rlabel metal1 9982 46512 9982 46512 0 rd_dout_muxed\[12\]
rlabel metal1 8045 43758 8045 43758 0 rd_dout_muxed\[13\]
rlabel metal1 8786 48518 8786 48518 0 rd_dout_muxed\[14\]
rlabel metal1 7130 37978 7130 37978 0 rd_dout_muxed\[15\]
rlabel metal1 7217 50966 7217 50966 0 rd_dout_muxed\[1\]
rlabel metal1 7309 52054 7309 52054 0 rd_dout_muxed\[2\]
rlabel metal1 7079 48110 7079 48110 0 rd_dout_muxed\[3\]
rlabel metal1 6936 52462 6936 52462 0 rd_dout_muxed\[4\]
rlabel metal1 7585 48790 7585 48790 0 rd_dout_muxed\[5\]
rlabel metal1 7539 49878 7539 49878 0 rd_dout_muxed\[6\]
rlabel metal1 4181 46954 4181 46954 0 rd_dout_muxed\[7\]
rlabel metal1 7820 40154 7820 40154 0 rd_dout_muxed\[8\]
rlabel metal1 6072 58310 6072 58310 0 rd_dout_muxed\[9\]
rlabel metal1 6716 57222 6716 57222 0 rd_dout_sel\[0\]
rlabel metal1 5566 59194 5566 59194 0 rd_dout_sel\[1\]
rlabel metal3 820 62492 820 62492 0 wr_addr[0]
rlabel metal3 1096 63444 1096 63444 0 wr_addr[1]
rlabel metal3 820 64396 820 64396 0 wr_addr[2]
rlabel metal3 820 65348 820 65348 0 wr_addr[3]
rlabel metal3 820 66300 820 66300 0 wr_addr[4]
rlabel metal3 751 67252 751 67252 0 wr_addr[5]
rlabel metal3 820 68204 820 68204 0 wr_addr[6]
rlabel metal3 820 69156 820 69156 0 wr_addr[7]
rlabel metal3 866 37740 866 37740 0 wr_data[0]
rlabel metal3 820 28220 820 28220 0 wr_data[10]
rlabel metal3 820 29172 820 29172 0 wr_data[11]
rlabel metal3 820 30124 820 30124 0 wr_data[12]
rlabel metal3 820 31076 820 31076 0 wr_data[13]
rlabel metal3 820 43452 820 43452 0 wr_data[14]
rlabel metal3 820 44404 820 44404 0 wr_data[15]
rlabel metal2 1426 70431 1426 70431 0 wr_data[16]
rlabel metal3 820 71060 820 71060 0 wr_data[17]
rlabel metal3 820 72012 820 72012 0 wr_data[18]
rlabel metal3 820 72964 820 72964 0 wr_data[19]
rlabel metal3 866 38692 866 38692 0 wr_data[1]
rlabel metal3 820 73916 820 73916 0 wr_data[20]
rlabel metal3 820 74868 820 74868 0 wr_data[21]
rlabel metal3 1096 75820 1096 75820 0 wr_data[22]
rlabel metal3 820 76772 820 76772 0 wr_data[23]
rlabel metal3 820 77724 820 77724 0 wr_data[24]
rlabel metal3 820 78676 820 78676 0 wr_data[25]
rlabel metal3 820 79628 820 79628 0 wr_data[26]
rlabel metal3 820 80580 820 80580 0 wr_data[27]
rlabel metal3 820 81532 820 81532 0 wr_data[28]
rlabel metal3 751 82484 751 82484 0 wr_data[29]
rlabel metal3 751 39644 751 39644 0 wr_data[2]
rlabel metal3 820 83436 820 83436 0 wr_data[30]
rlabel metal3 820 84388 820 84388 0 wr_data[31]
rlabel metal3 866 40596 866 40596 0 wr_data[3]
rlabel metal3 820 41548 820 41548 0 wr_data[4]
rlabel metal3 820 42500 820 42500 0 wr_data[5]
rlabel metal3 820 32028 820 32028 0 wr_data[6]
rlabel metal3 751 32980 751 32980 0 wr_data[7]
rlabel metal3 820 33932 820 33932 0 wr_data[8]
rlabel metal3 820 34884 820 34884 0 wr_data[9]
<< properties >>
string FIXED_BBOX 0 0 110000 88000
<< end >>
