magic
tech sky130A
magscale 1 2
timestamp 1734655017
<< viali >>
rect 1133 22729 1167 22763
rect 2053 22729 2087 22763
rect 3341 22729 3375 22763
rect 3893 22729 3927 22763
rect 4813 22729 4847 22763
rect 5917 22729 5951 22763
rect 6653 22729 6687 22763
rect 7573 22729 7607 22763
rect 8493 22729 8527 22763
rect 9413 22729 9447 22763
rect 10333 22729 10367 22763
rect 11253 22729 11287 22763
rect 12173 22729 12207 22763
rect 13093 22729 13127 22763
rect 13645 22729 13679 22763
rect 14013 22729 14047 22763
rect 14565 22729 14599 22763
rect 14933 22729 14967 22763
rect 15209 22729 15243 22763
rect 16221 22729 16255 22763
rect 16589 22729 16623 22763
rect 17693 22729 17727 22763
rect 18797 22729 18831 22763
rect 19349 22729 19383 22763
rect 20453 22729 20487 22763
rect 21373 22729 21407 22763
rect 21557 22729 21591 22763
rect 22293 22729 22327 22763
rect 23213 22729 23247 22763
rect 24133 22729 24167 22763
rect 24869 22729 24903 22763
rect 25421 22729 25455 22763
rect 25973 22729 26007 22763
rect 26893 22729 26927 22763
rect 27077 22729 27111 22763
rect 27905 22729 27939 22763
rect 29653 22729 29687 22763
rect 30573 22729 30607 22763
rect 31125 22729 31159 22763
rect 31493 22729 31527 22763
rect 33425 22729 33459 22763
rect 37013 22729 37047 22763
rect 37749 22729 37783 22763
rect 38485 22729 38519 22763
rect 40969 22729 41003 22763
rect 42809 22729 42843 22763
rect 29377 22661 29411 22695
rect 32413 22661 32447 22695
rect 949 22593 983 22627
rect 1869 22593 1903 22627
rect 3249 22593 3283 22627
rect 3709 22593 3743 22627
rect 4629 22593 4663 22627
rect 5825 22593 5859 22627
rect 6469 22593 6503 22627
rect 7389 22593 7423 22627
rect 8125 22593 8159 22627
rect 8401 22593 8435 22627
rect 9229 22593 9263 22627
rect 10149 22593 10183 22627
rect 11161 22593 11195 22627
rect 11989 22593 12023 22627
rect 12909 22593 12943 22627
rect 13921 22593 13955 22627
rect 14749 22593 14783 22627
rect 15393 22593 15427 22627
rect 15485 22593 15519 22627
rect 15669 22593 15703 22627
rect 16037 22593 16071 22627
rect 16497 22593 16531 22627
rect 17509 22593 17543 22627
rect 18613 22593 18647 22627
rect 19257 22593 19291 22627
rect 20269 22593 20303 22627
rect 21189 22593 21223 22627
rect 21749 22597 21783 22631
rect 22201 22593 22235 22627
rect 23029 22593 23063 22627
rect 23949 22593 23983 22627
rect 24777 22593 24811 22627
rect 25605 22593 25639 22627
rect 25789 22593 25823 22627
rect 26525 22593 26559 22627
rect 26709 22593 26743 22627
rect 27261 22593 27295 22627
rect 28457 22593 28491 22627
rect 29009 22593 29043 22627
rect 29561 22593 29595 22627
rect 30021 22593 30055 22627
rect 30481 22593 30515 22627
rect 30941 22593 30975 22627
rect 31861 22593 31895 22627
rect 33057 22593 33091 22627
rect 33333 22593 33367 22627
rect 33609 22593 33643 22627
rect 33885 22593 33919 22627
rect 34437 22593 34471 22627
rect 35081 22593 35115 22627
rect 35357 22593 35391 22627
rect 36001 22593 36035 22627
rect 36277 22593 36311 22627
rect 37657 22593 37691 22627
rect 37933 22593 37967 22627
rect 38393 22593 38427 22627
rect 39037 22593 39071 22627
rect 39405 22593 39439 22627
rect 39773 22593 39807 22627
rect 40693 22593 40727 22627
rect 41613 22593 41647 22627
rect 42533 22593 42567 22627
rect 43453 22593 43487 22627
rect 44557 22593 44591 22627
rect 45201 22593 45235 22627
rect 12817 22525 12851 22559
rect 27997 22525 28031 22559
rect 28089 22525 28123 22559
rect 31953 22525 31987 22559
rect 32137 22525 32171 22559
rect 34529 22525 34563 22559
rect 34621 22525 34655 22559
rect 37105 22525 37139 22559
rect 37197 22525 37231 22559
rect 38577 22525 38611 22559
rect 10057 22457 10091 22491
rect 20913 22457 20947 22491
rect 30205 22457 30239 22491
rect 32873 22457 32907 22491
rect 34897 22457 34931 22491
rect 40049 22457 40083 22491
rect 44833 22457 44867 22491
rect 7205 22389 7239 22423
rect 9137 22389 9171 22423
rect 11897 22389 11931 22423
rect 15853 22389 15887 22423
rect 17417 22389 17451 22423
rect 18429 22389 18463 22423
rect 20177 22389 20211 22423
rect 22845 22389 22879 22423
rect 24593 22389 24627 22423
rect 26341 22389 26375 22423
rect 27537 22389 27571 22423
rect 28641 22389 28675 22423
rect 32505 22389 32539 22423
rect 33149 22389 33183 22423
rect 33701 22389 33735 22423
rect 34069 22389 34103 22423
rect 35173 22389 35207 22423
rect 35725 22389 35759 22423
rect 35817 22389 35851 22423
rect 36093 22389 36127 22423
rect 36645 22389 36679 22423
rect 37473 22389 37507 22423
rect 38025 22389 38059 22423
rect 38853 22389 38887 22423
rect 39221 22389 39255 22423
rect 39589 22389 39623 22423
rect 40509 22389 40543 22423
rect 41429 22389 41463 22423
rect 42073 22389 42107 22423
rect 42349 22389 42383 22423
rect 43269 22389 43303 22423
rect 43821 22389 43855 22423
rect 44189 22389 44223 22423
rect 44373 22389 44407 22423
rect 45017 22389 45051 22423
rect 1409 22185 1443 22219
rect 2053 22185 2087 22219
rect 2789 22185 2823 22219
rect 3893 22185 3927 22219
rect 4629 22185 4663 22219
rect 5457 22185 5491 22219
rect 6009 22185 6043 22219
rect 6469 22185 6503 22219
rect 7297 22185 7331 22219
rect 8309 22185 8343 22219
rect 9413 22185 9447 22219
rect 10149 22185 10183 22219
rect 10885 22185 10919 22219
rect 11805 22185 11839 22219
rect 12817 22185 12851 22219
rect 13553 22185 13587 22219
rect 14105 22185 14139 22219
rect 16773 22185 16807 22219
rect 17233 22185 17267 22219
rect 17785 22185 17819 22219
rect 18245 22185 18279 22219
rect 19717 22185 19751 22219
rect 19993 22185 20027 22219
rect 22109 22185 22143 22219
rect 22753 22185 22787 22219
rect 23121 22185 23155 22219
rect 24961 22185 24995 22219
rect 29377 22185 29411 22219
rect 31020 22185 31054 22219
rect 36264 22185 36298 22219
rect 40969 22185 41003 22219
rect 41705 22185 41739 22219
rect 42441 22185 42475 22219
rect 32505 22117 32539 22151
rect 40141 22117 40175 22151
rect 9321 22049 9355 22083
rect 12357 22049 12391 22083
rect 20269 22049 20303 22083
rect 24777 22049 24811 22083
rect 27813 22049 27847 22083
rect 28549 22049 28583 22083
rect 30021 22049 30055 22083
rect 33149 22049 33183 22083
rect 34069 22049 34103 22083
rect 36001 22049 36035 22083
rect 38393 22049 38427 22083
rect 39773 22049 39807 22083
rect 44557 22049 44591 22083
rect 1593 21981 1627 22015
rect 1961 21981 1995 22015
rect 2237 21981 2271 22015
rect 2973 21981 3007 22015
rect 3341 21981 3375 22015
rect 4077 21981 4111 22015
rect 4445 21981 4479 22015
rect 4813 21981 4847 22015
rect 5089 21981 5123 22015
rect 5641 21981 5675 22015
rect 6653 21981 6687 22015
rect 7481 21981 7515 22015
rect 8493 21981 8527 22015
rect 9597 21981 9631 22015
rect 10333 21981 10367 22015
rect 11069 21981 11103 22015
rect 11989 21981 12023 22015
rect 13001 21981 13035 22015
rect 13737 21981 13771 22015
rect 14289 21981 14323 22015
rect 14381 21981 14415 22015
rect 14749 21981 14783 22015
rect 16175 21981 16209 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 16957 21981 16991 22015
rect 17417 21981 17451 22015
rect 18429 21981 18463 22015
rect 18613 21981 18647 22015
rect 18981 21981 19015 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 19901 21981 19935 22015
rect 20177 21981 20211 22015
rect 22293 21981 22327 22015
rect 22937 21981 22971 22015
rect 23305 21981 23339 22015
rect 23581 21981 23615 22015
rect 24041 21981 24075 22015
rect 25145 21981 25179 22015
rect 25329 21981 25363 22015
rect 27537 21981 27571 22015
rect 28917 21981 28951 22015
rect 29745 21981 29779 22015
rect 30205 21981 30239 22015
rect 30757 21981 30791 22015
rect 33609 21981 33643 22015
rect 33885 21981 33919 22015
rect 38209 21981 38243 22015
rect 39589 21981 39623 22015
rect 40325 21981 40359 22015
rect 44925 21981 44959 22015
rect 2605 21913 2639 21947
rect 10793 21913 10827 21947
rect 18797 21913 18831 21947
rect 18889 21913 18923 21947
rect 20545 21913 20579 21947
rect 24501 21913 24535 21947
rect 25605 21913 25639 21947
rect 28365 21913 28399 21947
rect 29837 21913 29871 21947
rect 32965 21913 32999 21947
rect 34345 21913 34379 21947
rect 43177 21913 43211 21947
rect 6377 21845 6411 21879
rect 7205 21845 7239 21879
rect 8033 21845 8067 21879
rect 8953 21845 8987 21879
rect 10057 21845 10091 21879
rect 11713 21845 11747 21879
rect 12725 21845 12759 21879
rect 16681 21845 16715 21879
rect 18153 21845 18187 21879
rect 19165 21845 19199 21879
rect 19349 21845 19383 21879
rect 22017 21845 22051 21879
rect 22661 21845 22695 21879
rect 23397 21845 23431 21879
rect 23857 21845 23891 21879
rect 24133 21845 24167 21879
rect 24593 21845 24627 21879
rect 27077 21845 27111 21879
rect 27169 21845 27203 21879
rect 27629 21845 27663 21879
rect 27997 21845 28031 21879
rect 28457 21845 28491 21879
rect 29101 21845 29135 21879
rect 30389 21845 30423 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 33701 21845 33735 21879
rect 35817 21845 35851 21879
rect 37749 21845 37783 21879
rect 37841 21845 37875 21879
rect 38301 21845 38335 21879
rect 38853 21845 38887 21879
rect 39221 21845 39255 21879
rect 39681 21845 39715 21879
rect 40601 21845 40635 21879
rect 41337 21845 41371 21879
rect 42165 21845 42199 21879
rect 42809 21845 42843 21879
rect 43545 21845 43579 21879
rect 43913 21845 43947 21879
rect 12265 21641 12299 21675
rect 16037 21641 16071 21675
rect 19441 21641 19475 21675
rect 19625 21641 19659 21675
rect 20361 21641 20395 21675
rect 21373 21641 21407 21675
rect 25421 21641 25455 21675
rect 25789 21641 25823 21675
rect 25881 21641 25915 21675
rect 28365 21641 28399 21675
rect 29561 21641 29595 21675
rect 30389 21641 30423 21675
rect 35173 21641 35207 21675
rect 36001 21641 36035 21675
rect 36277 21641 36311 21675
rect 40693 21641 40727 21675
rect 41337 21641 41371 21675
rect 41981 21641 42015 21675
rect 42349 21641 42383 21675
rect 43085 21641 43119 21675
rect 44189 21641 44223 21675
rect 44557 21641 44591 21675
rect 11161 21573 11195 21607
rect 16313 21573 16347 21607
rect 16405 21573 16439 21607
rect 16523 21573 16557 21607
rect 17141 21573 17175 21607
rect 17969 21573 18003 21607
rect 19993 21573 20027 21607
rect 26617 21573 26651 21607
rect 29101 21573 29135 21607
rect 36921 21573 36955 21607
rect 38761 21573 38795 21607
rect 42717 21573 42751 21607
rect 43821 21573 43855 21607
rect 13737 21505 13771 21539
rect 13829 21505 13863 21539
rect 15623 21505 15657 21539
rect 16221 21505 16255 21539
rect 16681 21505 16715 21539
rect 16957 21505 16991 21539
rect 17233 21505 17267 21539
rect 17325 21505 17359 21539
rect 17509 21505 17543 21539
rect 17693 21505 17727 21539
rect 19809 21505 19843 21539
rect 19901 21505 19935 21539
rect 20111 21505 20145 21539
rect 20545 21505 20579 21539
rect 20637 21505 20671 21539
rect 21189 21505 21223 21539
rect 21465 21505 21499 21539
rect 21741 21505 21775 21539
rect 26341 21505 26375 21539
rect 28181 21505 28215 21539
rect 29193 21505 29227 21539
rect 29929 21505 29963 21539
rect 30021 21505 30055 21539
rect 30757 21505 30791 21539
rect 30849 21505 30883 21539
rect 35541 21505 35575 21539
rect 36185 21505 36219 21539
rect 36461 21505 36495 21539
rect 6101 21437 6135 21471
rect 10149 21437 10183 21471
rect 14197 21437 14231 21471
rect 16773 21437 16807 21471
rect 20269 21437 20303 21471
rect 20913 21437 20947 21471
rect 21005 21437 21039 21471
rect 22017 21437 22051 21471
rect 23581 21437 23615 21471
rect 25329 21437 25363 21471
rect 26065 21437 26099 21471
rect 29285 21437 29319 21471
rect 30113 21437 30147 21471
rect 30941 21437 30975 21471
rect 31493 21437 31527 21471
rect 31769 21437 31803 21471
rect 33333 21437 33367 21471
rect 33609 21437 33643 21471
rect 35633 21437 35667 21471
rect 35725 21437 35759 21471
rect 36645 21437 36679 21471
rect 38485 21437 38519 21471
rect 40785 21437 40819 21471
rect 40877 21437 40911 21471
rect 7849 21369 7883 21403
rect 8217 21369 8251 21403
rect 8677 21369 8711 21403
rect 9321 21369 9355 21403
rect 11529 21369 11563 21403
rect 11897 21369 11931 21403
rect 17417 21369 17451 21403
rect 21189 21369 21223 21403
rect 23489 21369 23523 21403
rect 28733 21369 28767 21403
rect 40233 21369 40267 21403
rect 40325 21369 40359 21403
rect 6377 21301 6411 21335
rect 6837 21301 6871 21335
rect 7113 21301 7147 21335
rect 7481 21301 7515 21335
rect 9045 21301 9079 21335
rect 9781 21301 9815 21335
rect 10517 21301 10551 21335
rect 12633 21301 12667 21335
rect 13001 21301 13035 21335
rect 13369 21301 13403 21335
rect 23844 21301 23878 21335
rect 28089 21301 28123 21335
rect 33241 21301 33275 21335
rect 35081 21301 35115 21335
rect 38393 21301 38427 21335
rect 43453 21301 43487 21335
rect 44925 21301 44959 21335
rect 13737 21097 13771 21131
rect 14473 21097 14507 21131
rect 19349 21097 19383 21131
rect 23213 21097 23247 21131
rect 25513 21097 25547 21131
rect 26525 21097 26559 21131
rect 30757 21097 30791 21131
rect 32597 21097 32631 21131
rect 32873 21097 32907 21131
rect 35817 21097 35851 21131
rect 37749 21097 37783 21131
rect 40969 21097 41003 21131
rect 42901 21097 42935 21131
rect 44557 21097 44591 21131
rect 12541 21029 12575 21063
rect 18613 21029 18647 21063
rect 22845 21029 22879 21063
rect 27353 21029 27387 21063
rect 30665 21029 30699 21063
rect 37657 21029 37691 21063
rect 41061 21029 41095 21063
rect 8125 20961 8159 20995
rect 9229 20961 9263 20995
rect 15117 20961 15151 20995
rect 16681 20961 16715 20995
rect 16957 20961 16991 20995
rect 19165 20961 19199 20995
rect 19625 20961 19659 20995
rect 19809 20961 19843 20995
rect 20453 20961 20487 20995
rect 22385 20961 22419 20995
rect 24041 20961 24075 20995
rect 26341 20961 26375 20995
rect 26985 20961 27019 20995
rect 27169 20961 27203 20995
rect 27905 20961 27939 20995
rect 31401 20961 31435 20995
rect 32321 20961 32355 20995
rect 33609 20961 33643 20995
rect 33793 20961 33827 20995
rect 35909 20961 35943 20995
rect 36185 20961 36219 20995
rect 38209 20961 38243 20995
rect 38393 20961 38427 20995
rect 41521 20961 41555 20995
rect 41613 20961 41647 20995
rect 42441 20961 42475 20995
rect 949 20893 983 20927
rect 6377 20893 6411 20927
rect 8953 20893 8987 20927
rect 11069 20893 11103 20927
rect 11437 20893 11471 20927
rect 11805 20893 11839 20927
rect 12173 20893 12207 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 14841 20893 14875 20927
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 19533 20893 19567 20927
rect 19717 20893 19751 20927
rect 19993 20893 20027 20927
rect 22477 20893 22511 20927
rect 22937 20893 22971 20927
rect 23121 20893 23155 20927
rect 23397 20893 23431 20927
rect 23765 20893 23799 20927
rect 26065 20893 26099 20927
rect 26893 20893 26927 20927
rect 27721 20893 27755 20927
rect 28181 20893 28215 20927
rect 28549 20893 28583 20927
rect 28917 20893 28951 20927
rect 31125 20893 31159 20927
rect 32781 20893 32815 20927
rect 33057 20893 33091 20927
rect 34069 20893 34103 20927
rect 38761 20893 38795 20927
rect 39037 20893 39071 20927
rect 39221 20893 39255 20927
rect 42257 20893 42291 20927
rect 6193 20825 6227 20859
rect 6653 20825 6687 20859
rect 12909 20825 12943 20859
rect 13277 20825 13311 20859
rect 14105 20825 14139 20859
rect 19257 20825 19291 20859
rect 20177 20825 20211 20859
rect 20729 20825 20763 20859
rect 26157 20825 26191 20859
rect 28365 20825 28399 20859
rect 28457 20825 28491 20859
rect 29193 20825 29227 20859
rect 32137 20825 32171 20859
rect 32229 20825 32263 20859
rect 34345 20825 34379 20859
rect 39497 20825 39531 20859
rect 43361 20825 43395 20859
rect 44833 20825 44867 20859
rect 45201 20825 45235 20859
rect 765 20757 799 20791
rect 3709 20757 3743 20791
rect 5549 20757 5583 20791
rect 5917 20757 5951 20791
rect 8861 20757 8895 20791
rect 10701 20757 10735 20791
rect 14749 20757 14783 20791
rect 16589 20757 16623 20791
rect 18429 20757 18463 20791
rect 20361 20757 20395 20791
rect 22201 20757 22235 20791
rect 23029 20757 23063 20791
rect 25697 20757 25731 20791
rect 27813 20757 27847 20791
rect 28733 20757 28767 20791
rect 31217 20757 31251 20791
rect 31769 20757 31803 20791
rect 33149 20757 33183 20791
rect 33517 20757 33551 20791
rect 38117 20757 38151 20791
rect 38577 20757 38611 20791
rect 38853 20757 38887 20791
rect 41429 20757 41463 20791
rect 41889 20757 41923 20791
rect 42349 20757 42383 20791
rect 43637 20757 43671 20791
rect 44005 20757 44039 20791
rect 3617 20553 3651 20587
rect 5549 20553 5583 20587
rect 9229 20553 9263 20587
rect 9597 20553 9631 20587
rect 9965 20553 9999 20587
rect 11805 20553 11839 20587
rect 12541 20553 12575 20587
rect 13553 20553 13587 20587
rect 13921 20553 13955 20587
rect 16037 20553 16071 20587
rect 17141 20553 17175 20587
rect 17693 20553 17727 20587
rect 19533 20553 19567 20587
rect 20269 20553 20303 20587
rect 20453 20553 20487 20587
rect 22753 20553 22787 20587
rect 23489 20553 23523 20587
rect 23949 20553 23983 20587
rect 25605 20553 25639 20587
rect 29929 20553 29963 20587
rect 32045 20553 32079 20587
rect 33425 20553 33459 20587
rect 33701 20553 33735 20587
rect 34069 20553 34103 20587
rect 34161 20553 34195 20587
rect 34897 20553 34931 20587
rect 35725 20553 35759 20587
rect 36645 20553 36679 20587
rect 37105 20553 37139 20587
rect 39313 20553 39347 20587
rect 41429 20553 41463 20587
rect 42257 20553 42291 20587
rect 2145 20485 2179 20519
rect 4077 20485 4111 20519
rect 13277 20485 13311 20519
rect 14105 20485 14139 20519
rect 14473 20485 14507 20519
rect 15209 20485 15243 20519
rect 15301 20485 15335 20519
rect 15761 20485 15795 20519
rect 18889 20485 18923 20519
rect 21189 20485 21223 20519
rect 21557 20485 21591 20519
rect 22385 20485 22419 20519
rect 28457 20485 28491 20519
rect 31769 20485 31803 20519
rect 32965 20485 32999 20519
rect 34989 20485 35023 20519
rect 36093 20485 36127 20519
rect 37013 20485 37047 20519
rect 37841 20485 37875 20519
rect 39957 20485 39991 20519
rect 43085 20485 43119 20519
rect 43453 20485 43487 20519
rect 44557 20485 44591 20519
rect 44925 20485 44959 20519
rect 14703 20451 14737 20485
rect 14289 20417 14323 20451
rect 14381 20417 14415 20451
rect 15117 20417 15151 20451
rect 15439 20417 15473 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 16221 20417 16255 20451
rect 16313 20417 16347 20451
rect 16405 20417 16439 20451
rect 16523 20417 16557 20451
rect 16681 20417 16715 20451
rect 16773 20417 16807 20451
rect 17233 20417 17267 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 17601 20417 17635 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 18153 20417 18187 20451
rect 18245 20417 18279 20451
rect 18429 20417 18463 20451
rect 18521 20417 18555 20451
rect 18647 20417 18681 20451
rect 19165 20417 19199 20451
rect 19625 20417 19659 20451
rect 20183 20417 20217 20451
rect 20361 20417 20395 20451
rect 21373 20417 21407 20451
rect 21925 20417 21959 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22293 20417 22327 20451
rect 22569 20417 22603 20451
rect 23857 20417 23891 20451
rect 24777 20417 24811 20451
rect 25145 20417 25179 20451
rect 25789 20417 25823 20451
rect 26157 20417 26191 20451
rect 30205 20417 30239 20451
rect 30665 20417 30699 20451
rect 30757 20417 30791 20451
rect 31493 20417 31527 20451
rect 31677 20417 31711 20451
rect 31861 20417 31895 20451
rect 32137 20417 32171 20451
rect 33057 20417 33091 20451
rect 33609 20417 33643 20451
rect 36185 20417 36219 20451
rect 42165 20417 42199 20451
rect 42809 20417 42843 20451
rect 1869 20349 1903 20383
rect 3801 20349 3835 20383
rect 8033 20349 8067 20383
rect 15577 20349 15611 20383
rect 19257 20349 19291 20383
rect 19717 20349 19751 20383
rect 20637 20349 20671 20383
rect 20729 20349 20763 20383
rect 20821 20349 20855 20383
rect 20913 20349 20947 20383
rect 24133 20349 24167 20383
rect 26341 20349 26375 20383
rect 26617 20349 26651 20383
rect 28181 20349 28215 20383
rect 30941 20349 30975 20383
rect 33149 20349 33183 20383
rect 34253 20349 34287 20383
rect 35081 20349 35115 20383
rect 36369 20349 36403 20383
rect 37197 20349 37231 20383
rect 37565 20349 37599 20383
rect 39681 20349 39715 20383
rect 42349 20349 42383 20383
rect 6009 20281 6043 20315
rect 14105 20281 14139 20315
rect 14933 20281 14967 20315
rect 16911 20281 16945 20315
rect 17325 20281 17359 20315
rect 25973 20281 26007 20315
rect 30021 20281 30055 20315
rect 32321 20281 32355 20315
rect 32597 20281 32631 20315
rect 34529 20281 34563 20315
rect 43821 20281 43855 20315
rect 6285 20213 6319 20247
rect 6929 20213 6963 20247
rect 7297 20213 7331 20247
rect 7665 20213 7699 20247
rect 8401 20213 8435 20247
rect 8769 20213 8803 20247
rect 10241 20213 10275 20247
rect 10609 20213 10643 20247
rect 11345 20213 11379 20247
rect 12173 20213 12207 20247
rect 12909 20213 12943 20247
rect 14657 20213 14691 20247
rect 14841 20213 14875 20247
rect 17049 20213 17083 20247
rect 19809 20213 19843 20247
rect 19993 20213 20027 20247
rect 21649 20213 21683 20247
rect 23397 20213 23431 20247
rect 24593 20213 24627 20247
rect 24961 20213 24995 20247
rect 25329 20213 25363 20247
rect 28089 20213 28123 20247
rect 30297 20213 30331 20247
rect 35633 20213 35667 20247
rect 41797 20213 41831 20247
rect 42625 20213 42659 20247
rect 44281 20213 44315 20247
rect 3985 20009 4019 20043
rect 6929 20009 6963 20043
rect 7665 20009 7699 20043
rect 8769 20009 8803 20043
rect 9229 20009 9263 20043
rect 17693 20009 17727 20043
rect 18705 20009 18739 20043
rect 19717 20009 19751 20043
rect 21373 20009 21407 20043
rect 23765 20009 23799 20043
rect 27997 20009 28031 20043
rect 34253 20009 34287 20043
rect 36185 20009 36219 20043
rect 36645 20009 36679 20043
rect 44557 20009 44591 20043
rect 44925 20009 44959 20043
rect 12541 19941 12575 19975
rect 12817 19941 12851 19975
rect 14197 19941 14231 19975
rect 21557 19941 21591 19975
rect 23213 19941 23247 19975
rect 28641 19941 28675 19975
rect 30665 19941 30699 19975
rect 31309 19941 31343 19975
rect 32689 19941 32723 19975
rect 39405 19941 39439 19975
rect 5457 19873 5491 19907
rect 11621 19873 11655 19907
rect 13829 19873 13863 19907
rect 14749 19873 14783 19907
rect 15117 19873 15151 19907
rect 15485 19873 15519 19907
rect 17509 19873 17543 19907
rect 18061 19873 18095 19907
rect 19073 19873 19107 19907
rect 20637 19873 20671 19907
rect 20821 19873 20855 19907
rect 24317 19873 24351 19907
rect 25421 19873 25455 19907
rect 25973 19873 26007 19907
rect 26249 19873 26283 19907
rect 28917 19873 28951 19907
rect 29193 19873 29227 19907
rect 32137 19873 32171 19907
rect 33333 19873 33367 19907
rect 35725 19873 35759 19907
rect 37105 19873 37139 19907
rect 37197 19873 37231 19907
rect 38025 19873 38059 19907
rect 40141 19873 40175 19907
rect 42257 19873 42291 19907
rect 42533 19873 42567 19907
rect 9321 19805 9355 19839
rect 9505 19805 9539 19839
rect 9689 19805 9723 19839
rect 11713 19805 11747 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 14841 19805 14875 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 18153 19805 18187 19839
rect 18245 19805 18279 19839
rect 18429 19805 18463 19839
rect 18613 19805 18647 19839
rect 19349 19805 19383 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20269 19805 20303 19839
rect 20361 19805 20395 19839
rect 20729 19805 20763 19839
rect 20913 19805 20947 19839
rect 21557 19805 21591 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 21925 19805 21959 19839
rect 22109 19805 22143 19839
rect 24225 19805 24259 19839
rect 25329 19805 25363 19839
rect 28089 19805 28123 19839
rect 28457 19805 28491 19839
rect 30777 19805 30811 19839
rect 31029 19805 31063 19839
rect 31125 19805 31159 19839
rect 32321 19805 32355 19839
rect 33057 19805 33091 19839
rect 34897 19805 34931 19839
rect 35541 19805 35575 19839
rect 37013 19805 37047 19839
rect 37841 19805 37875 19839
rect 38485 19805 38519 19839
rect 38761 19805 38795 19839
rect 40049 19805 40083 19839
rect 40417 19805 40451 19839
rect 7297 19737 7331 19771
rect 9965 19737 9999 19771
rect 17233 19737 17267 19771
rect 19165 19737 19199 19771
rect 20085 19737 20119 19771
rect 23581 19737 23615 19771
rect 25237 19737 25271 19771
rect 26525 19737 26559 19771
rect 28273 19737 28307 19771
rect 28365 19737 28399 19771
rect 30941 19737 30975 19771
rect 31861 19737 31895 19771
rect 34161 19737 34195 19771
rect 40693 19737 40727 19771
rect 4721 19669 4755 19703
rect 5089 19669 5123 19703
rect 5825 19669 5859 19703
rect 6193 19669 6227 19703
rect 6653 19669 6687 19703
rect 8125 19669 8159 19703
rect 9413 19669 9447 19703
rect 11437 19669 11471 19703
rect 12081 19669 12115 19703
rect 13185 19669 13219 19703
rect 14381 19669 14415 19703
rect 16911 19669 16945 19703
rect 17877 19669 17911 19703
rect 18429 19669 18463 19703
rect 19533 19669 19567 19703
rect 20453 19669 20487 19703
rect 22017 19669 22051 19703
rect 22385 19669 22419 19703
rect 22845 19669 22879 19703
rect 24133 19669 24167 19703
rect 24869 19669 24903 19703
rect 31493 19669 31527 19703
rect 31953 19669 31987 19703
rect 32505 19669 32539 19703
rect 33149 19669 33183 19703
rect 33793 19669 33827 19703
rect 34713 19669 34747 19703
rect 35173 19669 35207 19703
rect 35633 19669 35667 19703
rect 37473 19669 37507 19703
rect 37933 19669 37967 19703
rect 38301 19669 38335 19703
rect 39589 19669 39623 19703
rect 39957 19669 39991 19703
rect 42165 19669 42199 19703
rect 44005 19669 44039 19703
rect 7757 19465 7791 19499
rect 8401 19465 8435 19499
rect 10333 19465 10367 19499
rect 12633 19465 12667 19499
rect 14841 19465 14875 19499
rect 18981 19465 19015 19499
rect 19165 19465 19199 19499
rect 21649 19465 21683 19499
rect 24593 19465 24627 19499
rect 25605 19465 25639 19499
rect 27905 19465 27939 19499
rect 28917 19465 28951 19499
rect 31677 19465 31711 19499
rect 33609 19465 33643 19499
rect 34529 19465 34563 19499
rect 41337 19465 41371 19499
rect 41797 19465 41831 19499
rect 42165 19465 42199 19499
rect 42257 19465 42291 19499
rect 43085 19465 43119 19499
rect 8861 19397 8895 19431
rect 15485 19397 15519 19431
rect 19901 19397 19935 19431
rect 21189 19397 21223 19431
rect 29653 19397 29687 19431
rect 30205 19397 30239 19431
rect 30297 19397 30331 19431
rect 37565 19397 37599 19431
rect 42993 19397 43027 19431
rect 44097 19397 44131 19431
rect 7021 19329 7055 19363
rect 7389 19329 7423 19363
rect 7573 19329 7607 19363
rect 7757 19329 7791 19363
rect 8125 19329 8159 19363
rect 8585 19329 8619 19363
rect 10425 19329 10459 19363
rect 10609 19329 10643 19363
rect 13185 19329 13219 19363
rect 15302 19329 15336 19363
rect 15669 19329 15703 19363
rect 15761 19329 15795 19363
rect 16037 19329 16071 19363
rect 16313 19329 16347 19363
rect 16681 19329 16715 19363
rect 16957 19329 16991 19363
rect 17509 19329 17543 19363
rect 17969 19329 18003 19363
rect 18245 19329 18279 19363
rect 18613 19329 18647 19363
rect 18797 19329 18831 19363
rect 19073 19329 19107 19363
rect 19257 19329 19291 19363
rect 19809 19329 19843 19363
rect 19993 19329 20027 19363
rect 20085 19329 20119 19363
rect 20269 19329 20303 19363
rect 20361 19329 20395 19363
rect 21481 19329 21515 19363
rect 25145 19329 25179 19363
rect 25789 19329 25823 19363
rect 27353 19329 27387 19363
rect 27537 19329 27571 19363
rect 27629 19329 27663 19363
rect 27721 19329 27755 19363
rect 28089 19329 28123 19363
rect 28733 19329 28767 19363
rect 29377 19329 29411 19363
rect 29561 19329 29595 19363
rect 29745 19329 29779 19363
rect 30021 19329 30055 19363
rect 30413 19329 30447 19363
rect 31493 19329 31527 19363
rect 33977 19329 34011 19363
rect 34897 19329 34931 19363
rect 34989 19329 35023 19363
rect 35725 19329 35759 19363
rect 36369 19329 36403 19363
rect 37197 19353 37231 19387
rect 41245 19329 41279 19363
rect 41521 19329 41555 19363
rect 6745 19261 6779 19295
rect 10885 19261 10919 19295
rect 12817 19261 12851 19295
rect 15025 19261 15059 19295
rect 15118 19261 15152 19295
rect 15209 19261 15243 19295
rect 16405 19261 16439 19295
rect 17693 19261 17727 19295
rect 20821 19261 20855 19295
rect 21373 19261 21407 19295
rect 22845 19261 22879 19295
rect 23121 19261 23155 19295
rect 25237 19261 25271 19295
rect 25329 19261 25363 19295
rect 30941 19261 30975 19295
rect 31033 19261 31067 19295
rect 31125 19261 31159 19295
rect 31217 19261 31251 19295
rect 31861 19261 31895 19295
rect 32137 19261 32171 19295
rect 33701 19261 33735 19295
rect 33885 19261 33919 19295
rect 34069 19261 34103 19295
rect 34161 19261 34195 19295
rect 35173 19261 35207 19295
rect 35817 19261 35851 19295
rect 35909 19261 35943 19295
rect 37289 19261 37323 19295
rect 39228 19261 39262 19295
rect 39497 19261 39531 19295
rect 42349 19261 42383 19295
rect 43177 19261 43211 19295
rect 44741 19261 44775 19295
rect 15485 19193 15519 19227
rect 16865 19193 16899 19227
rect 18061 19193 18095 19227
rect 19625 19193 19659 19227
rect 41061 19193 41095 19227
rect 42625 19193 42659 19227
rect 43637 19193 43671 19227
rect 44373 19193 44407 19227
rect 45109 19193 45143 19227
rect 5549 19125 5583 19159
rect 6009 19125 6043 19159
rect 6285 19125 6319 19159
rect 10517 19125 10551 19159
rect 11148 19125 11182 19159
rect 14611 19125 14645 19159
rect 18797 19125 18831 19159
rect 20637 19125 20671 19159
rect 21189 19125 21223 19159
rect 21925 19125 21959 19159
rect 22293 19125 22327 19159
rect 22753 19125 22787 19159
rect 24777 19125 24811 19159
rect 26157 19125 26191 19159
rect 26617 19125 26651 19159
rect 26893 19125 26927 19159
rect 28365 19125 28399 19159
rect 29929 19125 29963 19159
rect 30573 19125 30607 19159
rect 30757 19125 30791 19159
rect 35357 19125 35391 19159
rect 36185 19125 36219 19159
rect 36921 19125 36955 19159
rect 37013 19125 37047 19159
rect 39037 19125 39071 19159
rect 40969 19125 41003 19159
rect 5457 18921 5491 18955
rect 6469 18921 6503 18955
rect 8033 18921 8067 18955
rect 8750 18921 8784 18955
rect 10425 18921 10459 18955
rect 10977 18921 11011 18955
rect 13185 18921 13219 18955
rect 16681 18921 16715 18955
rect 18613 18921 18647 18955
rect 22845 18921 22879 18955
rect 23765 18921 23799 18955
rect 28181 18921 28215 18955
rect 29469 18921 29503 18955
rect 32229 18921 32263 18955
rect 38117 18921 38151 18955
rect 40969 18921 41003 18955
rect 41061 18921 41095 18955
rect 6009 18853 6043 18887
rect 18245 18853 18279 18887
rect 19901 18853 19935 18887
rect 28641 18853 28675 18887
rect 29193 18853 29227 18887
rect 32965 18853 32999 18887
rect 4445 18785 4479 18819
rect 7113 18785 7147 18819
rect 7665 18785 7699 18819
rect 10241 18785 10275 18819
rect 13461 18785 13495 18819
rect 13829 18785 13863 18819
rect 15761 18785 15795 18819
rect 19165 18785 19199 18819
rect 19441 18785 19475 18819
rect 20637 18785 20671 18819
rect 23489 18785 23523 18819
rect 24317 18785 24351 18819
rect 26709 18785 26743 18819
rect 30021 18785 30055 18819
rect 30481 18785 30515 18819
rect 32505 18785 32539 18819
rect 32597 18785 32631 18819
rect 33425 18785 33459 18819
rect 33517 18785 33551 18819
rect 34713 18785 34747 18819
rect 36553 18785 36587 18819
rect 38669 18785 38703 18819
rect 39221 18785 39255 18819
rect 41613 18785 41647 18819
rect 42441 18785 42475 18819
rect 4537 18717 4571 18751
rect 5549 18717 5583 18751
rect 5733 18717 5767 18751
rect 6561 18717 6595 18751
rect 6745 18717 6779 18751
rect 7021 18717 7055 18751
rect 7757 18717 7791 18751
rect 8493 18717 8527 18751
rect 10333 18717 10367 18751
rect 10517 18717 10551 18751
rect 10609 18717 10643 18751
rect 10793 18717 10827 18751
rect 11069 18717 11103 18751
rect 13093 18717 13127 18751
rect 15393 18717 15427 18751
rect 15878 18717 15912 18751
rect 16129 18717 16163 18751
rect 16313 18717 16347 18751
rect 16497 18717 16531 18751
rect 17049 18717 17083 18751
rect 17417 18717 17451 18751
rect 17969 18717 18003 18751
rect 18613 18717 18647 18751
rect 18797 18717 18831 18751
rect 19073 18717 19107 18751
rect 19257 18717 19291 18751
rect 19533 18717 19567 18751
rect 19993 18717 20027 18751
rect 20269 18717 20303 18751
rect 20361 18717 20395 18751
rect 22753 18717 22787 18751
rect 24133 18717 24167 18751
rect 24593 18717 24627 18751
rect 26433 18717 26467 18751
rect 28273 18717 28307 18751
rect 28457 18717 28491 18751
rect 29837 18717 29871 18751
rect 29929 18717 29963 18751
rect 32689 18717 32723 18751
rect 32781 18717 32815 18751
rect 34069 18717 34103 18751
rect 34437 18717 34471 18751
rect 36277 18717 36311 18751
rect 38485 18717 38519 18751
rect 38577 18717 38611 18751
rect 41429 18717 41463 18751
rect 41521 18717 41555 18751
rect 42901 18717 42935 18751
rect 11345 18649 11379 18683
rect 16405 18649 16439 18683
rect 20177 18649 20211 18683
rect 20913 18649 20947 18683
rect 23305 18649 23339 18683
rect 24869 18649 24903 18683
rect 30757 18649 30791 18683
rect 33333 18649 33367 18683
rect 39497 18649 39531 18683
rect 42349 18649 42383 18683
rect 4905 18581 4939 18615
rect 5641 18581 5675 18615
rect 6745 18581 6779 18615
rect 7389 18581 7423 18615
rect 12817 18581 12851 18615
rect 15255 18581 15289 18615
rect 15669 18581 15703 18615
rect 16037 18581 16071 18615
rect 20545 18581 20579 18615
rect 22385 18581 22419 18615
rect 22569 18581 22603 18615
rect 23213 18581 23247 18615
rect 24225 18581 24259 18615
rect 26341 18581 26375 18615
rect 32321 18581 32355 18615
rect 34253 18581 34287 18615
rect 36185 18581 36219 18615
rect 38025 18581 38059 18615
rect 41889 18581 41923 18615
rect 42257 18581 42291 18615
rect 42717 18581 42751 18615
rect 43269 18581 43303 18615
rect 43545 18581 43579 18615
rect 43913 18581 43947 18615
rect 44557 18581 44591 18615
rect 44925 18581 44959 18615
rect 5549 18377 5583 18411
rect 6101 18377 6135 18411
rect 8493 18377 8527 18411
rect 12449 18377 12483 18411
rect 13001 18377 13035 18411
rect 13553 18377 13587 18411
rect 17699 18377 17733 18411
rect 17785 18377 17819 18411
rect 21833 18377 21867 18411
rect 22477 18377 22511 18411
rect 24685 18377 24719 18411
rect 25513 18377 25547 18411
rect 28273 18377 28307 18411
rect 31493 18377 31527 18411
rect 34069 18377 34103 18411
rect 34529 18377 34563 18411
rect 36461 18377 36495 18411
rect 38761 18377 38795 18411
rect 39221 18377 39255 18411
rect 40049 18377 40083 18411
rect 41245 18377 41279 18411
rect 43545 18377 43579 18411
rect 44189 18377 44223 18411
rect 44925 18377 44959 18411
rect 4077 18309 4111 18343
rect 6285 18309 6319 18343
rect 7021 18309 7055 18343
rect 8861 18309 8895 18343
rect 11805 18309 11839 18343
rect 16221 18309 16255 18343
rect 16773 18309 16807 18343
rect 17141 18309 17175 18343
rect 17341 18309 17375 18343
rect 20545 18309 20579 18343
rect 21281 18309 21315 18343
rect 23121 18309 23155 18343
rect 27353 18309 27387 18343
rect 28825 18309 28859 18343
rect 29377 18309 29411 18343
rect 30941 18309 30975 18343
rect 31157 18309 31191 18343
rect 32597 18309 32631 18343
rect 34161 18309 34195 18343
rect 34361 18309 34395 18343
rect 37197 18309 37231 18343
rect 39129 18309 39163 18343
rect 42073 18309 42107 18343
rect 3801 18241 3835 18275
rect 5733 18241 5767 18275
rect 6193 18241 6227 18275
rect 6469 18241 6503 18275
rect 8585 18241 8619 18275
rect 11529 18241 11563 18275
rect 11897 18241 11931 18275
rect 12081 18241 12115 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 13737 18241 13771 18275
rect 13829 18241 13863 18275
rect 14197 18241 14231 18275
rect 16037 18241 16071 18275
rect 16313 18241 16347 18275
rect 16405 18241 16439 18275
rect 16680 18263 16714 18297
rect 16907 18241 16941 18275
rect 17049 18241 17083 18275
rect 17601 18241 17635 18275
rect 17877 18241 17911 18275
rect 17969 18241 18003 18275
rect 18153 18241 18187 18275
rect 20361 18241 20395 18275
rect 20453 18241 20487 18275
rect 20663 18241 20697 18275
rect 21189 18241 21223 18275
rect 21373 18241 21407 18275
rect 21465 18241 21499 18275
rect 21640 18241 21674 18275
rect 21765 18241 21799 18275
rect 21925 18241 21959 18275
rect 22753 18241 22787 18275
rect 22845 18241 22879 18275
rect 25053 18241 25087 18275
rect 25145 18241 25179 18275
rect 25697 18241 25731 18275
rect 26617 18241 26651 18275
rect 26893 18241 26927 18275
rect 28181 18241 28215 18275
rect 28641 18241 28675 18275
rect 29101 18241 29135 18275
rect 31677 18241 31711 18275
rect 31769 18241 31803 18275
rect 31861 18241 31895 18275
rect 34713 18241 34747 18275
rect 39957 18241 39991 18275
rect 40785 18241 40819 18275
rect 6745 18173 6779 18207
rect 10609 18173 10643 18207
rect 11805 18173 11839 18207
rect 18337 18173 18371 18207
rect 18613 18173 18647 18207
rect 20177 18173 20211 18207
rect 20821 18173 20855 18207
rect 24593 18173 24627 18207
rect 25237 18173 25271 18207
rect 27445 18173 27479 18207
rect 27629 18173 27663 18207
rect 28365 18173 28399 18207
rect 30849 18173 30883 18207
rect 31953 18173 31987 18207
rect 32321 18173 32355 18207
rect 34989 18173 35023 18207
rect 36921 18173 36955 18207
rect 39313 18173 39347 18207
rect 40141 18173 40175 18207
rect 41337 18173 41371 18207
rect 41429 18173 41463 18207
rect 41797 18173 41831 18207
rect 43821 18173 43855 18207
rect 44557 18173 44591 18207
rect 12265 18105 12299 18139
rect 16589 18105 16623 18139
rect 17049 18105 17083 18139
rect 18061 18105 18095 18139
rect 20085 18105 20119 18139
rect 22569 18105 22603 18139
rect 26065 18105 26099 18139
rect 26985 18105 27019 18139
rect 27813 18105 27847 18139
rect 31309 18105 31343 18139
rect 38669 18105 38703 18139
rect 40877 18105 40911 18139
rect 5871 18037 5905 18071
rect 6009 18037 6043 18071
rect 6653 18037 6687 18071
rect 10333 18037 10367 18071
rect 11345 18037 11379 18071
rect 11621 18037 11655 18071
rect 12081 18037 12115 18071
rect 13461 18037 13495 18071
rect 15623 18037 15657 18071
rect 17325 18037 17359 18071
rect 17509 18037 17543 18071
rect 21557 18037 21591 18071
rect 26433 18037 26467 18071
rect 26709 18037 26743 18071
rect 29009 18037 29043 18071
rect 31125 18037 31159 18071
rect 34345 18037 34379 18071
rect 39589 18037 39623 18071
rect 40601 18037 40635 18071
rect 3893 17833 3927 17867
rect 4445 17833 4479 17867
rect 8401 17833 8435 17867
rect 9321 17833 9355 17867
rect 9597 17833 9631 17867
rect 9873 17833 9907 17867
rect 10793 17833 10827 17867
rect 13185 17833 13219 17867
rect 15393 17833 15427 17867
rect 17049 17833 17083 17867
rect 17877 17833 17911 17867
rect 19073 17833 19107 17867
rect 20085 17833 20119 17867
rect 20821 17833 20855 17867
rect 22017 17833 22051 17867
rect 22845 17833 22879 17867
rect 28273 17833 28307 17867
rect 30665 17833 30699 17867
rect 31033 17833 31067 17867
rect 31217 17833 31251 17867
rect 33701 17833 33735 17867
rect 35081 17833 35115 17867
rect 35725 17833 35759 17867
rect 37105 17833 37139 17867
rect 37657 17833 37691 17867
rect 38393 17833 38427 17867
rect 40325 17833 40359 17867
rect 42441 17833 42475 17867
rect 8769 17765 8803 17799
rect 9229 17765 9263 17799
rect 15255 17765 15289 17799
rect 19257 17765 19291 17799
rect 20729 17765 20763 17799
rect 23765 17765 23799 17799
rect 28733 17765 28767 17799
rect 4813 17697 4847 17731
rect 8125 17697 8159 17731
rect 8493 17697 8527 17731
rect 9413 17697 9447 17731
rect 11437 17697 11471 17731
rect 12173 17697 12207 17731
rect 12541 17697 12575 17731
rect 13829 17697 13863 17731
rect 15853 17697 15887 17731
rect 16037 17697 16071 17731
rect 16497 17697 16531 17731
rect 17049 17697 17083 17731
rect 18981 17697 19015 17731
rect 20269 17697 20303 17731
rect 23305 17697 23339 17731
rect 23397 17697 23431 17731
rect 24317 17697 24351 17731
rect 25053 17697 25087 17731
rect 28917 17697 28951 17731
rect 29193 17697 29227 17731
rect 31493 17697 31527 17731
rect 31585 17697 31619 17731
rect 32229 17697 32263 17731
rect 34713 17697 34747 17731
rect 36369 17697 36403 17731
rect 38025 17697 38059 17731
rect 39773 17697 39807 17731
rect 40693 17697 40727 17731
rect 42993 17697 43027 17731
rect 43085 17697 43119 17731
rect 3525 17629 3559 17663
rect 3709 17629 3743 17663
rect 3801 17629 3835 17663
rect 3985 17629 4019 17663
rect 4537 17629 4571 17663
rect 6377 17629 6411 17663
rect 8585 17629 8619 17663
rect 9137 17629 9171 17663
rect 9505 17629 9539 17663
rect 9597 17629 9631 17663
rect 11253 17629 11287 17663
rect 12449 17629 12483 17663
rect 13461 17629 13495 17663
rect 16313 17629 16347 17663
rect 16405 17629 16439 17663
rect 16681 17629 16715 17663
rect 17141 17629 17175 17663
rect 17417 17629 17451 17663
rect 17785 17629 17819 17663
rect 18337 17629 18371 17663
rect 19073 17629 19107 17663
rect 19441 17629 19475 17663
rect 19625 17629 19659 17663
rect 19809 17629 19843 17663
rect 20085 17629 20119 17663
rect 20361 17629 20395 17663
rect 21005 17629 21039 17663
rect 21281 17629 21315 17663
rect 22753 17629 22787 17663
rect 24961 17629 24995 17663
rect 26893 17629 26927 17663
rect 27149 17629 27183 17663
rect 28365 17629 28399 17663
rect 31677 17629 31711 17663
rect 31769 17629 31803 17663
rect 31942 17629 31976 17663
rect 34989 17629 35023 17663
rect 35265 17629 35299 17663
rect 36093 17629 36127 17663
rect 36185 17629 36219 17663
rect 37841 17629 37875 17663
rect 38577 17629 38611 17663
rect 38853 17629 38887 17663
rect 42901 17629 42935 17663
rect 31079 17595 31113 17629
rect 4077 17561 4111 17595
rect 4261 17561 4295 17595
rect 6653 17561 6687 17595
rect 8309 17561 8343 17595
rect 10333 17561 10367 17595
rect 15761 17561 15795 17595
rect 16865 17561 16899 17595
rect 18613 17561 18647 17595
rect 19993 17561 20027 17595
rect 24225 17561 24259 17595
rect 25329 17561 25363 17595
rect 28549 17561 28583 17595
rect 30849 17561 30883 17595
rect 34345 17561 34379 17595
rect 37381 17561 37415 17595
rect 39589 17561 39623 17595
rect 40233 17561 40267 17595
rect 40969 17561 41003 17595
rect 3433 17493 3467 17527
rect 3709 17493 3743 17527
rect 6285 17493 6319 17527
rect 10885 17493 10919 17527
rect 11345 17493 11379 17527
rect 12817 17493 12851 17527
rect 16589 17493 16623 17527
rect 17325 17493 17359 17527
rect 17601 17493 17635 17527
rect 19533 17493 19567 17527
rect 21189 17493 21223 17527
rect 21649 17493 21683 17527
rect 22385 17493 22419 17527
rect 22569 17493 22603 17527
rect 23213 17493 23247 17527
rect 24133 17493 24167 17527
rect 24777 17493 24811 17527
rect 26801 17493 26835 17527
rect 31309 17493 31343 17527
rect 34805 17493 34839 17527
rect 35633 17493 35667 17527
rect 36737 17493 36771 17527
rect 38669 17493 38703 17527
rect 39221 17493 39255 17527
rect 39681 17493 39715 17527
rect 42533 17493 42567 17527
rect 43545 17493 43579 17527
rect 43913 17493 43947 17527
rect 44557 17493 44591 17527
rect 44925 17493 44959 17527
rect 5549 17289 5583 17323
rect 6193 17289 6227 17323
rect 7021 17289 7055 17323
rect 7665 17289 7699 17323
rect 8125 17289 8159 17323
rect 9781 17289 9815 17323
rect 9873 17289 9907 17323
rect 14473 17289 14507 17323
rect 15051 17289 15085 17323
rect 15761 17289 15795 17323
rect 16589 17289 16623 17323
rect 20453 17289 20487 17323
rect 20637 17289 20671 17323
rect 22385 17289 22419 17323
rect 24317 17289 24351 17323
rect 25053 17289 25087 17323
rect 25421 17289 25455 17323
rect 27905 17289 27939 17323
rect 29469 17289 29503 17323
rect 31309 17289 31343 17323
rect 31861 17289 31895 17323
rect 32889 17289 32923 17323
rect 33793 17289 33827 17323
rect 41245 17289 41279 17323
rect 42809 17289 42843 17323
rect 43913 17289 43947 17323
rect 44281 17289 44315 17323
rect 45017 17289 45051 17323
rect 3709 17221 3743 17255
rect 11161 17221 11195 17255
rect 13001 17221 13035 17255
rect 14841 17221 14875 17255
rect 18705 17221 18739 17255
rect 19073 17221 19107 17255
rect 19165 17221 19199 17255
rect 19809 17221 19843 17255
rect 22845 17221 22879 17255
rect 25513 17221 25547 17255
rect 26770 17221 26804 17255
rect 30941 17221 30975 17255
rect 31141 17221 31175 17255
rect 31585 17221 31619 17255
rect 32229 17221 32263 17255
rect 32689 17221 32723 17255
rect 34713 17221 34747 17255
rect 38209 17221 38243 17255
rect 40049 17221 40083 17255
rect 5733 17153 5767 17187
rect 6009 17153 6043 17187
rect 6929 17153 6963 17187
rect 7113 17153 7147 17187
rect 7389 17153 7423 17187
rect 9045 17153 9079 17187
rect 10057 17153 10091 17187
rect 10333 17153 10367 17187
rect 10701 17153 10735 17187
rect 10885 17153 10919 17187
rect 15301 17153 15335 17187
rect 15583 17153 15617 17187
rect 16405 17153 16439 17187
rect 16865 17153 16899 17187
rect 17049 17153 17083 17187
rect 17141 17153 17175 17187
rect 17233 17153 17267 17187
rect 17509 17153 17543 17187
rect 17693 17153 17727 17187
rect 18337 17153 18371 17187
rect 18521 17153 18555 17187
rect 18981 17153 19015 17187
rect 19283 17153 19317 17187
rect 19717 17153 19751 17187
rect 19902 17153 19936 17187
rect 20039 17153 20073 17187
rect 20269 17153 20303 17187
rect 20361 17153 20395 17187
rect 22569 17153 22603 17187
rect 24409 17153 24443 17187
rect 24961 17153 24995 17187
rect 27997 17153 28031 17187
rect 28264 17153 28298 17187
rect 29699 17153 29733 17187
rect 29837 17153 29871 17187
rect 29934 17153 29968 17187
rect 30113 17153 30147 17187
rect 30481 17153 30515 17187
rect 30573 17153 30607 17187
rect 30665 17153 30699 17187
rect 30849 17153 30883 17187
rect 31769 17153 31803 17187
rect 34161 17153 34195 17187
rect 34437 17153 34471 17187
rect 36829 17153 36863 17187
rect 37933 17153 37967 17187
rect 39957 17153 39991 17187
rect 40141 17153 40175 17187
rect 40785 17153 40819 17187
rect 41337 17153 41371 17187
rect 42165 17153 42199 17187
rect 42257 17153 42291 17187
rect 3801 17085 3835 17119
rect 4077 17085 4111 17119
rect 5825 17085 5859 17119
rect 7481 17085 7515 17119
rect 7665 17085 7699 17119
rect 9137 17085 9171 17119
rect 9321 17085 9355 17119
rect 12725 17085 12759 17119
rect 16313 17085 16347 17119
rect 16681 17085 16715 17119
rect 16773 17085 16807 17119
rect 19441 17085 19475 17119
rect 20177 17085 20211 17119
rect 20637 17085 20671 17119
rect 25605 17085 25639 17119
rect 26157 17085 26191 17119
rect 26525 17085 26559 17119
rect 32321 17085 32355 17119
rect 32505 17085 32539 17119
rect 41429 17085 41463 17119
rect 42349 17085 42383 17119
rect 15209 17017 15243 17051
rect 17509 17017 17543 17051
rect 18797 17017 18831 17051
rect 20913 17017 20947 17051
rect 22017 17017 22051 17051
rect 30205 17017 30239 17051
rect 33057 17017 33091 17051
rect 39773 17017 39807 17051
rect 40877 17017 40911 17051
rect 5733 16949 5767 16983
rect 6837 16949 6871 16983
rect 8493 16949 8527 16983
rect 8677 16949 8711 16983
rect 10149 16949 10183 16983
rect 10517 16949 10551 16983
rect 12633 16949 12667 16983
rect 15025 16949 15059 16983
rect 15393 16949 15427 16983
rect 16129 16949 16163 16983
rect 17417 16949 17451 16983
rect 18245 16949 18279 16983
rect 19533 16949 19567 16983
rect 21741 16949 21775 16983
rect 24593 16949 24627 16983
rect 24777 16949 24811 16983
rect 29377 16949 29411 16983
rect 31125 16949 31159 16983
rect 32873 16949 32907 16983
rect 33425 16949 33459 16983
rect 36185 16949 36219 16983
rect 36645 16949 36679 16983
rect 37197 16949 37231 16983
rect 37473 16949 37507 16983
rect 39681 16949 39715 16983
rect 40325 16949 40359 16983
rect 40601 16949 40635 16983
rect 41797 16949 41831 16983
rect 43177 16949 43211 16983
rect 43545 16949 43579 16983
rect 44649 16949 44683 16983
rect 7389 16745 7423 16779
rect 12357 16745 12391 16779
rect 14105 16745 14139 16779
rect 16405 16745 16439 16779
rect 20361 16745 20395 16779
rect 21189 16745 21223 16779
rect 24593 16745 24627 16779
rect 28549 16745 28583 16779
rect 30113 16745 30147 16779
rect 32597 16745 32631 16779
rect 35909 16745 35943 16779
rect 36737 16745 36771 16779
rect 37749 16745 37783 16779
rect 40969 16745 41003 16779
rect 43913 16745 43947 16779
rect 44925 16745 44959 16779
rect 21097 16677 21131 16711
rect 28917 16677 28951 16711
rect 33701 16677 33735 16711
rect 4721 16609 4755 16643
rect 9321 16609 9355 16643
rect 9505 16609 9539 16643
rect 9965 16609 9999 16643
rect 11989 16609 12023 16643
rect 12081 16609 12115 16643
rect 12909 16609 12943 16643
rect 14657 16609 14691 16643
rect 14933 16609 14967 16643
rect 16497 16609 16531 16643
rect 16865 16609 16899 16643
rect 18291 16609 18325 16643
rect 18889 16609 18923 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 23213 16609 23247 16643
rect 24409 16609 24443 16643
rect 25053 16609 25087 16643
rect 25237 16609 25271 16643
rect 25973 16609 26007 16643
rect 27169 16609 27203 16643
rect 29469 16609 29503 16643
rect 31125 16609 31159 16643
rect 33241 16609 33275 16643
rect 34345 16609 34379 16643
rect 36461 16609 36495 16643
rect 37289 16609 37323 16643
rect 38761 16609 38795 16643
rect 38853 16609 38887 16643
rect 39497 16609 39531 16643
rect 41337 16609 41371 16643
rect 43361 16609 43395 16643
rect 43453 16609 43487 16643
rect 44557 16609 44591 16643
rect 4813 16541 4847 16575
rect 8493 16541 8527 16575
rect 8769 16541 8803 16575
rect 9689 16541 9723 16575
rect 18613 16541 18647 16575
rect 20637 16541 20671 16575
rect 20729 16541 20763 16575
rect 20913 16541 20947 16575
rect 21005 16541 21039 16575
rect 21373 16541 21407 16575
rect 21557 16541 21591 16575
rect 22937 16541 22971 16575
rect 25789 16541 25823 16575
rect 28089 16541 28123 16575
rect 28181 16541 28215 16575
rect 28273 16541 28307 16575
rect 28457 16541 28491 16575
rect 28733 16541 28767 16575
rect 29285 16541 29319 16575
rect 29745 16541 29779 16575
rect 29929 16541 29963 16575
rect 30849 16541 30883 16575
rect 33517 16541 33551 16575
rect 34069 16541 34103 16575
rect 37933 16541 37967 16575
rect 38209 16541 38243 16575
rect 38669 16541 38703 16575
rect 39221 16541 39255 16575
rect 41061 16541 41095 16575
rect 43269 16541 43303 16575
rect 5089 16473 5123 16507
rect 12817 16473 12851 16507
rect 20453 16473 20487 16507
rect 21925 16473 21959 16507
rect 24225 16473 24259 16507
rect 25881 16473 25915 16507
rect 27353 16473 27387 16507
rect 27537 16473 27571 16507
rect 30481 16473 30515 16507
rect 33149 16473 33183 16507
rect 36369 16473 36403 16507
rect 37105 16473 37139 16507
rect 3525 16405 3559 16439
rect 3893 16405 3927 16439
rect 4261 16405 4295 16439
rect 6561 16405 6595 16439
rect 7021 16405 7055 16439
rect 7665 16405 7699 16439
rect 8125 16405 8159 16439
rect 8309 16405 8343 16439
rect 8585 16405 8619 16439
rect 8861 16405 8895 16439
rect 9229 16405 9263 16439
rect 11437 16405 11471 16439
rect 11529 16405 11563 16439
rect 11897 16405 11931 16439
rect 12725 16405 12759 16439
rect 13829 16405 13863 16439
rect 14565 16405 14599 16439
rect 22017 16405 22051 16439
rect 22385 16405 22419 16439
rect 23765 16405 23799 16439
rect 24133 16405 24167 16439
rect 24961 16405 24995 16439
rect 25421 16405 25455 16439
rect 26433 16405 26467 16439
rect 26893 16405 26927 16439
rect 27721 16405 27755 16439
rect 27813 16405 27847 16439
rect 29377 16405 29411 16439
rect 32689 16405 32723 16439
rect 33057 16405 33091 16439
rect 35817 16405 35851 16439
rect 36277 16405 36311 16439
rect 37197 16405 37231 16439
rect 38025 16405 38059 16439
rect 38301 16405 38335 16439
rect 42809 16405 42843 16439
rect 42901 16405 42935 16439
rect 4721 16201 4755 16235
rect 5365 16201 5399 16235
rect 6101 16201 6135 16235
rect 6561 16201 6595 16235
rect 7113 16201 7147 16235
rect 7389 16201 7423 16235
rect 7757 16201 7791 16235
rect 9965 16201 9999 16235
rect 15301 16201 15335 16235
rect 17049 16201 17083 16235
rect 17509 16201 17543 16235
rect 18061 16201 18095 16235
rect 20637 16201 20671 16235
rect 21557 16201 21591 16235
rect 24133 16201 24167 16235
rect 26893 16201 26927 16235
rect 28549 16201 28583 16235
rect 31217 16201 31251 16235
rect 36185 16201 36219 16235
rect 40693 16201 40727 16235
rect 43545 16201 43579 16235
rect 8217 16133 8251 16167
rect 17141 16133 17175 16167
rect 18429 16133 18463 16167
rect 20269 16133 20303 16167
rect 21373 16133 21407 16167
rect 24501 16133 24535 16167
rect 27414 16133 27448 16167
rect 35817 16133 35851 16167
rect 36921 16133 36955 16167
rect 42073 16133 42107 16167
rect 5273 16065 5307 16099
rect 5457 16065 5491 16099
rect 5733 16065 5767 16099
rect 6286 16087 6320 16121
rect 6377 16065 6411 16099
rect 7941 16065 7975 16099
rect 10333 16065 10367 16099
rect 12909 16065 12943 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 15761 16065 15795 16099
rect 16129 16065 16163 16099
rect 16313 16065 16347 16099
rect 16405 16065 16439 16099
rect 16681 16065 16715 16099
rect 16865 16065 16899 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 17785 16065 17819 16099
rect 17877 16065 17911 16099
rect 20085 16065 20119 16099
rect 20361 16065 20395 16099
rect 20453 16065 20487 16099
rect 21281 16065 21315 16099
rect 21925 16065 21959 16099
rect 27077 16065 27111 16099
rect 28641 16065 28675 16099
rect 28825 16065 28859 16099
rect 28917 16065 28951 16099
rect 29010 16055 29044 16089
rect 31493 16065 31527 16099
rect 33517 16065 33551 16099
rect 35725 16065 35759 16099
rect 36369 16065 36403 16099
rect 40785 16065 40819 16099
rect 41337 16065 41371 16099
rect 41613 16065 41647 16099
rect 3617 15997 3651 16031
rect 4353 15997 4387 16031
rect 5089 15997 5123 16031
rect 5825 15997 5859 16031
rect 6561 15997 6595 16031
rect 10425 15997 10459 16031
rect 10517 15997 10551 16031
rect 10885 15997 10919 16031
rect 11161 15997 11195 16031
rect 13185 15997 13219 16031
rect 14933 15997 14967 16031
rect 15669 15997 15703 16031
rect 18153 15997 18187 16031
rect 22017 15997 22051 16031
rect 22201 15997 22235 16031
rect 22385 15997 22419 16031
rect 22661 15997 22695 16031
rect 24225 15997 24259 16031
rect 27169 15997 27203 16031
rect 29469 15997 29503 16031
rect 29745 15997 29779 16031
rect 31769 15997 31803 16031
rect 33793 15997 33827 16031
rect 35909 15997 35943 16031
rect 36645 15997 36679 16031
rect 38393 15997 38427 16031
rect 38485 15997 38519 16031
rect 38761 15997 38795 16031
rect 40877 15997 40911 16031
rect 41797 15997 41831 16031
rect 16129 15929 16163 15963
rect 19901 15929 19935 15963
rect 25973 15929 26007 15963
rect 26525 15929 26559 15963
rect 29285 15929 29319 15963
rect 35357 15929 35391 15963
rect 40325 15929 40359 15963
rect 41429 15929 41463 15963
rect 44557 15929 44591 15963
rect 44925 15929 44959 15963
rect 3341 15861 3375 15895
rect 4077 15861 4111 15895
rect 5917 15861 5951 15895
rect 9689 15861 9723 15895
rect 12633 15861 12667 15895
rect 16865 15861 16899 15895
rect 20913 15861 20947 15895
rect 33241 15861 33275 15895
rect 35265 15861 35299 15895
rect 40233 15861 40267 15895
rect 41153 15861 41187 15895
rect 43913 15861 43947 15895
rect 44281 15861 44315 15895
rect 3985 15657 4019 15691
rect 6837 15657 6871 15691
rect 14197 15657 14231 15691
rect 17233 15657 17267 15691
rect 19809 15657 19843 15691
rect 20361 15657 20395 15691
rect 21097 15657 21131 15691
rect 21649 15657 21683 15691
rect 27721 15657 27755 15691
rect 30205 15657 30239 15691
rect 30665 15657 30699 15691
rect 30849 15657 30883 15691
rect 33701 15657 33735 15691
rect 37933 15657 37967 15691
rect 38301 15657 38335 15691
rect 40969 15657 41003 15691
rect 7389 15589 7423 15623
rect 13461 15589 13495 15623
rect 13553 15589 13587 15623
rect 16681 15589 16715 15623
rect 16865 15589 16899 15623
rect 17417 15589 17451 15623
rect 19349 15589 19383 15623
rect 22845 15589 22879 15623
rect 28549 15589 28583 15623
rect 4721 15521 4755 15555
rect 8033 15521 8067 15555
rect 12725 15521 12759 15555
rect 13183 15521 13217 15555
rect 13921 15521 13955 15555
rect 14933 15521 14967 15555
rect 15209 15521 15243 15555
rect 20177 15521 20211 15555
rect 21005 15521 21039 15555
rect 22385 15521 22419 15555
rect 23305 15521 23339 15555
rect 23397 15521 23431 15555
rect 25513 15521 25547 15555
rect 25881 15521 25915 15555
rect 28273 15521 28307 15555
rect 30941 15521 30975 15555
rect 31217 15521 31251 15555
rect 32781 15521 32815 15555
rect 32965 15521 32999 15555
rect 33149 15521 33183 15555
rect 35909 15521 35943 15555
rect 38853 15521 38887 15555
rect 39497 15521 39531 15555
rect 41889 15521 41923 15555
rect 42717 15521 42751 15555
rect 4629 15453 4663 15487
rect 5089 15453 5123 15487
rect 7297 15453 7331 15487
rect 7757 15453 7791 15487
rect 8309 15453 8343 15487
rect 10517 15453 10551 15487
rect 10609 15453 10643 15487
rect 12541 15453 12575 15487
rect 12817 15453 12851 15487
rect 13461 15453 13495 15487
rect 13829 15453 13863 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 14841 15453 14875 15487
rect 17693 15453 17727 15487
rect 17877 15453 17911 15487
rect 17969 15453 18003 15487
rect 19625 15453 19659 15487
rect 20085 15453 20119 15487
rect 20269 15453 20303 15487
rect 20361 15453 20395 15487
rect 20545 15453 20579 15487
rect 20821 15453 20855 15487
rect 21281 15453 21315 15487
rect 23213 15453 23247 15487
rect 23765 15453 23799 15487
rect 25605 15453 25639 15487
rect 28089 15453 28123 15487
rect 28181 15453 28215 15487
rect 28733 15453 28767 15487
rect 29193 15453 29227 15487
rect 29285 15453 29319 15487
rect 29377 15453 29411 15487
rect 29561 15453 29595 15487
rect 29653 15453 29687 15487
rect 30021 15453 30055 15487
rect 33057 15453 33091 15487
rect 33241 15453 33275 15487
rect 33609 15453 33643 15487
rect 33885 15453 33919 15487
rect 34069 15453 34103 15487
rect 38669 15453 38703 15487
rect 39221 15453 39255 15487
rect 41245 15453 41279 15487
rect 41705 15453 41739 15487
rect 43177 15453 43211 15487
rect 44925 15453 44959 15487
rect 5365 15385 5399 15419
rect 8585 15385 8619 15419
rect 10885 15385 10919 15419
rect 13737 15385 13771 15419
rect 17509 15385 17543 15419
rect 19441 15385 19475 15419
rect 21189 15385 21223 15419
rect 21465 15385 21499 15419
rect 22201 15385 22235 15419
rect 24041 15385 24075 15419
rect 28917 15385 28951 15419
rect 29837 15385 29871 15419
rect 29929 15385 29963 15419
rect 30481 15385 30515 15419
rect 34345 15385 34379 15419
rect 36185 15385 36219 15419
rect 37749 15385 37783 15419
rect 37965 15385 37999 15419
rect 41797 15385 41831 15419
rect 42533 15385 42567 15419
rect 3525 15317 3559 15351
rect 4261 15317 4295 15351
rect 4997 15317 5031 15351
rect 7113 15317 7147 15351
rect 7849 15317 7883 15351
rect 10057 15317 10091 15351
rect 10333 15317 10367 15351
rect 12357 15317 12391 15351
rect 13001 15317 13035 15351
rect 13093 15317 13127 15351
rect 14657 15317 14691 15351
rect 17233 15317 17267 15351
rect 18337 15317 18371 15351
rect 18889 15317 18923 15351
rect 21833 15317 21867 15351
rect 22293 15317 22327 15351
rect 27353 15317 27387 15351
rect 30691 15317 30725 15351
rect 32689 15317 32723 15351
rect 33425 15317 33459 15351
rect 35817 15317 35851 15351
rect 37657 15317 37691 15351
rect 38117 15317 38151 15351
rect 38761 15317 38795 15351
rect 41061 15317 41095 15351
rect 41337 15317 41371 15351
rect 42165 15317 42199 15351
rect 42625 15317 42659 15351
rect 42993 15317 43027 15351
rect 43453 15317 43487 15351
rect 43913 15317 43947 15351
rect 44557 15317 44591 15351
rect 3985 15113 4019 15147
rect 4353 15113 4387 15147
rect 4629 15113 4663 15147
rect 9965 15113 9999 15147
rect 14289 15113 14323 15147
rect 15117 15113 15151 15147
rect 15485 15113 15519 15147
rect 17325 15113 17359 15147
rect 20637 15113 20671 15147
rect 22937 15113 22971 15147
rect 23489 15113 23523 15147
rect 23857 15113 23891 15147
rect 24317 15113 24351 15147
rect 25513 15113 25547 15147
rect 26617 15113 26651 15147
rect 27629 15113 27663 15147
rect 30665 15113 30699 15147
rect 31861 15113 31895 15147
rect 32689 15113 32723 15147
rect 34345 15113 34379 15147
rect 34713 15113 34747 15147
rect 35173 15113 35207 15147
rect 35541 15113 35575 15147
rect 36277 15113 36311 15147
rect 37013 15113 37047 15147
rect 6009 15045 6043 15079
rect 8033 15045 8067 15079
rect 10609 15045 10643 15079
rect 16957 15045 16991 15079
rect 17157 15045 17191 15079
rect 17509 15045 17543 15079
rect 22569 15045 22603 15079
rect 22753 15045 22787 15079
rect 30205 15045 30239 15079
rect 30297 15045 30331 15079
rect 30941 15045 30975 15079
rect 31585 15045 31619 15079
rect 32229 15045 32263 15079
rect 32321 15045 32355 15079
rect 33609 15045 33643 15079
rect 34253 15045 34287 15079
rect 37105 15045 37139 15079
rect 38393 15045 38427 15079
rect 39405 15045 39439 15079
rect 40141 15045 40175 15079
rect 42073 15045 42107 15079
rect 31171 15011 31205 15045
rect 949 14977 983 15011
rect 4445 14977 4479 15011
rect 4629 14977 4663 15011
rect 4721 14977 4755 15011
rect 5089 14977 5123 15011
rect 5273 14977 5307 15011
rect 11253 14977 11287 15011
rect 11437 14977 11471 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 12449 14977 12483 15011
rect 13093 14977 13127 15011
rect 13185 14977 13219 15011
rect 13921 14977 13955 15011
rect 16129 14977 16163 15011
rect 16589 14977 16623 15011
rect 17417 14977 17451 15011
rect 19809 14977 19843 15011
rect 20361 14977 20395 15011
rect 20545 14977 20579 15011
rect 20821 14977 20855 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 21557 14977 21591 15011
rect 22109 14977 22143 15011
rect 22385 14977 22419 15011
rect 23121 14977 23155 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 24501 14977 24535 15011
rect 25053 14977 25087 15011
rect 26157 14977 26191 15011
rect 26525 14977 26559 15011
rect 26801 14977 26835 15011
rect 27077 14977 27111 15011
rect 27169 14977 27203 15011
rect 27353 14977 27387 15011
rect 27905 14977 27939 15011
rect 27997 14977 28031 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28632 14977 28666 15011
rect 29837 14977 29871 15011
rect 30021 14977 30055 15011
rect 30481 14977 30515 15011
rect 32873 14977 32907 15011
rect 32965 14977 32999 15011
rect 33149 14977 33183 15011
rect 33885 14977 33919 15011
rect 35633 14977 35667 15011
rect 36461 14977 36495 15011
rect 39313 14977 39347 15011
rect 39865 14977 39899 15011
rect 45201 14977 45235 15011
rect 4997 14909 5031 14943
rect 5733 14909 5767 14943
rect 7757 14909 7791 14943
rect 9505 14909 9539 14943
rect 10057 14909 10091 14943
rect 10149 14909 10183 14943
rect 12173 14909 12207 14943
rect 15577 14909 15611 14943
rect 15761 14909 15795 14943
rect 16313 14909 16347 14943
rect 16865 14909 16899 14943
rect 22293 14909 22327 14943
rect 23949 14909 23983 14943
rect 24041 14909 24075 14943
rect 25605 14909 25639 14943
rect 25697 14909 25731 14943
rect 28365 14909 28399 14943
rect 32505 14909 32539 14943
rect 33057 14909 33091 14943
rect 34805 14909 34839 14943
rect 34989 14909 35023 14943
rect 35725 14909 35759 14943
rect 37197 14909 37231 14943
rect 39497 14909 39531 14943
rect 41797 14909 41831 14943
rect 4905 14841 4939 14875
rect 16773 14841 16807 14875
rect 18613 14841 18647 14875
rect 18981 14841 19015 14875
rect 19717 14841 19751 14875
rect 21373 14841 21407 14875
rect 25145 14841 25179 14875
rect 31769 14841 31803 14875
rect 36645 14841 36679 14875
rect 765 14773 799 14807
rect 4813 14773 4847 14807
rect 5273 14773 5307 14807
rect 5457 14773 5491 14807
rect 7481 14773 7515 14807
rect 9597 14773 9631 14807
rect 13645 14773 13679 14807
rect 14565 14773 14599 14807
rect 14933 14773 14967 14807
rect 17141 14773 17175 14807
rect 18153 14773 18187 14807
rect 19349 14773 19383 14807
rect 19993 14773 20027 14807
rect 20177 14773 20211 14807
rect 20821 14773 20855 14807
rect 23305 14773 23339 14807
rect 24869 14773 24903 14807
rect 25973 14773 26007 14807
rect 26341 14773 26375 14807
rect 26893 14773 26927 14807
rect 27537 14773 27571 14807
rect 29745 14773 29779 14807
rect 31125 14773 31159 14807
rect 31309 14773 31343 14807
rect 37657 14773 37691 14807
rect 38025 14773 38059 14807
rect 38761 14773 38795 14807
rect 38945 14773 38979 14807
rect 41613 14773 41647 14807
rect 43545 14773 43579 14807
rect 43913 14773 43947 14807
rect 44189 14773 44223 14807
rect 44557 14773 44591 14807
rect 45017 14773 45051 14807
rect 4261 14569 4295 14603
rect 6745 14569 6779 14603
rect 12173 14569 12207 14603
rect 16865 14569 16899 14603
rect 19533 14569 19567 14603
rect 19809 14569 19843 14603
rect 21695 14569 21729 14603
rect 24593 14569 24627 14603
rect 27261 14569 27295 14603
rect 31401 14569 31435 14603
rect 32229 14569 32263 14603
rect 32597 14569 32631 14603
rect 36645 14569 36679 14603
rect 38301 14569 38335 14603
rect 41705 14569 41739 14603
rect 43913 14569 43947 14603
rect 7113 14501 7147 14535
rect 7573 14501 7607 14535
rect 13461 14501 13495 14535
rect 18337 14501 18371 14535
rect 23305 14501 23339 14535
rect 23765 14501 23799 14535
rect 31585 14501 31619 14535
rect 32965 14501 32999 14535
rect 33333 14501 33367 14535
rect 33609 14501 33643 14535
rect 36001 14501 36035 14535
rect 37013 14501 37047 14535
rect 4629 14433 4663 14467
rect 11345 14433 11379 14467
rect 11805 14433 11839 14467
rect 12014 14433 12048 14467
rect 13185 14433 13219 14467
rect 14105 14433 14139 14467
rect 15393 14433 15427 14467
rect 19533 14433 19567 14467
rect 25053 14433 25087 14467
rect 25145 14433 25179 14467
rect 25697 14433 25731 14467
rect 27813 14433 27847 14467
rect 28917 14433 28951 14467
rect 30757 14433 30791 14467
rect 30849 14433 30883 14467
rect 30941 14433 30975 14467
rect 31033 14433 31067 14467
rect 34621 14433 34655 14467
rect 35357 14433 35391 14467
rect 35725 14433 35759 14467
rect 38945 14433 38979 14467
rect 40969 14433 41003 14467
rect 42257 14433 42291 14467
rect 4537 14365 4571 14399
rect 4997 14365 5031 14399
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 11529 14365 11563 14399
rect 12449 14365 12483 14399
rect 14473 14365 14507 14399
rect 15117 14365 15151 14399
rect 18153 14365 18187 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 18797 14365 18831 14399
rect 18981 14365 19015 14399
rect 19625 14365 19659 14399
rect 19901 14365 19935 14399
rect 20269 14365 20303 14399
rect 21833 14365 21867 14399
rect 22569 14365 22603 14399
rect 22753 14365 22787 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 23397 14365 23431 14399
rect 23949 14365 23983 14399
rect 24041 14365 24075 14399
rect 24225 14365 24259 14399
rect 24317 14365 24351 14399
rect 25421 14365 25455 14399
rect 27629 14365 27663 14399
rect 28273 14365 28307 14399
rect 28365 14365 28399 14399
rect 29173 14365 29207 14399
rect 31953 14365 31987 14399
rect 33517 14365 33551 14399
rect 33793 14365 33827 14399
rect 34529 14365 34563 14399
rect 34897 14365 34931 14399
rect 35633 14365 35667 14399
rect 36277 14365 36311 14399
rect 37197 14365 37231 14399
rect 38025 14365 38059 14399
rect 39221 14365 39255 14399
rect 42165 14365 42199 14399
rect 5273 14297 5307 14331
rect 8585 14297 8619 14331
rect 10241 14297 10275 14331
rect 11069 14297 11103 14331
rect 11897 14297 11931 14331
rect 13829 14297 13863 14331
rect 18889 14297 18923 14331
rect 19349 14297 19383 14331
rect 22385 14297 22419 14331
rect 24961 14297 24995 14331
rect 31217 14297 31251 14331
rect 34437 14297 34471 14331
rect 35842 14297 35876 14331
rect 37289 14297 37323 14331
rect 38669 14297 38703 14331
rect 39497 14297 39531 14331
rect 3801 14229 3835 14263
rect 4905 14229 4939 14263
rect 7665 14229 7699 14263
rect 7941 14229 7975 14263
rect 10057 14229 10091 14263
rect 10333 14229 10367 14263
rect 10701 14229 10735 14263
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 12541 14229 12575 14263
rect 12909 14229 12943 14263
rect 13001 14229 13035 14263
rect 13921 14229 13955 14263
rect 14289 14229 14323 14263
rect 14933 14229 14967 14263
rect 17417 14229 17451 14263
rect 17785 14229 17819 14263
rect 17969 14229 18003 14263
rect 19165 14229 19199 14263
rect 22017 14229 22051 14263
rect 27169 14229 27203 14263
rect 27721 14229 27755 14263
rect 28089 14229 28123 14263
rect 28549 14229 28583 14263
rect 30297 14229 30331 14263
rect 30573 14229 30607 14263
rect 31417 14229 31451 14263
rect 34069 14229 34103 14263
rect 35081 14229 35115 14263
rect 36093 14229 36127 14263
rect 37381 14229 37415 14263
rect 37565 14229 37599 14263
rect 37841 14229 37875 14263
rect 38761 14229 38795 14263
rect 41245 14229 41279 14263
rect 42073 14229 42107 14263
rect 42809 14229 42843 14263
rect 43085 14229 43119 14263
rect 43453 14229 43487 14263
rect 44557 14229 44591 14263
rect 44925 14229 44959 14263
rect 3525 14025 3559 14059
rect 6929 14025 6963 14059
rect 7205 14025 7239 14059
rect 7389 14025 7423 14059
rect 12817 14025 12851 14059
rect 15209 14025 15243 14059
rect 20085 14025 20119 14059
rect 20377 14025 20411 14059
rect 20545 14025 20579 14059
rect 21649 14025 21683 14059
rect 26065 14025 26099 14059
rect 27721 14025 27755 14059
rect 27813 14025 27847 14059
rect 28181 14025 28215 14059
rect 28273 14025 28307 14059
rect 28641 14025 28675 14059
rect 29009 14025 29043 14059
rect 29101 14025 29135 14059
rect 31585 14025 31619 14059
rect 32689 14025 32723 14059
rect 34713 14025 34747 14059
rect 35725 14025 35759 14059
rect 36185 14025 36219 14059
rect 41153 14025 41187 14059
rect 41797 14025 41831 14059
rect 42257 14025 42291 14059
rect 4077 13957 4111 13991
rect 7757 13957 7791 13991
rect 8493 13957 8527 13991
rect 15117 13957 15151 13991
rect 17877 13957 17911 13991
rect 17969 13957 18003 13991
rect 18613 13957 18647 13991
rect 20177 13957 20211 13991
rect 20637 13957 20671 13991
rect 20837 13957 20871 13991
rect 21373 13957 21407 13991
rect 22569 13957 22603 13991
rect 25237 13957 25271 13991
rect 25329 13957 25363 13991
rect 26608 13957 26642 13991
rect 33149 13957 33183 13991
rect 36093 13957 36127 13991
rect 37749 13957 37783 13991
rect 1777 13889 1811 13923
rect 7849 13889 7883 13923
rect 8217 13889 8251 13923
rect 10241 13889 10275 13923
rect 10701 13889 10735 13923
rect 15761 13889 15795 13923
rect 16773 13889 16807 13923
rect 17693 13889 17727 13923
rect 18061 13889 18095 13923
rect 18337 13889 18371 13923
rect 22017 13889 22051 13923
rect 22201 13889 22235 13923
rect 22661 13889 22695 13923
rect 23121 13889 23155 13923
rect 23397 13889 23431 13923
rect 23857 13889 23891 13923
rect 24225 13889 24259 13923
rect 24869 13889 24903 13923
rect 25513 13889 25547 13923
rect 25605 13889 25639 13923
rect 25789 13889 25823 13923
rect 29561 13889 29595 13923
rect 31953 13889 31987 13923
rect 35081 13889 35115 13923
rect 36737 13889 36771 13923
rect 37197 13889 37231 13923
rect 37473 13889 37507 13923
rect 41337 13889 41371 13923
rect 42165 13889 42199 13923
rect 2053 13821 2087 13855
rect 3801 13821 3835 13855
rect 8033 13821 8067 13855
rect 9965 13821 9999 13855
rect 11069 13821 11103 13855
rect 12909 13821 12943 13855
rect 14657 13821 14691 13855
rect 15301 13821 15335 13855
rect 16589 13821 16623 13855
rect 16865 13821 16899 13855
rect 16957 13821 16991 13855
rect 17049 13821 17083 13855
rect 24685 13821 24719 13855
rect 26341 13821 26375 13855
rect 28365 13821 28399 13855
rect 29193 13821 29227 13855
rect 31309 13821 31343 13855
rect 32045 13821 32079 13855
rect 32137 13821 32171 13855
rect 32873 13821 32907 13855
rect 35173 13821 35207 13855
rect 35265 13821 35299 13855
rect 36369 13821 36403 13855
rect 37105 13821 37139 13855
rect 39313 13821 39347 13855
rect 39589 13821 39623 13855
rect 41061 13821 41095 13855
rect 42349 13821 42383 13855
rect 42809 13821 42843 13855
rect 14749 13753 14783 13787
rect 21005 13753 21039 13787
rect 22201 13753 22235 13787
rect 43545 13753 43579 13787
rect 43913 13753 43947 13787
rect 44741 13753 44775 13787
rect 5549 13685 5583 13719
rect 6193 13685 6227 13719
rect 6469 13685 6503 13719
rect 10057 13685 10091 13719
rect 10517 13685 10551 13719
rect 11332 13685 11366 13719
rect 13172 13685 13206 13719
rect 15577 13685 15611 13719
rect 16497 13685 16531 13719
rect 17509 13685 17543 13719
rect 18245 13685 18279 13719
rect 20361 13685 20395 13719
rect 20821 13685 20855 13719
rect 24501 13685 24535 13719
rect 25145 13685 25179 13719
rect 25329 13685 25363 13719
rect 29824 13685 29858 13719
rect 34621 13685 34655 13719
rect 37197 13685 37231 13719
rect 37381 13685 37415 13719
rect 39221 13685 39255 13719
rect 43177 13685 43211 13719
rect 44281 13685 44315 13719
rect 45109 13685 45143 13719
rect 3893 13481 3927 13515
rect 4721 13481 4755 13515
rect 5549 13481 5583 13515
rect 8769 13481 8803 13515
rect 11345 13481 11379 13515
rect 13185 13481 13219 13515
rect 16497 13481 16531 13515
rect 18429 13481 18463 13515
rect 19349 13481 19383 13515
rect 19717 13481 19751 13515
rect 20164 13481 20198 13515
rect 22845 13481 22879 13515
rect 23305 13481 23339 13515
rect 24317 13481 24351 13515
rect 26617 13481 26651 13515
rect 26893 13481 26927 13515
rect 27077 13481 27111 13515
rect 29653 13481 29687 13515
rect 30113 13481 30147 13515
rect 32597 13481 32631 13515
rect 37749 13481 37783 13515
rect 38117 13481 38151 13515
rect 41337 13481 41371 13515
rect 5733 13413 5767 13447
rect 19165 13413 19199 13447
rect 24501 13413 24535 13447
rect 30573 13413 30607 13447
rect 41613 13413 41647 13447
rect 42349 13413 42383 13447
rect 43085 13413 43119 13447
rect 43453 13413 43487 13447
rect 5917 13345 5951 13379
rect 9413 13345 9447 13379
rect 9873 13345 9907 13379
rect 13737 13345 13771 13379
rect 16037 13345 16071 13379
rect 16957 13345 16991 13379
rect 21925 13345 21959 13379
rect 22109 13345 22143 13379
rect 22661 13345 22695 13379
rect 25145 13345 25179 13379
rect 27353 13345 27387 13379
rect 33149 13345 33183 13379
rect 33241 13345 33275 13379
rect 34069 13345 34103 13379
rect 35909 13345 35943 13379
rect 36185 13345 36219 13379
rect 37657 13345 37691 13379
rect 38761 13345 38795 13379
rect 5641 13277 5675 13311
rect 6285 13277 6319 13311
rect 8677 13277 8711 13311
rect 9597 13277 9631 13311
rect 11437 13277 11471 13311
rect 13461 13277 13495 13311
rect 15301 13277 15335 13311
rect 15945 13277 15979 13311
rect 16405 13277 16439 13311
rect 16681 13277 16715 13311
rect 18613 13277 18647 13311
rect 18797 13277 18831 13311
rect 18889 13277 18923 13311
rect 18981 13277 19015 13311
rect 19441 13277 19475 13311
rect 19533 13277 19567 13311
rect 19901 13277 19935 13311
rect 22017 13277 22051 13311
rect 22195 13277 22229 13311
rect 22315 13277 22349 13311
rect 22937 13277 22971 13311
rect 23305 13277 23339 13311
rect 23489 13277 23523 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 24317 13277 24351 13311
rect 24869 13277 24903 13311
rect 27620 13277 27654 13311
rect 29193 13277 29227 13311
rect 29285 13277 29319 13311
rect 29377 13277 29411 13311
rect 29561 13277 29595 13311
rect 29837 13277 29871 13311
rect 30757 13277 30791 13311
rect 30849 13277 30883 13311
rect 33701 13277 33735 13311
rect 37749 13277 37783 13311
rect 37933 13277 37967 13311
rect 39221 13277 39255 13311
rect 6561 13209 6595 13243
rect 11713 13209 11747 13243
rect 19257 13209 19291 13243
rect 26709 13209 26743 13243
rect 31125 13209 31159 13243
rect 34345 13209 34379 13243
rect 38485 13209 38519 13243
rect 39497 13209 39531 13243
rect 45017 13209 45051 13243
rect 3433 13141 3467 13175
rect 4353 13141 4387 13175
rect 5089 13141 5123 13175
rect 5917 13141 5951 13175
rect 8033 13141 8067 13175
rect 8493 13141 8527 13175
rect 9137 13141 9171 13175
rect 9229 13141 9263 13175
rect 15209 13141 15243 13175
rect 22477 13141 22511 13175
rect 23121 13141 23155 13175
rect 26909 13141 26943 13175
rect 28733 13141 28767 13175
rect 28917 13141 28951 13175
rect 32689 13141 32723 13175
rect 33057 13141 33091 13175
rect 33517 13141 33551 13175
rect 35817 13141 35851 13175
rect 38577 13141 38611 13175
rect 40969 13141 41003 13175
rect 41981 13141 42015 13175
rect 42717 13141 42751 13175
rect 43821 13141 43855 13175
rect 44557 13141 44591 13175
rect 7481 12937 7515 12971
rect 11437 12937 11471 12971
rect 12173 12937 12207 12971
rect 12265 12937 12299 12971
rect 13553 12937 13587 12971
rect 13645 12937 13679 12971
rect 17831 12937 17865 12971
rect 20269 12937 20303 12971
rect 20729 12937 20763 12971
rect 20821 12937 20855 12971
rect 22937 12937 22971 12971
rect 23121 12937 23155 12971
rect 24501 12937 24535 12971
rect 25697 12937 25731 12971
rect 27813 12937 27847 12971
rect 28273 12937 28307 12971
rect 29009 12937 29043 12971
rect 31125 12937 31159 12971
rect 35081 12937 35115 12971
rect 35265 12937 35299 12971
rect 35909 12937 35943 12971
rect 38393 12937 38427 12971
rect 40049 12937 40083 12971
rect 42441 12937 42475 12971
rect 4813 12869 4847 12903
rect 6009 12869 6043 12903
rect 9045 12869 9079 12903
rect 10977 12869 11011 12903
rect 11713 12869 11747 12903
rect 13369 12869 13403 12903
rect 13737 12869 13771 12903
rect 18245 12869 18279 12903
rect 20361 12869 20395 12903
rect 20577 12869 20611 12903
rect 25789 12869 25823 12903
rect 26341 12869 26375 12903
rect 26557 12869 26591 12903
rect 28181 12869 28215 12903
rect 29193 12869 29227 12903
rect 30113 12869 30147 12903
rect 30665 12869 30699 12903
rect 31769 12869 31803 12903
rect 33609 12869 33643 12903
rect 36001 12869 36035 12903
rect 39221 12869 39255 12903
rect 39681 12869 39715 12903
rect 39773 12869 39807 12903
rect 39957 12869 39991 12903
rect 4721 12801 4755 12835
rect 4905 12801 4939 12835
rect 5181 12801 5215 12835
rect 8769 12801 8803 12835
rect 12817 12801 12851 12835
rect 17969 12801 18003 12835
rect 19809 12801 19843 12835
rect 20085 12801 20119 12835
rect 21005 12801 21039 12835
rect 23489 12801 23523 12835
rect 23581 12801 23615 12835
rect 23765 12801 23799 12835
rect 23857 12801 23891 12835
rect 24317 12801 24351 12835
rect 24869 12781 24903 12815
rect 27261 12801 27295 12835
rect 27353 12801 27387 12835
rect 27445 12801 27479 12835
rect 27629 12801 27663 12835
rect 28641 12801 28675 12835
rect 28825 12801 28859 12835
rect 29101 12801 29135 12835
rect 29745 12801 29779 12835
rect 30297 12801 30331 12835
rect 30389 12801 30423 12835
rect 31309 12801 31343 12835
rect 33333 12801 33367 12835
rect 35449 12801 35483 12835
rect 36645 12801 36679 12835
rect 39037 12801 39071 12835
rect 40233 12801 40267 12835
rect 5273 12733 5307 12767
rect 5733 12733 5767 12767
rect 8585 12733 8619 12767
rect 10517 12733 10551 12767
rect 11529 12733 11563 12767
rect 12357 12733 12391 12767
rect 13001 12733 13035 12767
rect 14013 12733 14047 12767
rect 14289 12733 14323 12767
rect 16037 12733 16071 12767
rect 16405 12733 16439 12767
rect 19901 12733 19935 12767
rect 21189 12733 21223 12767
rect 21465 12733 21499 12767
rect 24133 12733 24167 12767
rect 24778 12733 24812 12767
rect 25145 12733 25179 12767
rect 25237 12733 25271 12767
rect 25973 12733 26007 12767
rect 28365 12733 28399 12767
rect 29561 12733 29595 12767
rect 31493 12733 31527 12767
rect 36093 12733 36127 12767
rect 36921 12733 36955 12767
rect 41981 12733 42015 12767
rect 42717 12733 42751 12767
rect 43453 12733 43487 12767
rect 43821 12733 43855 12767
rect 44189 12733 44223 12767
rect 44557 12733 44591 12767
rect 8309 12665 8343 12699
rect 10977 12665 11011 12699
rect 26985 12665 27019 12699
rect 35541 12665 35575 12699
rect 38853 12665 38887 12699
rect 39221 12665 39255 12699
rect 40601 12665 40635 12699
rect 41245 12665 41279 12699
rect 5457 12597 5491 12631
rect 7849 12597 7883 12631
rect 11805 12597 11839 12631
rect 13921 12597 13955 12631
rect 15761 12597 15795 12631
rect 19717 12597 19751 12631
rect 20085 12597 20119 12631
rect 20545 12597 20579 12631
rect 24133 12597 24167 12631
rect 24593 12597 24627 12631
rect 25329 12597 25363 12631
rect 26525 12597 26559 12631
rect 26709 12597 26743 12631
rect 29929 12597 29963 12631
rect 30113 12597 30147 12631
rect 33241 12597 33275 12631
rect 38761 12597 38795 12631
rect 40877 12597 40911 12631
rect 43085 12597 43119 12631
rect 44925 12597 44959 12631
rect 5181 12393 5215 12427
rect 7021 12393 7055 12427
rect 7113 12393 7147 12427
rect 8033 12393 8067 12427
rect 11345 12393 11379 12427
rect 11621 12393 11655 12427
rect 12449 12393 12483 12427
rect 15393 12393 15427 12427
rect 17693 12393 17727 12427
rect 19349 12393 19383 12427
rect 19809 12393 19843 12427
rect 23397 12393 23431 12427
rect 23581 12393 23615 12427
rect 24593 12393 24627 12427
rect 25053 12393 25087 12427
rect 26893 12393 26927 12427
rect 30941 12393 30975 12427
rect 33241 12393 33275 12427
rect 33885 12393 33919 12427
rect 34069 12393 34103 12427
rect 34897 12393 34931 12427
rect 37197 12393 37231 12427
rect 43545 12393 43579 12427
rect 7573 12325 7607 12359
rect 8769 12325 8803 12359
rect 16865 12325 16899 12359
rect 17417 12325 17451 12359
rect 19257 12325 19291 12359
rect 19993 12325 20027 12359
rect 22845 12325 22879 12359
rect 23765 12325 23799 12359
rect 28365 12325 28399 12359
rect 41429 12325 41463 12359
rect 5273 12257 5307 12291
rect 7297 12257 7331 12291
rect 9873 12257 9907 12291
rect 14749 12257 14783 12291
rect 24777 12257 24811 12291
rect 25421 12257 25455 12291
rect 27905 12257 27939 12291
rect 29009 12257 29043 12291
rect 32597 12257 32631 12291
rect 33333 12257 33367 12291
rect 34621 12257 34655 12291
rect 34989 12257 35023 12291
rect 35449 12257 35483 12291
rect 35725 12257 35759 12291
rect 37749 12257 37783 12291
rect 37933 12257 37967 12291
rect 38577 12257 38611 12291
rect 38669 12257 38703 12291
rect 39773 12257 39807 12291
rect 40325 12257 40359 12291
rect 40969 12257 41003 12291
rect 7389 12189 7423 12223
rect 9597 12189 9631 12223
rect 11805 12189 11839 12223
rect 12633 12189 12667 12223
rect 13737 12189 13771 12223
rect 14013 12189 14047 12223
rect 14933 12189 14967 12223
rect 15485 12189 15519 12223
rect 15741 12189 15775 12223
rect 17877 12189 17911 12223
rect 18153 12189 18187 12223
rect 18245 12189 18279 12223
rect 18613 12189 18647 12223
rect 18761 12189 18795 12223
rect 18981 12189 19015 12223
rect 19078 12189 19112 12223
rect 19349 12189 19383 12223
rect 19533 12189 19567 12223
rect 20177 12189 20211 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 20545 12189 20579 12223
rect 20729 12189 20763 12223
rect 21097 12189 21131 12223
rect 23121 12189 23155 12223
rect 24041 12189 24075 12223
rect 24133 12189 24167 12223
rect 24225 12189 24259 12223
rect 24409 12189 24443 12223
rect 24501 12189 24535 12223
rect 25145 12189 25179 12223
rect 27169 12189 27203 12223
rect 31125 12189 31159 12223
rect 31585 12189 31619 12223
rect 32505 12189 32539 12223
rect 33701 12189 33735 12223
rect 34437 12189 34471 12223
rect 35173 12189 35207 12223
rect 37657 12189 37691 12223
rect 38485 12189 38519 12223
rect 4813 12121 4847 12155
rect 4997 12121 5031 12155
rect 5549 12121 5583 12155
rect 7113 12121 7147 12155
rect 18061 12121 18095 12155
rect 18889 12121 18923 12155
rect 19625 12121 19659 12155
rect 19825 12121 19859 12155
rect 21373 12121 21407 12155
rect 27721 12121 27755 12155
rect 29285 12121 29319 12155
rect 34897 12121 34931 12155
rect 39589 12121 39623 12155
rect 42533 12121 42567 12155
rect 43177 12121 43211 12155
rect 9045 12053 9079 12087
rect 9413 12053 9447 12087
rect 12265 12053 12299 12087
rect 13185 12053 13219 12087
rect 13829 12053 13863 12087
rect 18429 12053 18463 12087
rect 20637 12053 20671 12087
rect 26985 12053 27019 12087
rect 27353 12053 27387 12087
rect 27813 12053 27847 12087
rect 30757 12053 30791 12087
rect 31953 12053 31987 12087
rect 32873 12053 32907 12087
rect 33517 12053 33551 12087
rect 34529 12053 34563 12087
rect 35357 12053 35391 12087
rect 37289 12053 37323 12087
rect 38117 12053 38151 12087
rect 39221 12053 39255 12087
rect 39681 12053 39715 12087
rect 40693 12053 40727 12087
rect 41797 12053 41831 12087
rect 42073 12053 42107 12087
rect 42809 12053 42843 12087
rect 43913 12053 43947 12087
rect 44557 12053 44591 12087
rect 44925 12053 44959 12087
rect 4905 11849 4939 11883
rect 8217 11849 8251 11883
rect 8953 11849 8987 11883
rect 9505 11849 9539 11883
rect 9965 11849 9999 11883
rect 11161 11849 11195 11883
rect 16037 11849 16071 11883
rect 16405 11849 16439 11883
rect 19441 11849 19475 11883
rect 20453 11849 20487 11883
rect 21189 11849 21223 11883
rect 28089 11849 28123 11883
rect 31033 11849 31067 11883
rect 31677 11849 31711 11883
rect 32505 11849 32539 11883
rect 33625 11849 33659 11883
rect 33793 11849 33827 11883
rect 35633 11849 35667 11883
rect 38393 11849 38427 11883
rect 40785 11849 40819 11883
rect 41521 11849 41555 11883
rect 42349 11849 42383 11883
rect 42717 11849 42751 11883
rect 5181 11781 5215 11815
rect 6009 11781 6043 11815
rect 9873 11781 9907 11815
rect 14381 11781 14415 11815
rect 16497 11781 16531 11815
rect 17325 11781 17359 11815
rect 17785 11781 17819 11815
rect 19625 11781 19659 11815
rect 23673 11781 23707 11815
rect 24409 11781 24443 11815
rect 26617 11781 26651 11815
rect 28457 11781 28491 11815
rect 32781 11781 32815 11815
rect 33425 11781 33459 11815
rect 34345 11781 34379 11815
rect 5089 11713 5123 11747
rect 5281 11713 5315 11747
rect 5371 11713 5405 11747
rect 5549 11711 5583 11745
rect 11529 11713 11563 11747
rect 16957 11713 16991 11747
rect 17233 11713 17267 11747
rect 19341 11719 19375 11753
rect 19855 11747 19889 11781
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 20637 11713 20671 11747
rect 20729 11713 20763 11747
rect 21005 11713 21039 11747
rect 21373 11713 21407 11747
rect 30021 11713 30055 11747
rect 30573 11713 30607 11747
rect 31493 11713 31527 11747
rect 31769 11713 31803 11747
rect 31953 11713 31987 11747
rect 33333 11713 33367 11747
rect 34253 11713 34287 11747
rect 34713 11713 34747 11747
rect 35265 11713 35299 11747
rect 36093 11713 36127 11747
rect 36369 11713 36403 11747
rect 40325 11713 40359 11747
rect 40601 11713 40635 11747
rect 43085 11713 43119 11747
rect 43453 11713 43487 11747
rect 5457 11645 5491 11679
rect 5733 11645 5767 11679
rect 7481 11645 7515 11679
rect 10149 11645 10183 11679
rect 11345 11645 11379 11679
rect 12265 11645 12299 11679
rect 12541 11645 12575 11679
rect 14105 11645 14139 11679
rect 16589 11645 16623 11679
rect 17509 11645 17543 11679
rect 19257 11645 19291 11679
rect 21741 11645 21775 11679
rect 22017 11645 22051 11679
rect 24133 11645 24167 11679
rect 26157 11645 26191 11679
rect 26341 11645 26375 11679
rect 28181 11645 28215 11679
rect 29929 11645 29963 11679
rect 30481 11645 30515 11679
rect 34437 11645 34471 11679
rect 36645 11645 36679 11679
rect 36921 11645 36955 11679
rect 38485 11645 38519 11679
rect 38761 11645 38795 11679
rect 40417 11645 40451 11679
rect 42073 11645 42107 11679
rect 44833 11645 44867 11679
rect 10609 11577 10643 11611
rect 12081 11577 12115 11611
rect 19993 11577 20027 11611
rect 20177 11577 20211 11611
rect 23489 11577 23523 11611
rect 31493 11577 31527 11611
rect 34897 11577 34931 11611
rect 35909 11577 35943 11611
rect 7849 11509 7883 11543
rect 8585 11509 8619 11543
rect 9321 11509 9355 11543
rect 11713 11509 11747 11543
rect 14013 11509 14047 11543
rect 15853 11509 15887 11543
rect 17049 11509 17083 11543
rect 19809 11509 19843 11543
rect 20913 11509 20947 11543
rect 23765 11509 23799 11543
rect 30113 11509 30147 11543
rect 30849 11509 30883 11543
rect 32045 11509 32079 11543
rect 33149 11509 33183 11543
rect 33609 11509 33643 11543
rect 33885 11509 33919 11543
rect 35081 11509 35115 11543
rect 36185 11509 36219 11543
rect 40233 11509 40267 11543
rect 40325 11509 40359 11543
rect 41061 11509 41095 11543
rect 5457 11305 5491 11339
rect 7021 11305 7055 11339
rect 7757 11305 7791 11339
rect 8125 11305 8159 11339
rect 8861 11305 8895 11339
rect 10149 11305 10183 11339
rect 13461 11305 13495 11339
rect 14105 11305 14139 11339
rect 18245 11305 18279 11339
rect 18797 11305 18831 11339
rect 19533 11305 19567 11339
rect 20729 11305 20763 11339
rect 21005 11305 21039 11339
rect 21189 11305 21223 11339
rect 22017 11305 22051 11339
rect 23305 11305 23339 11339
rect 24961 11305 24995 11339
rect 27905 11305 27939 11339
rect 27997 11305 28031 11339
rect 32413 11305 32447 11339
rect 32873 11305 32907 11339
rect 37197 11305 37231 11339
rect 42625 11305 42659 11339
rect 43361 11305 43395 11339
rect 11437 11237 11471 11271
rect 12817 11237 12851 11271
rect 13185 11237 13219 11271
rect 14657 11237 14691 11271
rect 17601 11237 17635 11271
rect 25329 11237 25363 11271
rect 32597 11237 32631 11271
rect 33057 11237 33091 11271
rect 33149 11237 33183 11271
rect 38301 11237 38335 11271
rect 41153 11237 41187 11271
rect 43637 11237 43671 11271
rect 5089 11169 5123 11203
rect 11989 11169 12023 11203
rect 12449 11169 12483 11203
rect 20085 11169 20119 11203
rect 21741 11169 21775 11203
rect 22477 11169 22511 11203
rect 24225 11169 24259 11203
rect 26157 11169 26191 11203
rect 26433 11169 26467 11203
rect 29285 11169 29319 11203
rect 30113 11169 30147 11203
rect 32137 11169 32171 11203
rect 33609 11169 33643 11203
rect 33793 11169 33827 11203
rect 34437 11169 34471 11203
rect 38025 11169 38059 11203
rect 38761 11169 38795 11203
rect 38853 11169 38887 11203
rect 41797 11169 41831 11203
rect 4813 11101 4847 11135
rect 4905 11101 4939 11135
rect 9413 11101 9447 11135
rect 9597 11101 9631 11135
rect 10425 11101 10459 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10701 11101 10735 11135
rect 11253 11101 11287 11135
rect 11345 11101 11379 11135
rect 11529 11101 11563 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 13645 11101 13679 11135
rect 13921 11101 13955 11135
rect 14013 11101 14047 11135
rect 14105 11101 14139 11135
rect 14473 11101 14507 11135
rect 15117 11101 15151 11135
rect 17785 11101 17819 11135
rect 17877 11101 17911 11135
rect 18705 11101 18739 11135
rect 19993 11101 20027 11135
rect 20177 11101 20211 11135
rect 20913 11101 20947 11135
rect 22201 11101 22235 11135
rect 22293 11101 22327 11135
rect 22569 11101 22603 11135
rect 22937 11101 22971 11135
rect 24041 11101 24075 11135
rect 24685 11101 24719 11135
rect 28181 11101 28215 11135
rect 28549 11101 28583 11135
rect 29009 11101 29043 11135
rect 34253 11101 34287 11135
rect 36553 11101 36587 11135
rect 37381 11101 37415 11135
rect 38669 11101 38703 11135
rect 39221 11101 39255 11135
rect 41521 11101 41555 11135
rect 42257 11101 42291 11135
rect 8953 11033 8987 11067
rect 9137 11033 9171 11067
rect 9505 11033 9539 11067
rect 13829 11033 13863 11067
rect 15393 11033 15427 11067
rect 17509 11033 17543 11067
rect 18061 11033 18095 11067
rect 23121 11033 23155 11067
rect 29561 11033 29595 11067
rect 30389 11033 30423 11067
rect 32229 11033 32263 11067
rect 32689 11033 32723 11067
rect 33517 11033 33551 11067
rect 34713 11033 34747 11067
rect 37841 11033 37875 11067
rect 39497 11033 39531 11067
rect 44097 11033 44131 11067
rect 5089 10965 5123 10999
rect 5733 10965 5767 10999
rect 6193 10965 6227 10999
rect 6561 10965 6595 10999
rect 7297 10965 7331 10999
rect 9321 10965 9355 10999
rect 10241 10965 10275 10999
rect 11069 10965 11103 10999
rect 11713 10965 11747 10999
rect 14381 10965 14415 10999
rect 16865 10965 16899 10999
rect 19901 10965 19935 10999
rect 21557 10965 21591 10999
rect 21649 10965 21683 10999
rect 25697 10965 25731 10999
rect 28641 10965 28675 10999
rect 29653 10965 29687 10999
rect 32434 10965 32468 10999
rect 32899 10965 32933 10999
rect 34069 10965 34103 10999
rect 36185 10965 36219 10999
rect 36829 10965 36863 10999
rect 37473 10965 37507 10999
rect 37933 10965 37967 10999
rect 40969 10965 41003 10999
rect 41613 10965 41647 10999
rect 42993 10965 43027 10999
rect 44557 10965 44591 10999
rect 44925 10965 44959 10999
rect 7113 10761 7147 10795
rect 8493 10761 8527 10795
rect 10609 10761 10643 10795
rect 12633 10761 12667 10795
rect 17141 10761 17175 10795
rect 18981 10761 19015 10795
rect 21833 10761 21867 10795
rect 22385 10761 22419 10795
rect 22569 10761 22603 10795
rect 25329 10761 25363 10795
rect 25697 10761 25731 10795
rect 28273 10761 28307 10795
rect 29393 10761 29427 10795
rect 30021 10761 30055 10795
rect 30757 10761 30791 10795
rect 35081 10761 35115 10795
rect 35541 10761 35575 10795
rect 36461 10761 36495 10795
rect 36645 10761 36679 10795
rect 37565 10761 37599 10795
rect 39589 10761 39623 10795
rect 41429 10761 41463 10795
rect 42349 10761 42383 10795
rect 43085 10761 43119 10795
rect 43821 10761 43855 10795
rect 6101 10693 6135 10727
rect 11161 10693 11195 10727
rect 14841 10693 14875 10727
rect 15025 10693 15059 10727
rect 16037 10693 16071 10727
rect 21649 10693 21683 10727
rect 29193 10693 29227 10727
rect 30113 10693 30147 10727
rect 31769 10693 31803 10727
rect 33609 10693 33643 10727
rect 37105 10693 37139 10727
rect 38117 10693 38151 10727
rect 42717 10693 42751 10727
rect 43453 10693 43487 10727
rect 44189 10693 44223 10727
rect 30343 10659 30377 10693
rect 5089 10625 5123 10659
rect 5733 10625 5767 10659
rect 5917 10625 5951 10659
rect 6009 10625 6043 10659
rect 6193 10625 6227 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8585 10625 8619 10659
rect 10517 10625 10551 10659
rect 10701 10625 10735 10659
rect 12725 10625 12759 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 15209 10625 15243 10659
rect 16773 10625 16807 10659
rect 19533 10625 19567 10659
rect 21925 10625 21959 10659
rect 22477 10625 22511 10659
rect 25053 10625 25087 10659
rect 26341 10625 26375 10659
rect 28273 10625 28307 10659
rect 28641 10625 28675 10659
rect 29745 10625 29779 10659
rect 29837 10625 29871 10659
rect 31125 10625 31159 10659
rect 31493 10625 31527 10659
rect 33333 10625 33367 10659
rect 36001 10625 36035 10659
rect 36277 10625 36311 10659
rect 36829 10625 36863 10659
rect 37749 10625 37783 10659
rect 41981 10625 42015 10659
rect 3065 10557 3099 10591
rect 3341 10557 3375 10591
rect 4813 10557 4847 10591
rect 5181 10557 5215 10591
rect 8125 10557 8159 10591
rect 8677 10557 8711 10591
rect 8953 10557 8987 10591
rect 10885 10557 10919 10591
rect 13277 10557 13311 10591
rect 16497 10557 16531 10591
rect 17233 10557 17267 10591
rect 17509 10557 17543 10591
rect 19165 10557 19199 10591
rect 22937 10557 22971 10591
rect 23213 10557 23247 10591
rect 24685 10557 24719 10591
rect 26617 10557 26651 10591
rect 30941 10557 30975 10591
rect 31033 10557 31067 10591
rect 31217 10557 31251 10591
rect 35633 10557 35667 10591
rect 35725 10557 35759 10591
rect 36093 10557 36127 10591
rect 37841 10557 37875 10591
rect 39681 10557 39715 10591
rect 39957 10557 39991 10591
rect 5457 10489 5491 10523
rect 6745 10489 6779 10523
rect 7481 10489 7515 10523
rect 7849 10489 7883 10523
rect 16313 10489 16347 10523
rect 21281 10489 21315 10523
rect 22201 10489 22235 10523
rect 33241 10489 33275 10523
rect 35173 10489 35207 10523
rect 5089 10421 5123 10455
rect 5825 10421 5859 10455
rect 8309 10421 8343 10455
rect 10425 10421 10459 10455
rect 12817 10421 12851 10455
rect 14749 10421 14783 10455
rect 15853 10421 15887 10455
rect 16589 10421 16623 10455
rect 20913 10421 20947 10455
rect 21649 10421 21683 10455
rect 24869 10421 24903 10455
rect 26065 10421 26099 10455
rect 28089 10421 28123 10455
rect 29377 10421 29411 10455
rect 29561 10421 29595 10455
rect 30297 10421 30331 10455
rect 30481 10421 30515 10455
rect 36093 10421 36127 10455
rect 41797 10421 41831 10455
rect 44557 10421 44591 10455
rect 44833 10421 44867 10455
rect 3433 10217 3467 10251
rect 10057 10217 10091 10251
rect 10241 10217 10275 10251
rect 12265 10217 12299 10251
rect 12633 10217 12667 10251
rect 13461 10217 13495 10251
rect 14013 10217 14047 10251
rect 14289 10217 14323 10251
rect 17693 10217 17727 10251
rect 20177 10217 20211 10251
rect 20361 10217 20395 10251
rect 21281 10217 21315 10251
rect 23029 10217 23063 10251
rect 24298 10217 24332 10251
rect 28549 10217 28583 10251
rect 29009 10217 29043 10251
rect 33609 10217 33643 10251
rect 35817 10217 35851 10251
rect 35909 10217 35943 10251
rect 38853 10217 38887 10251
rect 42257 10217 42291 10251
rect 42625 10217 42659 10251
rect 42993 10217 43027 10251
rect 43729 10217 43763 10251
rect 44557 10217 44591 10251
rect 13001 10149 13035 10183
rect 19625 10149 19659 10183
rect 20453 10149 20487 10183
rect 29745 10149 29779 10183
rect 30113 10149 30147 10183
rect 37565 10149 37599 10183
rect 38577 10149 38611 10183
rect 39221 10149 39255 10183
rect 43269 10149 43303 10183
rect 44005 10149 44039 10183
rect 44925 10149 44959 10183
rect 4169 10081 4203 10115
rect 4813 10081 4847 10115
rect 6377 10081 6411 10115
rect 10701 10081 10735 10115
rect 15393 10081 15427 10115
rect 17417 10081 17451 10115
rect 19257 10081 19291 10115
rect 21005 10081 21039 10115
rect 21833 10081 21867 10115
rect 22845 10081 22879 10115
rect 23489 10081 23523 10115
rect 23857 10081 23891 10115
rect 26433 10081 26467 10115
rect 28733 10081 28767 10115
rect 30297 10081 30331 10115
rect 31033 10081 31067 10115
rect 32505 10081 32539 10115
rect 33057 10081 33091 10115
rect 33149 10081 33183 10115
rect 34345 10081 34379 10115
rect 36461 10081 36495 10115
rect 38209 10081 38243 10115
rect 39681 10081 39715 10115
rect 39773 10081 39807 10115
rect 40785 10081 40819 10115
rect 3341 10013 3375 10047
rect 3617 10013 3651 10047
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 4537 10013 4571 10047
rect 8309 10013 8343 10047
rect 10149 10013 10183 10047
rect 10425 10013 10459 10047
rect 12265 10013 12299 10047
rect 12357 10013 12391 10047
rect 13001 10013 13035 10047
rect 13277 10013 13311 10047
rect 13737 10013 13771 10047
rect 13829 10013 13863 10047
rect 14565 10013 14599 10047
rect 15117 10013 15151 10047
rect 17141 10013 17175 10047
rect 17233 10013 17267 10047
rect 17509 10013 17543 10047
rect 17877 10013 17911 10047
rect 18153 10013 18187 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 19073 10013 19107 10047
rect 19533 10013 19567 10047
rect 19809 10013 19843 10047
rect 20913 10013 20947 10047
rect 22109 10013 22143 10047
rect 22293 10013 22327 10047
rect 22569 10013 22603 10047
rect 22661 10013 22695 10047
rect 22937 10013 22971 10047
rect 23214 10013 23248 10047
rect 23305 10013 23339 10047
rect 23581 10013 23615 10047
rect 23765 10013 23799 10047
rect 24041 10013 24075 10047
rect 26065 10013 26099 10047
rect 26157 10013 26191 10047
rect 28457 10013 28491 10047
rect 29193 10013 29227 10047
rect 29469 10013 29503 10047
rect 30021 10013 30055 10047
rect 30389 10013 30423 10047
rect 30481 10013 30515 10047
rect 30573 10013 30607 10047
rect 30757 10013 30791 10047
rect 34069 10013 34103 10047
rect 36277 10013 36311 10047
rect 36921 10013 36955 10047
rect 37197 10013 37231 10047
rect 37473 10013 37507 10047
rect 38761 10013 38795 10047
rect 39037 10013 39071 10047
rect 39589 10013 39623 10047
rect 40509 10013 40543 10047
rect 6653 9945 6687 9979
rect 8585 9945 8619 9979
rect 13461 9945 13495 9979
rect 14381 9945 14415 9979
rect 20177 9945 20211 9979
rect 21649 9945 21683 9979
rect 28181 9945 28215 9979
rect 29745 9945 29779 9979
rect 29929 9945 29963 9979
rect 33425 9945 33459 9979
rect 33625 9945 33659 9979
rect 3801 9877 3835 9911
rect 4445 9877 4479 9911
rect 6285 9877 6319 9911
rect 8125 9877 8159 9911
rect 12173 9877 12207 9911
rect 13185 9877 13219 9911
rect 13645 9877 13679 9911
rect 14749 9877 14783 9911
rect 16865 9877 16899 9911
rect 16957 9877 16991 9911
rect 17969 9877 18003 9911
rect 18705 9877 18739 9911
rect 19165 9877 19199 9911
rect 20821 9877 20855 9911
rect 21741 9877 21775 9911
rect 22201 9877 22235 9911
rect 22385 9877 22419 9911
rect 28733 9877 28767 9911
rect 32597 9877 32631 9911
rect 32965 9877 32999 9911
rect 33793 9877 33827 9911
rect 36369 9877 36403 9911
rect 36737 9877 36771 9911
rect 37013 9877 37047 9911
rect 37289 9877 37323 9911
rect 37933 9877 37967 9911
rect 38025 9877 38059 9911
rect 40233 9877 40267 9911
rect 6193 9673 6227 9707
rect 9597 9673 9631 9707
rect 10149 9673 10183 9707
rect 13001 9673 13035 9707
rect 22385 9673 22419 9707
rect 22845 9673 22879 9707
rect 24409 9673 24443 9707
rect 31703 9673 31737 9707
rect 32505 9673 32539 9707
rect 32965 9673 32999 9707
rect 34161 9673 34195 9707
rect 36277 9673 36311 9707
rect 38945 9673 38979 9707
rect 40785 9673 40819 9707
rect 42993 9673 43027 9707
rect 4077 9605 4111 9639
rect 5733 9605 5767 9639
rect 6653 9605 6687 9639
rect 7389 9605 7423 9639
rect 8125 9605 8159 9639
rect 10701 9605 10735 9639
rect 11345 9605 11379 9639
rect 12449 9605 12483 9639
rect 13369 9605 13403 9639
rect 16304 9605 16338 9639
rect 17785 9605 17819 9639
rect 19809 9605 19843 9639
rect 20361 9605 20395 9639
rect 22477 9605 22511 9639
rect 24501 9605 24535 9639
rect 25605 9605 25639 9639
rect 25973 9605 26007 9639
rect 26525 9605 26559 9639
rect 30389 9605 30423 9639
rect 30589 9605 30623 9639
rect 30849 9605 30883 9639
rect 31493 9605 31527 9639
rect 33793 9605 33827 9639
rect 33993 9605 34027 9639
rect 34805 9605 34839 9639
rect 36645 9605 36679 9639
rect 36845 9605 36879 9639
rect 37381 9605 37415 9639
rect 39313 9605 39347 9639
rect 40141 9605 40175 9639
rect 42625 9605 42659 9639
rect 3801 9537 3835 9571
rect 6009 9537 6043 9571
rect 9689 9537 9723 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 10425 9537 10459 9571
rect 10517 9537 10551 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 12817 9537 12851 9571
rect 13001 9537 13035 9571
rect 13100 9537 13134 9571
rect 15485 9537 15519 9571
rect 16037 9537 16071 9571
rect 17509 9537 17543 9571
rect 19717 9537 19751 9571
rect 20637 9537 20671 9571
rect 20729 9537 20763 9571
rect 20821 9537 20855 9571
rect 21005 9537 21039 9571
rect 21465 9537 21499 9571
rect 21554 9543 21588 9577
rect 21649 9540 21683 9574
rect 31079 9571 31113 9605
rect 21833 9537 21867 9571
rect 23213 9537 23247 9571
rect 23765 9537 23799 9571
rect 24961 9537 24995 9571
rect 26985 9537 27019 9571
rect 27997 9537 28031 9571
rect 29837 9537 29871 9571
rect 30113 9537 30147 9571
rect 32413 9537 32447 9571
rect 33333 9537 33367 9571
rect 33425 9537 33459 9571
rect 37105 9537 37139 9571
rect 41153 9537 41187 9571
rect 41797 9537 41831 9571
rect 43453 9537 43487 9571
rect 5917 9469 5951 9503
rect 7849 9469 7883 9503
rect 15577 9469 15611 9503
rect 19257 9469 19291 9503
rect 19901 9469 19935 9503
rect 22569 9469 22603 9503
rect 23305 9469 23339 9503
rect 23397 9469 23431 9503
rect 24593 9469 24627 9503
rect 26709 9469 26743 9503
rect 27629 9469 27663 9503
rect 32689 9469 32723 9503
rect 33609 9469 33643 9503
rect 34529 9469 34563 9503
rect 38853 9469 38887 9503
rect 39405 9469 39439 9503
rect 39589 9469 39623 9503
rect 40233 9469 40267 9503
rect 40325 9469 40359 9503
rect 41429 9469 41463 9503
rect 41981 9469 42015 9503
rect 15117 9401 15151 9435
rect 19349 9401 19383 9435
rect 21189 9401 21223 9435
rect 30757 9401 30791 9435
rect 31217 9401 31251 9435
rect 44741 9401 44775 9435
rect 5549 9333 5583 9367
rect 5733 9333 5767 9367
rect 7021 9333 7055 9367
rect 7757 9333 7791 9367
rect 9689 9333 9723 9367
rect 11253 9333 11287 9367
rect 11713 9333 11747 9367
rect 12081 9333 12115 9367
rect 12633 9333 12667 9367
rect 14841 9333 14875 9367
rect 15853 9333 15887 9367
rect 17417 9333 17451 9367
rect 22017 9333 22051 9367
rect 23857 9333 23891 9367
rect 24041 9333 24075 9367
rect 25053 9333 25087 9367
rect 29377 9333 29411 9367
rect 29653 9333 29687 9367
rect 30573 9333 30607 9367
rect 31033 9333 31067 9367
rect 31677 9333 31711 9367
rect 31861 9333 31895 9367
rect 32045 9333 32079 9367
rect 33977 9333 34011 9367
rect 36829 9333 36863 9367
rect 37013 9333 37047 9367
rect 39773 9333 39807 9367
rect 43361 9333 43395 9367
rect 6101 9129 6135 9163
rect 6653 9129 6687 9163
rect 7757 9129 7791 9163
rect 8861 9129 8895 9163
rect 9597 9129 9631 9163
rect 11069 9129 11103 9163
rect 12909 9129 12943 9163
rect 13461 9129 13495 9163
rect 15301 9129 15335 9163
rect 21557 9129 21591 9163
rect 22661 9129 22695 9163
rect 23121 9129 23155 9163
rect 23489 9129 23523 9163
rect 24133 9129 24167 9163
rect 24777 9129 24811 9163
rect 26157 9129 26191 9163
rect 29193 9129 29227 9163
rect 29377 9129 29411 9163
rect 29732 9129 29766 9163
rect 33609 9129 33643 9163
rect 35909 9129 35943 9163
rect 36093 9129 36127 9163
rect 36369 9129 36403 9163
rect 38485 9129 38519 9163
rect 43177 9129 43211 9163
rect 43729 9129 43763 9163
rect 8585 9061 8619 9095
rect 9965 9061 9999 9095
rect 10609 9061 10643 9095
rect 13001 9061 13035 9095
rect 14197 9061 14231 9095
rect 23305 9061 23339 9095
rect 34897 9061 34931 9095
rect 36553 9061 36587 9095
rect 38577 9061 38611 9095
rect 16405 8993 16439 9027
rect 16957 8993 16991 9027
rect 19165 8993 19199 9027
rect 19257 8993 19291 9027
rect 20085 8993 20119 9027
rect 22293 8993 22327 9027
rect 23765 8993 23799 9027
rect 24409 8993 24443 9027
rect 25513 8993 25547 9027
rect 26801 8993 26835 9027
rect 31953 8993 31987 9027
rect 32689 8993 32723 9027
rect 32873 8993 32907 9027
rect 32965 8993 32999 9027
rect 34713 8993 34747 9027
rect 35541 8993 35575 9027
rect 37013 8993 37047 9027
rect 765 8925 799 8959
rect 4353 8925 4387 8959
rect 8585 8925 8619 8959
rect 8769 8925 8803 8959
rect 9045 8925 9079 8959
rect 9137 8925 9171 8959
rect 10241 8925 10275 8959
rect 11161 8925 11195 8959
rect 13277 8925 13311 8959
rect 13737 8925 13771 8959
rect 14013 8925 14047 8959
rect 16681 8925 16715 8959
rect 19533 8925 19567 8959
rect 19717 8925 19751 8959
rect 19809 8925 19843 8959
rect 22017 8925 22051 8959
rect 22109 8925 22143 8959
rect 22753 8925 22787 8959
rect 23397 8925 23431 8959
rect 25237 8925 25271 8959
rect 25329 8925 25363 8959
rect 25605 8925 25639 8959
rect 26617 8925 26651 8959
rect 28917 8925 28951 8959
rect 29469 8925 29503 8959
rect 31677 8925 31711 8959
rect 32229 8925 32263 8959
rect 32781 8925 32815 8959
rect 33517 8925 33551 8959
rect 35357 8925 35391 8959
rect 36737 8925 36771 8959
rect 38761 8925 38795 8959
rect 39037 8925 39071 8959
rect 39773 8925 39807 8959
rect 39865 8925 39899 8959
rect 8861 8891 8895 8925
rect 4629 8857 4663 8891
rect 9229 8857 9263 8891
rect 9413 8857 9447 8891
rect 9965 8857 9999 8891
rect 11437 8857 11471 8891
rect 13001 8857 13035 8891
rect 13185 8857 13219 8891
rect 13461 8857 13495 8891
rect 13645 8857 13679 8891
rect 13829 8857 13863 8891
rect 16313 8857 16347 8891
rect 19073 8857 19107 8891
rect 21649 8857 21683 8891
rect 23121 8857 23155 8891
rect 25053 8857 25087 8891
rect 26525 8857 26559 8891
rect 26985 8857 27019 8891
rect 31769 8857 31803 8891
rect 35725 8857 35759 8891
rect 35941 8857 35975 8891
rect 36185 8857 36219 8891
rect 36401 8857 36435 8891
rect 40141 8857 40175 8891
rect 41705 8857 41739 8891
rect 949 8789 983 8823
rect 6929 8789 6963 8823
rect 7297 8789 7331 8823
rect 8125 8789 8159 8823
rect 10149 8789 10183 8823
rect 14565 8789 14599 8823
rect 14933 8789 14967 8823
rect 15669 8789 15703 8823
rect 15853 8789 15887 8823
rect 16221 8789 16255 8823
rect 18429 8789 18463 8823
rect 18705 8789 18739 8823
rect 19717 8789 19751 8823
rect 24133 8789 24167 8823
rect 24317 8789 24351 8823
rect 24777 8789 24811 8823
rect 24961 8789 24995 8823
rect 25973 8789 26007 8823
rect 28457 8789 28491 8823
rect 31217 8789 31251 8823
rect 31309 8789 31343 8823
rect 32321 8789 32355 8823
rect 32505 8789 32539 8823
rect 34069 8789 34103 8823
rect 34437 8789 34471 8823
rect 34529 8789 34563 8823
rect 35265 8789 35299 8823
rect 38853 8789 38887 8823
rect 39405 8789 39439 8823
rect 39589 8789 39623 8823
rect 41613 8789 41647 8823
rect 44189 8789 44223 8823
rect 44557 8789 44591 8823
rect 44925 8789 44959 8823
rect 6009 8585 6043 8619
rect 6469 8585 6503 8619
rect 7665 8585 7699 8619
rect 8125 8585 8159 8619
rect 8769 8585 8803 8619
rect 11069 8585 11103 8619
rect 15117 8585 15151 8619
rect 17325 8585 17359 8619
rect 19165 8585 19199 8619
rect 21833 8585 21867 8619
rect 26525 8585 26559 8619
rect 27261 8585 27295 8619
rect 30113 8585 30147 8619
rect 30957 8585 30991 8619
rect 34253 8585 34287 8619
rect 34345 8585 34379 8619
rect 36369 8585 36403 8619
rect 40877 8585 40911 8619
rect 41245 8585 41279 8619
rect 9229 8517 9263 8551
rect 11345 8517 11379 8551
rect 13192 8517 13226 8551
rect 15761 8517 15795 8551
rect 17693 8517 17727 8551
rect 19533 8517 19567 8551
rect 20729 8517 20763 8551
rect 21649 8517 21683 8551
rect 22385 8517 22419 8551
rect 26433 8517 26467 8551
rect 27997 8517 28031 8551
rect 30757 8517 30791 8551
rect 31585 8517 31619 8551
rect 32781 8517 32815 8551
rect 34897 8517 34931 8551
rect 42073 8517 42107 8551
rect 10885 8449 10919 8483
rect 11161 8449 11195 8483
rect 11253 8449 11287 8483
rect 11437 8449 11471 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 12449 8449 12483 8483
rect 12633 8449 12667 8483
rect 12817 8449 12851 8483
rect 14749 8449 14783 8483
rect 16313 8449 16347 8483
rect 16497 8449 16531 8483
rect 16957 8449 16991 8483
rect 17417 8449 17451 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 20637 8449 20671 8483
rect 22293 8449 22327 8483
rect 22937 8449 22971 8483
rect 23397 8449 23431 8483
rect 23857 8449 23891 8483
rect 27353 8449 27387 8483
rect 27721 8449 27755 8483
rect 29745 8449 29779 8483
rect 30389 8449 30423 8483
rect 30573 8449 30607 8483
rect 32045 8449 32079 8483
rect 32505 8449 32539 8483
rect 34529 8449 34563 8483
rect 34621 8449 34655 8483
rect 36645 8449 36679 8483
rect 38485 8449 38519 8483
rect 40785 8449 40819 8483
rect 41429 8449 41463 8483
rect 41797 8449 41831 8483
rect 5549 8381 5583 8415
rect 6837 8381 6871 8415
rect 7389 8381 7423 8415
rect 8493 8381 8527 8415
rect 8953 8381 8987 8415
rect 12909 8381 12943 8415
rect 14841 8381 14875 8415
rect 19901 8381 19935 8415
rect 19993 8381 20027 8415
rect 20913 8381 20947 8415
rect 22477 8381 22511 8415
rect 23489 8381 23523 8415
rect 23673 8381 23707 8415
rect 24133 8381 24167 8415
rect 24409 8381 24443 8415
rect 26157 8381 26191 8415
rect 27445 8381 27479 8415
rect 30297 8381 30331 8415
rect 30481 8381 30515 8415
rect 31769 8381 31803 8415
rect 32137 8381 32171 8415
rect 32229 8381 32263 8415
rect 32321 8381 32355 8415
rect 40233 8381 40267 8415
rect 40969 8381 41003 8415
rect 43821 8381 43855 8415
rect 44189 8381 44223 8415
rect 44925 8381 44959 8415
rect 10701 8313 10735 8347
rect 11989 8313 12023 8347
rect 14657 8313 14691 8347
rect 21281 8313 21315 8347
rect 21925 8313 21959 8347
rect 22753 8313 22787 8347
rect 31125 8313 31159 8347
rect 40417 8313 40451 8347
rect 10885 8245 10919 8279
rect 11897 8245 11931 8279
rect 14933 8245 14967 8279
rect 15393 8245 15427 8279
rect 16405 8245 16439 8279
rect 16773 8245 16807 8279
rect 19349 8245 19383 8279
rect 20177 8245 20211 8279
rect 20269 8245 20303 8279
rect 21649 8245 21683 8279
rect 23029 8245 23063 8279
rect 23949 8245 23983 8279
rect 26893 8245 26927 8279
rect 30941 8245 30975 8279
rect 31861 8245 31895 8279
rect 36908 8245 36942 8279
rect 38393 8245 38427 8279
rect 38748 8245 38782 8279
rect 43545 8245 43579 8279
rect 44649 8245 44683 8279
rect 8125 8041 8159 8075
rect 8769 8041 8803 8075
rect 9965 8041 9999 8075
rect 12817 8041 12851 8075
rect 13185 8041 13219 8075
rect 15209 8041 15243 8075
rect 18245 8041 18279 8075
rect 23857 8041 23891 8075
rect 27997 8041 28031 8075
rect 31493 8041 31527 8075
rect 33885 8041 33919 8075
rect 37013 8041 37047 8075
rect 38025 8041 38059 8075
rect 38393 8041 38427 8075
rect 41521 8041 41555 8075
rect 43361 8041 43395 8075
rect 22477 7973 22511 8007
rect 22569 7973 22603 8007
rect 22845 7973 22879 8007
rect 42349 7973 42383 8007
rect 8585 7905 8619 7939
rect 10333 7905 10367 7939
rect 13093 7905 13127 7939
rect 13277 7905 13311 7939
rect 16129 7905 16163 7939
rect 16405 7905 16439 7939
rect 18613 7905 18647 7939
rect 21005 7905 21039 7939
rect 23397 7905 23431 7939
rect 24133 7905 24167 7939
rect 24409 7905 24443 7939
rect 26157 7905 26191 7939
rect 26525 7905 26559 7939
rect 28089 7905 28123 7939
rect 28365 7905 28399 7939
rect 28549 7905 28583 7939
rect 29101 7905 29135 7939
rect 29377 7905 29411 7939
rect 30021 7905 30055 7939
rect 30941 7905 30975 7939
rect 31033 7905 31067 7939
rect 32137 7905 32171 7939
rect 32413 7905 32447 7939
rect 35449 7905 35483 7939
rect 37657 7905 37691 7939
rect 41429 7905 41463 7939
rect 42073 7905 42107 7939
rect 42809 7905 42843 7939
rect 42901 7905 42935 7939
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9045 7837 9079 7871
rect 9137 7837 9171 7871
rect 9321 7837 9355 7871
rect 10057 7837 10091 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 13461 7837 13495 7871
rect 16037 7837 16071 7871
rect 18429 7837 18463 7871
rect 20729 7837 20763 7871
rect 22753 7837 22787 7871
rect 23765 7837 23799 7871
rect 26249 7837 26283 7871
rect 28273 7837 28307 7871
rect 28457 7837 28491 7871
rect 29193 7837 29227 7871
rect 29285 7837 29319 7871
rect 29745 7837 29779 7871
rect 29837 7837 29871 7871
rect 29929 7837 29963 7871
rect 30757 7837 30791 7871
rect 30849 7837 30883 7871
rect 31677 7837 31711 7871
rect 31769 7837 31803 7871
rect 31861 7837 31895 7871
rect 31954 7837 31988 7871
rect 34069 7837 34103 7871
rect 34345 7837 34379 7871
rect 35173 7837 35207 7871
rect 37381 7837 37415 7871
rect 39589 7837 39623 7871
rect 39681 7837 39715 7871
rect 41889 7837 41923 7871
rect 41981 7837 42015 7871
rect 8769 7769 8803 7803
rect 9597 7769 9631 7803
rect 9781 7769 9815 7803
rect 13737 7769 13771 7803
rect 15761 7769 15795 7803
rect 18889 7769 18923 7803
rect 20637 7769 20671 7803
rect 23213 7769 23247 7803
rect 30297 7769 30331 7803
rect 38853 7769 38887 7803
rect 39957 7769 39991 7803
rect 7757 7701 7791 7735
rect 8953 7701 8987 7735
rect 9505 7701 9539 7735
rect 11805 7701 11839 7735
rect 12265 7701 12299 7735
rect 12541 7701 12575 7735
rect 15669 7701 15703 7735
rect 15859 7701 15893 7735
rect 15945 7701 15979 7735
rect 17877 7701 17911 7735
rect 23305 7701 23339 7735
rect 28917 7701 28951 7735
rect 29561 7701 29595 7735
rect 30389 7701 30423 7735
rect 30573 7701 30607 7735
rect 36921 7701 36955 7735
rect 37473 7701 37507 7735
rect 39405 7701 39439 7735
rect 42717 7701 42751 7735
rect 43729 7701 43763 7735
rect 44189 7701 44223 7735
rect 44557 7701 44591 7735
rect 44925 7701 44959 7735
rect 7665 7497 7699 7531
rect 8493 7497 8527 7531
rect 10701 7497 10735 7531
rect 11345 7497 11379 7531
rect 11805 7497 11839 7531
rect 12081 7497 12115 7531
rect 13645 7497 13679 7531
rect 14381 7497 14415 7531
rect 17785 7497 17819 7531
rect 18429 7497 18463 7531
rect 20821 7497 20855 7531
rect 21741 7497 21775 7531
rect 24317 7497 24351 7531
rect 24409 7497 24443 7531
rect 25329 7497 25363 7531
rect 26525 7497 26559 7531
rect 28365 7497 28399 7531
rect 33333 7497 33367 7531
rect 33701 7497 33735 7531
rect 34161 7497 34195 7531
rect 35541 7497 35575 7531
rect 36001 7497 36035 7531
rect 36829 7497 36863 7531
rect 38669 7497 38703 7531
rect 40141 7497 40175 7531
rect 40601 7497 40635 7531
rect 42165 7497 42199 7531
rect 43177 7497 43211 7531
rect 44005 7497 44039 7531
rect 44649 7497 44683 7531
rect 8769 7429 8803 7463
rect 10885 7429 10919 7463
rect 15669 7429 15703 7463
rect 16313 7429 16347 7463
rect 18981 7429 19015 7463
rect 19349 7429 19383 7463
rect 21465 7429 21499 7463
rect 21649 7429 21683 7463
rect 22845 7429 22879 7463
rect 28733 7429 28767 7463
rect 31861 7429 31895 7463
rect 34989 7429 35023 7463
rect 35909 7429 35943 7463
rect 39497 7429 39531 7463
rect 40509 7429 40543 7463
rect 45017 7429 45051 7463
rect 8033 7361 8067 7395
rect 8953 7361 8987 7395
rect 11161 7361 11195 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 15117 7361 15151 7395
rect 15301 7361 15335 7395
rect 15393 7361 15427 7395
rect 15485 7361 15519 7395
rect 16037 7361 16071 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 18337 7361 18371 7395
rect 18521 7361 18555 7395
rect 19073 7361 19107 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 24593 7361 24627 7395
rect 24685 7361 24719 7395
rect 24943 7361 24977 7395
rect 26341 7361 26375 7395
rect 31585 7361 31619 7395
rect 34069 7361 34103 7395
rect 34897 7361 34931 7395
rect 37197 7361 37231 7395
rect 38025 7361 38059 7395
rect 38577 7361 38611 7395
rect 39405 7361 39439 7395
rect 40049 7361 40083 7395
rect 41245 7361 41279 7395
rect 41521 7361 41555 7395
rect 42257 7361 42291 7395
rect 9229 7293 9263 7327
rect 10977 7293 11011 7327
rect 14933 7293 14967 7327
rect 22385 7293 22419 7327
rect 22569 7293 22603 7327
rect 25697 7293 25731 7327
rect 26157 7293 26191 7327
rect 26617 7293 26651 7327
rect 26893 7293 26927 7327
rect 28457 7293 28491 7327
rect 30297 7293 30331 7327
rect 30573 7293 30607 7327
rect 34345 7293 34379 7327
rect 35173 7293 35207 7327
rect 36093 7293 36127 7327
rect 37289 7293 37323 7327
rect 37473 7293 37507 7327
rect 39589 7293 39623 7327
rect 40693 7293 40727 7327
rect 42349 7293 42383 7327
rect 13277 7225 13311 7259
rect 13921 7225 13955 7259
rect 14749 7225 14783 7259
rect 39037 7225 39071 7259
rect 10885 7157 10919 7191
rect 12541 7157 12575 7191
rect 12817 7157 12851 7191
rect 15117 7157 15151 7191
rect 15853 7157 15887 7191
rect 18245 7157 18279 7191
rect 24869 7157 24903 7191
rect 30205 7157 30239 7191
rect 34529 7157 34563 7191
rect 38117 7157 38151 7191
rect 39865 7157 39899 7191
rect 41061 7157 41095 7191
rect 41337 7157 41371 7191
rect 41797 7157 41831 7191
rect 42809 7157 42843 7191
rect 43545 7157 43579 7191
rect 44281 7157 44315 7191
rect 7021 6953 7055 6987
rect 10149 6953 10183 6987
rect 11069 6953 11103 6987
rect 11345 6953 11379 6987
rect 15104 6953 15138 6987
rect 16589 6953 16623 6987
rect 17049 6953 17083 6987
rect 17969 6953 18003 6987
rect 19533 6953 19567 6987
rect 20637 6953 20671 6987
rect 22845 6953 22879 6987
rect 26801 6953 26835 6987
rect 27997 6953 28031 6987
rect 33701 6953 33735 6987
rect 34253 6953 34287 6987
rect 34437 6953 34471 6987
rect 39484 6953 39518 6987
rect 40969 6953 41003 6987
rect 41324 6953 41358 6987
rect 43913 6953 43947 6987
rect 44557 6953 44591 6987
rect 44925 6953 44959 6987
rect 8125 6885 8159 6919
rect 9229 6885 9263 6919
rect 16681 6885 16715 6919
rect 19165 6885 19199 6919
rect 7297 6817 7331 6851
rect 9505 6817 9539 6851
rect 9965 6817 9999 6851
rect 10333 6817 10367 6851
rect 17693 6817 17727 6851
rect 21005 6817 21039 6851
rect 22753 6817 22787 6851
rect 23305 6817 23339 6851
rect 23397 6817 23431 6851
rect 24685 6817 24719 6851
rect 25145 6817 25179 6851
rect 26433 6817 26467 6851
rect 27169 6817 27203 6851
rect 28181 6817 28215 6851
rect 29193 6817 29227 6851
rect 31033 6817 31067 6851
rect 31125 6817 31159 6851
rect 31217 6817 31251 6851
rect 31769 6817 31803 6851
rect 32045 6817 32079 6851
rect 33149 6817 33183 6851
rect 33333 6817 33367 6851
rect 35357 6817 35391 6851
rect 36185 6817 36219 6851
rect 36921 6817 36955 6851
rect 37933 6817 37967 6851
rect 38669 6817 38703 6851
rect 39221 6817 39255 6851
rect 41061 6817 41095 6851
rect 42809 6817 42843 6851
rect 43361 6817 43395 6851
rect 43545 6817 43579 6851
rect 7757 6749 7791 6783
rect 10057 6749 10091 6783
rect 14841 6749 14875 6783
rect 17509 6749 17543 6783
rect 19349 6749 19383 6783
rect 19442 6749 19476 6783
rect 19809 6749 19843 6783
rect 19993 6749 20027 6783
rect 20085 6749 20119 6783
rect 20269 6749 20303 6783
rect 20821 6749 20855 6783
rect 23213 6749 23247 6783
rect 25973 6749 26007 6783
rect 27445 6749 27479 6783
rect 28365 6749 28399 6783
rect 28457 6749 28491 6783
rect 28549 6749 28583 6783
rect 28641 6749 28675 6783
rect 28917 6749 28951 6783
rect 30941 6749 30975 6783
rect 35909 6749 35943 6783
rect 36737 6749 36771 6783
rect 37473 6749 37507 6783
rect 38485 6749 38519 6783
rect 33747 6715 33781 6749
rect 12817 6681 12851 6715
rect 13921 6681 13955 6715
rect 14289 6681 14323 6715
rect 14657 6681 14691 6715
rect 17049 6681 17083 6715
rect 17325 6681 17359 6715
rect 21281 6681 21315 6715
rect 24317 6681 24351 6715
rect 25421 6681 25455 6715
rect 25697 6681 25731 6715
rect 33517 6681 33551 6715
rect 34069 6681 34103 6715
rect 34285 6681 34319 6715
rect 35173 6681 35207 6715
rect 37657 6681 37691 6715
rect 8769 6613 8803 6647
rect 10333 6613 10367 6647
rect 10609 6613 10643 6647
rect 11713 6613 11747 6647
rect 12081 6613 12115 6647
rect 12449 6613 12483 6647
rect 13185 6613 13219 6647
rect 17233 6613 17267 6647
rect 18337 6613 18371 6647
rect 18797 6613 18831 6647
rect 19993 6613 20027 6647
rect 20177 6613 20211 6647
rect 23949 6613 23983 6647
rect 25789 6613 25823 6647
rect 26157 6613 26191 6647
rect 27629 6613 27663 6647
rect 30665 6613 30699 6647
rect 30757 6613 30791 6647
rect 31677 6613 31711 6647
rect 32689 6613 32723 6647
rect 33057 6613 33091 6647
rect 33885 6613 33919 6647
rect 34713 6613 34747 6647
rect 35081 6613 35115 6647
rect 35541 6613 35575 6647
rect 36001 6613 36035 6647
rect 36369 6613 36403 6647
rect 36829 6613 36863 6647
rect 37289 6613 37323 6647
rect 38117 6613 38151 6647
rect 38577 6613 38611 6647
rect 42901 6613 42935 6647
rect 43269 6613 43303 6647
rect 16405 6409 16439 6443
rect 18061 6409 18095 6443
rect 18521 6409 18555 6443
rect 21373 6409 21407 6443
rect 21557 6409 21591 6443
rect 24133 6409 24167 6443
rect 25145 6409 25179 6443
rect 25697 6409 25731 6443
rect 27721 6409 27755 6443
rect 28181 6409 28215 6443
rect 28549 6409 28583 6443
rect 29009 6409 29043 6443
rect 31309 6409 31343 6443
rect 36093 6409 36127 6443
rect 38853 6409 38887 6443
rect 40693 6409 40727 6443
rect 41245 6409 41279 6443
rect 41797 6409 41831 6443
rect 42257 6409 42291 6443
rect 43085 6409 43119 6443
rect 43637 6409 43671 6443
rect 44373 6409 44407 6443
rect 44741 6409 44775 6443
rect 7665 6341 7699 6375
rect 8125 6341 8159 6375
rect 9505 6341 9539 6375
rect 10609 6341 10643 6375
rect 17141 6341 17175 6375
rect 22661 6341 22695 6375
rect 25329 6341 25363 6375
rect 25605 6341 25639 6375
rect 26433 6341 26467 6375
rect 29837 6341 29871 6375
rect 33609 6341 33643 6375
rect 37381 6341 37415 6375
rect 42165 6341 42199 6375
rect 7021 6273 7055 6307
rect 9229 6273 9263 6307
rect 16037 6273 16071 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 16773 6273 16807 6307
rect 16865 6273 16899 6307
rect 16957 6273 16991 6307
rect 17233 6273 17267 6307
rect 20453 6273 20487 6307
rect 20637 6273 20671 6307
rect 21189 6273 21223 6307
rect 21741 6273 21775 6307
rect 22385 6273 22419 6307
rect 25513 6273 25547 6307
rect 26617 6273 26651 6307
rect 26893 6273 26927 6307
rect 28089 6273 28123 6307
rect 28917 6273 28951 6307
rect 29561 6273 29595 6307
rect 31677 6273 31711 6307
rect 36369 6273 36403 6307
rect 37013 6273 37047 6307
rect 38945 6273 38979 6307
rect 41153 6273 41187 6307
rect 42993 6273 43027 6307
rect 5273 6205 5307 6239
rect 6653 6205 6687 6239
rect 14105 6205 14139 6239
rect 14381 6205 14415 6239
rect 16129 6205 16163 6239
rect 17141 6205 17175 6239
rect 17509 6205 17543 6239
rect 18613 6205 18647 6239
rect 18889 6205 18923 6239
rect 26801 6205 26835 6239
rect 27077 6205 27111 6239
rect 28365 6205 28399 6239
rect 29101 6205 29135 6239
rect 31953 6205 31987 6239
rect 34345 6205 34379 6239
rect 34621 6205 34655 6239
rect 37105 6205 37139 6239
rect 39221 6205 39255 6239
rect 41337 6205 41371 6239
rect 42349 6205 42383 6239
rect 43269 6205 43303 6239
rect 8401 6137 8435 6171
rect 8769 6137 8803 6171
rect 9873 6137 9907 6171
rect 12449 6137 12483 6171
rect 12817 6137 12851 6171
rect 13645 6137 13679 6171
rect 16497 6137 16531 6171
rect 17325 6137 17359 6171
rect 20361 6137 20395 6171
rect 26709 6137 26743 6171
rect 27353 6137 27387 6171
rect 40785 6137 40819 6171
rect 42625 6137 42659 6171
rect 7297 6069 7331 6103
rect 10333 6069 10367 6103
rect 11345 6069 11379 6103
rect 11713 6069 11747 6103
rect 12081 6069 12115 6103
rect 13277 6069 13311 6103
rect 14013 6069 14047 6103
rect 15853 6069 15887 6103
rect 16221 6069 16255 6103
rect 17417 6069 17451 6103
rect 20821 6069 20855 6103
rect 22201 6069 22235 6103
rect 24501 6069 24535 6103
rect 24869 6069 24903 6103
rect 25881 6069 25915 6103
rect 27537 6069 27571 6103
rect 33425 6069 33459 6103
rect 33701 6069 33735 6103
rect 36185 6069 36219 6103
rect 36829 6069 36863 6103
rect 44005 6069 44039 6103
rect 45109 6069 45143 6103
rect 1685 5865 1719 5899
rect 4537 5865 4571 5899
rect 6745 5865 6779 5899
rect 8769 5865 8803 5899
rect 9229 5865 9263 5899
rect 13185 5865 13219 5899
rect 14841 5865 14875 5899
rect 16037 5865 16071 5899
rect 17693 5865 17727 5899
rect 21281 5865 21315 5899
rect 21373 5865 21407 5899
rect 24225 5865 24259 5899
rect 25145 5865 25179 5899
rect 27169 5865 27203 5899
rect 28089 5865 28123 5899
rect 32505 5865 32539 5899
rect 33241 5865 33275 5899
rect 34897 5865 34931 5899
rect 37013 5865 37047 5899
rect 38117 5865 38151 5899
rect 42809 5865 42843 5899
rect 43453 5865 43487 5899
rect 43821 5865 43855 5899
rect 44557 5865 44591 5899
rect 44925 5865 44959 5899
rect 6377 5797 6411 5831
rect 10701 5797 10735 5831
rect 14105 5797 14139 5831
rect 17877 5797 17911 5831
rect 17969 5797 18003 5831
rect 18613 5797 18647 5831
rect 30665 5797 30699 5831
rect 5089 5729 5123 5763
rect 5825 5729 5859 5763
rect 14657 5729 14691 5763
rect 19533 5729 19567 5763
rect 19809 5729 19843 5763
rect 21465 5729 21499 5763
rect 23857 5729 23891 5763
rect 25421 5729 25455 5763
rect 28917 5729 28951 5763
rect 30757 5729 30791 5763
rect 31033 5729 31067 5763
rect 33057 5729 33091 5763
rect 33421 5729 33455 5763
rect 34069 5729 34103 5763
rect 34529 5729 34563 5763
rect 35541 5729 35575 5763
rect 37749 5729 37783 5763
rect 38669 5729 38703 5763
rect 41337 5729 41371 5763
rect 2973 5661 3007 5695
rect 10333 5661 10367 5695
rect 12909 5661 12943 5695
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 15117 5671 15151 5705
rect 15393 5661 15427 5695
rect 16405 5661 16439 5695
rect 16589 5661 16623 5695
rect 16681 5661 16715 5695
rect 16865 5661 16899 5695
rect 17141 5661 17175 5695
rect 17417 5661 17451 5695
rect 17509 5661 17543 5695
rect 17693 5661 17727 5695
rect 18245 5661 18279 5695
rect 18797 5661 18831 5695
rect 18889 5661 18923 5695
rect 18981 5661 19015 5695
rect 19165 5661 19199 5695
rect 19441 5661 19475 5695
rect 21373 5661 21407 5695
rect 22385 5661 22419 5695
rect 22661 5661 22695 5695
rect 23213 5661 23247 5695
rect 23397 5661 23431 5695
rect 23949 5661 23983 5695
rect 24317 5661 24351 5695
rect 24685 5661 24719 5695
rect 24961 5661 24995 5695
rect 25145 5661 25179 5695
rect 27353 5661 27387 5695
rect 27629 5661 27663 5695
rect 32781 5661 32815 5695
rect 32873 5661 32907 5695
rect 32965 5661 32999 5695
rect 33506 5661 33540 5695
rect 33609 5661 33643 5695
rect 33701 5661 33735 5695
rect 34253 5661 34287 5695
rect 34345 5661 34379 5695
rect 34437 5661 34471 5695
rect 35081 5661 35115 5695
rect 35265 5661 35299 5695
rect 37473 5661 37507 5695
rect 39221 5661 39255 5695
rect 41061 5661 41095 5695
rect 7481 5593 7515 5627
rect 9597 5593 9631 5627
rect 14473 5593 14507 5627
rect 14841 5593 14875 5627
rect 15227 5593 15261 5627
rect 15669 5593 15703 5627
rect 15853 5593 15887 5627
rect 16773 5593 16807 5627
rect 17969 5593 18003 5627
rect 18613 5593 18647 5627
rect 23029 5593 23063 5627
rect 25697 5593 25731 5627
rect 27537 5593 27571 5627
rect 27905 5593 27939 5627
rect 28110 5593 28144 5627
rect 28549 5593 28583 5627
rect 29193 5593 29227 5627
rect 37565 5593 37599 5627
rect 39497 5593 39531 5627
rect 1317 5525 1351 5559
rect 3341 5525 3375 5559
rect 3985 5525 4019 5559
rect 5457 5525 5491 5559
rect 7113 5525 7147 5559
rect 8125 5525 8159 5559
rect 9965 5525 9999 5559
rect 11069 5525 11103 5559
rect 11437 5525 11471 5559
rect 11805 5525 11839 5559
rect 12173 5525 12207 5559
rect 12541 5525 12575 5559
rect 13737 5525 13771 5559
rect 15025 5525 15059 5559
rect 15577 5525 15611 5559
rect 16497 5525 16531 5559
rect 16957 5525 16991 5559
rect 17325 5525 17359 5559
rect 18153 5525 18187 5559
rect 19349 5525 19383 5559
rect 21741 5525 21775 5559
rect 22477 5525 22511 5559
rect 23305 5525 23339 5559
rect 23581 5525 23615 5559
rect 24501 5525 24535 5559
rect 25329 5525 25363 5559
rect 28273 5525 28307 5559
rect 28641 5525 28675 5559
rect 32597 5525 32631 5559
rect 37105 5525 37139 5559
rect 38485 5525 38519 5559
rect 38577 5525 38611 5559
rect 40969 5525 41003 5559
rect 43085 5525 43119 5559
rect 2329 5321 2363 5355
rect 3433 5321 3467 5355
rect 4261 5321 4295 5355
rect 4721 5321 4755 5355
rect 5089 5321 5123 5355
rect 6285 5321 6319 5355
rect 7297 5321 7331 5355
rect 8033 5321 8067 5355
rect 8769 5321 8803 5355
rect 9965 5321 9999 5355
rect 10701 5321 10735 5355
rect 18613 5321 18647 5355
rect 25605 5321 25639 5355
rect 29101 5321 29135 5355
rect 29561 5321 29595 5355
rect 29929 5321 29963 5355
rect 30389 5321 30423 5355
rect 33793 5321 33827 5355
rect 36461 5321 36495 5355
rect 39497 5321 39531 5355
rect 40049 5321 40083 5355
rect 41429 5321 41463 5355
rect 42349 5321 42383 5355
rect 43085 5321 43119 5355
rect 43453 5321 43487 5355
rect 43821 5321 43855 5355
rect 44557 5321 44591 5355
rect 9137 5253 9171 5287
rect 11529 5253 11563 5287
rect 11897 5253 11931 5287
rect 14381 5253 14415 5287
rect 16037 5253 16071 5287
rect 16587 5253 16621 5287
rect 17141 5253 17175 5287
rect 18889 5253 18923 5287
rect 19441 5253 19475 5287
rect 22109 5253 22143 5287
rect 24593 5253 24627 5287
rect 28135 5253 28169 5287
rect 28825 5253 28859 5287
rect 31769 5253 31803 5287
rect 33701 5253 33735 5287
rect 42809 5253 42843 5287
rect 1869 5185 1903 5219
rect 4537 5185 4571 5219
rect 5181 5185 5215 5219
rect 6377 5185 6411 5219
rect 12265 5185 12299 5219
rect 12909 5185 12943 5219
rect 13645 5185 13679 5219
rect 14105 5185 14139 5219
rect 16221 5185 16255 5219
rect 16313 5185 16347 5219
rect 16405 5185 16439 5219
rect 18705 5185 18739 5219
rect 21741 5185 21775 5219
rect 22937 5185 22971 5219
rect 23305 5185 23339 5219
rect 23673 5185 23707 5219
rect 23765 5185 23799 5219
rect 24133 5185 24167 5219
rect 24961 5185 24995 5219
rect 25329 5185 25363 5219
rect 25789 5185 25823 5219
rect 26341 5185 26375 5219
rect 26709 5185 26743 5219
rect 28273 5185 28307 5219
rect 28365 5185 28399 5219
rect 29469 5185 29503 5219
rect 30297 5185 30331 5219
rect 31033 5185 31067 5219
rect 31217 5185 31251 5219
rect 31493 5185 31527 5219
rect 34621 5185 34655 5219
rect 36829 5185 36863 5219
rect 37749 5185 37783 5219
rect 39957 5185 39991 5219
rect 40785 5185 40819 5219
rect 2421 5117 2455 5151
rect 2605 5117 2639 5151
rect 5273 5117 5307 5151
rect 6561 5117 6595 5151
rect 10333 5117 10367 5151
rect 15853 5117 15887 5151
rect 16773 5117 16807 5151
rect 16865 5117 16899 5151
rect 19165 5117 19199 5151
rect 22477 5117 22511 5151
rect 22845 5117 22879 5151
rect 24869 5117 24903 5151
rect 29009 5117 29043 5151
rect 29653 5117 29687 5151
rect 30481 5117 30515 5151
rect 30941 5117 30975 5151
rect 31125 5117 31159 5151
rect 33977 5117 34011 5151
rect 34713 5117 34747 5151
rect 34989 5117 35023 5151
rect 37473 5117 37507 5151
rect 38025 5117 38059 5151
rect 40141 5117 40175 5151
rect 40877 5117 40911 5151
rect 40969 5117 41003 5151
rect 1961 5049 1995 5083
rect 7021 5049 7055 5083
rect 11253 5049 11287 5083
rect 13277 5049 13311 5083
rect 14013 5049 14047 5083
rect 28641 5049 28675 5083
rect 36645 5049 36679 5083
rect 40417 5049 40451 5083
rect 44925 5049 44959 5083
rect 1133 4981 1167 5015
rect 1501 4981 1535 5015
rect 1685 4981 1719 5015
rect 3065 4981 3099 5015
rect 3893 4981 3927 5015
rect 4353 4981 4387 5015
rect 5917 4981 5951 5015
rect 7757 4981 7791 5015
rect 8493 4981 8527 5015
rect 9505 4981 9539 5015
rect 12081 4981 12115 5015
rect 16037 4981 16071 5015
rect 19073 4981 19107 5015
rect 20913 4981 20947 5015
rect 23213 4981 23247 5015
rect 23489 4981 23523 5015
rect 24133 4981 24167 5015
rect 24317 4981 24351 5015
rect 25237 4981 25271 5015
rect 25513 4981 25547 5015
rect 26065 4981 26099 5015
rect 28273 4981 28307 5015
rect 30757 4981 30791 5015
rect 33241 4981 33275 5015
rect 33333 4981 33367 5015
rect 34437 4981 34471 5015
rect 37105 4981 37139 5015
rect 39589 4981 39623 5015
rect 41981 4981 42015 5015
rect 44189 4981 44223 5015
rect 3157 4777 3191 4811
rect 11621 4777 11655 4811
rect 12541 4777 12575 4811
rect 14013 4777 14047 4811
rect 15853 4777 15887 4811
rect 18337 4777 18371 4811
rect 19441 4777 19475 4811
rect 19717 4777 19751 4811
rect 20729 4777 20763 4811
rect 21465 4777 21499 4811
rect 23765 4777 23799 4811
rect 25421 4777 25455 4811
rect 33793 4777 33827 4811
rect 36737 4777 36771 4811
rect 38209 4777 38243 4811
rect 38669 4777 38703 4811
rect 38853 4777 38887 4811
rect 41797 4777 41831 4811
rect 42257 4777 42291 4811
rect 42901 4777 42935 4811
rect 44557 4777 44591 4811
rect 9505 4709 9539 4743
rect 10057 4709 10091 4743
rect 15945 4709 15979 4743
rect 18153 4709 18187 4743
rect 19993 4709 20027 4743
rect 24777 4709 24811 4743
rect 30021 4709 30055 4743
rect 35909 4709 35943 4743
rect 41153 4709 41187 4743
rect 43269 4709 43303 4743
rect 43637 4709 43671 4743
rect 44005 4709 44039 4743
rect 1501 4641 1535 4675
rect 3801 4641 3835 4675
rect 4813 4641 4847 4675
rect 8125 4641 8159 4675
rect 8953 4641 8987 4675
rect 10609 4641 10643 4675
rect 12265 4641 12299 4675
rect 13093 4641 13127 4675
rect 21097 4641 21131 4675
rect 22109 4641 22143 4675
rect 24317 4641 24351 4675
rect 25053 4641 25087 4675
rect 27537 4641 27571 4675
rect 28273 4641 28307 4675
rect 30665 4641 30699 4675
rect 31493 4641 31527 4675
rect 32045 4641 32079 4675
rect 32321 4641 32355 4675
rect 34345 4641 34379 4675
rect 36369 4641 36403 4675
rect 36553 4641 36587 4675
rect 37289 4641 37323 4675
rect 39773 4641 39807 4675
rect 40601 4641 40635 4675
rect 44925 4641 44959 4675
rect 1133 4573 1167 4607
rect 1225 4573 1259 4607
rect 3525 4573 3559 4607
rect 4537 4573 4571 4607
rect 4997 4573 5031 4607
rect 7297 4573 7331 4607
rect 8677 4573 8711 4607
rect 9781 4573 9815 4607
rect 14105 4573 14139 4607
rect 16129 4573 16163 4607
rect 16221 4573 16255 4607
rect 16405 4573 16439 4607
rect 18245 4573 18279 4607
rect 18429 4573 18463 4607
rect 19625 4573 19659 4607
rect 19809 4573 19843 4607
rect 19901 4573 19935 4607
rect 20085 4573 20119 4607
rect 21741 4573 21775 4607
rect 21833 4573 21867 4607
rect 25145 4573 25179 4607
rect 25513 4573 25547 4607
rect 25789 4573 25823 4607
rect 27721 4573 27755 4607
rect 27813 4573 27847 4607
rect 28135 4573 28169 4607
rect 28917 4573 28951 4607
rect 29101 4573 29135 4607
rect 29285 4573 29319 4607
rect 34069 4573 34103 4607
rect 36277 4573 36311 4607
rect 37105 4573 37139 4607
rect 38393 4573 38427 4607
rect 39037 4573 39071 4607
rect 39589 4573 39623 4607
rect 40417 4573 40451 4607
rect 3617 4505 3651 4539
rect 5273 4505 5307 4539
rect 8769 4505 8803 4539
rect 14381 4505 14415 4539
rect 15945 4505 15979 4539
rect 16681 4505 16715 4539
rect 24225 4505 24259 4539
rect 26065 4505 26099 4539
rect 29009 4505 29043 4539
rect 29837 4505 29871 4539
rect 30481 4505 30515 4539
rect 30573 4505 30607 4539
rect 37749 4505 37783 4539
rect 39681 4505 39715 4539
rect 41521 4505 41555 4539
rect 42533 4505 42567 4539
rect 949 4437 983 4471
rect 2973 4437 3007 4471
rect 4169 4437 4203 4471
rect 4629 4437 4663 4471
rect 6745 4437 6779 4471
rect 7113 4437 7147 4471
rect 7757 4437 7791 4471
rect 8309 4437 8343 4471
rect 9597 4437 9631 4471
rect 10425 4437 10459 4471
rect 10517 4437 10551 4471
rect 11253 4437 11287 4471
rect 11713 4437 11747 4471
rect 12081 4437 12115 4471
rect 12173 4437 12207 4471
rect 12909 4437 12943 4471
rect 13001 4437 13035 4471
rect 19073 4437 19107 4471
rect 21557 4437 21591 4471
rect 23581 4437 23615 4471
rect 24133 4437 24167 4471
rect 25697 4437 25731 4471
rect 28549 4437 28583 4471
rect 29377 4437 29411 4471
rect 30113 4437 30147 4471
rect 30941 4437 30975 4471
rect 31309 4437 31343 4471
rect 31401 4437 31435 4471
rect 35817 4437 35851 4471
rect 37197 4437 37231 4471
rect 39221 4437 39255 4471
rect 40049 4437 40083 4471
rect 40509 4437 40543 4471
rect 5733 4233 5767 4267
rect 14105 4233 14139 4267
rect 15025 4233 15059 4267
rect 23121 4233 23155 4267
rect 24317 4233 24351 4267
rect 31033 4233 31067 4267
rect 39865 4233 39899 4267
rect 40417 4233 40451 4267
rect 41245 4233 41279 4267
rect 41981 4233 42015 4267
rect 43085 4233 43119 4267
rect 43453 4233 43487 4267
rect 43913 4233 43947 4267
rect 44557 4233 44591 4267
rect 44925 4233 44959 4267
rect 4077 4165 4111 4199
rect 9229 4165 9263 4199
rect 11805 4165 11839 4199
rect 20177 4165 20211 4199
rect 25329 4165 25363 4199
rect 27471 4165 27505 4199
rect 27721 4165 27755 4199
rect 27937 4165 27971 4199
rect 29009 4165 29043 4199
rect 30757 4165 30791 4199
rect 31677 4165 31711 4199
rect 33241 4165 33275 4199
rect 33793 4165 33827 4199
rect 41153 4165 41187 4199
rect 42349 4165 42383 4199
rect 42717 4165 42751 4199
rect 44189 4165 44223 4199
rect 1225 4097 1259 4131
rect 5917 4097 5951 4131
rect 6469 4097 6503 4131
rect 6561 4097 6595 4131
rect 8861 4097 8895 4131
rect 8953 4097 8987 4131
rect 11437 4097 11471 4131
rect 13553 4097 13587 4131
rect 14197 4097 14231 4131
rect 14933 4097 14967 4131
rect 15117 4097 15151 4131
rect 15853 4097 15887 4131
rect 16405 4097 16439 4131
rect 19257 4097 19291 4131
rect 20269 4097 20303 4131
rect 21005 4097 21039 4131
rect 21281 4097 21315 4131
rect 23489 4097 23523 4131
rect 24593 4097 24627 4131
rect 25053 4097 25087 4131
rect 25697 4097 25731 4131
rect 25789 4097 25823 4131
rect 26525 4097 26559 4131
rect 26709 4097 26743 4131
rect 26801 4097 26835 4131
rect 27169 4097 27203 4131
rect 27261 4097 27295 4131
rect 27353 4097 27387 4131
rect 28457 4097 28491 4131
rect 28825 4097 28859 4131
rect 29285 4097 29319 4131
rect 29745 4097 29779 4131
rect 29837 4097 29871 4131
rect 30113 4097 30147 4131
rect 30205 4097 30239 4131
rect 31217 4097 31251 4131
rect 32229 4097 32263 4131
rect 33333 4097 33367 4131
rect 36185 4097 36219 4131
rect 38117 4097 38151 4131
rect 40325 4097 40359 4131
rect 1501 4029 1535 4063
rect 3617 4029 3651 4063
rect 3801 4029 3835 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 11161 4029 11195 4063
rect 11529 4029 11563 4063
rect 14289 4029 14323 4063
rect 16313 4029 16347 4063
rect 16681 4029 16715 4063
rect 18153 4029 18187 4063
rect 19073 4029 19107 4063
rect 19533 4029 19567 4063
rect 20361 4029 20395 4063
rect 21557 4029 21591 4063
rect 23581 4029 23615 4063
rect 23765 4029 23799 4063
rect 24869 4029 24903 4063
rect 26341 4029 26375 4063
rect 26985 4029 27019 4063
rect 27629 4029 27663 4063
rect 28733 4029 28767 4063
rect 29193 4029 29227 4063
rect 30297 4029 30331 4063
rect 31953 4029 31987 4063
rect 33517 4029 33551 4063
rect 34161 4029 34195 4063
rect 34437 4029 34471 4063
rect 37197 4029 37231 4063
rect 38393 4029 38427 4063
rect 40509 4029 40543 4063
rect 41337 4029 41371 4063
rect 3341 3961 3375 3995
rect 13737 3961 13771 3995
rect 18705 3961 18739 3995
rect 25237 3961 25271 3995
rect 28089 3961 28123 3995
rect 28273 3961 28307 3995
rect 31861 3961 31895 3995
rect 32873 3961 32907 3995
rect 33977 3961 34011 3995
rect 36829 3961 36863 3995
rect 40785 3961 40819 3995
rect 1133 3893 1167 3927
rect 2973 3893 3007 3927
rect 8309 3893 8343 3927
rect 8677 3893 8711 3927
rect 10701 3893 10735 3927
rect 11253 3893 11287 3927
rect 13277 3893 13311 3927
rect 13369 3893 13403 3927
rect 14841 3893 14875 3927
rect 15485 3893 15519 3927
rect 19809 3893 19843 3927
rect 23029 3893 23063 3927
rect 24869 3893 24903 3927
rect 25421 3893 25455 3927
rect 25973 3893 26007 3927
rect 27905 3893 27939 3927
rect 28641 3893 28675 3927
rect 29377 3893 29411 3927
rect 29561 3893 29595 3927
rect 30021 3893 30055 3927
rect 30389 3893 30423 3927
rect 30573 3893 30607 3927
rect 30849 3893 30883 3927
rect 35909 3893 35943 3927
rect 37565 3893 37599 3927
rect 37933 3893 37967 3927
rect 39957 3893 39991 3927
rect 5089 3689 5123 3723
rect 5549 3689 5583 3723
rect 5917 3689 5951 3723
rect 8033 3689 8067 3723
rect 10149 3689 10183 3723
rect 13093 3689 13127 3723
rect 14841 3689 14875 3723
rect 27445 3689 27479 3723
rect 28089 3689 28123 3723
rect 31125 3689 31159 3723
rect 32413 3689 32447 3723
rect 34253 3689 34287 3723
rect 34713 3689 34747 3723
rect 38485 3689 38519 3723
rect 40969 3689 41003 3723
rect 41705 3689 41739 3723
rect 42717 3689 42751 3723
rect 43085 3689 43119 3723
rect 43913 3689 43947 3723
rect 44925 3689 44959 3723
rect 1501 3621 1535 3655
rect 2605 3621 2639 3655
rect 30941 3621 30975 3655
rect 41245 3621 41279 3655
rect 42073 3621 42107 3655
rect 42441 3621 42475 3655
rect 43453 3621 43487 3655
rect 44649 3621 44683 3655
rect 2973 3553 3007 3587
rect 3341 3553 3375 3587
rect 7389 3553 7423 3587
rect 10701 3553 10735 3587
rect 11621 3553 11655 3587
rect 14105 3553 14139 3587
rect 17417 3553 17451 3587
rect 18061 3553 18095 3587
rect 19349 3553 19383 3587
rect 20177 3553 20211 3587
rect 22661 3553 22695 3587
rect 22753 3553 22787 3587
rect 24317 3553 24351 3587
rect 25605 3553 25639 3587
rect 26433 3553 26467 3587
rect 28181 3553 28215 3587
rect 29193 3553 29227 3587
rect 29469 3553 29503 3587
rect 32873 3553 32907 3587
rect 33057 3553 33091 3587
rect 35541 3553 35575 3587
rect 35725 3553 35759 3587
rect 36369 3553 36403 3587
rect 36553 3553 36587 3587
rect 37381 3553 37415 3587
rect 38209 3553 38243 3587
rect 1133 3485 1167 3519
rect 1869 3485 1903 3519
rect 6193 3485 6227 3519
rect 6561 3485 6595 3519
rect 7113 3485 7147 3519
rect 8309 3485 8343 3519
rect 10517 3485 10551 3519
rect 11345 3485 11379 3519
rect 13921 3485 13955 3519
rect 15025 3485 15059 3519
rect 17233 3485 17267 3519
rect 17785 3485 17819 3519
rect 18429 3485 18463 3519
rect 19073 3485 19107 3519
rect 19901 3485 19935 3519
rect 20361 3485 20395 3519
rect 23213 3485 23247 3519
rect 23581 3485 23615 3519
rect 24133 3485 24167 3519
rect 24869 3485 24903 3519
rect 26249 3485 26283 3519
rect 26709 3485 26743 3519
rect 27905 3485 27939 3519
rect 27997 3485 28031 3519
rect 28457 3485 28491 3519
rect 28549 3485 28583 3519
rect 28733 3485 28767 3519
rect 28917 3485 28951 3519
rect 29101 3485 29135 3519
rect 31131 3485 31165 3519
rect 31309 3485 31343 3519
rect 31539 3485 31573 3519
rect 31861 3485 31895 3519
rect 32137 3485 32171 3519
rect 32321 3485 32355 3519
rect 33425 3485 33459 3519
rect 34621 3485 34655 3519
rect 34897 3485 34931 3519
rect 38669 3485 38703 3519
rect 39037 3485 39071 3519
rect 39221 3485 39255 3519
rect 3617 3417 3651 3451
rect 8585 3417 8619 3451
rect 15301 3417 15335 3451
rect 17325 3417 17359 3451
rect 19165 3417 19199 3451
rect 20637 3417 20671 3451
rect 22569 3417 22603 3451
rect 26985 3417 27019 3451
rect 27261 3417 27295 3451
rect 27477 3417 27511 3451
rect 31677 3417 31711 3451
rect 31769 3417 31803 3451
rect 33701 3417 33735 3451
rect 35449 3417 35483 3451
rect 37197 3417 37231 3451
rect 39497 3417 39531 3451
rect 2237 3349 2271 3383
rect 6377 3349 6411 3383
rect 6745 3349 6779 3383
rect 7205 3349 7239 3383
rect 10057 3349 10091 3383
rect 10609 3349 10643 3383
rect 11253 3349 11287 3383
rect 13553 3349 13587 3383
rect 14013 3349 14047 3383
rect 16773 3349 16807 3383
rect 16865 3349 16899 3383
rect 18245 3349 18279 3383
rect 18705 3349 18739 3383
rect 19533 3349 19567 3383
rect 19993 3349 20027 3383
rect 22109 3349 22143 3383
rect 22201 3349 22235 3383
rect 23029 3349 23063 3383
rect 23765 3349 23799 3383
rect 24225 3349 24259 3383
rect 24685 3349 24719 3383
rect 25053 3349 25087 3383
rect 25421 3349 25455 3383
rect 25513 3349 25547 3383
rect 25881 3349 25915 3383
rect 26341 3349 26375 3383
rect 27629 3349 27663 3383
rect 28273 3349 28307 3383
rect 28641 3349 28675 3383
rect 29009 3349 29043 3383
rect 32045 3349 32079 3383
rect 32321 3349 32355 3383
rect 32781 3349 32815 3383
rect 33241 3349 33275 3383
rect 34437 3349 34471 3383
rect 35081 3349 35115 3383
rect 35909 3349 35943 3383
rect 36277 3349 36311 3383
rect 36829 3349 36863 3383
rect 37289 3349 37323 3383
rect 37657 3349 37691 3383
rect 38025 3349 38059 3383
rect 38117 3349 38151 3383
rect 38853 3349 38887 3383
rect 949 3145 983 3179
rect 4445 3145 4479 3179
rect 5549 3145 5583 3179
rect 7665 3145 7699 3179
rect 8401 3145 8435 3179
rect 10425 3145 10459 3179
rect 14473 3145 14507 3179
rect 15669 3145 15703 3179
rect 20821 3145 20855 3179
rect 25881 3145 25915 3179
rect 26065 3145 26099 3179
rect 29653 3145 29687 3179
rect 29745 3145 29779 3179
rect 33609 3145 33643 3179
rect 34989 3145 35023 3179
rect 35357 3145 35391 3179
rect 40233 3145 40267 3179
rect 41981 3145 42015 3179
rect 42717 3145 42751 3179
rect 43085 3145 43119 3179
rect 44741 3145 44775 3179
rect 3985 3077 4019 3111
rect 6193 3077 6227 3111
rect 11437 3077 11471 3111
rect 17325 3077 17359 3111
rect 19165 3077 19199 3111
rect 21465 3077 21499 3111
rect 23765 3077 23799 3111
rect 24409 3077 24443 3111
rect 28917 3077 28951 3111
rect 31953 3077 31987 3111
rect 34529 3077 34563 3111
rect 35449 3077 35483 3111
rect 41337 3077 41371 3111
rect 42349 3077 42383 3111
rect 765 3009 799 3043
rect 1501 3009 1535 3043
rect 4629 3009 4663 3043
rect 5181 3009 5215 3043
rect 5917 3009 5951 3043
rect 8585 3009 8619 3043
rect 11345 3009 11379 3043
rect 12633 3009 12667 3043
rect 15025 3009 15059 3043
rect 15853 3009 15887 3043
rect 16405 3009 16439 3043
rect 17049 3009 17083 3043
rect 21005 3009 21039 3043
rect 23213 3009 23247 3043
rect 23673 3009 23707 3043
rect 24133 3009 24167 3043
rect 25973 3009 26007 3043
rect 26157 3009 26191 3043
rect 26525 3009 26559 3043
rect 28733 3009 28767 3043
rect 30021 3009 30055 3043
rect 30113 3009 30147 3043
rect 30205 3009 30239 3043
rect 30389 3009 30423 3043
rect 30665 3009 30699 3043
rect 33517 3009 33551 3043
rect 33701 3009 33735 3043
rect 34069 3009 34103 3043
rect 34621 3009 34655 3043
rect 36001 3009 36035 3043
rect 36461 3009 36495 3043
rect 38485 3009 38519 3043
rect 40693 3009 40727 3043
rect 43453 3009 43487 3043
rect 1777 2941 1811 2975
rect 4077 2941 4111 2975
rect 4169 2941 4203 2975
rect 8677 2941 8711 2975
rect 8953 2941 8987 2975
rect 11529 2941 11563 2975
rect 12725 2941 12759 2975
rect 13001 2941 13035 2975
rect 16497 2941 16531 2975
rect 16589 2941 16623 2975
rect 18889 2941 18923 2975
rect 20637 2941 20671 2975
rect 21189 2941 21223 2975
rect 23857 2941 23891 2975
rect 26617 2941 26651 2975
rect 26893 2941 26927 2975
rect 29377 2941 29411 2975
rect 29469 2941 29503 2975
rect 30757 2941 30791 2975
rect 31677 2941 31711 2975
rect 34805 2941 34839 2975
rect 35541 2941 35575 2975
rect 36645 2941 36679 2975
rect 36921 2941 36955 2975
rect 38761 2941 38795 2975
rect 40785 2941 40819 2975
rect 40877 2941 40911 2975
rect 8309 2873 8343 2907
rect 16037 2873 16071 2907
rect 18797 2873 18831 2907
rect 23305 2873 23339 2907
rect 28917 2873 28951 2907
rect 34161 2873 34195 2907
rect 36277 2873 36311 2907
rect 38393 2873 38427 2907
rect 40325 2873 40359 2907
rect 1409 2805 1443 2839
rect 3249 2805 3283 2839
rect 3617 2805 3651 2839
rect 10977 2805 11011 2839
rect 12357 2805 12391 2839
rect 12449 2805 12483 2839
rect 14841 2805 14875 2839
rect 15393 2805 15427 2839
rect 22937 2805 22971 2839
rect 23029 2805 23063 2839
rect 26341 2805 26375 2839
rect 28365 2805 28399 2839
rect 28549 2805 28583 2839
rect 30665 2805 30699 2839
rect 31033 2805 31067 2839
rect 33425 2805 33459 2839
rect 33885 2805 33919 2839
rect 35817 2805 35851 2839
rect 1501 2601 1535 2635
rect 1961 2601 1995 2635
rect 9137 2601 9171 2635
rect 11805 2601 11839 2635
rect 12173 2601 12207 2635
rect 13277 2601 13311 2635
rect 16037 2601 16071 2635
rect 19441 2601 19475 2635
rect 23581 2601 23615 2635
rect 27353 2601 27387 2635
rect 27537 2601 27571 2635
rect 28273 2601 28307 2635
rect 29745 2601 29779 2635
rect 30757 2601 30791 2635
rect 35817 2601 35851 2635
rect 37657 2601 37691 2635
rect 38853 2601 38887 2635
rect 42349 2601 42383 2635
rect 43085 2601 43119 2635
rect 43361 2601 43395 2635
rect 43729 2601 43763 2635
rect 44189 2601 44223 2635
rect 45017 2601 45051 2635
rect 1593 2533 1627 2567
rect 7021 2533 7055 2567
rect 12909 2533 12943 2567
rect 27813 2533 27847 2567
rect 29377 2533 29411 2567
rect 29469 2533 29503 2567
rect 30113 2533 30147 2567
rect 38577 2533 38611 2567
rect 39221 2533 39255 2567
rect 41981 2533 42015 2567
rect 42625 2533 42659 2567
rect 2789 2465 2823 2499
rect 3157 2465 3191 2499
rect 5457 2465 5491 2499
rect 9689 2465 9723 2499
rect 14289 2465 14323 2499
rect 16497 2465 16531 2499
rect 16681 2465 16715 2499
rect 18429 2465 18463 2499
rect 19073 2465 19107 2499
rect 19257 2465 19291 2499
rect 19901 2465 19935 2499
rect 21833 2465 21867 2499
rect 25605 2465 25639 2499
rect 25881 2465 25915 2499
rect 27721 2465 27755 2499
rect 28733 2465 28767 2499
rect 30021 2465 30055 2499
rect 31217 2465 31251 2499
rect 31401 2465 31435 2499
rect 31861 2465 31895 2499
rect 34345 2465 34379 2499
rect 36185 2465 36219 2499
rect 38209 2465 38243 2499
rect 38301 2465 38335 2499
rect 39681 2465 39715 2499
rect 39773 2465 39807 2499
rect 40601 2465 40635 2499
rect 41429 2465 41463 2499
rect 44557 2465 44591 2499
rect 1777 2397 1811 2431
rect 2145 2397 2179 2431
rect 2605 2397 2639 2431
rect 2697 2397 2731 2431
rect 7205 2397 7239 2431
rect 9505 2397 9539 2431
rect 9597 2397 9631 2431
rect 10057 2397 10091 2431
rect 13921 2397 13955 2431
rect 19625 2397 19659 2431
rect 23765 2397 23799 2431
rect 27445 2397 27479 2431
rect 27997 2397 28031 2431
rect 28457 2397 28491 2431
rect 28641 2397 28675 2431
rect 29101 2397 29135 2431
rect 29285 2397 29319 2431
rect 29561 2397 29595 2431
rect 29929 2397 29963 2431
rect 30205 2397 30239 2431
rect 30389 2397 30423 2431
rect 31585 2397 31619 2431
rect 33701 2397 33735 2431
rect 34069 2397 34103 2431
rect 35909 2397 35943 2431
rect 38761 2397 38795 2431
rect 39037 2397 39071 2431
rect 39589 2397 39623 2431
rect 40417 2397 40451 2431
rect 3433 2329 3467 2363
rect 6929 2329 6963 2363
rect 9045 2329 9079 2363
rect 10333 2329 10367 2363
rect 12449 2329 12483 2363
rect 14565 2329 14599 2363
rect 16957 2329 16991 2363
rect 18981 2329 19015 2363
rect 20177 2329 20211 2363
rect 22109 2329 22143 2363
rect 24041 2329 24075 2363
rect 27721 2329 27755 2363
rect 31125 2329 31159 2363
rect 38117 2329 38151 2363
rect 40509 2329 40543 2363
rect 41337 2329 41371 2363
rect 1133 2261 1167 2295
rect 2237 2261 2271 2295
rect 4905 2261 4939 2295
rect 5733 2261 5767 2295
rect 6101 2261 6135 2295
rect 6561 2261 6595 2295
rect 7757 2261 7791 2295
rect 8125 2261 8159 2295
rect 8585 2261 8619 2295
rect 13737 2261 13771 2295
rect 18613 2261 18647 2295
rect 21649 2261 21683 2295
rect 25513 2261 25547 2295
rect 30573 2261 30607 2295
rect 33333 2261 33367 2295
rect 33517 2261 33551 2295
rect 37749 2261 37783 2295
rect 40049 2261 40083 2295
rect 40877 2261 40911 2295
rect 41245 2261 41279 2295
rect 1685 2057 1719 2091
rect 2053 2057 2087 2091
rect 3341 2057 3375 2091
rect 4445 2057 4479 2091
rect 10149 2057 10183 2091
rect 10885 2057 10919 2091
rect 11897 2057 11931 2091
rect 14289 2057 14323 2091
rect 17785 2057 17819 2091
rect 19257 2057 19291 2091
rect 19625 2057 19659 2091
rect 20453 2057 20487 2091
rect 21189 2057 21223 2091
rect 21649 2057 21683 2091
rect 22477 2057 22511 2091
rect 25145 2057 25179 2091
rect 29929 2057 29963 2091
rect 31125 2057 31159 2091
rect 35725 2057 35759 2091
rect 36093 2057 36127 2091
rect 40601 2057 40635 2091
rect 40693 2057 40727 2091
rect 42073 2057 42107 2091
rect 42717 2057 42751 2091
rect 43821 2057 43855 2091
rect 44189 2057 44223 2091
rect 44557 2057 44591 2091
rect 44925 2057 44959 2091
rect 12817 1989 12851 2023
rect 16865 1989 16899 2023
rect 23029 1989 23063 2023
rect 34161 1989 34195 2023
rect 41521 1989 41555 2023
rect 42441 1989 42475 2023
rect 43085 1989 43119 2023
rect 43453 1989 43487 2023
rect 2329 1921 2363 1955
rect 2881 1921 2915 1955
rect 3525 1921 3559 1955
rect 3985 1921 4019 1955
rect 4721 1921 4755 1955
rect 5365 1921 5399 1955
rect 6377 1921 6411 1955
rect 7941 1921 7975 1955
rect 9137 1921 9171 1955
rect 9873 1921 9907 1955
rect 10517 1921 10551 1955
rect 11069 1921 11103 1955
rect 11345 1921 11379 1955
rect 12173 1921 12207 1955
rect 12449 1921 12483 1955
rect 12541 1921 12575 1955
rect 14565 1921 14599 1955
rect 15577 1921 15611 1955
rect 16405 1921 16439 1955
rect 17233 1921 17267 1955
rect 17417 1921 17451 1955
rect 17969 1921 18003 1955
rect 18521 1921 18555 1955
rect 18889 1921 18923 1955
rect 19901 1921 19935 1955
rect 20361 1921 20395 1955
rect 20637 1921 20671 1955
rect 21005 1921 21039 1955
rect 21557 1921 21591 1955
rect 22385 1921 22419 1955
rect 22661 1921 22695 1955
rect 22753 1921 22787 1955
rect 24685 1921 24719 1955
rect 25329 1921 25363 1955
rect 25421 1921 25455 1955
rect 25605 1921 25639 1955
rect 26065 1921 26099 1955
rect 26341 1921 26375 1955
rect 28181 1921 28215 1955
rect 30021 1921 30055 1955
rect 30573 1921 30607 1955
rect 31309 1921 31343 1955
rect 31493 1921 31527 1955
rect 31953 1921 31987 1955
rect 36645 1921 36679 1955
rect 38669 1921 38703 1955
rect 38853 1921 38887 1955
rect 40877 1921 40911 1955
rect 41153 1921 41187 1955
rect 3249 1853 3283 1887
rect 5089 1853 5123 1887
rect 6101 1853 6135 1887
rect 6929 1853 6963 1887
rect 7665 1853 7699 1887
rect 8493 1853 8527 1887
rect 8861 1853 8895 1887
rect 15209 1853 15243 1887
rect 18245 1853 18279 1887
rect 21833 1853 21867 1887
rect 26617 1853 26651 1887
rect 28457 1853 28491 1887
rect 31033 1853 31067 1887
rect 32229 1853 32263 1887
rect 33885 1853 33919 1887
rect 35633 1853 35667 1887
rect 36185 1853 36219 1887
rect 36369 1853 36403 1887
rect 39129 1853 39163 1887
rect 7297 1785 7331 1819
rect 9597 1785 9631 1819
rect 24869 1785 24903 1819
rect 25789 1785 25823 1819
rect 38393 1785 38427 1819
rect 38485 1785 38519 1819
rect 40969 1785 41003 1819
rect 1225 1717 1259 1751
rect 2145 1717 2179 1751
rect 2697 1717 2731 1751
rect 3801 1717 3835 1751
rect 4537 1717 4571 1751
rect 5181 1717 5215 1751
rect 6193 1717 6227 1751
rect 7757 1717 7791 1751
rect 8953 1717 8987 1751
rect 9689 1717 9723 1751
rect 10333 1717 10367 1751
rect 11161 1717 11195 1751
rect 11989 1717 12023 1751
rect 12265 1717 12299 1751
rect 14381 1717 14415 1751
rect 14933 1717 14967 1751
rect 15393 1717 15427 1751
rect 16221 1717 16255 1751
rect 17601 1717 17635 1751
rect 18337 1717 18371 1751
rect 18705 1717 18739 1751
rect 19717 1717 19751 1751
rect 20177 1717 20211 1751
rect 20821 1717 20855 1751
rect 22201 1717 22235 1751
rect 24501 1717 24535 1751
rect 25881 1717 25915 1751
rect 28089 1717 28123 1751
rect 30113 1717 30147 1751
rect 30481 1717 30515 1751
rect 30757 1717 30791 1751
rect 31677 1717 31711 1751
rect 33701 1717 33735 1751
rect 36908 1717 36942 1751
rect 3341 1513 3375 1547
rect 5181 1513 5215 1547
rect 6009 1513 6043 1547
rect 6929 1513 6963 1547
rect 7665 1513 7699 1547
rect 9229 1513 9263 1547
rect 11069 1513 11103 1547
rect 15209 1513 15243 1547
rect 16681 1513 16715 1547
rect 17693 1513 17727 1547
rect 17969 1513 18003 1547
rect 19349 1513 19383 1547
rect 25973 1513 26007 1547
rect 26525 1513 26559 1547
rect 27077 1513 27111 1547
rect 27813 1513 27847 1547
rect 28641 1513 28675 1547
rect 29193 1513 29227 1547
rect 29653 1513 29687 1547
rect 29929 1513 29963 1547
rect 30389 1513 30423 1547
rect 32689 1513 32723 1547
rect 40049 1513 40083 1547
rect 40601 1513 40635 1547
rect 41153 1513 41187 1547
rect 42993 1513 43027 1547
rect 43913 1513 43947 1547
rect 1041 1445 1075 1479
rect 1869 1445 1903 1479
rect 2973 1445 3007 1479
rect 11713 1445 11747 1479
rect 12541 1445 12575 1479
rect 15853 1445 15887 1479
rect 31125 1445 31159 1479
rect 32045 1445 32079 1479
rect 33149 1445 33183 1479
rect 36185 1445 36219 1479
rect 40325 1445 40359 1479
rect 24501 1377 24535 1411
rect 31585 1377 31619 1411
rect 33425 1377 33459 1411
rect 33609 1377 33643 1411
rect 35357 1377 35391 1411
rect 37289 1377 37323 1411
rect 37565 1377 37599 1411
rect 39865 1377 39899 1411
rect 1133 1309 1167 1343
rect 1961 1309 1995 1343
rect 3249 1309 3283 1343
rect 3709 1309 3743 1343
rect 4445 1309 4479 1343
rect 5273 1309 5307 1343
rect 6101 1309 6135 1343
rect 6837 1309 6871 1343
rect 7757 1309 7791 1343
rect 8585 1309 8619 1343
rect 9413 1309 9447 1343
rect 10241 1309 10275 1343
rect 10977 1309 11011 1343
rect 11897 1309 11931 1343
rect 12725 1309 12759 1343
rect 13553 1309 13587 1343
rect 14381 1309 14415 1343
rect 15117 1309 15151 1343
rect 16037 1309 16071 1343
rect 16865 1309 16899 1343
rect 18613 1309 18647 1343
rect 19257 1309 19291 1343
rect 20177 1309 20211 1343
rect 21189 1309 21223 1343
rect 21741 1309 21775 1343
rect 21833 1309 21867 1343
rect 22569 1309 22603 1343
rect 22661 1309 22695 1343
rect 23949 1309 23983 1343
rect 24225 1309 24259 1343
rect 26433 1309 26467 1343
rect 26985 1309 27019 1343
rect 27721 1309 27755 1343
rect 28181 1309 28215 1343
rect 28549 1309 28583 1343
rect 28733 1309 28767 1343
rect 28917 1309 28951 1343
rect 29469 1309 29503 1343
rect 30757 1309 30791 1343
rect 31309 1309 31343 1343
rect 31677 1309 31711 1343
rect 32137 1309 32171 1343
rect 32505 1309 32539 1343
rect 33333 1309 33367 1343
rect 33885 1309 33919 1343
rect 34253 1309 34287 1343
rect 34529 1309 34563 1343
rect 35173 1309 35207 1343
rect 35265 1309 35299 1343
rect 35817 1309 35851 1343
rect 36093 1309 36127 1343
rect 36369 1309 36403 1343
rect 36829 1309 36863 1343
rect 37105 1309 37139 1343
rect 39589 1309 39623 1343
rect 39681 1309 39715 1343
rect 40233 1309 40267 1343
rect 40509 1309 40543 1343
rect 40785 1309 40819 1343
rect 41061 1309 41095 1343
rect 41337 1309 41371 1343
rect 41613 1309 41647 1343
rect 41981 1309 42015 1343
rect 42257 1309 42291 1343
rect 42717 1309 42751 1343
rect 43545 1309 43579 1343
rect 44557 1309 44591 1343
rect 44833 1309 44867 1343
rect 45201 1309 45235 1343
rect 2605 1241 2639 1275
rect 4261 1241 4295 1275
rect 10149 1241 10183 1275
rect 20913 1241 20947 1275
rect 23213 1241 23247 1275
rect 30297 1241 30331 1275
rect 32321 1241 32355 1275
rect 32413 1241 32447 1275
rect 32855 1241 32889 1275
rect 1317 1173 1351 1207
rect 2145 1173 2179 1207
rect 3893 1173 3927 1207
rect 4629 1173 4663 1207
rect 5457 1173 5491 1207
rect 6285 1173 6319 1207
rect 7941 1173 7975 1207
rect 8769 1173 8803 1207
rect 9597 1173 9631 1207
rect 10425 1173 10459 1207
rect 12081 1173 12115 1207
rect 12909 1173 12943 1207
rect 13737 1173 13771 1207
rect 14197 1173 14231 1207
rect 14565 1173 14599 1207
rect 16221 1173 16255 1207
rect 17049 1173 17083 1207
rect 18337 1173 18371 1207
rect 18797 1173 18831 1207
rect 20085 1173 20119 1207
rect 20361 1173 20395 1207
rect 21373 1173 21407 1207
rect 21557 1173 21591 1207
rect 22017 1173 22051 1207
rect 22385 1173 22419 1207
rect 22845 1173 22879 1207
rect 23305 1173 23339 1207
rect 23765 1173 23799 1207
rect 28365 1173 28399 1207
rect 29377 1173 29411 1207
rect 30941 1173 30975 1207
rect 33609 1173 33643 1207
rect 33701 1173 33735 1207
rect 34069 1173 34103 1207
rect 34345 1173 34379 1207
rect 34805 1173 34839 1207
rect 35633 1173 35667 1207
rect 35909 1173 35943 1207
rect 36645 1173 36679 1207
rect 36921 1173 36955 1207
rect 39037 1173 39071 1207
rect 39221 1173 39255 1207
rect 40877 1173 40911 1207
rect 41429 1173 41463 1207
rect 41797 1173 41831 1207
rect 42073 1173 42107 1207
rect 42533 1173 42567 1207
rect 43361 1173 43395 1207
rect 44373 1173 44407 1207
rect 45017 1173 45051 1207
<< metal1 >>
rect 17954 23508 17960 23520
rect 12406 23480 17960 23508
rect 11698 23264 11704 23316
rect 11756 23304 11762 23316
rect 12406 23304 12434 23480
rect 17954 23468 17960 23480
rect 18012 23468 18018 23520
rect 22830 23440 22836 23452
rect 11756 23276 12434 23304
rect 12544 23412 22836 23440
rect 11756 23264 11762 23276
rect 12544 23236 12572 23412
rect 22830 23400 22836 23412
rect 22888 23400 22894 23452
rect 14918 23332 14924 23384
rect 14976 23372 14982 23384
rect 23474 23372 23480 23384
rect 14976 23344 23480 23372
rect 14976 23332 14982 23344
rect 23474 23332 23480 23344
rect 23532 23332 23538 23384
rect 15102 23264 15108 23316
rect 15160 23304 15166 23316
rect 24026 23304 24032 23316
rect 15160 23276 24032 23304
rect 15160 23264 15166 23276
rect 24026 23264 24032 23276
rect 24084 23264 24090 23316
rect 8266 23208 12572 23236
rect 5994 22992 6000 23044
rect 6052 23032 6058 23044
rect 8266 23032 8294 23208
rect 14550 23196 14556 23248
rect 14608 23236 14614 23248
rect 22370 23236 22376 23248
rect 14608 23208 22376 23236
rect 14608 23196 14614 23208
rect 22370 23196 22376 23208
rect 22428 23196 22434 23248
rect 27430 23196 27436 23248
rect 27488 23236 27494 23248
rect 27488 23208 28304 23236
rect 27488 23196 27494 23208
rect 23290 23128 23296 23180
rect 23348 23168 23354 23180
rect 28166 23168 28172 23180
rect 23348 23140 28172 23168
rect 23348 23128 23354 23140
rect 28166 23128 28172 23140
rect 28224 23128 28230 23180
rect 28276 23168 28304 23208
rect 31294 23196 31300 23248
rect 31352 23236 31358 23248
rect 33594 23236 33600 23248
rect 31352 23208 33600 23236
rect 31352 23196 31358 23208
rect 33594 23196 33600 23208
rect 33652 23196 33658 23248
rect 34054 23196 34060 23248
rect 34112 23236 34118 23248
rect 35066 23236 35072 23248
rect 34112 23208 35072 23236
rect 34112 23196 34118 23208
rect 35066 23196 35072 23208
rect 35124 23196 35130 23248
rect 28276 23140 41000 23168
rect 12710 23060 12716 23112
rect 12768 23100 12774 23112
rect 22278 23100 22284 23112
rect 12768 23072 22284 23100
rect 12768 23060 12774 23072
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 28074 23060 28080 23112
rect 28132 23100 28138 23112
rect 32858 23100 32864 23112
rect 28132 23072 32864 23100
rect 28132 23060 28138 23072
rect 32858 23060 32864 23072
rect 32916 23100 32922 23112
rect 34606 23100 34612 23112
rect 32916 23072 34612 23100
rect 32916 23060 32922 23072
rect 34606 23060 34612 23072
rect 34664 23060 34670 23112
rect 40972 23044 41000 23140
rect 6052 23004 8294 23032
rect 6052 22992 6058 23004
rect 13630 22992 13636 23044
rect 13688 23032 13694 23044
rect 24854 23032 24860 23044
rect 13688 23004 24860 23032
rect 13688 22992 13694 23004
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 27890 22992 27896 23044
rect 27948 23032 27954 23044
rect 33410 23032 33416 23044
rect 27948 23004 33416 23032
rect 27948 22992 27954 23004
rect 33410 22992 33416 23004
rect 33468 22992 33474 23044
rect 40954 22992 40960 23044
rect 41012 22992 41018 23044
rect 8294 22924 8300 22976
rect 8352 22964 8358 22976
rect 30650 22964 30656 22976
rect 8352 22936 30656 22964
rect 8352 22924 8358 22936
rect 30650 22924 30656 22936
rect 30708 22924 30714 22976
rect 32398 22924 32404 22976
rect 32456 22964 32462 22976
rect 42794 22964 42800 22976
rect 32456 22936 42800 22964
rect 32456 22924 32462 22936
rect 42794 22924 42800 22936
rect 42852 22924 42858 22976
rect 460 22874 45540 22896
rect 460 22822 6070 22874
rect 6122 22822 6134 22874
rect 6186 22822 6198 22874
rect 6250 22822 6262 22874
rect 6314 22822 6326 22874
rect 6378 22822 11070 22874
rect 11122 22822 11134 22874
rect 11186 22822 11198 22874
rect 11250 22822 11262 22874
rect 11314 22822 11326 22874
rect 11378 22822 16070 22874
rect 16122 22822 16134 22874
rect 16186 22822 16198 22874
rect 16250 22822 16262 22874
rect 16314 22822 16326 22874
rect 16378 22822 21070 22874
rect 21122 22822 21134 22874
rect 21186 22822 21198 22874
rect 21250 22822 21262 22874
rect 21314 22822 21326 22874
rect 21378 22822 26070 22874
rect 26122 22822 26134 22874
rect 26186 22822 26198 22874
rect 26250 22822 26262 22874
rect 26314 22822 26326 22874
rect 26378 22822 31070 22874
rect 31122 22822 31134 22874
rect 31186 22822 31198 22874
rect 31250 22822 31262 22874
rect 31314 22822 31326 22874
rect 31378 22822 36070 22874
rect 36122 22822 36134 22874
rect 36186 22822 36198 22874
rect 36250 22822 36262 22874
rect 36314 22822 36326 22874
rect 36378 22822 41070 22874
rect 41122 22822 41134 22874
rect 41186 22822 41198 22874
rect 41250 22822 41262 22874
rect 41314 22822 41326 22874
rect 41378 22822 45540 22874
rect 460 22800 45540 22822
rect 842 22720 848 22772
rect 900 22760 906 22772
rect 1121 22763 1179 22769
rect 1121 22760 1133 22763
rect 900 22732 1133 22760
rect 900 22720 906 22732
rect 1121 22729 1133 22732
rect 1167 22729 1179 22763
rect 1121 22723 1179 22729
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1820 22732 2053 22760
rect 1820 22720 1826 22732
rect 2041 22729 2053 22732
rect 2087 22729 2099 22763
rect 2041 22723 2099 22729
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3329 22763 3387 22769
rect 3329 22760 3341 22763
rect 2832 22732 3341 22760
rect 2832 22720 2838 22732
rect 3329 22729 3341 22732
rect 3375 22729 3387 22763
rect 3329 22723 3387 22729
rect 3602 22720 3608 22772
rect 3660 22760 3666 22772
rect 3881 22763 3939 22769
rect 3881 22760 3893 22763
rect 3660 22732 3893 22760
rect 3660 22720 3666 22732
rect 3881 22729 3893 22732
rect 3927 22729 3939 22763
rect 3881 22723 3939 22729
rect 4522 22720 4528 22772
rect 4580 22760 4586 22772
rect 4801 22763 4859 22769
rect 4801 22760 4813 22763
rect 4580 22732 4813 22760
rect 4580 22720 4586 22732
rect 4801 22729 4813 22732
rect 4847 22729 4859 22763
rect 4801 22723 4859 22729
rect 5442 22720 5448 22772
rect 5500 22760 5506 22772
rect 5905 22763 5963 22769
rect 5905 22760 5917 22763
rect 5500 22732 5917 22760
rect 5500 22720 5506 22732
rect 5905 22729 5917 22732
rect 5951 22729 5963 22763
rect 5905 22723 5963 22729
rect 6454 22720 6460 22772
rect 6512 22760 6518 22772
rect 6641 22763 6699 22769
rect 6641 22760 6653 22763
rect 6512 22732 6653 22760
rect 6512 22720 6518 22732
rect 6641 22729 6653 22732
rect 6687 22729 6699 22763
rect 6641 22723 6699 22729
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7561 22763 7619 22769
rect 7561 22760 7573 22763
rect 7340 22732 7573 22760
rect 7340 22720 7346 22732
rect 7561 22729 7573 22732
rect 7607 22729 7619 22763
rect 7561 22723 7619 22729
rect 8202 22720 8208 22772
rect 8260 22760 8266 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 8260 22732 8493 22760
rect 8260 22720 8266 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 8481 22723 8539 22729
rect 9122 22720 9128 22772
rect 9180 22760 9186 22772
rect 9401 22763 9459 22769
rect 9401 22760 9413 22763
rect 9180 22732 9413 22760
rect 9180 22720 9186 22732
rect 9401 22729 9413 22732
rect 9447 22729 9459 22763
rect 9401 22723 9459 22729
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 10321 22763 10379 22769
rect 10321 22760 10333 22763
rect 10100 22732 10333 22760
rect 10100 22720 10106 22732
rect 10321 22729 10333 22732
rect 10367 22729 10379 22763
rect 10321 22723 10379 22729
rect 10962 22720 10968 22772
rect 11020 22760 11026 22772
rect 11241 22763 11299 22769
rect 11241 22760 11253 22763
rect 11020 22732 11253 22760
rect 11020 22720 11026 22732
rect 11241 22729 11253 22732
rect 11287 22729 11299 22763
rect 11241 22723 11299 22729
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 12161 22763 12219 22769
rect 12161 22760 12173 22763
rect 11940 22732 12173 22760
rect 11940 22720 11946 22732
rect 12161 22729 12173 22732
rect 12207 22729 12219 22763
rect 12161 22723 12219 22729
rect 12802 22720 12808 22772
rect 12860 22760 12866 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12860 22732 13093 22760
rect 12860 22720 12866 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13630 22720 13636 22772
rect 13688 22720 13694 22772
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 14001 22763 14059 22769
rect 14001 22760 14013 22763
rect 13872 22732 14013 22760
rect 13872 22720 13878 22732
rect 14001 22729 14013 22732
rect 14047 22729 14059 22763
rect 14001 22723 14059 22729
rect 14550 22720 14556 22772
rect 14608 22720 14614 22772
rect 14642 22720 14648 22772
rect 14700 22760 14706 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14700 22732 14933 22760
rect 14700 22720 14706 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 14921 22723 14979 22729
rect 15102 22720 15108 22772
rect 15160 22720 15166 22772
rect 15197 22763 15255 22769
rect 15197 22729 15209 22763
rect 15243 22729 15255 22763
rect 15197 22723 15255 22729
rect 1946 22652 1952 22704
rect 2004 22692 2010 22704
rect 15120 22692 15148 22720
rect 2004 22664 15148 22692
rect 15212 22692 15240 22723
rect 15562 22720 15568 22772
rect 15620 22760 15626 22772
rect 16209 22763 16267 22769
rect 16209 22760 16221 22763
rect 15620 22732 16221 22760
rect 15620 22720 15626 22732
rect 16209 22729 16221 22732
rect 16255 22729 16267 22763
rect 16209 22723 16267 22729
rect 16482 22720 16488 22772
rect 16540 22760 16546 22772
rect 16577 22763 16635 22769
rect 16577 22760 16589 22763
rect 16540 22732 16589 22760
rect 16540 22720 16546 22732
rect 16577 22729 16589 22732
rect 16623 22729 16635 22763
rect 16577 22723 16635 22729
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 17460 22732 17693 22760
rect 17460 22720 17466 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 17681 22723 17739 22729
rect 18322 22720 18328 22772
rect 18380 22760 18386 22772
rect 18785 22763 18843 22769
rect 18785 22760 18797 22763
rect 18380 22732 18797 22760
rect 18380 22720 18386 22732
rect 18785 22729 18797 22732
rect 18831 22729 18843 22763
rect 18785 22723 18843 22729
rect 19242 22720 19248 22772
rect 19300 22760 19306 22772
rect 19337 22763 19395 22769
rect 19337 22760 19349 22763
rect 19300 22732 19349 22760
rect 19300 22720 19306 22732
rect 19337 22729 19349 22732
rect 19383 22729 19395 22763
rect 19337 22723 19395 22729
rect 20162 22720 20168 22772
rect 20220 22760 20226 22772
rect 20441 22763 20499 22769
rect 20441 22760 20453 22763
rect 20220 22732 20453 22760
rect 20220 22720 20226 22732
rect 20441 22729 20453 22732
rect 20487 22729 20499 22763
rect 20441 22723 20499 22729
rect 20990 22720 20996 22772
rect 21048 22760 21054 22772
rect 21361 22763 21419 22769
rect 21361 22760 21373 22763
rect 21048 22732 21373 22760
rect 21048 22720 21054 22732
rect 21361 22729 21373 22732
rect 21407 22729 21419 22763
rect 21361 22723 21419 22729
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22729 21603 22763
rect 21545 22723 21603 22729
rect 15212 22664 16068 22692
rect 2004 22652 2010 22664
rect 934 22584 940 22636
rect 992 22584 998 22636
rect 1854 22584 1860 22636
rect 1912 22584 1918 22636
rect 3234 22584 3240 22636
rect 3292 22584 3298 22636
rect 3697 22627 3755 22633
rect 3697 22593 3709 22627
rect 3743 22624 3755 22627
rect 3970 22624 3976 22636
rect 3743 22596 3976 22624
rect 3743 22593 3755 22596
rect 3697 22587 3755 22593
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 4614 22584 4620 22636
rect 4672 22584 4678 22636
rect 5810 22584 5816 22636
rect 5868 22584 5874 22636
rect 6454 22584 6460 22636
rect 6512 22584 6518 22636
rect 7374 22584 7380 22636
rect 7432 22584 7438 22636
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22624 8171 22627
rect 8294 22624 8300 22636
rect 8159 22596 8300 22624
rect 8159 22593 8171 22596
rect 8113 22587 8171 22593
rect 8294 22584 8300 22596
rect 8352 22584 8358 22636
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 9214 22584 9220 22636
rect 9272 22584 9278 22636
rect 10134 22584 10140 22636
rect 10192 22584 10198 22636
rect 11146 22584 11152 22636
rect 11204 22584 11210 22636
rect 11698 22584 11704 22636
rect 11756 22584 11762 22636
rect 11974 22584 11980 22636
rect 12032 22584 12038 22636
rect 12894 22584 12900 22636
rect 12952 22584 12958 22636
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13909 22627 13967 22633
rect 13909 22624 13921 22627
rect 13504 22596 13921 22624
rect 13504 22584 13510 22596
rect 13909 22593 13921 22596
rect 13955 22593 13967 22627
rect 13909 22587 13967 22593
rect 14734 22584 14740 22636
rect 14792 22584 14798 22636
rect 15378 22584 15384 22636
rect 15436 22584 15442 22636
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15654 22584 15660 22636
rect 15712 22584 15718 22636
rect 16040 22633 16068 22664
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22593 16083 22627
rect 16025 22587 16083 22593
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 16758 22624 16764 22636
rect 16531 22596 16764 22624
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 17494 22584 17500 22636
rect 17552 22584 17558 22636
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18601 22627 18659 22633
rect 18601 22624 18613 22627
rect 18288 22596 18613 22624
rect 18288 22584 18294 22596
rect 18601 22593 18613 22596
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 19245 22627 19303 22633
rect 19245 22593 19257 22627
rect 19291 22624 19303 22627
rect 19702 22624 19708 22636
rect 19291 22596 19708 22624
rect 19291 22593 19303 22596
rect 19245 22587 19303 22593
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 20254 22584 20260 22636
rect 20312 22584 20318 22636
rect 21177 22627 21235 22633
rect 21177 22593 21189 22627
rect 21223 22624 21235 22627
rect 21560 22624 21588 22723
rect 22002 22720 22008 22772
rect 22060 22760 22066 22772
rect 22281 22763 22339 22769
rect 22281 22760 22293 22763
rect 22060 22732 22293 22760
rect 22060 22720 22066 22732
rect 22281 22729 22293 22732
rect 22327 22729 22339 22763
rect 22281 22723 22339 22729
rect 22922 22720 22928 22772
rect 22980 22760 22986 22772
rect 23201 22763 23259 22769
rect 23201 22760 23213 22763
rect 22980 22732 23213 22760
rect 22980 22720 22986 22732
rect 23201 22729 23213 22732
rect 23247 22729 23259 22763
rect 23201 22723 23259 22729
rect 23842 22720 23848 22772
rect 23900 22760 23906 22772
rect 24121 22763 24179 22769
rect 24121 22760 24133 22763
rect 23900 22732 24133 22760
rect 23900 22720 23906 22732
rect 24121 22729 24133 22732
rect 24167 22729 24179 22763
rect 24121 22723 24179 22729
rect 24762 22720 24768 22772
rect 24820 22760 24826 22772
rect 24857 22763 24915 22769
rect 24857 22760 24869 22763
rect 24820 22732 24869 22760
rect 24820 22720 24826 22732
rect 24857 22729 24869 22732
rect 24903 22729 24915 22763
rect 24857 22723 24915 22729
rect 25409 22763 25467 22769
rect 25409 22729 25421 22763
rect 25455 22729 25467 22763
rect 25409 22723 25467 22729
rect 25424 22692 25452 22723
rect 25682 22720 25688 22772
rect 25740 22760 25746 22772
rect 25961 22763 26019 22769
rect 25961 22760 25973 22763
rect 25740 22732 25973 22760
rect 25740 22720 25746 22732
rect 25961 22729 25973 22732
rect 26007 22729 26019 22763
rect 25961 22723 26019 22729
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 26881 22763 26939 22769
rect 26881 22760 26893 22763
rect 26660 22732 26893 22760
rect 26660 22720 26666 22732
rect 26881 22729 26893 22732
rect 26927 22729 26939 22763
rect 26881 22723 26939 22729
rect 27065 22763 27123 22769
rect 27065 22729 27077 22763
rect 27111 22729 27123 22763
rect 27065 22723 27123 22729
rect 25424 22664 25820 22692
rect 21223 22596 21588 22624
rect 21737 22631 21795 22637
rect 21737 22597 21749 22631
rect 21783 22624 21795 22631
rect 21783 22597 21864 22624
rect 21737 22596 21864 22597
rect 21223 22593 21235 22596
rect 21177 22587 21235 22593
rect 21737 22591 21795 22596
rect 3050 22516 3056 22568
rect 3108 22556 3114 22568
rect 11716 22556 11744 22584
rect 3108 22528 11744 22556
rect 3108 22516 3114 22528
rect 12802 22516 12808 22568
rect 12860 22516 12866 22568
rect 17126 22516 17132 22568
rect 17184 22556 17190 22568
rect 21836 22556 21864 22596
rect 22186 22584 22192 22636
rect 22244 22584 22250 22636
rect 23014 22584 23020 22636
rect 23072 22584 23078 22636
rect 23106 22584 23112 22636
rect 23164 22624 23170 22636
rect 23937 22627 23995 22633
rect 23937 22624 23949 22627
rect 23164 22596 23949 22624
rect 23164 22584 23170 22596
rect 23937 22593 23949 22596
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 25590 22584 25596 22636
rect 25648 22584 25654 22636
rect 25792 22633 25820 22664
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22593 25835 22627
rect 25777 22587 25835 22593
rect 26510 22584 26516 22636
rect 26568 22584 26574 22636
rect 26697 22627 26755 22633
rect 26697 22593 26709 22627
rect 26743 22624 26755 22627
rect 27080 22624 27108 22723
rect 27890 22720 27896 22772
rect 27948 22720 27954 22772
rect 28626 22720 28632 22772
rect 28684 22760 28690 22772
rect 29641 22763 29699 22769
rect 29641 22760 29653 22763
rect 28684 22732 29653 22760
rect 28684 22720 28690 22732
rect 29641 22729 29653 22732
rect 29687 22729 29699 22763
rect 29641 22723 29699 22729
rect 29730 22720 29736 22772
rect 29788 22760 29794 22772
rect 30561 22763 30619 22769
rect 30561 22760 30573 22763
rect 29788 22732 30573 22760
rect 29788 22720 29794 22732
rect 30561 22729 30573 22732
rect 30607 22729 30619 22763
rect 30561 22723 30619 22729
rect 30650 22720 30656 22772
rect 30708 22760 30714 22772
rect 31113 22763 31171 22769
rect 31113 22760 31125 22763
rect 30708 22732 31125 22760
rect 30708 22720 30714 22732
rect 31113 22729 31125 22732
rect 31159 22729 31171 22763
rect 31113 22723 31171 22729
rect 31481 22763 31539 22769
rect 31481 22729 31493 22763
rect 31527 22760 31539 22763
rect 31527 22732 33364 22760
rect 31527 22729 31539 22732
rect 31481 22723 31539 22729
rect 27430 22652 27436 22704
rect 27488 22652 27494 22704
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 29365 22695 29423 22701
rect 29365 22692 29377 22695
rect 27672 22664 29377 22692
rect 27672 22652 27678 22664
rect 29365 22661 29377 22664
rect 29411 22661 29423 22695
rect 29365 22655 29423 22661
rect 32398 22652 32404 22704
rect 32456 22652 32462 22704
rect 26743 22596 27108 22624
rect 27249 22627 27307 22633
rect 26743 22593 26755 22596
rect 26697 22587 26755 22593
rect 27249 22593 27261 22627
rect 27295 22624 27307 22627
rect 27448 22624 27476 22652
rect 27295 22596 27476 22624
rect 27295 22593 27307 22596
rect 27249 22587 27307 22593
rect 28166 22584 28172 22636
rect 28224 22584 28230 22636
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22593 28503 22627
rect 28445 22587 28503 22593
rect 17184 22528 21864 22556
rect 17184 22516 17190 22528
rect 21836 22500 21864 22528
rect 25866 22516 25872 22568
rect 25924 22556 25930 22568
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 25924 22528 27997 22556
rect 25924 22516 25930 22528
rect 27985 22525 27997 22528
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 28074 22516 28080 22568
rect 28132 22516 28138 22568
rect 10045 22491 10103 22497
rect 10045 22457 10057 22491
rect 10091 22488 10103 22491
rect 10594 22488 10600 22500
rect 10091 22460 10600 22488
rect 10091 22457 10103 22460
rect 10045 22451 10103 22457
rect 10594 22448 10600 22460
rect 10652 22488 10658 22500
rect 15378 22488 15384 22500
rect 10652 22460 15384 22488
rect 10652 22448 10658 22460
rect 15378 22448 15384 22460
rect 15436 22448 15442 22500
rect 20070 22488 20076 22500
rect 15488 22460 20076 22488
rect 7190 22380 7196 22432
rect 7248 22380 7254 22432
rect 9125 22423 9183 22429
rect 9125 22389 9137 22423
rect 9171 22420 9183 22423
rect 9582 22420 9588 22432
rect 9171 22392 9588 22420
rect 9171 22389 9183 22392
rect 9125 22383 9183 22389
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 11882 22380 11888 22432
rect 11940 22380 11946 22432
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 15488 22420 15516 22460
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 20901 22491 20959 22497
rect 20901 22457 20913 22491
rect 20947 22488 20959 22491
rect 21542 22488 21548 22500
rect 20947 22460 21548 22488
rect 20947 22457 20959 22460
rect 20901 22451 20959 22457
rect 21542 22448 21548 22460
rect 21600 22448 21606 22500
rect 21818 22448 21824 22500
rect 21876 22448 21882 22500
rect 28184 22488 28212 22584
rect 28460 22556 28488 22587
rect 28994 22584 29000 22636
rect 29052 22584 29058 22636
rect 29549 22627 29607 22633
rect 29549 22593 29561 22627
rect 29595 22593 29607 22627
rect 29549 22587 29607 22593
rect 30009 22627 30067 22633
rect 30009 22593 30021 22627
rect 30055 22624 30067 22627
rect 30374 22624 30380 22636
rect 30055 22596 30380 22624
rect 30055 22593 30067 22596
rect 30009 22587 30067 22593
rect 29362 22556 29368 22568
rect 28460 22528 29368 22556
rect 29362 22516 29368 22528
rect 29420 22516 29426 22568
rect 29564 22556 29592 22587
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30466 22584 30472 22636
rect 30524 22584 30530 22636
rect 30926 22584 30932 22636
rect 30984 22584 30990 22636
rect 31846 22584 31852 22636
rect 31904 22584 31910 22636
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 33336 22633 33364 22732
rect 33410 22720 33416 22772
rect 33468 22720 33474 22772
rect 37001 22763 37059 22769
rect 37001 22729 37013 22763
rect 37047 22760 37059 22763
rect 37737 22763 37795 22769
rect 37737 22760 37749 22763
rect 37047 22732 37749 22760
rect 37047 22729 37059 22732
rect 37001 22723 37059 22729
rect 37737 22729 37749 22732
rect 37783 22729 37795 22763
rect 37737 22723 37795 22729
rect 38473 22763 38531 22769
rect 38473 22729 38485 22763
rect 38519 22760 38531 22763
rect 39666 22760 39672 22772
rect 38519 22732 39672 22760
rect 38519 22729 38531 22732
rect 38473 22723 38531 22729
rect 39666 22720 39672 22732
rect 39724 22720 39730 22772
rect 40954 22720 40960 22772
rect 41012 22720 41018 22772
rect 42794 22720 42800 22772
rect 42852 22720 42858 22772
rect 34882 22652 34888 22704
rect 34940 22692 34946 22704
rect 34940 22664 35388 22692
rect 34940 22652 34946 22664
rect 33045 22627 33103 22633
rect 33045 22624 33057 22627
rect 33008 22596 33057 22624
rect 33008 22584 33014 22596
rect 33045 22593 33057 22596
rect 33091 22593 33103 22627
rect 33045 22587 33103 22593
rect 33321 22627 33379 22633
rect 33321 22593 33333 22627
rect 33367 22593 33379 22627
rect 33321 22587 33379 22593
rect 33594 22584 33600 22636
rect 33652 22584 33658 22636
rect 33873 22627 33931 22633
rect 33873 22593 33885 22627
rect 33919 22593 33931 22627
rect 33873 22587 33931 22593
rect 34425 22627 34483 22633
rect 34425 22593 34437 22627
rect 34471 22624 34483 22627
rect 34471 22596 34928 22624
rect 34471 22593 34483 22596
rect 34425 22587 34483 22593
rect 31941 22559 31999 22565
rect 29564 22528 31892 22556
rect 30193 22491 30251 22497
rect 30193 22488 30205 22491
rect 28184 22460 30205 22488
rect 30193 22457 30205 22460
rect 30239 22457 30251 22491
rect 30193 22451 30251 22457
rect 30282 22448 30288 22500
rect 30340 22488 30346 22500
rect 31864 22488 31892 22528
rect 31941 22525 31953 22559
rect 31987 22556 31999 22559
rect 32030 22556 32036 22568
rect 31987 22528 32036 22556
rect 31987 22525 31999 22528
rect 31941 22519 31999 22525
rect 32030 22516 32036 22528
rect 32088 22516 32094 22568
rect 32122 22516 32128 22568
rect 32180 22516 32186 22568
rect 32582 22516 32588 22568
rect 32640 22556 32646 22568
rect 33888 22556 33916 22587
rect 32640 22528 33916 22556
rect 32640 22516 32646 22528
rect 34054 22516 34060 22568
rect 34112 22556 34118 22568
rect 34517 22559 34575 22565
rect 34517 22556 34529 22559
rect 34112 22528 34529 22556
rect 34112 22516 34118 22528
rect 34517 22525 34529 22528
rect 34563 22525 34575 22559
rect 34517 22519 34575 22525
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 34664 22528 34836 22556
rect 34664 22516 34670 22528
rect 32861 22491 32919 22497
rect 32861 22488 32873 22491
rect 30340 22460 31754 22488
rect 31864 22460 32873 22488
rect 30340 22448 30346 22460
rect 13412 22392 15516 22420
rect 13412 22380 13418 22392
rect 15838 22380 15844 22432
rect 15896 22380 15902 22432
rect 17405 22423 17463 22429
rect 17405 22389 17417 22423
rect 17451 22420 17463 22423
rect 17678 22420 17684 22432
rect 17451 22392 17684 22420
rect 17451 22389 17463 22392
rect 17405 22383 17463 22389
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 18417 22423 18475 22429
rect 18417 22389 18429 22423
rect 18463 22420 18475 22423
rect 19518 22420 19524 22432
rect 18463 22392 19524 22420
rect 18463 22389 18475 22392
rect 18417 22383 18475 22389
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 20165 22423 20223 22429
rect 20165 22389 20177 22423
rect 20211 22420 20223 22423
rect 21634 22420 21640 22432
rect 20211 22392 21640 22420
rect 20211 22389 20223 22392
rect 20165 22383 20223 22389
rect 21634 22380 21640 22392
rect 21692 22420 21698 22432
rect 22833 22423 22891 22429
rect 22833 22420 22845 22423
rect 21692 22392 22845 22420
rect 21692 22380 21698 22392
rect 22833 22389 22845 22392
rect 22879 22389 22891 22423
rect 22833 22383 22891 22389
rect 24302 22380 24308 22432
rect 24360 22420 24366 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 24360 22392 24593 22420
rect 24360 22380 24366 22392
rect 24581 22389 24593 22392
rect 24627 22420 24639 22423
rect 25314 22420 25320 22432
rect 24627 22392 25320 22420
rect 24627 22389 24639 22392
rect 24581 22383 24639 22389
rect 25314 22380 25320 22392
rect 25372 22380 25378 22432
rect 26329 22423 26387 22429
rect 26329 22389 26341 22423
rect 26375 22420 26387 22423
rect 26602 22420 26608 22432
rect 26375 22392 26608 22420
rect 26375 22389 26387 22392
rect 26329 22383 26387 22389
rect 26602 22380 26608 22392
rect 26660 22380 26666 22432
rect 27522 22380 27528 22432
rect 27580 22380 27586 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 28629 22423 28687 22429
rect 28629 22420 28641 22423
rect 27672 22392 28641 22420
rect 27672 22380 27678 22392
rect 28629 22389 28641 22392
rect 28675 22389 28687 22423
rect 31726 22420 31754 22460
rect 32861 22457 32873 22460
rect 32907 22457 32919 22491
rect 32861 22451 32919 22457
rect 32493 22423 32551 22429
rect 32493 22420 32505 22423
rect 31726 22392 32505 22420
rect 28629 22383 28687 22389
rect 32493 22389 32505 22392
rect 32539 22389 32551 22423
rect 32493 22383 32551 22389
rect 33134 22380 33140 22432
rect 33192 22380 33198 22432
rect 33502 22380 33508 22432
rect 33560 22420 33566 22432
rect 33689 22423 33747 22429
rect 33689 22420 33701 22423
rect 33560 22392 33701 22420
rect 33560 22380 33566 22392
rect 33689 22389 33701 22392
rect 33735 22389 33747 22423
rect 33689 22383 33747 22389
rect 33962 22380 33968 22432
rect 34020 22420 34026 22432
rect 34057 22423 34115 22429
rect 34057 22420 34069 22423
rect 34020 22392 34069 22420
rect 34020 22380 34026 22392
rect 34057 22389 34069 22392
rect 34103 22389 34115 22423
rect 34808 22420 34836 22528
rect 34900 22497 34928 22596
rect 35066 22584 35072 22636
rect 35124 22584 35130 22636
rect 35360 22633 35388 22664
rect 36906 22652 36912 22704
rect 36964 22692 36970 22704
rect 36964 22664 37964 22692
rect 36964 22652 36970 22664
rect 35345 22627 35403 22633
rect 35345 22593 35357 22627
rect 35391 22593 35403 22627
rect 35345 22587 35403 22593
rect 35986 22584 35992 22636
rect 36044 22584 36050 22636
rect 36265 22627 36323 22633
rect 36265 22593 36277 22627
rect 36311 22624 36323 22627
rect 37274 22624 37280 22636
rect 36311 22596 37280 22624
rect 36311 22593 36323 22596
rect 36265 22587 36323 22593
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 37642 22584 37648 22636
rect 37700 22584 37706 22636
rect 37936 22633 37964 22664
rect 38286 22652 38292 22704
rect 38344 22692 38350 22704
rect 38344 22664 38608 22692
rect 38344 22652 38350 22664
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22593 37979 22627
rect 37921 22587 37979 22593
rect 38378 22584 38384 22636
rect 38436 22584 38442 22636
rect 38580 22624 38608 22664
rect 38654 22652 38660 22704
rect 38712 22692 38718 22704
rect 38712 22664 39436 22692
rect 38712 22652 38718 22664
rect 39408 22633 39436 22664
rect 39025 22627 39083 22633
rect 39025 22624 39037 22627
rect 38580 22596 39037 22624
rect 39025 22593 39037 22596
rect 39071 22593 39083 22627
rect 39025 22587 39083 22593
rect 39393 22627 39451 22633
rect 39393 22593 39405 22627
rect 39439 22593 39451 22627
rect 39393 22587 39451 22593
rect 39482 22584 39488 22636
rect 39540 22624 39546 22636
rect 39761 22627 39819 22633
rect 39761 22624 39773 22627
rect 39540 22596 39773 22624
rect 39540 22584 39546 22596
rect 39761 22593 39773 22596
rect 39807 22593 39819 22627
rect 39761 22587 39819 22593
rect 40402 22584 40408 22636
rect 40460 22624 40466 22636
rect 40681 22627 40739 22633
rect 40681 22624 40693 22627
rect 40460 22596 40693 22624
rect 40460 22584 40466 22596
rect 40681 22593 40693 22596
rect 40727 22593 40739 22627
rect 40681 22587 40739 22593
rect 41598 22584 41604 22636
rect 41656 22584 41662 22636
rect 42242 22584 42248 22636
rect 42300 22624 42306 22636
rect 42521 22627 42579 22633
rect 42521 22624 42533 22627
rect 42300 22596 42533 22624
rect 42300 22584 42306 22596
rect 42521 22593 42533 22596
rect 42567 22593 42579 22627
rect 42521 22587 42579 22593
rect 43162 22584 43168 22636
rect 43220 22624 43226 22636
rect 43441 22627 43499 22633
rect 43441 22624 43453 22627
rect 43220 22596 43453 22624
rect 43220 22584 43226 22596
rect 43441 22593 43453 22596
rect 43487 22593 43499 22627
rect 43441 22587 43499 22593
rect 44266 22584 44272 22636
rect 44324 22624 44330 22636
rect 44545 22627 44603 22633
rect 44545 22624 44557 22627
rect 44324 22596 44557 22624
rect 44324 22584 44330 22596
rect 44545 22593 44557 22596
rect 44591 22593 44603 22627
rect 44545 22587 44603 22593
rect 45186 22584 45192 22636
rect 45244 22584 45250 22636
rect 37090 22516 37096 22568
rect 37148 22516 37154 22568
rect 37185 22559 37243 22565
rect 37185 22525 37197 22559
rect 37231 22525 37243 22559
rect 37185 22519 37243 22525
rect 34885 22491 34943 22497
rect 34885 22457 34897 22491
rect 34931 22457 34943 22491
rect 37200 22488 37228 22519
rect 37550 22516 37556 22568
rect 37608 22556 37614 22568
rect 38565 22559 38623 22565
rect 37608 22528 38056 22556
rect 37608 22516 37614 22528
rect 37366 22488 37372 22500
rect 34885 22451 34943 22457
rect 35084 22460 37372 22488
rect 35084 22420 35112 22460
rect 37366 22448 37372 22460
rect 37424 22448 37430 22500
rect 37918 22488 37924 22500
rect 37476 22460 37924 22488
rect 34808 22392 35112 22420
rect 34057 22383 34115 22389
rect 35158 22380 35164 22432
rect 35216 22380 35222 22432
rect 35710 22380 35716 22432
rect 35768 22380 35774 22432
rect 35802 22380 35808 22432
rect 35860 22380 35866 22432
rect 36078 22380 36084 22432
rect 36136 22380 36142 22432
rect 36630 22380 36636 22432
rect 36688 22380 36694 22432
rect 37476 22429 37504 22460
rect 37918 22448 37924 22460
rect 37976 22448 37982 22500
rect 38028 22488 38056 22528
rect 38565 22525 38577 22559
rect 38611 22525 38623 22559
rect 38565 22519 38623 22525
rect 38580 22488 38608 22519
rect 40037 22491 40095 22497
rect 40037 22488 40049 22491
rect 38028 22460 38608 22488
rect 38764 22460 40049 22488
rect 37461 22423 37519 22429
rect 37461 22389 37473 22423
rect 37507 22389 37519 22423
rect 37461 22383 37519 22389
rect 38010 22380 38016 22432
rect 38068 22380 38074 22432
rect 38286 22380 38292 22432
rect 38344 22420 38350 22432
rect 38764 22420 38792 22460
rect 40037 22457 40049 22460
rect 40083 22488 40095 22491
rect 40954 22488 40960 22500
rect 40083 22460 40960 22488
rect 40083 22457 40095 22460
rect 40037 22451 40095 22457
rect 40954 22448 40960 22460
rect 41012 22448 41018 22500
rect 44821 22491 44879 22497
rect 44821 22488 44833 22491
rect 44192 22460 44833 22488
rect 44192 22432 44220 22460
rect 44821 22457 44833 22460
rect 44867 22457 44879 22491
rect 44821 22451 44879 22457
rect 38344 22392 38792 22420
rect 38344 22380 38350 22392
rect 38838 22380 38844 22432
rect 38896 22380 38902 22432
rect 39206 22380 39212 22432
rect 39264 22380 39270 22432
rect 39298 22380 39304 22432
rect 39356 22420 39362 22432
rect 39577 22423 39635 22429
rect 39577 22420 39589 22423
rect 39356 22392 39589 22420
rect 39356 22380 39362 22392
rect 39577 22389 39589 22392
rect 39623 22389 39635 22423
rect 39577 22383 39635 22389
rect 40494 22380 40500 22432
rect 40552 22380 40558 22432
rect 41414 22380 41420 22432
rect 41472 22380 41478 22432
rect 42061 22423 42119 22429
rect 42061 22389 42073 22423
rect 42107 22420 42119 22423
rect 42150 22420 42156 22432
rect 42107 22392 42156 22420
rect 42107 22389 42119 22392
rect 42061 22383 42119 22389
rect 42150 22380 42156 22392
rect 42208 22380 42214 22432
rect 42337 22423 42395 22429
rect 42337 22389 42349 22423
rect 42383 22420 42395 22423
rect 42702 22420 42708 22432
rect 42383 22392 42708 22420
rect 42383 22389 42395 22392
rect 42337 22383 42395 22389
rect 42702 22380 42708 22392
rect 42760 22380 42766 22432
rect 43254 22380 43260 22432
rect 43312 22380 43318 22432
rect 43809 22423 43867 22429
rect 43809 22389 43821 22423
rect 43855 22420 43867 22423
rect 43898 22420 43904 22432
rect 43855 22392 43904 22420
rect 43855 22389 43867 22392
rect 43809 22383 43867 22389
rect 43898 22380 43904 22392
rect 43956 22380 43962 22432
rect 44174 22380 44180 22432
rect 44232 22380 44238 22432
rect 44358 22380 44364 22432
rect 44416 22380 44422 22432
rect 45002 22380 45008 22432
rect 45060 22380 45066 22432
rect 460 22330 45540 22352
rect 460 22278 3570 22330
rect 3622 22278 3634 22330
rect 3686 22278 3698 22330
rect 3750 22278 3762 22330
rect 3814 22278 3826 22330
rect 3878 22278 8570 22330
rect 8622 22278 8634 22330
rect 8686 22278 8698 22330
rect 8750 22278 8762 22330
rect 8814 22278 8826 22330
rect 8878 22278 13570 22330
rect 13622 22278 13634 22330
rect 13686 22278 13698 22330
rect 13750 22278 13762 22330
rect 13814 22278 13826 22330
rect 13878 22278 18570 22330
rect 18622 22278 18634 22330
rect 18686 22278 18698 22330
rect 18750 22278 18762 22330
rect 18814 22278 18826 22330
rect 18878 22278 23570 22330
rect 23622 22278 23634 22330
rect 23686 22278 23698 22330
rect 23750 22278 23762 22330
rect 23814 22278 23826 22330
rect 23878 22278 28570 22330
rect 28622 22278 28634 22330
rect 28686 22278 28698 22330
rect 28750 22278 28762 22330
rect 28814 22278 28826 22330
rect 28878 22278 33570 22330
rect 33622 22278 33634 22330
rect 33686 22278 33698 22330
rect 33750 22278 33762 22330
rect 33814 22278 33826 22330
rect 33878 22278 38570 22330
rect 38622 22278 38634 22330
rect 38686 22278 38698 22330
rect 38750 22278 38762 22330
rect 38814 22278 38826 22330
rect 38878 22278 43570 22330
rect 43622 22278 43634 22330
rect 43686 22278 43698 22330
rect 43750 22278 43762 22330
rect 43814 22278 43826 22330
rect 43878 22278 45540 22330
rect 460 22256 45540 22278
rect 934 22176 940 22228
rect 992 22216 998 22228
rect 1397 22219 1455 22225
rect 1397 22216 1409 22219
rect 992 22188 1409 22216
rect 992 22176 998 22188
rect 1397 22185 1409 22188
rect 1443 22185 1455 22219
rect 1397 22179 1455 22185
rect 1854 22176 1860 22228
rect 1912 22216 1918 22228
rect 2041 22219 2099 22225
rect 2041 22216 2053 22219
rect 1912 22188 2053 22216
rect 1912 22176 1918 22188
rect 2041 22185 2053 22188
rect 2087 22185 2099 22219
rect 2041 22179 2099 22185
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 3234 22216 3240 22228
rect 2823 22188 3240 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 3881 22219 3939 22225
rect 3881 22185 3893 22219
rect 3927 22216 3939 22219
rect 3970 22216 3976 22228
rect 3927 22188 3976 22216
rect 3927 22185 3939 22188
rect 3881 22179 3939 22185
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 4614 22176 4620 22228
rect 4672 22176 4678 22228
rect 5445 22219 5503 22225
rect 5445 22185 5457 22219
rect 5491 22216 5503 22219
rect 5810 22216 5816 22228
rect 5491 22188 5816 22216
rect 5491 22185 5503 22188
rect 5445 22179 5503 22185
rect 5810 22176 5816 22188
rect 5868 22176 5874 22228
rect 5994 22176 6000 22228
rect 6052 22176 6058 22228
rect 6454 22176 6460 22228
rect 6512 22176 6518 22228
rect 7285 22219 7343 22225
rect 7285 22185 7297 22219
rect 7331 22216 7343 22219
rect 7374 22216 7380 22228
rect 7331 22188 7380 22216
rect 7331 22185 7343 22188
rect 7285 22179 7343 22185
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8386 22216 8392 22228
rect 8343 22188 8392 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8386 22176 8392 22188
rect 8444 22176 8450 22228
rect 9214 22176 9220 22228
rect 9272 22216 9278 22228
rect 9401 22219 9459 22225
rect 9401 22216 9413 22219
rect 9272 22188 9413 22216
rect 9272 22176 9278 22188
rect 9401 22185 9413 22188
rect 9447 22185 9459 22219
rect 9401 22179 9459 22185
rect 10134 22176 10140 22228
rect 10192 22176 10198 22228
rect 10873 22219 10931 22225
rect 10873 22185 10885 22219
rect 10919 22216 10931 22219
rect 11146 22216 11152 22228
rect 10919 22188 11152 22216
rect 10919 22185 10931 22188
rect 10873 22179 10931 22185
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11793 22219 11851 22225
rect 11793 22185 11805 22219
rect 11839 22216 11851 22219
rect 11974 22216 11980 22228
rect 11839 22188 11980 22216
rect 11839 22185 11851 22188
rect 11793 22179 11851 22185
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12805 22219 12863 22225
rect 12805 22185 12817 22219
rect 12851 22216 12863 22219
rect 12894 22216 12900 22228
rect 12851 22188 12900 22216
rect 12851 22185 12863 22188
rect 12805 22179 12863 22185
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13446 22176 13452 22228
rect 13504 22216 13510 22228
rect 13541 22219 13599 22225
rect 13541 22216 13553 22219
rect 13504 22188 13553 22216
rect 13504 22176 13510 22188
rect 13541 22185 13553 22188
rect 13587 22185 13599 22219
rect 13541 22179 13599 22185
rect 13998 22176 14004 22228
rect 14056 22176 14062 22228
rect 14093 22219 14151 22225
rect 14093 22185 14105 22219
rect 14139 22216 14151 22219
rect 14734 22216 14740 22228
rect 14139 22188 14740 22216
rect 14139 22185 14151 22188
rect 14093 22179 14151 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 16758 22176 16764 22228
rect 16816 22176 16822 22228
rect 17221 22219 17279 22225
rect 17221 22185 17233 22219
rect 17267 22216 17279 22219
rect 17494 22216 17500 22228
rect 17267 22188 17500 22216
rect 17267 22185 17279 22188
rect 17221 22179 17279 22185
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 17678 22176 17684 22228
rect 17736 22216 17742 22228
rect 17773 22219 17831 22225
rect 17773 22216 17785 22219
rect 17736 22188 17785 22216
rect 17736 22176 17742 22188
rect 17773 22185 17785 22188
rect 17819 22216 17831 22219
rect 17819 22188 18184 22216
rect 17819 22185 17831 22188
rect 17773 22179 17831 22185
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 1946 22012 1952 22024
rect 1627 21984 1952 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 1946 21972 1952 21984
rect 2004 21972 2010 22024
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 2961 22015 3019 22021
rect 2961 21981 2973 22015
rect 3007 22012 3019 22015
rect 3050 22012 3056 22024
rect 3007 21984 3056 22012
rect 3007 21981 3019 21984
rect 2961 21975 3019 21981
rect 2240 21944 2268 21975
rect 3050 21972 3056 21984
rect 3108 22012 3114 22024
rect 3329 22015 3387 22021
rect 3329 22012 3341 22015
rect 3108 21984 3341 22012
rect 3108 21972 3114 21984
rect 3329 21981 3341 21984
rect 3375 21981 3387 22015
rect 3329 21975 3387 21981
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4430 22012 4436 22024
rect 4111 21984 4436 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 4430 21972 4436 21984
rect 4488 21972 4494 22024
rect 4801 22015 4859 22021
rect 4801 21981 4813 22015
rect 4847 22012 4859 22015
rect 5074 22012 5080 22024
rect 4847 21984 5080 22012
rect 4847 21981 4859 21984
rect 4801 21975 4859 21981
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 22012 5687 22015
rect 6012 22012 6040 22176
rect 14016 22148 14044 22176
rect 7484 22120 14044 22148
rect 7484 22021 7512 22120
rect 16298 22108 16304 22160
rect 16356 22148 16362 22160
rect 18156 22148 18184 22188
rect 18230 22176 18236 22228
rect 18288 22176 18294 22228
rect 19702 22176 19708 22228
rect 19760 22176 19766 22228
rect 19981 22219 20039 22225
rect 19981 22185 19993 22219
rect 20027 22216 20039 22219
rect 20254 22216 20260 22228
rect 20027 22188 20260 22216
rect 20027 22185 20039 22188
rect 19981 22179 20039 22185
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 22097 22219 22155 22225
rect 20364 22188 21588 22216
rect 16356 22120 17954 22148
rect 18156 22120 19472 22148
rect 16356 22108 16362 22120
rect 9309 22083 9367 22089
rect 9309 22049 9321 22083
rect 9355 22080 9367 22083
rect 12345 22083 12403 22089
rect 9355 22052 12204 22080
rect 9355 22049 9367 22052
rect 9309 22043 9367 22049
rect 6641 22015 6699 22021
rect 6641 22012 6653 22015
rect 5675 21984 6040 22012
rect 6472 21984 6653 22012
rect 5675 21981 5687 21984
rect 5629 21975 5687 21981
rect 2593 21947 2651 21953
rect 2593 21944 2605 21947
rect 2240 21916 2605 21944
rect 2593 21913 2605 21916
rect 2639 21944 2651 21947
rect 5442 21944 5448 21956
rect 2639 21916 5448 21944
rect 2639 21913 2651 21916
rect 2593 21907 2651 21913
rect 5442 21904 5448 21916
rect 5500 21904 5506 21956
rect 6472 21888 6500 21984
rect 6641 21981 6653 21984
rect 6687 21981 6699 22015
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 6641 21975 6699 21981
rect 7208 21984 7481 22012
rect 7208 21888 7236 21984
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 9582 21972 9588 22024
rect 9640 21972 9646 22024
rect 11072 22021 11100 22052
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 21981 11115 22015
rect 11057 21975 11115 21981
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12066 22012 12072 22024
rect 12023 21984 12072 22012
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 10336 21944 10364 21975
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12176 22012 12204 22052
rect 12345 22049 12357 22083
rect 12391 22080 12403 22083
rect 17926 22080 17954 22120
rect 19444 22080 19472 22120
rect 19518 22108 19524 22160
rect 19576 22148 19582 22160
rect 20364 22148 20392 22188
rect 19576 22120 20392 22148
rect 21560 22148 21588 22188
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22186 22216 22192 22228
rect 22143 22188 22192 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 22741 22219 22799 22225
rect 22741 22185 22753 22219
rect 22787 22216 22799 22219
rect 23014 22216 23020 22228
rect 22787 22188 23020 22216
rect 22787 22185 22799 22188
rect 22741 22179 22799 22185
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 23106 22176 23112 22228
rect 23164 22176 23170 22228
rect 24762 22176 24768 22228
rect 24820 22216 24826 22228
rect 24949 22219 25007 22225
rect 24949 22216 24961 22219
rect 24820 22188 24961 22216
rect 24820 22176 24826 22188
rect 24949 22185 24961 22188
rect 24995 22185 25007 22219
rect 24949 22179 25007 22185
rect 29362 22176 29368 22228
rect 29420 22176 29426 22228
rect 31008 22219 31066 22225
rect 31008 22185 31020 22219
rect 31054 22216 31066 22219
rect 33134 22216 33140 22228
rect 31054 22188 33140 22216
rect 31054 22185 31066 22188
rect 31008 22179 31066 22185
rect 33134 22176 33140 22188
rect 33192 22176 33198 22228
rect 33962 22176 33968 22228
rect 34020 22176 34026 22228
rect 36252 22219 36310 22225
rect 36252 22185 36264 22219
rect 36298 22216 36310 22219
rect 36446 22216 36452 22228
rect 36298 22188 36452 22216
rect 36298 22185 36310 22188
rect 36252 22179 36310 22185
rect 36446 22176 36452 22188
rect 36504 22176 36510 22228
rect 40954 22176 40960 22228
rect 41012 22216 41018 22228
rect 41693 22219 41751 22225
rect 41693 22216 41705 22219
rect 41012 22188 41705 22216
rect 41012 22176 41018 22188
rect 41693 22185 41705 22188
rect 41739 22216 41751 22219
rect 42429 22219 42487 22225
rect 42429 22216 42441 22219
rect 41739 22188 42441 22216
rect 41739 22185 41751 22188
rect 41693 22179 41751 22185
rect 42429 22185 42441 22188
rect 42475 22185 42487 22219
rect 42429 22179 42487 22185
rect 21560 22120 22508 22148
rect 19576 22108 19582 22120
rect 20257 22083 20315 22089
rect 20257 22080 20269 22083
rect 12391 22052 16896 22080
rect 17926 22052 18552 22080
rect 12391 22049 12403 22052
rect 12345 22043 12403 22049
rect 12710 22012 12716 22024
rect 12176 21984 12716 22012
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12989 22015 13047 22021
rect 12989 21981 13001 22015
rect 13035 22012 13047 22015
rect 13078 22012 13084 22024
rect 13035 21984 13084 22012
rect 13035 21981 13047 21984
rect 12989 21975 13047 21981
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13725 22015 13783 22021
rect 13188 21984 13676 22012
rect 8956 21916 10364 21944
rect 8956 21888 8984 21916
rect 6365 21879 6423 21885
rect 6365 21845 6377 21879
rect 6411 21876 6423 21879
rect 6454 21876 6460 21888
rect 6411 21848 6460 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 7190 21836 7196 21888
rect 7248 21836 7254 21888
rect 7282 21836 7288 21888
rect 7340 21876 7346 21888
rect 8021 21879 8079 21885
rect 8021 21876 8033 21879
rect 7340 21848 8033 21876
rect 7340 21836 7346 21848
rect 8021 21845 8033 21848
rect 8067 21845 8079 21879
rect 8021 21839 8079 21845
rect 8938 21836 8944 21888
rect 8996 21836 9002 21888
rect 10042 21836 10048 21888
rect 10100 21836 10106 21888
rect 10336 21876 10364 21916
rect 10781 21947 10839 21953
rect 10781 21913 10793 21947
rect 10827 21944 10839 21947
rect 13188 21944 13216 21984
rect 10827 21916 13216 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 11606 21876 11612 21888
rect 10336 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 11698 21836 11704 21888
rect 11756 21836 11762 21888
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21876 12771 21879
rect 13446 21876 13452 21888
rect 12759 21848 13452 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 13648 21876 13676 21984
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 13725 21975 13783 21981
rect 14108 21984 14289 22012
rect 13748 21944 13776 21975
rect 13906 21944 13912 21956
rect 13748 21916 13912 21944
rect 13906 21904 13912 21916
rect 13964 21904 13970 21956
rect 14108 21888 14136 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 22012 14427 22015
rect 14458 22012 14464 22024
rect 14415 21984 14464 22012
rect 14415 21981 14427 21984
rect 14369 21975 14427 21981
rect 14458 21972 14464 21984
rect 14516 21972 14522 22024
rect 14734 21972 14740 22024
rect 14792 21972 14798 22024
rect 15654 21972 15660 22024
rect 15712 22012 15718 22024
rect 16163 22015 16221 22021
rect 16163 22012 16175 22015
rect 15712 21984 16175 22012
rect 15712 21972 15718 21984
rect 16163 21981 16175 21984
rect 16209 22012 16221 22015
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 16209 21984 16313 22012
rect 16209 21981 16221 21984
rect 16163 21975 16221 21981
rect 16301 21981 16313 21984
rect 16347 22012 16359 22015
rect 16390 22012 16396 22024
rect 16347 21984 16396 22012
rect 16347 21981 16359 21984
rect 16301 21975 16359 21981
rect 16390 21972 16396 21984
rect 16448 21972 16454 22024
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 15930 21944 15936 21956
rect 15778 21916 15936 21944
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 16500 21944 16528 21975
rect 16758 21944 16764 21956
rect 16500 21916 16764 21944
rect 14090 21876 14096 21888
rect 13648 21848 14096 21876
rect 14090 21836 14096 21848
rect 14148 21836 14154 21888
rect 15654 21836 15660 21888
rect 15712 21876 15718 21888
rect 16500 21876 16528 21916
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 16868 21944 16896 22052
rect 16945 22015 17003 22021
rect 16945 21981 16957 22015
rect 16991 22012 17003 22015
rect 17310 22012 17316 22024
rect 16991 21984 17316 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 17494 22012 17500 22024
rect 17451 21984 17500 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 17920 21984 18429 22012
rect 17920 21972 17926 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 18322 21944 18328 21956
rect 16868 21916 18328 21944
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 18524 21944 18552 22052
rect 18616 22052 19196 22080
rect 19444 22052 20269 22080
rect 18616 22021 18644 22052
rect 19168 22024 19196 22052
rect 20257 22049 20269 22052
rect 20303 22080 20315 22083
rect 20303 22052 21588 22080
rect 20303 22049 20315 22052
rect 20257 22043 20315 22049
rect 21560 22024 21588 22052
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 21981 18659 22015
rect 18601 21975 18659 21981
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 18969 22015 19027 22021
rect 18969 22012 18981 22015
rect 18748 21984 18981 22012
rect 18748 21972 18754 21984
rect 18969 21981 18981 21984
rect 19015 22012 19027 22015
rect 19058 22012 19064 22024
rect 19015 21984 19064 22012
rect 19015 21981 19027 21984
rect 18969 21975 19027 21981
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 19150 21972 19156 22024
rect 19208 21972 19214 22024
rect 19242 21972 19248 22024
rect 19300 21972 19306 22024
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 22012 19487 22015
rect 19889 22015 19947 22021
rect 19889 22012 19901 22015
rect 19475 21984 19748 22012
rect 19475 21981 19487 21984
rect 19429 21975 19487 21981
rect 18782 21944 18788 21956
rect 18524 21916 18788 21944
rect 18782 21904 18788 21916
rect 18840 21904 18846 21956
rect 18877 21947 18935 21953
rect 18877 21913 18889 21947
rect 18923 21944 18935 21947
rect 18923 21916 19472 21944
rect 18923 21913 18935 21916
rect 18877 21907 18935 21913
rect 19444 21888 19472 21916
rect 19720 21888 19748 21984
rect 19812 21984 19901 22012
rect 19812 21888 19840 21984
rect 19889 21981 19901 21984
rect 19935 21981 19947 22015
rect 19889 21975 19947 21981
rect 20162 21972 20168 22024
rect 20220 21972 20226 22024
rect 21542 21972 21548 22024
rect 21600 21972 21606 22024
rect 21634 21972 21640 22024
rect 21692 21972 21698 22024
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22370 22012 22376 22024
rect 22327 21984 22376 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 22480 22012 22508 22120
rect 32030 22108 32036 22160
rect 32088 22148 32094 22160
rect 32490 22148 32496 22160
rect 32088 22120 32496 22148
rect 32088 22108 32094 22120
rect 32490 22108 32496 22120
rect 32548 22108 32554 22160
rect 32674 22108 32680 22160
rect 32732 22148 32738 22160
rect 33980 22148 34008 22176
rect 32732 22120 34008 22148
rect 32732 22108 32738 22120
rect 35434 22108 35440 22160
rect 35492 22148 35498 22160
rect 35492 22120 36124 22148
rect 35492 22108 35498 22120
rect 24762 22040 24768 22092
rect 24820 22040 24826 22092
rect 27798 22040 27804 22092
rect 27856 22040 27862 22092
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28442 22080 28448 22092
rect 28132 22052 28448 22080
rect 28132 22040 28138 22052
rect 28442 22040 28448 22052
rect 28500 22080 28506 22092
rect 28537 22083 28595 22089
rect 28537 22080 28549 22083
rect 28500 22052 28549 22080
rect 28500 22040 28506 22052
rect 28537 22049 28549 22052
rect 28583 22049 28595 22083
rect 28537 22043 28595 22049
rect 30006 22040 30012 22092
rect 30064 22040 30070 22092
rect 30116 22052 32352 22080
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22480 21984 22937 22012
rect 22925 21981 22937 21984
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 22012 23351 22015
rect 23382 22012 23388 22024
rect 23339 21984 23388 22012
rect 23339 21981 23351 21984
rect 23293 21975 23351 21981
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 23566 21972 23572 22024
rect 23624 21972 23630 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 20533 21947 20591 21953
rect 20533 21944 20545 21947
rect 19904 21916 20545 21944
rect 19904 21888 19932 21916
rect 20533 21913 20545 21916
rect 20579 21913 20591 21947
rect 20533 21907 20591 21913
rect 15712 21848 16528 21876
rect 16669 21879 16727 21885
rect 15712 21836 15718 21848
rect 16669 21845 16681 21879
rect 16715 21876 16727 21879
rect 17034 21876 17040 21888
rect 16715 21848 17040 21876
rect 16715 21845 16727 21848
rect 16669 21839 16727 21845
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 18138 21836 18144 21888
rect 18196 21836 18202 21888
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 19153 21879 19211 21885
rect 19153 21876 19165 21879
rect 18288 21848 19165 21876
rect 18288 21836 18294 21848
rect 19153 21845 19165 21848
rect 19199 21845 19211 21879
rect 19153 21839 19211 21845
rect 19334 21836 19340 21888
rect 19392 21836 19398 21888
rect 19426 21836 19432 21888
rect 19484 21836 19490 21888
rect 19702 21836 19708 21888
rect 19760 21836 19766 21888
rect 19794 21836 19800 21888
rect 19852 21836 19858 21888
rect 19886 21836 19892 21888
rect 19944 21836 19950 21888
rect 20438 21836 20444 21888
rect 20496 21876 20502 21888
rect 22005 21879 22063 21885
rect 22005 21876 22017 21879
rect 20496 21848 22017 21876
rect 20496 21836 20502 21848
rect 22005 21845 22017 21848
rect 22051 21876 22063 21879
rect 22186 21876 22192 21888
rect 22051 21848 22192 21876
rect 22051 21845 22063 21848
rect 22005 21839 22063 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22336 21848 22661 21876
rect 22336 21836 22342 21848
rect 22649 21845 22661 21848
rect 22695 21876 22707 21879
rect 23198 21876 23204 21888
rect 22695 21848 23204 21876
rect 22695 21845 22707 21848
rect 22649 21839 22707 21845
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 23385 21879 23443 21885
rect 23385 21845 23397 21879
rect 23431 21876 23443 21879
rect 23474 21876 23480 21888
rect 23431 21848 23480 21876
rect 23431 21845 23443 21848
rect 23385 21839 23443 21845
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23842 21836 23848 21888
rect 23900 21836 23906 21888
rect 24044 21876 24072 21975
rect 25130 21972 25136 22024
rect 25188 21972 25194 22024
rect 25314 21972 25320 22024
rect 25372 21972 25378 22024
rect 26726 21984 27292 22012
rect 24486 21904 24492 21956
rect 24544 21944 24550 21956
rect 24544 21916 25452 21944
rect 24544 21904 24550 21916
rect 24121 21879 24179 21885
rect 24121 21876 24133 21879
rect 24044 21848 24133 21876
rect 24121 21845 24133 21848
rect 24167 21845 24179 21879
rect 24121 21839 24179 21845
rect 24581 21879 24639 21885
rect 24581 21845 24593 21879
rect 24627 21876 24639 21879
rect 25314 21876 25320 21888
rect 24627 21848 25320 21876
rect 24627 21845 24639 21848
rect 24581 21839 24639 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 25424 21876 25452 21916
rect 25590 21904 25596 21956
rect 25648 21904 25654 21956
rect 27264 21944 27292 21984
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 28902 21972 28908 22024
rect 28960 21972 28966 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 22012 29791 22015
rect 30116 22012 30144 22052
rect 29779 21984 30144 22012
rect 29779 21981 29791 21984
rect 29733 21975 29791 21981
rect 30190 21972 30196 22024
rect 30248 21972 30254 22024
rect 30282 21972 30288 22024
rect 30340 22012 30346 22024
rect 30745 22015 30803 22021
rect 30340 21984 30696 22012
rect 30340 21972 30346 21984
rect 27890 21944 27896 21956
rect 26988 21916 27200 21944
rect 27264 21916 27896 21944
rect 25774 21876 25780 21888
rect 25424 21848 25780 21876
rect 25774 21836 25780 21848
rect 25832 21836 25838 21888
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 26988 21876 27016 21916
rect 26016 21848 27016 21876
rect 26016 21836 26022 21848
rect 27062 21836 27068 21888
rect 27120 21836 27126 21888
rect 27172 21885 27200 21916
rect 27890 21904 27896 21916
rect 27948 21904 27954 21956
rect 28350 21904 28356 21956
rect 28408 21904 28414 21956
rect 29825 21947 29883 21953
rect 29825 21913 29837 21947
rect 29871 21944 29883 21947
rect 30558 21944 30564 21956
rect 29871 21916 30564 21944
rect 29871 21913 29883 21916
rect 29825 21907 29883 21913
rect 30558 21904 30564 21916
rect 30616 21904 30622 21956
rect 27157 21879 27215 21885
rect 27157 21845 27169 21879
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 27522 21836 27528 21888
rect 27580 21876 27586 21888
rect 27617 21879 27675 21885
rect 27617 21876 27629 21879
rect 27580 21848 27629 21876
rect 27580 21836 27586 21848
rect 27617 21845 27629 21848
rect 27663 21845 27675 21879
rect 27617 21839 27675 21845
rect 27982 21836 27988 21888
rect 28040 21836 28046 21888
rect 28074 21836 28080 21888
rect 28132 21876 28138 21888
rect 28445 21879 28503 21885
rect 28445 21876 28457 21879
rect 28132 21848 28457 21876
rect 28132 21836 28138 21848
rect 28445 21845 28457 21848
rect 28491 21845 28503 21879
rect 28445 21839 28503 21845
rect 29086 21836 29092 21888
rect 29144 21836 29150 21888
rect 30006 21836 30012 21888
rect 30064 21876 30070 21888
rect 30377 21879 30435 21885
rect 30377 21876 30389 21879
rect 30064 21848 30389 21876
rect 30064 21836 30070 21848
rect 30377 21845 30389 21848
rect 30423 21845 30435 21879
rect 30668 21876 30696 21984
rect 30745 21981 30757 22015
rect 30791 21981 30803 22015
rect 30745 21975 30803 21981
rect 30760 21944 30788 21975
rect 30926 21944 30932 21956
rect 30760 21916 30932 21944
rect 30926 21904 30932 21916
rect 30984 21904 30990 21956
rect 32140 21876 32168 21998
rect 32324 21944 32352 22052
rect 32858 22040 32864 22092
rect 32916 22080 32922 22092
rect 33137 22083 33195 22089
rect 33137 22080 33149 22083
rect 32916 22052 33149 22080
rect 32916 22040 32922 22052
rect 33137 22049 33149 22052
rect 33183 22049 33195 22083
rect 33137 22043 33195 22049
rect 33318 22040 33324 22092
rect 33376 22080 33382 22092
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 33376 22052 34069 22080
rect 33376 22040 33382 22052
rect 34057 22049 34069 22052
rect 34103 22080 34115 22083
rect 35989 22083 36047 22089
rect 35989 22080 36001 22083
rect 34103 22052 36001 22080
rect 34103 22049 34115 22052
rect 34057 22043 34115 22049
rect 35989 22049 36001 22052
rect 36035 22049 36047 22083
rect 36096 22080 36124 22120
rect 37366 22108 37372 22160
rect 37424 22148 37430 22160
rect 38194 22148 38200 22160
rect 37424 22120 38200 22148
rect 37424 22108 37430 22120
rect 38194 22108 38200 22120
rect 38252 22148 38258 22160
rect 40129 22151 40187 22157
rect 38252 22120 39804 22148
rect 38252 22108 38258 22120
rect 38396 22089 38424 22120
rect 39776 22089 39804 22120
rect 40129 22117 40141 22151
rect 40175 22148 40187 22151
rect 40175 22120 40209 22148
rect 40175 22117 40187 22120
rect 40129 22111 40187 22117
rect 38381 22083 38439 22089
rect 36096 22052 37596 22080
rect 35989 22043 36047 22049
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 32548 21984 32904 22012
rect 32548 21972 32554 21984
rect 32674 21944 32680 21956
rect 32324 21916 32680 21944
rect 32674 21904 32680 21916
rect 32732 21904 32738 21956
rect 32306 21876 32312 21888
rect 30668 21848 32312 21876
rect 30377 21839 30435 21845
rect 32306 21836 32312 21848
rect 32364 21836 32370 21888
rect 32582 21836 32588 21888
rect 32640 21836 32646 21888
rect 32876 21876 32904 21984
rect 33042 21972 33048 22024
rect 33100 22012 33106 22024
rect 33597 22015 33655 22021
rect 33597 22012 33609 22015
rect 33100 21984 33609 22012
rect 33100 21972 33106 21984
rect 33597 21981 33609 21984
rect 33643 21981 33655 22015
rect 33597 21975 33655 21981
rect 33870 21972 33876 22024
rect 33928 21972 33934 22024
rect 35434 21972 35440 22024
rect 35492 21972 35498 22024
rect 32953 21947 33011 21953
rect 32953 21913 32965 21947
rect 32999 21944 33011 21947
rect 34333 21947 34391 21953
rect 34333 21944 34345 21947
rect 32999 21916 33456 21944
rect 32999 21913 33011 21916
rect 32953 21907 33011 21913
rect 33428 21885 33456 21916
rect 33704 21916 34345 21944
rect 33704 21885 33732 21916
rect 34333 21913 34345 21916
rect 34379 21913 34391 21947
rect 36004 21944 36032 22043
rect 37366 21972 37372 22024
rect 37424 21972 37430 22024
rect 36538 21944 36544 21956
rect 36004 21916 36544 21944
rect 34333 21907 34391 21913
rect 36538 21904 36544 21916
rect 36596 21904 36602 21956
rect 37568 21944 37596 22052
rect 38381 22049 38393 22083
rect 38427 22080 38439 22083
rect 39761 22083 39819 22089
rect 38427 22052 38461 22080
rect 38427 22049 38439 22052
rect 38381 22043 38439 22049
rect 39761 22049 39773 22083
rect 39807 22080 39819 22083
rect 39807 22052 39841 22080
rect 39807 22049 39819 22052
rect 39761 22043 39819 22049
rect 40034 22040 40040 22092
rect 40092 22080 40098 22092
rect 40144 22080 40172 22111
rect 40092 22052 40172 22080
rect 40092 22040 40098 22052
rect 43162 22040 43168 22092
rect 43220 22080 43226 22092
rect 44545 22083 44603 22089
rect 44545 22080 44557 22083
rect 43220 22052 44557 22080
rect 43220 22040 43226 22052
rect 44545 22049 44557 22052
rect 44591 22049 44603 22083
rect 44545 22043 44603 22049
rect 38197 22015 38255 22021
rect 38197 21981 38209 22015
rect 38243 22012 38255 22015
rect 38930 22012 38936 22024
rect 38243 21984 38936 22012
rect 38243 21981 38255 21984
rect 38197 21975 38255 21981
rect 38930 21972 38936 21984
rect 38988 21972 38994 22024
rect 39206 21972 39212 22024
rect 39264 22012 39270 22024
rect 39577 22015 39635 22021
rect 39577 22012 39589 22015
rect 39264 21984 39589 22012
rect 39264 21972 39270 21984
rect 39577 21981 39589 21984
rect 39623 21981 39635 22015
rect 39577 21975 39635 21981
rect 40313 22015 40371 22021
rect 40313 21981 40325 22015
rect 40359 22012 40371 22015
rect 41690 22012 41696 22024
rect 40359 21984 41696 22012
rect 40359 21981 40371 21984
rect 40313 21975 40371 21981
rect 41690 21972 41696 21984
rect 41748 21972 41754 22024
rect 43898 21972 43904 22024
rect 43956 22012 43962 22024
rect 44913 22015 44971 22021
rect 44913 22012 44925 22015
rect 43956 21984 44925 22012
rect 43956 21972 43962 21984
rect 44913 21981 44925 21984
rect 44959 21981 44971 22015
rect 44913 21975 44971 21981
rect 43165 21947 43223 21953
rect 43165 21944 43177 21947
rect 37568 21916 43177 21944
rect 43165 21913 43177 21916
rect 43211 21913 43223 21947
rect 43165 21907 43223 21913
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32876 21848 33057 21876
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33413 21879 33471 21885
rect 33413 21845 33425 21879
rect 33459 21845 33471 21879
rect 33413 21839 33471 21845
rect 33689 21879 33747 21885
rect 33689 21845 33701 21879
rect 33735 21845 33747 21879
rect 33689 21839 33747 21845
rect 35618 21836 35624 21888
rect 35676 21876 35682 21888
rect 35805 21879 35863 21885
rect 35805 21876 35817 21879
rect 35676 21848 35817 21876
rect 35676 21836 35682 21848
rect 35805 21845 35817 21848
rect 35851 21845 35863 21879
rect 35805 21839 35863 21845
rect 37734 21836 37740 21888
rect 37792 21836 37798 21888
rect 37826 21836 37832 21888
rect 37884 21836 37890 21888
rect 38286 21836 38292 21888
rect 38344 21836 38350 21888
rect 38378 21836 38384 21888
rect 38436 21876 38442 21888
rect 38841 21879 38899 21885
rect 38841 21876 38853 21879
rect 38436 21848 38853 21876
rect 38436 21836 38442 21848
rect 38841 21845 38853 21848
rect 38887 21845 38899 21879
rect 38841 21839 38899 21845
rect 38930 21836 38936 21888
rect 38988 21876 38994 21888
rect 39209 21879 39267 21885
rect 39209 21876 39221 21879
rect 38988 21848 39221 21876
rect 38988 21836 38994 21848
rect 39209 21845 39221 21848
rect 39255 21845 39267 21879
rect 39209 21839 39267 21845
rect 39666 21836 39672 21888
rect 39724 21836 39730 21888
rect 39758 21836 39764 21888
rect 39816 21876 39822 21888
rect 40589 21879 40647 21885
rect 40589 21876 40601 21879
rect 39816 21848 40601 21876
rect 39816 21836 39822 21848
rect 40589 21845 40601 21848
rect 40635 21876 40647 21879
rect 41325 21879 41383 21885
rect 41325 21876 41337 21879
rect 40635 21848 41337 21876
rect 40635 21845 40647 21848
rect 40589 21839 40647 21845
rect 41325 21845 41337 21848
rect 41371 21876 41383 21879
rect 41966 21876 41972 21888
rect 41371 21848 41972 21876
rect 41371 21845 41383 21848
rect 41325 21839 41383 21845
rect 41966 21836 41972 21848
rect 42024 21836 42030 21888
rect 42150 21836 42156 21888
rect 42208 21836 42214 21888
rect 42794 21836 42800 21888
rect 42852 21876 42858 21888
rect 43533 21879 43591 21885
rect 43533 21876 43545 21879
rect 42852 21848 43545 21876
rect 42852 21836 42858 21848
rect 43533 21845 43545 21848
rect 43579 21876 43591 21879
rect 43901 21879 43959 21885
rect 43901 21876 43913 21879
rect 43579 21848 43913 21876
rect 43579 21845 43591 21848
rect 43533 21839 43591 21845
rect 43901 21845 43913 21848
rect 43947 21845 43959 21879
rect 43901 21839 43959 21845
rect 460 21786 45540 21808
rect 460 21734 6070 21786
rect 6122 21734 6134 21786
rect 6186 21734 6198 21786
rect 6250 21734 6262 21786
rect 6314 21734 6326 21786
rect 6378 21734 11070 21786
rect 11122 21734 11134 21786
rect 11186 21734 11198 21786
rect 11250 21734 11262 21786
rect 11314 21734 11326 21786
rect 11378 21734 16070 21786
rect 16122 21734 16134 21786
rect 16186 21734 16198 21786
rect 16250 21734 16262 21786
rect 16314 21734 16326 21786
rect 16378 21734 21070 21786
rect 21122 21734 21134 21786
rect 21186 21734 21198 21786
rect 21250 21734 21262 21786
rect 21314 21734 21326 21786
rect 21378 21734 26070 21786
rect 26122 21734 26134 21786
rect 26186 21734 26198 21786
rect 26250 21734 26262 21786
rect 26314 21734 26326 21786
rect 26378 21734 31070 21786
rect 31122 21734 31134 21786
rect 31186 21734 31198 21786
rect 31250 21734 31262 21786
rect 31314 21734 31326 21786
rect 31378 21734 36070 21786
rect 36122 21734 36134 21786
rect 36186 21734 36198 21786
rect 36250 21734 36262 21786
rect 36314 21734 36326 21786
rect 36378 21734 41070 21786
rect 41122 21734 41134 21786
rect 41186 21734 41198 21786
rect 41250 21734 41262 21786
rect 41314 21734 41326 21786
rect 41378 21734 45540 21786
rect 460 21712 45540 21734
rect 10042 21632 10048 21684
rect 10100 21632 10106 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 14274 21672 14280 21684
rect 12299 21644 14280 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 16025 21675 16083 21681
rect 16025 21672 16037 21675
rect 14792 21644 16037 21672
rect 14792 21632 14798 21644
rect 16025 21641 16037 21644
rect 16071 21641 16083 21675
rect 18690 21672 18696 21684
rect 16025 21635 16083 21641
rect 16500 21644 18696 21672
rect 10060 21536 10088 21632
rect 11149 21607 11207 21613
rect 11149 21573 11161 21607
rect 11195 21604 11207 21607
rect 13906 21604 13912 21616
rect 11195 21576 13912 21604
rect 11195 21573 11207 21576
rect 11149 21567 11207 21573
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 15226 21590 15792 21604
rect 15212 21576 15792 21590
rect 13078 21536 13084 21548
rect 10060 21508 13084 21536
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 13817 21539 13875 21545
rect 13817 21536 13829 21539
rect 13771 21508 13829 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 13817 21505 13829 21508
rect 13863 21536 13875 21539
rect 13863 21508 14320 21536
rect 13863 21505 13875 21508
rect 13817 21499 13875 21505
rect 6089 21471 6147 21477
rect 6089 21437 6101 21471
rect 6135 21468 6147 21471
rect 6730 21468 6736 21480
rect 6135 21440 6736 21468
rect 6135 21437 6147 21440
rect 6089 21431 6147 21437
rect 6730 21428 6736 21440
rect 6788 21468 6794 21480
rect 7098 21468 7104 21480
rect 6788 21440 7104 21468
rect 6788 21428 6794 21440
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 10137 21471 10195 21477
rect 10137 21437 10149 21471
rect 10183 21468 10195 21471
rect 12066 21468 12072 21480
rect 10183 21440 12072 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 12066 21428 12072 21440
rect 12124 21428 12130 21480
rect 14182 21428 14188 21480
rect 14240 21428 14246 21480
rect 14292 21468 14320 21508
rect 14458 21468 14464 21480
rect 14292 21440 14464 21468
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 14550 21428 14556 21480
rect 14608 21468 14614 21480
rect 15212 21468 15240 21576
rect 15611 21539 15669 21545
rect 15611 21505 15623 21539
rect 15657 21505 15669 21539
rect 15764 21536 15792 21576
rect 15838 21564 15844 21616
rect 15896 21604 15902 21616
rect 16301 21607 16359 21613
rect 16301 21604 16313 21607
rect 15896 21576 16313 21604
rect 15896 21564 15902 21576
rect 16301 21573 16313 21576
rect 16347 21573 16359 21607
rect 16301 21567 16359 21573
rect 16390 21564 16396 21616
rect 16448 21564 16454 21616
rect 16500 21613 16528 21644
rect 18690 21632 18696 21644
rect 18748 21632 18754 21684
rect 18782 21632 18788 21684
rect 18840 21672 18846 21684
rect 18840 21644 19288 21672
rect 18840 21632 18846 21644
rect 16500 21607 16569 21613
rect 16500 21576 16523 21607
rect 16511 21573 16523 21576
rect 16557 21573 16569 21607
rect 17129 21607 17187 21613
rect 17129 21604 17141 21607
rect 16511 21567 16569 21573
rect 16776 21576 17141 21604
rect 15930 21536 15936 21548
rect 15764 21508 15936 21536
rect 15611 21499 15669 21505
rect 14608 21440 15240 21468
rect 15626 21468 15654 21499
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21505 16267 21539
rect 16209 21499 16267 21505
rect 15626 21440 15700 21468
rect 14608 21428 14614 21440
rect 15672 21412 15700 21440
rect 7837 21403 7895 21409
rect 7837 21400 7849 21403
rect 7116 21372 7849 21400
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 6365 21335 6423 21341
rect 6365 21332 6377 21335
rect 5960 21304 6377 21332
rect 5960 21292 5966 21304
rect 6365 21301 6377 21304
rect 6411 21301 6423 21335
rect 6365 21295 6423 21301
rect 6822 21292 6828 21344
rect 6880 21332 6886 21344
rect 7116 21341 7144 21372
rect 7837 21369 7849 21372
rect 7883 21400 7895 21403
rect 8205 21403 8263 21409
rect 8205 21400 8217 21403
rect 7883 21372 8217 21400
rect 7883 21369 7895 21372
rect 7837 21363 7895 21369
rect 8205 21369 8217 21372
rect 8251 21400 8263 21403
rect 8665 21403 8723 21409
rect 8665 21400 8677 21403
rect 8251 21372 8677 21400
rect 8251 21369 8263 21372
rect 8205 21363 8263 21369
rect 8665 21369 8677 21372
rect 8711 21400 8723 21403
rect 9306 21400 9312 21412
rect 8711 21372 9312 21400
rect 8711 21369 8723 21372
rect 8665 21363 8723 21369
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 11517 21403 11575 21409
rect 11517 21400 11529 21403
rect 9692 21372 11529 21400
rect 7101 21335 7159 21341
rect 7101 21332 7113 21335
rect 6880 21304 7113 21332
rect 6880 21292 6886 21304
rect 7101 21301 7113 21304
rect 7147 21301 7159 21335
rect 7101 21295 7159 21301
rect 7282 21292 7288 21344
rect 7340 21332 7346 21344
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 7340 21304 7481 21332
rect 7340 21292 7346 21304
rect 7469 21301 7481 21304
rect 7515 21332 7527 21335
rect 9033 21335 9091 21341
rect 9033 21332 9045 21335
rect 7515 21304 9045 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 9033 21301 9045 21304
rect 9079 21332 9091 21335
rect 9692 21332 9720 21372
rect 11517 21369 11529 21372
rect 11563 21400 11575 21403
rect 11885 21403 11943 21409
rect 11885 21400 11897 21403
rect 11563 21372 11897 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 11885 21369 11897 21372
rect 11931 21400 11943 21403
rect 11931 21372 13032 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 9079 21304 9720 21332
rect 9769 21335 9827 21341
rect 9079 21301 9091 21304
rect 9033 21295 9091 21301
rect 9769 21301 9781 21335
rect 9815 21332 9827 21335
rect 10226 21332 10232 21344
rect 9815 21304 10232 21332
rect 9815 21301 9827 21304
rect 9769 21295 9827 21301
rect 10226 21292 10232 21304
rect 10284 21292 10290 21344
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 11054 21332 11060 21344
rect 10551 21304 11060 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 12618 21292 12624 21344
rect 12676 21292 12682 21344
rect 13004 21341 13032 21372
rect 15470 21360 15476 21412
rect 15528 21360 15534 21412
rect 15654 21360 15660 21412
rect 15712 21360 15718 21412
rect 16224 21400 16252 21499
rect 16666 21496 16672 21548
rect 16724 21536 16730 21548
rect 16776 21536 16804 21576
rect 17129 21573 17141 21576
rect 17175 21604 17187 21607
rect 17957 21607 18015 21613
rect 17175 21576 17540 21604
rect 17175 21573 17187 21576
rect 17129 21567 17187 21573
rect 16724 21508 16804 21536
rect 16724 21496 16730 21508
rect 16850 21496 16856 21548
rect 16908 21536 16914 21548
rect 17512 21545 17540 21576
rect 17957 21573 17969 21607
rect 18003 21604 18015 21607
rect 18230 21604 18236 21616
rect 18003 21576 18236 21604
rect 18003 21573 18015 21576
rect 17957 21567 18015 21573
rect 18230 21564 18236 21576
rect 18288 21564 18294 21616
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16908 21508 16957 21536
rect 16908 21496 16914 21508
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21536 17279 21539
rect 17313 21539 17371 21545
rect 17313 21536 17325 21539
rect 17267 21508 17325 21536
rect 17267 21505 17279 21508
rect 17221 21499 17279 21505
rect 17313 21505 17325 21508
rect 17359 21505 17371 21539
rect 17313 21499 17371 21505
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 16298 21428 16304 21480
rect 16356 21468 16362 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 16356 21440 16773 21468
rect 16356 21428 16362 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 17328 21468 17356 21499
rect 17678 21496 17684 21548
rect 17736 21496 17742 21548
rect 17328 21440 17540 21468
rect 16761 21431 16819 21437
rect 17405 21403 17463 21409
rect 17405 21400 17417 21403
rect 16224 21372 17417 21400
rect 17405 21369 17417 21372
rect 17451 21369 17463 21403
rect 17405 21363 17463 21369
rect 12989 21335 13047 21341
rect 12989 21301 13001 21335
rect 13035 21332 13047 21335
rect 13354 21332 13360 21344
rect 13035 21304 13360 21332
rect 13035 21301 13047 21304
rect 12989 21295 13047 21301
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 15488 21332 15516 21360
rect 17512 21332 17540 21440
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18966 21468 18972 21480
rect 18104 21440 18972 21468
rect 18104 21428 18110 21440
rect 18966 21428 18972 21440
rect 19024 21468 19030 21480
rect 19076 21468 19104 21522
rect 19024 21440 19104 21468
rect 19260 21468 19288 21644
rect 19426 21632 19432 21684
rect 19484 21632 19490 21684
rect 19613 21675 19671 21681
rect 19613 21641 19625 21675
rect 19659 21672 19671 21675
rect 19886 21672 19892 21684
rect 19659 21644 19892 21672
rect 19659 21641 19671 21644
rect 19613 21635 19671 21641
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 20162 21632 20168 21684
rect 20220 21632 20226 21684
rect 20349 21675 20407 21681
rect 20349 21641 20361 21675
rect 20395 21672 20407 21675
rect 20622 21672 20628 21684
rect 20395 21644 20628 21672
rect 20395 21641 20407 21644
rect 20349 21635 20407 21641
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 21361 21675 21419 21681
rect 21361 21672 21373 21675
rect 20864 21644 21373 21672
rect 20864 21632 20870 21644
rect 21361 21641 21373 21644
rect 21407 21641 21419 21675
rect 21361 21635 21419 21641
rect 21652 21644 23336 21672
rect 19981 21607 20039 21613
rect 19981 21604 19993 21607
rect 19628 21576 19993 21604
rect 19628 21480 19656 21576
rect 19981 21573 19993 21576
rect 20027 21573 20039 21607
rect 20180 21604 20208 21632
rect 21652 21616 21680 21644
rect 20714 21604 20720 21616
rect 20180 21576 20720 21604
rect 19981 21567 20039 21573
rect 20714 21564 20720 21576
rect 20772 21604 20778 21616
rect 20772 21576 21496 21604
rect 20772 21564 20778 21576
rect 21468 21548 21496 21576
rect 21634 21564 21640 21616
rect 21692 21564 21698 21616
rect 22278 21604 22284 21616
rect 21744 21576 22284 21604
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19610 21468 19616 21480
rect 19260 21440 19616 21468
rect 19024 21428 19030 21440
rect 19610 21428 19616 21440
rect 19668 21428 19674 21480
rect 19812 21400 19840 21499
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20099 21539 20157 21545
rect 20099 21505 20111 21539
rect 20145 21505 20157 21539
rect 20099 21499 20157 21505
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20114 21468 20142 21499
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 20622 21496 20628 21548
rect 20680 21496 20686 21548
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21536 21235 21539
rect 21223 21508 21312 21536
rect 21223 21505 21235 21508
rect 21177 21499 21235 21505
rect 20036 21440 20142 21468
rect 20257 21471 20315 21477
rect 20036 21428 20042 21440
rect 20257 21437 20269 21471
rect 20303 21468 20315 21471
rect 20438 21468 20444 21480
rect 20303 21440 20444 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 20162 21400 20168 21412
rect 19812 21372 20168 21400
rect 20162 21360 20168 21372
rect 20220 21360 20226 21412
rect 20916 21400 20944 21431
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 20456 21372 20944 21400
rect 17954 21332 17960 21344
rect 15488 21304 17960 21332
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 20346 21332 20352 21344
rect 20036 21304 20352 21332
rect 20036 21292 20042 21304
rect 20346 21292 20352 21304
rect 20404 21332 20410 21344
rect 20456 21332 20484 21372
rect 21082 21360 21088 21412
rect 21140 21400 21146 21412
rect 21177 21403 21235 21409
rect 21177 21400 21189 21403
rect 21140 21372 21189 21400
rect 21140 21360 21146 21372
rect 21177 21369 21189 21372
rect 21223 21369 21235 21403
rect 21177 21363 21235 21369
rect 21284 21400 21312 21508
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 21744 21545 21772 21576
rect 22278 21564 22284 21576
rect 22336 21564 22342 21616
rect 22388 21604 22416 21644
rect 23308 21604 23336 21644
rect 23566 21632 23572 21684
rect 23624 21672 23630 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 23624 21644 25421 21672
rect 23624 21632 23630 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 25409 21635 25467 21641
rect 25774 21632 25780 21684
rect 25832 21632 25838 21684
rect 25866 21632 25872 21684
rect 25924 21632 25930 21684
rect 27614 21632 27620 21684
rect 27672 21672 27678 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27672 21644 28365 21672
rect 27672 21632 27678 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 28902 21632 28908 21684
rect 28960 21672 28966 21684
rect 29549 21675 29607 21681
rect 29549 21672 29561 21675
rect 28960 21644 29561 21672
rect 28960 21632 28966 21644
rect 29549 21641 29561 21644
rect 29595 21641 29607 21675
rect 29549 21635 29607 21641
rect 30374 21632 30380 21684
rect 30432 21632 30438 21684
rect 32582 21672 32588 21684
rect 31726 21644 32588 21672
rect 24118 21604 24124 21616
rect 22388 21576 22494 21604
rect 23308 21576 24124 21604
rect 24118 21564 24124 21576
rect 24176 21604 24182 21616
rect 24176 21576 24334 21604
rect 24176 21564 24182 21576
rect 25314 21564 25320 21616
rect 25372 21564 25378 21616
rect 25498 21564 25504 21616
rect 25556 21604 25562 21616
rect 26050 21604 26056 21616
rect 25556 21576 26056 21604
rect 25556 21564 25562 21576
rect 26050 21564 26056 21576
rect 26108 21604 26114 21616
rect 26108 21576 26234 21604
rect 26108 21564 26114 21576
rect 21729 21539 21787 21545
rect 21729 21536 21741 21539
rect 21600 21508 21741 21536
rect 21600 21496 21606 21508
rect 21729 21505 21741 21508
rect 21775 21505 21787 21539
rect 21729 21499 21787 21505
rect 22002 21428 22008 21480
rect 22060 21428 22066 21480
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 23569 21471 23627 21477
rect 23569 21468 23581 21471
rect 23256 21440 23581 21468
rect 23256 21428 23262 21440
rect 23569 21437 23581 21440
rect 23615 21437 23627 21471
rect 23934 21468 23940 21480
rect 23569 21431 23627 21437
rect 23676 21440 23940 21468
rect 23477 21403 23535 21409
rect 21284 21372 21772 21400
rect 20404 21304 20484 21332
rect 20404 21292 20410 21304
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 21284 21332 21312 21372
rect 21744 21344 21772 21372
rect 23477 21369 23489 21403
rect 23523 21400 23535 21403
rect 23676 21400 23704 21440
rect 23934 21428 23940 21440
rect 23992 21468 23998 21480
rect 24486 21468 24492 21480
rect 23992 21440 24492 21468
rect 23992 21428 23998 21440
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 25332 21477 25360 21564
rect 26206 21536 26234 21576
rect 26602 21564 26608 21616
rect 26660 21564 26666 21616
rect 29089 21607 29147 21613
rect 29089 21573 29101 21607
rect 29135 21604 29147 21607
rect 31726 21604 31754 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 33870 21632 33876 21684
rect 33928 21672 33934 21684
rect 35161 21675 35219 21681
rect 35161 21672 35173 21675
rect 33928 21644 35173 21672
rect 33928 21632 33934 21644
rect 35161 21641 35173 21644
rect 35207 21641 35219 21675
rect 35161 21635 35219 21641
rect 35989 21675 36047 21681
rect 35989 21641 36001 21675
rect 36035 21641 36047 21675
rect 35989 21635 36047 21641
rect 36265 21675 36323 21681
rect 36265 21641 36277 21675
rect 36311 21672 36323 21675
rect 36446 21672 36452 21684
rect 36311 21644 36452 21672
rect 36311 21641 36323 21644
rect 36265 21635 36323 21641
rect 34054 21604 34060 21616
rect 29135 21576 31754 21604
rect 32982 21590 34060 21604
rect 32968 21576 34060 21590
rect 29135 21573 29147 21576
rect 29089 21567 29147 21573
rect 26329 21539 26387 21545
rect 26329 21536 26341 21539
rect 26206 21508 26341 21536
rect 26329 21505 26341 21508
rect 26375 21505 26387 21539
rect 28169 21539 28227 21545
rect 26329 21499 26387 21505
rect 25317 21471 25375 21477
rect 25317 21437 25329 21471
rect 25363 21437 25375 21471
rect 25317 21431 25375 21437
rect 26053 21471 26111 21477
rect 26053 21437 26065 21471
rect 26099 21437 26111 21471
rect 27154 21468 27160 21480
rect 26053 21431 26111 21437
rect 26436 21440 27160 21468
rect 23523 21372 23704 21400
rect 26068 21400 26096 21431
rect 26436 21400 26464 21440
rect 27154 21428 27160 21440
rect 27212 21428 27218 21480
rect 27724 21468 27752 21522
rect 28169 21505 28181 21539
rect 28215 21536 28227 21539
rect 29181 21539 29239 21545
rect 28215 21508 28764 21536
rect 28215 21505 28227 21508
rect 28169 21499 28227 21505
rect 27890 21468 27896 21480
rect 27724 21440 27896 21468
rect 27890 21428 27896 21440
rect 27948 21468 27954 21480
rect 27948 21440 28304 21468
rect 27948 21428 27954 21440
rect 28276 21412 28304 21440
rect 26068 21372 26464 21400
rect 23523 21369 23535 21372
rect 23477 21363 23535 21369
rect 27798 21360 27804 21412
rect 27856 21400 27862 21412
rect 27856 21372 28212 21400
rect 27856 21360 27862 21372
rect 20588 21304 21312 21332
rect 20588 21292 20594 21304
rect 21726 21292 21732 21344
rect 21784 21292 21790 21344
rect 23842 21341 23848 21344
rect 23832 21335 23848 21341
rect 23832 21301 23844 21335
rect 23832 21295 23848 21301
rect 23842 21292 23848 21295
rect 23900 21292 23906 21344
rect 26970 21292 26976 21344
rect 27028 21332 27034 21344
rect 28074 21332 28080 21344
rect 27028 21304 28080 21332
rect 27028 21292 27034 21304
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 28184 21332 28212 21372
rect 28258 21360 28264 21412
rect 28316 21360 28322 21412
rect 28736 21409 28764 21508
rect 29181 21505 29193 21539
rect 29227 21536 29239 21539
rect 29362 21536 29368 21548
rect 29227 21508 29368 21536
rect 29227 21505 29239 21508
rect 29181 21499 29239 21505
rect 29362 21496 29368 21508
rect 29420 21496 29426 21548
rect 29914 21496 29920 21548
rect 29972 21496 29978 21548
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 30650 21536 30656 21548
rect 30055 21508 30656 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30742 21496 30748 21548
rect 30800 21496 30806 21548
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21536 30895 21539
rect 31018 21536 31024 21548
rect 30883 21508 31024 21536
rect 30883 21505 30895 21508
rect 30837 21499 30895 21505
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 29273 21471 29331 21477
rect 29273 21468 29285 21471
rect 28966 21440 29285 21468
rect 28721 21403 28779 21409
rect 28721 21369 28733 21403
rect 28767 21369 28779 21403
rect 28721 21363 28779 21369
rect 28966 21332 28994 21440
rect 29273 21437 29285 21440
rect 29319 21468 29331 21471
rect 30098 21468 30104 21480
rect 29319 21440 30104 21468
rect 29319 21437 29331 21440
rect 29273 21431 29331 21437
rect 30098 21428 30104 21440
rect 30156 21468 30162 21480
rect 30929 21471 30987 21477
rect 30929 21468 30941 21471
rect 30156 21440 30941 21468
rect 30156 21428 30162 21440
rect 30929 21437 30941 21440
rect 30975 21468 30987 21471
rect 31386 21468 31392 21480
rect 30975 21440 31392 21468
rect 30975 21437 30987 21440
rect 30929 21431 30987 21437
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 31481 21471 31539 21477
rect 31481 21437 31493 21471
rect 31527 21437 31539 21471
rect 31481 21431 31539 21437
rect 31757 21471 31815 21477
rect 31757 21437 31769 21471
rect 31803 21468 31815 21471
rect 32214 21468 32220 21480
rect 31803 21440 32220 21468
rect 31803 21437 31815 21440
rect 31757 21431 31815 21437
rect 30190 21360 30196 21412
rect 30248 21400 30254 21412
rect 30742 21400 30748 21412
rect 30248 21372 30748 21400
rect 30248 21360 30254 21372
rect 30742 21360 30748 21372
rect 30800 21360 30806 21412
rect 28184 21304 28994 21332
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31496 21332 31524 21431
rect 32214 21428 32220 21440
rect 32272 21428 32278 21480
rect 32306 21428 32312 21480
rect 32364 21468 32370 21480
rect 32968 21468 32996 21576
rect 34054 21564 34060 21576
rect 34112 21564 34118 21616
rect 36004 21604 36032 21635
rect 36446 21632 36452 21644
rect 36504 21632 36510 21684
rect 37918 21632 37924 21684
rect 37976 21672 37982 21684
rect 37976 21644 38240 21672
rect 37976 21632 37982 21644
rect 36909 21607 36967 21613
rect 36909 21604 36921 21607
rect 36004 21576 36921 21604
rect 36909 21573 36921 21576
rect 36955 21573 36967 21607
rect 38212 21604 38240 21644
rect 40494 21632 40500 21684
rect 40552 21672 40558 21684
rect 40681 21675 40739 21681
rect 40681 21672 40693 21675
rect 40552 21644 40693 21672
rect 40552 21632 40558 21644
rect 40681 21641 40693 21644
rect 40727 21641 40739 21675
rect 40681 21635 40739 21641
rect 40954 21632 40960 21684
rect 41012 21672 41018 21684
rect 41325 21675 41383 21681
rect 41325 21672 41337 21675
rect 41012 21644 41337 21672
rect 41012 21632 41018 21644
rect 41325 21641 41337 21644
rect 41371 21641 41383 21675
rect 41325 21635 41383 21641
rect 38749 21607 38807 21613
rect 38749 21604 38761 21607
rect 38212 21576 38761 21604
rect 36909 21567 36967 21573
rect 38749 21573 38761 21576
rect 38795 21573 38807 21607
rect 41340 21604 41368 21635
rect 41966 21632 41972 21684
rect 42024 21672 42030 21684
rect 42337 21675 42395 21681
rect 42337 21672 42349 21675
rect 42024 21644 42349 21672
rect 42024 21632 42030 21644
rect 42337 21641 42349 21644
rect 42383 21672 42395 21675
rect 42794 21672 42800 21684
rect 42383 21644 42800 21672
rect 42383 21641 42395 21644
rect 42337 21635 42395 21641
rect 42794 21632 42800 21644
rect 42852 21672 42858 21684
rect 43073 21675 43131 21681
rect 43073 21672 43085 21675
rect 42852 21644 43085 21672
rect 42852 21632 42858 21644
rect 43073 21641 43085 21644
rect 43119 21672 43131 21675
rect 44174 21672 44180 21684
rect 43119 21644 44180 21672
rect 43119 21641 43131 21644
rect 43073 21635 43131 21641
rect 44174 21632 44180 21644
rect 44232 21672 44238 21684
rect 44542 21672 44548 21684
rect 44232 21644 44548 21672
rect 44232 21632 44238 21644
rect 44542 21632 44548 21644
rect 44600 21632 44606 21684
rect 42705 21607 42763 21613
rect 42705 21604 42717 21607
rect 41340 21576 42717 21604
rect 38749 21567 38807 21573
rect 42705 21573 42717 21576
rect 42751 21604 42763 21607
rect 43809 21607 43867 21613
rect 43809 21604 43821 21607
rect 42751 21576 43821 21604
rect 42751 21573 42763 21576
rect 42705 21567 42763 21573
rect 43809 21573 43821 21576
rect 43855 21604 43867 21607
rect 43898 21604 43904 21616
rect 43855 21576 43904 21604
rect 43855 21573 43867 21576
rect 43809 21567 43867 21573
rect 43898 21564 43904 21576
rect 43956 21564 43962 21616
rect 35434 21536 35440 21548
rect 34730 21522 35440 21536
rect 34716 21508 35440 21522
rect 32364 21440 32996 21468
rect 32364 21428 32370 21440
rect 33134 21428 33140 21480
rect 33192 21468 33198 21480
rect 33318 21468 33324 21480
rect 33192 21440 33324 21468
rect 33192 21428 33198 21440
rect 33318 21428 33324 21440
rect 33376 21428 33382 21480
rect 33597 21471 33655 21477
rect 33597 21468 33609 21471
rect 33428 21440 33609 21468
rect 32858 21360 32864 21412
rect 32916 21400 32922 21412
rect 33428 21400 33456 21440
rect 33597 21437 33609 21440
rect 33643 21437 33655 21471
rect 33597 21431 33655 21437
rect 34054 21428 34060 21480
rect 34112 21468 34118 21480
rect 34716 21468 34744 21508
rect 35434 21496 35440 21508
rect 35492 21496 35498 21548
rect 35526 21496 35532 21548
rect 35584 21496 35590 21548
rect 35894 21496 35900 21548
rect 35952 21536 35958 21548
rect 36173 21539 36231 21545
rect 36173 21536 36185 21539
rect 35952 21508 36185 21536
rect 35952 21496 35958 21508
rect 36173 21505 36185 21508
rect 36219 21505 36231 21539
rect 36173 21499 36231 21505
rect 36446 21496 36452 21548
rect 36504 21496 36510 21548
rect 36538 21496 36544 21548
rect 36596 21496 36602 21548
rect 37918 21496 37924 21548
rect 37976 21536 37982 21548
rect 37976 21508 38042 21536
rect 37976 21496 37982 21508
rect 39758 21496 39764 21548
rect 39816 21536 39822 21548
rect 39816 21508 39882 21536
rect 39816 21496 39822 21508
rect 34112 21440 34744 21468
rect 34112 21428 34118 21440
rect 34974 21428 34980 21480
rect 35032 21468 35038 21480
rect 35618 21468 35624 21480
rect 35032 21440 35624 21468
rect 35032 21428 35038 21440
rect 35618 21428 35624 21440
rect 35676 21428 35682 21480
rect 35710 21428 35716 21480
rect 35768 21428 35774 21480
rect 36556 21468 36584 21496
rect 36633 21471 36691 21477
rect 36633 21468 36645 21471
rect 36556 21440 36645 21468
rect 36633 21437 36645 21440
rect 36679 21437 36691 21471
rect 36633 21431 36691 21437
rect 37458 21428 37464 21480
rect 37516 21468 37522 21480
rect 38378 21468 38384 21480
rect 37516 21440 38384 21468
rect 37516 21428 37522 21440
rect 38378 21428 38384 21440
rect 38436 21468 38442 21480
rect 38473 21471 38531 21477
rect 38473 21468 38485 21471
rect 38436 21440 38485 21468
rect 38436 21428 38442 21440
rect 38473 21437 38485 21440
rect 38519 21437 38531 21471
rect 38473 21431 38531 21437
rect 38580 21440 40356 21468
rect 32916 21372 33456 21400
rect 32916 21360 32922 21372
rect 38010 21360 38016 21412
rect 38068 21400 38074 21412
rect 38580 21400 38608 21440
rect 40328 21409 40356 21440
rect 40770 21428 40776 21480
rect 40828 21428 40834 21480
rect 40862 21428 40868 21480
rect 40920 21428 40926 21480
rect 38068 21372 38608 21400
rect 40221 21403 40279 21409
rect 38068 21360 38074 21372
rect 40221 21369 40233 21403
rect 40267 21369 40279 21403
rect 40221 21363 40279 21369
rect 40313 21403 40371 21409
rect 40313 21369 40325 21403
rect 40359 21369 40371 21403
rect 40313 21363 40371 21369
rect 31938 21332 31944 21344
rect 30984 21304 31944 21332
rect 30984 21292 30990 21304
rect 31938 21292 31944 21304
rect 31996 21292 32002 21344
rect 32122 21292 32128 21344
rect 32180 21332 32186 21344
rect 33042 21332 33048 21344
rect 32180 21304 33048 21332
rect 32180 21292 32186 21304
rect 33042 21292 33048 21304
rect 33100 21292 33106 21344
rect 33226 21292 33232 21344
rect 33284 21292 33290 21344
rect 33410 21292 33416 21344
rect 33468 21332 33474 21344
rect 33686 21332 33692 21344
rect 33468 21304 33692 21332
rect 33468 21292 33474 21304
rect 33686 21292 33692 21304
rect 33744 21332 33750 21344
rect 35069 21335 35127 21341
rect 35069 21332 35081 21335
rect 33744 21304 35081 21332
rect 33744 21292 33750 21304
rect 35069 21301 35081 21304
rect 35115 21301 35127 21335
rect 35069 21295 35127 21301
rect 36906 21292 36912 21344
rect 36964 21332 36970 21344
rect 38381 21335 38439 21341
rect 38381 21332 38393 21335
rect 36964 21304 38393 21332
rect 36964 21292 36970 21304
rect 38381 21301 38393 21304
rect 38427 21301 38439 21335
rect 38381 21295 38439 21301
rect 38470 21292 38476 21344
rect 38528 21332 38534 21344
rect 40236 21332 40264 21363
rect 40494 21360 40500 21412
rect 40552 21400 40558 21412
rect 40552 21372 42196 21400
rect 40552 21360 40558 21372
rect 42168 21344 42196 21372
rect 38528 21304 40264 21332
rect 38528 21292 38534 21304
rect 42150 21292 42156 21344
rect 42208 21332 42214 21344
rect 43441 21335 43499 21341
rect 43441 21332 43453 21335
rect 42208 21304 43453 21332
rect 42208 21292 42214 21304
rect 43441 21301 43453 21304
rect 43487 21332 43499 21335
rect 44266 21332 44272 21344
rect 43487 21304 44272 21332
rect 43487 21301 43499 21304
rect 43441 21295 43499 21301
rect 44266 21292 44272 21304
rect 44324 21292 44330 21344
rect 44910 21292 44916 21344
rect 44968 21292 44974 21344
rect 460 21242 45540 21264
rect 460 21190 3570 21242
rect 3622 21190 3634 21242
rect 3686 21190 3698 21242
rect 3750 21190 3762 21242
rect 3814 21190 3826 21242
rect 3878 21190 8570 21242
rect 8622 21190 8634 21242
rect 8686 21190 8698 21242
rect 8750 21190 8762 21242
rect 8814 21190 8826 21242
rect 8878 21190 13570 21242
rect 13622 21190 13634 21242
rect 13686 21190 13698 21242
rect 13750 21190 13762 21242
rect 13814 21190 13826 21242
rect 13878 21190 18570 21242
rect 18622 21190 18634 21242
rect 18686 21190 18698 21242
rect 18750 21190 18762 21242
rect 18814 21190 18826 21242
rect 18878 21190 23570 21242
rect 23622 21190 23634 21242
rect 23686 21190 23698 21242
rect 23750 21190 23762 21242
rect 23814 21190 23826 21242
rect 23878 21190 28570 21242
rect 28622 21190 28634 21242
rect 28686 21190 28698 21242
rect 28750 21190 28762 21242
rect 28814 21190 28826 21242
rect 28878 21190 33570 21242
rect 33622 21190 33634 21242
rect 33686 21190 33698 21242
rect 33750 21190 33762 21242
rect 33814 21190 33826 21242
rect 33878 21190 38570 21242
rect 38622 21190 38634 21242
rect 38686 21190 38698 21242
rect 38750 21190 38762 21242
rect 38814 21190 38826 21242
rect 38878 21190 43570 21242
rect 43622 21190 43634 21242
rect 43686 21190 43698 21242
rect 43750 21190 43762 21242
rect 43814 21190 43826 21242
rect 43878 21190 45540 21242
rect 460 21168 45540 21190
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 13725 21131 13783 21137
rect 13725 21128 13737 21131
rect 12768 21100 13737 21128
rect 12768 21088 12774 21100
rect 13725 21097 13737 21100
rect 13771 21128 13783 21131
rect 13998 21128 14004 21140
rect 13771 21100 14004 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 14461 21131 14519 21137
rect 14461 21097 14473 21131
rect 14507 21128 14519 21131
rect 14550 21128 14556 21140
rect 14507 21100 14556 21128
rect 14507 21097 14519 21100
rect 14461 21091 14519 21097
rect 12529 21063 12587 21069
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 13354 21060 13360 21072
rect 12575 21032 13360 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 13354 21020 13360 21032
rect 13412 21060 13418 21072
rect 13814 21060 13820 21072
rect 13412 21032 13820 21060
rect 13412 21020 13418 21032
rect 13814 21020 13820 21032
rect 13872 21060 13878 21072
rect 14476 21060 14504 21091
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 15470 21128 15476 21140
rect 14936 21100 15476 21128
rect 13872 21032 14504 21060
rect 13872 21020 13878 21032
rect 8113 20995 8171 21001
rect 8113 20961 8125 20995
rect 8159 20992 8171 20995
rect 9217 20995 9275 21001
rect 9217 20992 9229 20995
rect 8159 20964 9229 20992
rect 8159 20961 8171 20964
rect 8113 20955 8171 20961
rect 9217 20961 9229 20964
rect 9263 20961 9275 20995
rect 14936 20992 14964 21100
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 17678 21128 17684 21140
rect 15620 21100 17684 21128
rect 15620 21088 15626 21100
rect 16684 21001 16712 21100
rect 17678 21088 17684 21100
rect 17736 21088 17742 21140
rect 19337 21131 19395 21137
rect 19337 21128 19349 21131
rect 18984 21100 19349 21128
rect 18601 21063 18659 21069
rect 18601 21029 18613 21063
rect 18647 21029 18659 21063
rect 18601 21023 18659 21029
rect 9217 20955 9275 20961
rect 14568 20964 14964 20992
rect 15105 20995 15163 21001
rect 934 20884 940 20936
rect 992 20884 998 20936
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 6196 20896 6377 20924
rect 6196 20865 6224 20896
rect 6365 20893 6377 20896
rect 6411 20893 6423 20927
rect 6365 20887 6423 20893
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 6181 20859 6239 20865
rect 6181 20856 6193 20859
rect 5644 20828 6193 20856
rect 5644 20800 5672 20828
rect 6181 20825 6193 20828
rect 6227 20825 6239 20859
rect 6181 20819 6239 20825
rect 6638 20816 6644 20868
rect 6696 20816 6702 20868
rect 7926 20856 7932 20868
rect 7866 20828 7932 20856
rect 7926 20816 7932 20828
rect 7984 20816 7990 20868
rect 8956 20856 8984 20887
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 11112 20896 11437 20924
rect 11112 20884 11118 20896
rect 11425 20893 11437 20896
rect 11471 20924 11483 20927
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11471 20896 11805 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 11793 20893 11805 20896
rect 11839 20924 11851 20927
rect 11882 20924 11888 20936
rect 11839 20896 11888 20924
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 11882 20884 11888 20896
rect 11940 20924 11946 20936
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 11940 20896 12173 20924
rect 11940 20884 11946 20896
rect 12161 20893 12173 20896
rect 12207 20924 12219 20927
rect 12207 20896 12940 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 9306 20856 9312 20868
rect 8956 20828 9312 20856
rect 9306 20816 9312 20828
rect 9364 20816 9370 20868
rect 10226 20816 10232 20868
rect 10284 20816 10290 20868
rect 12912 20865 12940 20896
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 14568 20933 14596 20964
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 16669 20995 16727 21001
rect 15151 20964 16620 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 14424 20896 14565 20924
rect 14424 20884 14430 20896
rect 14553 20893 14565 20896
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 14734 20884 14740 20936
rect 14792 20884 14798 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 12897 20859 12955 20865
rect 10612 20828 12756 20856
rect 750 20748 756 20800
rect 808 20748 814 20800
rect 3142 20748 3148 20800
rect 3200 20788 3206 20800
rect 3697 20791 3755 20797
rect 3697 20788 3709 20791
rect 3200 20760 3709 20788
rect 3200 20748 3206 20760
rect 3697 20757 3709 20760
rect 3743 20788 3755 20791
rect 3786 20788 3792 20800
rect 3743 20760 3792 20788
rect 3743 20757 3755 20760
rect 3697 20751 3755 20757
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 5534 20748 5540 20800
rect 5592 20748 5598 20800
rect 5626 20748 5632 20800
rect 5684 20748 5690 20800
rect 5902 20748 5908 20800
rect 5960 20748 5966 20800
rect 8849 20791 8907 20797
rect 8849 20757 8861 20791
rect 8895 20788 8907 20791
rect 10612 20788 10640 20828
rect 12728 20800 12756 20828
rect 12897 20825 12909 20859
rect 12943 20856 12955 20859
rect 13265 20859 13323 20865
rect 13265 20856 13277 20859
rect 12943 20828 13277 20856
rect 12943 20825 12955 20828
rect 12897 20819 12955 20825
rect 13265 20825 13277 20828
rect 13311 20856 13323 20859
rect 13538 20856 13544 20868
rect 13311 20828 13544 20856
rect 13311 20825 13323 20828
rect 13265 20819 13323 20825
rect 13538 20816 13544 20828
rect 13596 20856 13602 20868
rect 14093 20859 14151 20865
rect 14093 20856 14105 20859
rect 13596 20828 14105 20856
rect 13596 20816 13602 20828
rect 14093 20825 14105 20828
rect 14139 20856 14151 20859
rect 14458 20856 14464 20868
rect 14139 20828 14464 20856
rect 14139 20825 14151 20828
rect 14093 20819 14151 20825
rect 14458 20816 14464 20828
rect 14516 20856 14522 20868
rect 14844 20856 14872 20887
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16482 20924 16488 20936
rect 16172 20896 16488 20924
rect 16172 20884 16178 20896
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 15378 20856 15384 20868
rect 14516 20828 15384 20856
rect 14516 20816 14522 20828
rect 15378 20816 15384 20828
rect 15436 20816 15442 20868
rect 16592 20856 16620 20964
rect 16669 20961 16681 20995
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20992 17003 20995
rect 18616 20992 18644 21023
rect 18984 20992 19012 21100
rect 19337 21097 19349 21100
rect 19383 21097 19395 21131
rect 19337 21091 19395 21097
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 23201 21131 23259 21137
rect 23201 21128 23213 21131
rect 22060 21100 23213 21128
rect 22060 21088 22066 21100
rect 23201 21097 23213 21100
rect 23247 21097 23259 21131
rect 23201 21091 23259 21097
rect 25501 21131 25559 21137
rect 25501 21097 25513 21131
rect 25547 21128 25559 21131
rect 25866 21128 25872 21140
rect 25547 21100 25872 21128
rect 25547 21097 25559 21100
rect 25501 21091 25559 21097
rect 25866 21088 25872 21100
rect 25924 21088 25930 21140
rect 26510 21088 26516 21140
rect 26568 21088 26574 21140
rect 26712 21100 30512 21128
rect 19518 21060 19524 21072
rect 19168 21032 19524 21060
rect 19168 21001 19196 21032
rect 19518 21020 19524 21032
rect 19576 21060 19582 21072
rect 19978 21060 19984 21072
rect 19576 21032 19984 21060
rect 19576 21020 19582 21032
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 21726 21020 21732 21072
rect 21784 21060 21790 21072
rect 22833 21063 22891 21069
rect 22833 21060 22845 21063
rect 21784 21032 22845 21060
rect 21784 21020 21790 21032
rect 22833 21029 22845 21032
rect 22879 21029 22891 21063
rect 22833 21023 22891 21029
rect 16991 20964 18644 20992
rect 18892 20964 19012 20992
rect 19153 20995 19211 21001
rect 16991 20961 17003 20964
rect 16945 20955 17003 20961
rect 18892 20933 18920 20964
rect 19153 20961 19165 20995
rect 19199 20961 19211 20995
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19153 20955 19211 20961
rect 19444 20964 19625 20992
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 16850 20856 16856 20868
rect 16592 20828 16856 20856
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 17402 20816 17408 20868
rect 17460 20816 17466 20868
rect 18800 20856 18828 20887
rect 18966 20884 18972 20936
rect 19024 20924 19030 20936
rect 19444 20924 19472 20964
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 19613 20955 19671 20961
rect 19797 20995 19855 21001
rect 19797 20961 19809 20995
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 20441 20995 20499 21001
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 20487 20964 21772 20992
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 19024 20896 19472 20924
rect 19024 20884 19030 20896
rect 19518 20884 19524 20936
rect 19576 20884 19582 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19245 20859 19303 20865
rect 19245 20856 19257 20859
rect 18248 20828 18828 20856
rect 18892 20828 19257 20856
rect 8895 20760 10640 20788
rect 10689 20791 10747 20797
rect 8895 20757 8907 20760
rect 8849 20751 8907 20757
rect 10689 20757 10701 20791
rect 10735 20788 10747 20791
rect 11422 20788 11428 20800
rect 10735 20760 11428 20788
rect 10735 20757 10747 20760
rect 10689 20751 10747 20757
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 12710 20748 12716 20800
rect 12768 20748 12774 20800
rect 14737 20791 14795 20797
rect 14737 20757 14749 20791
rect 14783 20788 14795 20791
rect 15102 20788 15108 20800
rect 14783 20760 15108 20788
rect 14783 20757 14795 20760
rect 14737 20751 14795 20757
rect 15102 20748 15108 20760
rect 15160 20748 15166 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16390 20788 16396 20800
rect 15988 20760 16396 20788
rect 15988 20748 15994 20760
rect 16390 20748 16396 20760
rect 16448 20748 16454 20800
rect 16574 20748 16580 20800
rect 16632 20748 16638 20800
rect 17770 20748 17776 20800
rect 17828 20788 17834 20800
rect 18248 20788 18276 20828
rect 17828 20760 18276 20788
rect 17828 20748 17834 20760
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18417 20791 18475 20797
rect 18417 20788 18429 20791
rect 18380 20760 18429 20788
rect 18380 20748 18386 20760
rect 18417 20757 18429 20760
rect 18463 20788 18475 20791
rect 18892 20788 18920 20828
rect 19245 20825 19257 20828
rect 19291 20825 19303 20859
rect 19245 20819 19303 20825
rect 18463 20760 18920 20788
rect 18463 20757 18475 20760
rect 18417 20751 18475 20757
rect 19058 20748 19064 20800
rect 19116 20788 19122 20800
rect 19720 20788 19748 20887
rect 19812 20856 19840 20955
rect 21744 20936 21772 20964
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 22060 20964 22385 20992
rect 22060 20952 22066 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 23474 20952 23480 21004
rect 23532 20992 23538 21004
rect 24029 20995 24087 21001
rect 24029 20992 24041 20995
rect 23532 20964 24041 20992
rect 23532 20952 23538 20964
rect 24029 20961 24041 20964
rect 24075 20961 24087 20995
rect 24029 20955 24087 20961
rect 24762 20952 24768 21004
rect 24820 20992 24826 21004
rect 26329 20995 26387 21001
rect 26329 20992 26341 20995
rect 24820 20964 26341 20992
rect 24820 20952 24826 20964
rect 26329 20961 26341 20964
rect 26375 20992 26387 20995
rect 26712 20992 26740 21100
rect 27338 21020 27344 21072
rect 27396 21020 27402 21072
rect 28350 21020 28356 21072
rect 28408 21060 28414 21072
rect 28902 21060 28908 21072
rect 28408 21032 28908 21060
rect 28408 21020 28414 21032
rect 28902 21020 28908 21032
rect 28960 21020 28966 21072
rect 26375 20964 26740 20992
rect 26375 20961 26387 20964
rect 26329 20955 26387 20961
rect 26970 20952 26976 21004
rect 27028 20952 27034 21004
rect 27154 20952 27160 21004
rect 27212 20952 27218 21004
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 27893 20995 27951 21001
rect 27893 20992 27905 20995
rect 27856 20964 27905 20992
rect 27856 20952 27862 20964
rect 27893 20961 27905 20964
rect 27939 20961 27951 20995
rect 30484 20992 30512 21100
rect 30742 21088 30748 21140
rect 30800 21088 30806 21140
rect 31938 21088 31944 21140
rect 31996 21088 32002 21140
rect 32214 21088 32220 21140
rect 32272 21128 32278 21140
rect 32585 21131 32643 21137
rect 32585 21128 32597 21131
rect 32272 21100 32597 21128
rect 32272 21088 32278 21100
rect 32585 21097 32597 21100
rect 32631 21097 32643 21131
rect 32585 21091 32643 21097
rect 32858 21088 32864 21140
rect 32916 21088 32922 21140
rect 33042 21088 33048 21140
rect 33100 21128 33106 21140
rect 33100 21100 33824 21128
rect 33100 21088 33106 21100
rect 30558 21020 30564 21072
rect 30616 21060 30622 21072
rect 30653 21063 30711 21069
rect 30653 21060 30665 21063
rect 30616 21032 30665 21060
rect 30616 21020 30622 21032
rect 30653 21029 30665 21032
rect 30699 21029 30711 21063
rect 31956 21060 31984 21088
rect 33134 21060 33140 21072
rect 30653 21023 30711 21029
rect 31312 21032 31892 21060
rect 31956 21032 33140 21060
rect 31312 20992 31340 21032
rect 27893 20955 27951 20961
rect 28276 20964 30420 20992
rect 30484 20964 31340 20992
rect 31389 20995 31447 21001
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20180 20924 20392 20934
rect 20027 20906 20484 20924
rect 20027 20896 20208 20906
rect 20364 20896 20484 20906
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20070 20856 20076 20868
rect 19812 20828 20076 20856
rect 20070 20816 20076 20828
rect 20128 20816 20134 20868
rect 20162 20816 20168 20868
rect 20220 20816 20226 20868
rect 20456 20856 20484 20896
rect 21726 20884 21732 20936
rect 21784 20884 21790 20936
rect 22462 20884 22468 20936
rect 22520 20884 22526 20936
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 22612 20896 22937 20924
rect 22612 20884 22618 20896
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23106 20884 23112 20936
rect 23164 20884 23170 20936
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 23753 20927 23811 20933
rect 23753 20893 23765 20927
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 20717 20859 20775 20865
rect 20456 20828 20576 20856
rect 20548 20800 20576 20828
rect 20717 20825 20729 20859
rect 20763 20825 20775 20859
rect 20717 20819 20775 20825
rect 19116 20760 19748 20788
rect 19116 20748 19122 20760
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 20254 20788 20260 20800
rect 20036 20760 20260 20788
rect 20036 20748 20042 20760
rect 20254 20748 20260 20760
rect 20312 20788 20318 20800
rect 20349 20791 20407 20797
rect 20349 20788 20361 20791
rect 20312 20760 20361 20788
rect 20312 20748 20318 20760
rect 20349 20757 20361 20760
rect 20395 20757 20407 20791
rect 20349 20751 20407 20757
rect 20530 20748 20536 20800
rect 20588 20748 20594 20800
rect 20732 20788 20760 20819
rect 20990 20816 20996 20868
rect 21048 20816 21054 20868
rect 21174 20816 21180 20868
rect 21232 20816 21238 20868
rect 23198 20816 23204 20868
rect 23256 20856 23262 20868
rect 23768 20856 23796 20887
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 25372 20896 26065 20924
rect 25372 20884 25378 20896
rect 26053 20893 26065 20896
rect 26099 20924 26111 20927
rect 26881 20927 26939 20933
rect 26881 20924 26893 20927
rect 26099 20896 26893 20924
rect 26099 20893 26111 20896
rect 26053 20887 26111 20893
rect 26881 20893 26893 20896
rect 26927 20893 26939 20927
rect 26881 20887 26939 20893
rect 27709 20927 27767 20933
rect 27709 20893 27721 20927
rect 27755 20924 27767 20927
rect 27982 20924 27988 20936
rect 27755 20896 27988 20924
rect 27755 20893 27767 20896
rect 27709 20887 27767 20893
rect 27982 20884 27988 20896
rect 28040 20884 28046 20936
rect 28166 20884 28172 20936
rect 28224 20884 28230 20936
rect 24302 20856 24308 20868
rect 23256 20828 24308 20856
rect 23256 20816 23262 20828
rect 24302 20816 24308 20828
rect 24360 20816 24366 20868
rect 26145 20859 26203 20865
rect 24412 20828 24518 20856
rect 25608 20828 25820 20856
rect 20898 20788 20904 20800
rect 20732 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21008 20788 21036 20816
rect 21726 20788 21732 20800
rect 21008 20760 21732 20788
rect 21726 20748 21732 20760
rect 21784 20788 21790 20800
rect 22189 20791 22247 20797
rect 22189 20788 22201 20791
rect 21784 20760 22201 20788
rect 21784 20748 21790 20760
rect 22189 20757 22201 20760
rect 22235 20788 22247 20791
rect 22462 20788 22468 20800
rect 22235 20760 22468 20788
rect 22235 20757 22247 20760
rect 22189 20751 22247 20757
rect 22462 20748 22468 20760
rect 22520 20748 22526 20800
rect 23014 20748 23020 20800
rect 23072 20748 23078 20800
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 24412 20788 24440 20828
rect 25608 20788 25636 20828
rect 24176 20760 25636 20788
rect 24176 20748 24182 20760
rect 25682 20748 25688 20800
rect 25740 20748 25746 20800
rect 25792 20788 25820 20828
rect 26145 20825 26157 20859
rect 26191 20856 26203 20859
rect 27062 20856 27068 20868
rect 26191 20828 27068 20856
rect 26191 20825 26203 20828
rect 26145 20819 26203 20825
rect 27062 20816 27068 20828
rect 27120 20856 27126 20868
rect 28276 20856 28304 20964
rect 28537 20927 28595 20933
rect 28537 20893 28549 20927
rect 28583 20924 28595 20927
rect 28810 20924 28816 20936
rect 28583 20896 28816 20924
rect 28583 20893 28595 20896
rect 28537 20887 28595 20893
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 28902 20884 28908 20936
rect 28960 20884 28966 20936
rect 30282 20884 30288 20936
rect 30340 20884 30346 20936
rect 30392 20924 30420 20964
rect 31389 20961 31401 20995
rect 31435 20992 31447 20995
rect 31478 20992 31484 21004
rect 31435 20964 31484 20992
rect 31435 20961 31447 20964
rect 31389 20955 31447 20961
rect 31478 20952 31484 20964
rect 31536 20952 31542 21004
rect 31864 20992 31892 21032
rect 33134 21020 33140 21032
rect 33192 21060 33198 21072
rect 33192 21032 33732 21060
rect 33192 21020 33198 21032
rect 32309 20995 32367 21001
rect 32309 20992 32321 20995
rect 31864 20964 32321 20992
rect 32309 20961 32321 20964
rect 32355 20992 32367 20995
rect 33318 20992 33324 21004
rect 32355 20964 33324 20992
rect 32355 20961 32367 20964
rect 32309 20955 32367 20961
rect 33318 20952 33324 20964
rect 33376 20952 33382 21004
rect 33410 20952 33416 21004
rect 33468 20992 33474 21004
rect 33597 20995 33655 21001
rect 33597 20992 33609 20995
rect 33468 20964 33609 20992
rect 33468 20952 33474 20964
rect 33597 20961 33609 20964
rect 33643 20961 33655 20995
rect 33597 20955 33655 20961
rect 30392 20896 30512 20924
rect 27120 20828 28304 20856
rect 27120 20816 27126 20828
rect 28350 20816 28356 20868
rect 28408 20816 28414 20868
rect 28445 20859 28503 20865
rect 28445 20825 28457 20859
rect 28491 20856 28503 20859
rect 28491 20828 29132 20856
rect 28491 20825 28503 20828
rect 28445 20819 28503 20825
rect 27614 20788 27620 20800
rect 25792 20760 27620 20788
rect 27614 20748 27620 20760
rect 27672 20748 27678 20800
rect 27801 20791 27859 20797
rect 27801 20757 27813 20791
rect 27847 20788 27859 20791
rect 28074 20788 28080 20800
rect 27847 20760 28080 20788
rect 27847 20757 27859 20760
rect 27801 20751 27859 20757
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 29104 20788 29132 20828
rect 29178 20816 29184 20868
rect 29236 20816 29242 20868
rect 30484 20856 30512 20896
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 32769 20927 32827 20933
rect 32769 20924 32781 20927
rect 31812 20896 32781 20924
rect 31812 20884 31818 20896
rect 32769 20893 32781 20896
rect 32815 20893 32827 20927
rect 32769 20887 32827 20893
rect 33045 20927 33103 20933
rect 33045 20893 33057 20927
rect 33091 20924 33103 20927
rect 33704 20924 33732 21032
rect 33796 21001 33824 21100
rect 34514 21088 34520 21140
rect 34572 21128 34578 21140
rect 35526 21128 35532 21140
rect 34572 21100 35532 21128
rect 34572 21088 34578 21100
rect 35526 21088 35532 21100
rect 35584 21128 35590 21140
rect 35805 21131 35863 21137
rect 35805 21128 35817 21131
rect 35584 21100 35817 21128
rect 35584 21088 35590 21100
rect 35805 21097 35817 21100
rect 35851 21097 35863 21131
rect 35805 21091 35863 21097
rect 37274 21088 37280 21140
rect 37332 21128 37338 21140
rect 37737 21131 37795 21137
rect 37737 21128 37749 21131
rect 37332 21100 37749 21128
rect 37332 21088 37338 21100
rect 37737 21097 37749 21100
rect 37783 21097 37795 21131
rect 37737 21091 37795 21097
rect 38286 21088 38292 21140
rect 38344 21088 38350 21140
rect 40494 21128 40500 21140
rect 38396 21100 40500 21128
rect 37645 21063 37703 21069
rect 37645 21029 37657 21063
rect 37691 21060 37703 21063
rect 38304 21060 38332 21088
rect 37691 21032 38332 21060
rect 37691 21029 37703 21032
rect 37645 21023 37703 21029
rect 33781 20995 33839 21001
rect 33781 20961 33793 20995
rect 33827 20992 33839 20995
rect 33962 20992 33968 21004
rect 33827 20964 33968 20992
rect 33827 20961 33839 20964
rect 33781 20955 33839 20961
rect 33962 20952 33968 20964
rect 34020 20952 34026 21004
rect 35897 20995 35955 21001
rect 35897 20992 35909 20995
rect 34072 20964 35909 20992
rect 34072 20933 34100 20964
rect 35897 20961 35909 20964
rect 35943 20961 35955 20995
rect 35897 20955 35955 20961
rect 36170 20952 36176 21004
rect 36228 20952 36234 21004
rect 37366 20992 37372 21004
rect 37200 20964 37372 20992
rect 34057 20927 34115 20933
rect 34057 20924 34069 20927
rect 33091 20896 33180 20924
rect 33704 20896 34069 20924
rect 33091 20893 33103 20896
rect 33045 20887 33103 20893
rect 31846 20856 31852 20868
rect 30484 20828 31852 20856
rect 31846 20816 31852 20828
rect 31904 20856 31910 20868
rect 32125 20859 32183 20865
rect 32125 20856 32137 20859
rect 31904 20828 32137 20856
rect 31904 20816 31910 20828
rect 32125 20825 32137 20828
rect 32171 20825 32183 20859
rect 32125 20819 32183 20825
rect 32217 20859 32275 20865
rect 32217 20825 32229 20859
rect 32263 20856 32275 20859
rect 32582 20856 32588 20868
rect 32263 20828 32588 20856
rect 32263 20825 32275 20828
rect 32217 20819 32275 20825
rect 32582 20816 32588 20828
rect 32640 20816 32646 20868
rect 29362 20788 29368 20800
rect 29104 20760 29368 20788
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 30098 20748 30104 20800
rect 30156 20788 30162 20800
rect 31205 20791 31263 20797
rect 31205 20788 31217 20791
rect 30156 20760 31217 20788
rect 30156 20748 30162 20760
rect 31205 20757 31217 20760
rect 31251 20757 31263 20791
rect 31205 20751 31263 20757
rect 31754 20748 31760 20800
rect 31812 20748 31818 20800
rect 33152 20797 33180 20896
rect 34057 20893 34069 20896
rect 34103 20893 34115 20927
rect 34057 20887 34115 20893
rect 35434 20884 35440 20936
rect 35492 20884 35498 20936
rect 33410 20816 33416 20868
rect 33468 20856 33474 20868
rect 34333 20859 34391 20865
rect 34333 20856 34345 20859
rect 33468 20828 34345 20856
rect 33468 20816 33474 20828
rect 34333 20825 34345 20828
rect 34379 20825 34391 20859
rect 34333 20819 34391 20825
rect 33137 20791 33195 20797
rect 33137 20757 33149 20791
rect 33183 20757 33195 20791
rect 33137 20751 33195 20757
rect 33226 20748 33232 20800
rect 33284 20788 33290 20800
rect 33505 20791 33563 20797
rect 33505 20788 33517 20791
rect 33284 20760 33517 20788
rect 33284 20748 33290 20760
rect 33505 20757 33517 20760
rect 33551 20788 33563 20791
rect 34054 20788 34060 20800
rect 33551 20760 34060 20788
rect 33551 20757 33563 20760
rect 33505 20751 33563 20757
rect 34054 20748 34060 20760
rect 34112 20748 34118 20800
rect 35452 20788 35480 20884
rect 35986 20788 35992 20800
rect 35452 20760 35992 20788
rect 35986 20748 35992 20760
rect 36044 20788 36050 20800
rect 37200 20788 37228 20964
rect 37292 20910 37320 20964
rect 37366 20952 37372 20964
rect 37424 20992 37430 21004
rect 38212 21001 38240 21032
rect 38396 21004 38424 21100
rect 40494 21088 40500 21100
rect 40552 21088 40558 21140
rect 40770 21088 40776 21140
rect 40828 21128 40834 21140
rect 40957 21131 41015 21137
rect 40957 21128 40969 21131
rect 40828 21100 40969 21128
rect 40828 21088 40834 21100
rect 40957 21097 40969 21100
rect 41003 21128 41015 21131
rect 41003 21100 41414 21128
rect 41003 21097 41015 21100
rect 40957 21091 41015 21097
rect 41049 21063 41107 21069
rect 41049 21029 41061 21063
rect 41095 21029 41107 21063
rect 41049 21023 41107 21029
rect 38197 20995 38255 21001
rect 37424 20964 37964 20992
rect 37424 20952 37430 20964
rect 37936 20936 37964 20964
rect 38197 20961 38209 20995
rect 38243 20961 38255 20995
rect 38197 20955 38255 20961
rect 38378 20952 38384 21004
rect 38436 20952 38442 21004
rect 41064 20992 41092 21023
rect 38626 20964 38792 20992
rect 37734 20884 37740 20936
rect 37792 20884 37798 20936
rect 37918 20884 37924 20936
rect 37976 20884 37982 20936
rect 38102 20884 38108 20936
rect 38160 20924 38166 20936
rect 38626 20924 38654 20964
rect 38764 20933 38792 20964
rect 39040 20964 41092 20992
rect 41386 20992 41414 21100
rect 42794 21088 42800 21140
rect 42852 21128 42858 21140
rect 42889 21131 42947 21137
rect 42889 21128 42901 21131
rect 42852 21100 42901 21128
rect 42852 21088 42858 21100
rect 42889 21097 42901 21100
rect 42935 21097 42947 21131
rect 42889 21091 42947 21097
rect 44542 21088 44548 21140
rect 44600 21088 44606 21140
rect 41509 20995 41567 21001
rect 41509 20992 41521 20995
rect 41386 20964 41521 20992
rect 39040 20933 39068 20964
rect 41509 20961 41521 20964
rect 41555 20961 41567 20995
rect 41509 20955 41567 20961
rect 41598 20952 41604 21004
rect 41656 20952 41662 21004
rect 42429 20995 42487 21001
rect 42429 20961 42441 20995
rect 42475 20961 42487 20995
rect 42429 20955 42487 20961
rect 38160 20896 38654 20924
rect 38749 20927 38807 20933
rect 38160 20884 38166 20896
rect 38749 20893 38761 20927
rect 38795 20893 38807 20927
rect 38749 20887 38807 20893
rect 39025 20927 39083 20933
rect 39025 20893 39037 20927
rect 39071 20893 39083 20927
rect 39025 20887 39083 20893
rect 39206 20884 39212 20936
rect 39264 20884 39270 20936
rect 41414 20884 41420 20936
rect 41472 20924 41478 20936
rect 42245 20927 42303 20933
rect 42245 20924 42257 20927
rect 41472 20896 42257 20924
rect 41472 20884 41478 20896
rect 42245 20893 42257 20896
rect 42291 20893 42303 20927
rect 42245 20887 42303 20893
rect 36044 20760 37228 20788
rect 37752 20788 37780 20884
rect 37826 20816 37832 20868
rect 37884 20856 37890 20868
rect 38654 20856 38660 20868
rect 37884 20828 38660 20856
rect 37884 20816 37890 20828
rect 38654 20816 38660 20828
rect 38712 20816 38718 20868
rect 39485 20859 39543 20865
rect 39485 20856 39497 20859
rect 38856 20828 39497 20856
rect 38105 20791 38163 20797
rect 38105 20788 38117 20791
rect 37752 20760 38117 20788
rect 36044 20748 36050 20760
rect 38105 20757 38117 20760
rect 38151 20757 38163 20791
rect 38105 20751 38163 20757
rect 38562 20748 38568 20800
rect 38620 20748 38626 20800
rect 38856 20797 38884 20828
rect 39485 20825 39497 20828
rect 39531 20825 39543 20859
rect 39485 20819 39543 20825
rect 39758 20816 39764 20868
rect 39816 20856 39822 20868
rect 40862 20856 40868 20868
rect 39816 20828 39974 20856
rect 40788 20828 40868 20856
rect 39816 20816 39822 20828
rect 38841 20791 38899 20797
rect 38841 20757 38853 20791
rect 38887 20757 38899 20791
rect 38841 20751 38899 20757
rect 39022 20748 39028 20800
rect 39080 20788 39086 20800
rect 40788 20788 40816 20828
rect 40862 20816 40868 20828
rect 40920 20856 40926 20868
rect 42444 20856 42472 20955
rect 43162 20856 43168 20868
rect 40920 20828 43168 20856
rect 40920 20816 40926 20828
rect 43162 20816 43168 20828
rect 43220 20816 43226 20868
rect 43349 20859 43407 20865
rect 43349 20825 43361 20859
rect 43395 20856 43407 20859
rect 43395 20828 44128 20856
rect 43395 20825 43407 20828
rect 43349 20819 43407 20825
rect 39080 20760 40816 20788
rect 39080 20748 39086 20760
rect 40954 20748 40960 20800
rect 41012 20788 41018 20800
rect 41417 20791 41475 20797
rect 41417 20788 41429 20791
rect 41012 20760 41429 20788
rect 41012 20748 41018 20760
rect 41417 20757 41429 20760
rect 41463 20757 41475 20791
rect 41417 20751 41475 20757
rect 41874 20748 41880 20800
rect 41932 20748 41938 20800
rect 42334 20748 42340 20800
rect 42392 20748 42398 20800
rect 43438 20748 43444 20800
rect 43496 20788 43502 20800
rect 43625 20791 43683 20797
rect 43625 20788 43637 20791
rect 43496 20760 43637 20788
rect 43496 20748 43502 20760
rect 43625 20757 43637 20760
rect 43671 20788 43683 20791
rect 43993 20791 44051 20797
rect 43993 20788 44005 20791
rect 43671 20760 44005 20788
rect 43671 20757 43683 20760
rect 43625 20751 43683 20757
rect 43993 20757 44005 20760
rect 44039 20757 44051 20791
rect 44100 20788 44128 20828
rect 44174 20816 44180 20868
rect 44232 20856 44238 20868
rect 44821 20859 44879 20865
rect 44821 20856 44833 20859
rect 44232 20828 44833 20856
rect 44232 20816 44238 20828
rect 44821 20825 44833 20828
rect 44867 20825 44879 20859
rect 44821 20819 44879 20825
rect 45186 20816 45192 20868
rect 45244 20816 45250 20868
rect 44266 20788 44272 20800
rect 44100 20760 44272 20788
rect 43993 20751 44051 20757
rect 44266 20748 44272 20760
rect 44324 20788 44330 20800
rect 44726 20788 44732 20800
rect 44324 20760 44732 20788
rect 44324 20748 44330 20760
rect 44726 20748 44732 20760
rect 44784 20748 44790 20800
rect 460 20698 45540 20720
rect 460 20646 6070 20698
rect 6122 20646 6134 20698
rect 6186 20646 6198 20698
rect 6250 20646 6262 20698
rect 6314 20646 6326 20698
rect 6378 20646 11070 20698
rect 11122 20646 11134 20698
rect 11186 20646 11198 20698
rect 11250 20646 11262 20698
rect 11314 20646 11326 20698
rect 11378 20646 16070 20698
rect 16122 20646 16134 20698
rect 16186 20646 16198 20698
rect 16250 20646 16262 20698
rect 16314 20646 16326 20698
rect 16378 20646 21070 20698
rect 21122 20646 21134 20698
rect 21186 20646 21198 20698
rect 21250 20646 21262 20698
rect 21314 20646 21326 20698
rect 21378 20646 26070 20698
rect 26122 20646 26134 20698
rect 26186 20646 26198 20698
rect 26250 20646 26262 20698
rect 26314 20646 26326 20698
rect 26378 20646 31070 20698
rect 31122 20646 31134 20698
rect 31186 20646 31198 20698
rect 31250 20646 31262 20698
rect 31314 20646 31326 20698
rect 31378 20646 36070 20698
rect 36122 20646 36134 20698
rect 36186 20646 36198 20698
rect 36250 20646 36262 20698
rect 36314 20646 36326 20698
rect 36378 20646 41070 20698
rect 41122 20646 41134 20698
rect 41186 20646 41198 20698
rect 41250 20646 41262 20698
rect 41314 20646 41326 20698
rect 41378 20646 45540 20698
rect 460 20624 45540 20646
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20553 3663 20587
rect 3605 20547 3663 20553
rect 5537 20587 5595 20593
rect 5537 20553 5549 20587
rect 5583 20584 5595 20587
rect 6638 20584 6644 20596
rect 5583 20556 6644 20584
rect 5583 20553 5595 20556
rect 5537 20547 5595 20553
rect 750 20476 756 20528
rect 808 20516 814 20528
rect 2133 20519 2191 20525
rect 2133 20516 2145 20519
rect 808 20488 2145 20516
rect 808 20476 814 20488
rect 2133 20485 2145 20488
rect 2179 20485 2191 20519
rect 3620 20516 3648 20547
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 9217 20587 9275 20593
rect 9217 20553 9229 20587
rect 9263 20584 9275 20587
rect 9306 20584 9312 20596
rect 9263 20556 9312 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 9306 20544 9312 20556
rect 9364 20584 9370 20596
rect 9585 20587 9643 20593
rect 9585 20584 9597 20587
rect 9364 20556 9597 20584
rect 9364 20544 9370 20556
rect 9585 20553 9597 20556
rect 9631 20584 9643 20587
rect 9674 20584 9680 20596
rect 9631 20556 9680 20584
rect 9631 20553 9643 20556
rect 9585 20547 9643 20553
rect 9674 20544 9680 20556
rect 9732 20584 9738 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 9732 20556 9965 20584
rect 9732 20544 9738 20556
rect 9953 20553 9965 20556
rect 9999 20584 10011 20587
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 9999 20556 11805 20584
rect 9999 20553 10011 20556
rect 9953 20547 10011 20553
rect 11793 20553 11805 20556
rect 11839 20584 11851 20587
rect 12526 20584 12532 20596
rect 11839 20556 12532 20584
rect 11839 20553 11851 20556
rect 11793 20547 11851 20553
rect 12526 20544 12532 20556
rect 12584 20584 12590 20596
rect 13538 20584 13544 20596
rect 12584 20556 13544 20584
rect 12584 20544 12590 20556
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 13814 20584 13820 20596
rect 13648 20556 13820 20584
rect 4065 20519 4123 20525
rect 4065 20516 4077 20519
rect 3620 20488 4077 20516
rect 2133 20479 2191 20485
rect 4065 20485 4077 20488
rect 4111 20485 4123 20519
rect 4065 20479 4123 20485
rect 13265 20519 13323 20525
rect 13265 20485 13277 20519
rect 13311 20516 13323 20519
rect 13354 20516 13360 20528
rect 13311 20488 13360 20516
rect 13311 20485 13323 20488
rect 13265 20479 13323 20485
rect 13354 20476 13360 20488
rect 13412 20516 13418 20528
rect 13648 20516 13676 20556
rect 13814 20544 13820 20556
rect 13872 20584 13878 20596
rect 13909 20587 13967 20593
rect 13909 20584 13921 20587
rect 13872 20556 13921 20584
rect 13872 20544 13878 20556
rect 13909 20553 13921 20556
rect 13955 20553 13967 20587
rect 14274 20584 14280 20596
rect 13909 20547 13967 20553
rect 14108 20556 14280 20584
rect 14108 20525 14136 20556
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 15102 20544 15108 20596
rect 15160 20544 15166 20596
rect 15930 20584 15936 20596
rect 15304 20556 15936 20584
rect 13412 20488 13676 20516
rect 14093 20519 14151 20525
rect 13412 20476 13418 20488
rect 14093 20485 14105 20519
rect 14139 20485 14151 20519
rect 14093 20479 14151 20485
rect 14458 20476 14464 20528
rect 14516 20476 14522 20528
rect 14691 20485 14749 20491
rect 14691 20482 14703 20485
rect 3266 20420 3372 20448
rect 3344 20392 3372 20420
rect 5166 20408 5172 20460
rect 5224 20448 5230 20460
rect 14277 20451 14335 20457
rect 5224 20420 6040 20448
rect 5224 20408 5230 20420
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 3142 20380 3148 20392
rect 1903 20352 3148 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 3786 20340 3792 20392
rect 3844 20340 3850 20392
rect 6012 20321 6040 20420
rect 14277 20417 14289 20451
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 6822 20340 6828 20392
rect 6880 20380 6886 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 6880 20352 8033 20380
rect 6880 20340 6886 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 14292 20380 14320 20411
rect 14366 20408 14372 20460
rect 14424 20446 14430 20460
rect 14676 20451 14703 20482
rect 14737 20451 14749 20485
rect 15120 20457 15148 20544
rect 15304 20528 15332 20556
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 16132 20556 16528 20584
rect 15194 20476 15200 20528
rect 15252 20476 15258 20528
rect 15286 20476 15292 20528
rect 15344 20476 15350 20528
rect 15749 20519 15807 20525
rect 15442 20488 15700 20516
rect 15442 20457 15470 20488
rect 15672 20457 15700 20488
rect 15749 20485 15761 20519
rect 15795 20516 15807 20519
rect 16132 20516 16160 20556
rect 15795 20488 16160 20516
rect 16500 20516 16528 20556
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17129 20587 17187 20593
rect 17129 20584 17141 20587
rect 16908 20556 17141 20584
rect 16908 20544 16914 20556
rect 17129 20553 17141 20556
rect 17175 20553 17187 20587
rect 17129 20547 17187 20553
rect 17681 20587 17739 20593
rect 17681 20553 17693 20587
rect 17727 20584 17739 20587
rect 18782 20584 18788 20596
rect 17727 20556 18788 20584
rect 17727 20553 17739 20556
rect 17681 20547 17739 20553
rect 17696 20516 17724 20547
rect 18782 20544 18788 20556
rect 18840 20544 18846 20596
rect 19058 20584 19064 20596
rect 18984 20556 19064 20584
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 16500 20488 17264 20516
rect 15795 20485 15807 20488
rect 15749 20479 15807 20485
rect 14676 20448 14749 20451
rect 14660 20446 14749 20448
rect 14424 20445 14749 20446
rect 15105 20451 15163 20457
rect 14424 20420 14704 20445
rect 14424 20418 14688 20420
rect 14424 20408 14430 20418
rect 15105 20417 15117 20451
rect 15151 20417 15163 20451
rect 15105 20411 15163 20417
rect 15427 20451 15485 20457
rect 15427 20417 15439 20451
rect 15473 20417 15485 20451
rect 15427 20411 15485 20417
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15657 20411 15715 20417
rect 15764 20420 15853 20448
rect 14734 20380 14740 20392
rect 14292 20352 14740 20380
rect 8021 20343 8079 20349
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 15442 20380 15470 20411
rect 15764 20392 15792 20420
rect 15841 20417 15853 20420
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 15988 20420 16068 20448
rect 15988 20408 15994 20420
rect 15565 20383 15623 20389
rect 15442 20352 15516 20380
rect 15488 20324 15516 20352
rect 15565 20349 15577 20383
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 5997 20315 6055 20321
rect 5997 20281 6009 20315
rect 6043 20312 6055 20315
rect 14093 20315 14151 20321
rect 6043 20284 7972 20312
rect 6043 20281 6055 20284
rect 5997 20275 6055 20281
rect 7944 20256 7972 20284
rect 14093 20281 14105 20315
rect 14139 20281 14151 20315
rect 14093 20275 14151 20281
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 6273 20247 6331 20253
rect 6273 20244 6285 20247
rect 5684 20216 6285 20244
rect 5684 20204 5690 20216
rect 6273 20213 6285 20216
rect 6319 20244 6331 20247
rect 6822 20244 6828 20256
rect 6319 20216 6828 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 6822 20204 6828 20216
rect 6880 20244 6886 20256
rect 6917 20247 6975 20253
rect 6917 20244 6929 20247
rect 6880 20216 6929 20244
rect 6880 20204 6886 20216
rect 6917 20213 6929 20216
rect 6963 20213 6975 20247
rect 6917 20207 6975 20213
rect 7282 20204 7288 20256
rect 7340 20244 7346 20256
rect 7653 20247 7711 20253
rect 7653 20244 7665 20247
rect 7340 20216 7665 20244
rect 7340 20204 7346 20216
rect 7653 20213 7665 20216
rect 7699 20213 7711 20247
rect 7653 20207 7711 20213
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8386 20244 8392 20256
rect 7984 20216 8392 20244
rect 7984 20204 7990 20216
rect 8386 20204 8392 20216
rect 8444 20244 8450 20256
rect 8757 20247 8815 20253
rect 8757 20244 8769 20247
rect 8444 20216 8769 20244
rect 8444 20204 8450 20216
rect 8757 20213 8769 20216
rect 8803 20244 8815 20247
rect 10226 20244 10232 20256
rect 8803 20216 10232 20244
rect 8803 20213 8815 20216
rect 8757 20207 8815 20213
rect 10226 20204 10232 20216
rect 10284 20244 10290 20256
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 10284 20216 10609 20244
rect 10284 20204 10290 20216
rect 10597 20213 10609 20216
rect 10643 20244 10655 20247
rect 10962 20244 10968 20256
rect 10643 20216 10968 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10962 20204 10968 20216
rect 11020 20244 11026 20256
rect 11333 20247 11391 20253
rect 11333 20244 11345 20247
rect 11020 20216 11345 20244
rect 11020 20204 11026 20216
rect 11333 20213 11345 20216
rect 11379 20244 11391 20247
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11379 20216 12173 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 12161 20213 12173 20216
rect 12207 20244 12219 20247
rect 12897 20247 12955 20253
rect 12897 20244 12909 20247
rect 12207 20216 12909 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12897 20213 12909 20216
rect 12943 20244 12955 20247
rect 13906 20244 13912 20256
rect 12943 20216 13912 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14108 20244 14136 20275
rect 14366 20272 14372 20324
rect 14424 20312 14430 20324
rect 14921 20315 14979 20321
rect 14921 20312 14933 20315
rect 14424 20284 14933 20312
rect 14424 20272 14430 20284
rect 14921 20281 14933 20284
rect 14967 20281 14979 20315
rect 14921 20275 14979 20281
rect 15470 20272 15476 20324
rect 15528 20272 15534 20324
rect 15580 20312 15608 20343
rect 15746 20340 15752 20392
rect 15804 20340 15810 20392
rect 16040 20380 16068 20420
rect 16114 20408 16120 20460
rect 16172 20446 16178 20460
rect 16209 20451 16267 20457
rect 16209 20446 16221 20451
rect 16172 20418 16221 20446
rect 16172 20408 16178 20418
rect 16209 20417 16221 20418
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 16298 20408 16304 20460
rect 16356 20408 16362 20460
rect 16393 20451 16451 20457
rect 16393 20417 16405 20451
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 16408 20380 16436 20411
rect 16482 20408 16488 20460
rect 16540 20457 16546 20460
rect 16540 20451 16569 20457
rect 16557 20417 16569 20451
rect 16540 20411 16569 20417
rect 16540 20408 16546 20411
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 16761 20451 16819 20457
rect 16761 20417 16773 20451
rect 16807 20448 16819 20451
rect 16942 20448 16948 20460
rect 16807 20420 16948 20448
rect 16807 20417 16819 20420
rect 16761 20411 16819 20417
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17236 20457 17264 20488
rect 17604 20488 17724 20516
rect 17788 20488 18889 20516
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17402 20448 17408 20460
rect 17359 20420 17408 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17604 20457 17632 20488
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20417 17647 20451
rect 17788 20448 17816 20488
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 18877 20479 18935 20485
rect 18984 20460 19012 20556
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19208 20556 19533 20584
rect 19208 20544 19214 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 19521 20547 19579 20553
rect 19886 20544 19892 20596
rect 19944 20584 19950 20596
rect 20257 20587 20315 20593
rect 20257 20584 20269 20587
rect 19944 20556 20269 20584
rect 19944 20544 19950 20556
rect 20257 20553 20269 20556
rect 20303 20553 20315 20587
rect 20257 20547 20315 20553
rect 20441 20587 20499 20593
rect 20441 20553 20453 20587
rect 20487 20584 20499 20587
rect 20622 20584 20628 20596
rect 20487 20556 20628 20584
rect 20487 20553 20499 20556
rect 20441 20547 20499 20553
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 22741 20587 22799 20593
rect 21192 20556 22508 20584
rect 19702 20516 19708 20528
rect 19081 20488 19708 20516
rect 17589 20411 17647 20417
rect 17696 20420 17816 20448
rect 17865 20451 17923 20457
rect 17512 20380 17540 20411
rect 17696 20392 17724 20420
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 16040 20352 16436 20380
rect 17236 20352 17540 20380
rect 15654 20312 15660 20324
rect 15580 20284 15660 20312
rect 15654 20272 15660 20284
rect 15712 20272 15718 20324
rect 16666 20272 16672 20324
rect 16724 20312 16730 20324
rect 16899 20315 16957 20321
rect 16899 20312 16911 20315
rect 16724 20284 16911 20312
rect 16724 20272 16730 20284
rect 16899 20281 16911 20284
rect 16945 20281 16957 20315
rect 16899 20275 16957 20281
rect 14182 20244 14188 20256
rect 14108 20216 14188 20244
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 14734 20244 14740 20256
rect 14691 20216 14740 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 14829 20247 14887 20253
rect 14829 20213 14841 20247
rect 14875 20244 14887 20247
rect 16298 20244 16304 20256
rect 14875 20216 16304 20244
rect 14875 20213 14887 20216
rect 14829 20207 14887 20213
rect 16298 20204 16304 20216
rect 16356 20244 16362 20256
rect 17037 20247 17095 20253
rect 17037 20244 17049 20247
rect 16356 20216 17049 20244
rect 16356 20204 16362 20216
rect 17037 20213 17049 20216
rect 17083 20213 17095 20247
rect 17236 20244 17264 20352
rect 17678 20340 17684 20392
rect 17736 20340 17742 20392
rect 17770 20340 17776 20392
rect 17828 20340 17834 20392
rect 17313 20315 17371 20321
rect 17313 20281 17325 20315
rect 17359 20312 17371 20315
rect 17788 20312 17816 20340
rect 17359 20284 17816 20312
rect 17880 20312 17908 20411
rect 18064 20380 18092 20411
rect 18138 20408 18144 20460
rect 18196 20408 18202 20460
rect 18230 20408 18236 20460
rect 18288 20408 18294 20460
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 18417 20451 18475 20457
rect 18417 20448 18429 20451
rect 18380 20420 18429 20448
rect 18380 20408 18386 20420
rect 18417 20417 18429 20420
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 18635 20451 18693 20457
rect 18635 20417 18647 20451
rect 18681 20448 18693 20451
rect 18966 20448 18972 20460
rect 18681 20420 18972 20448
rect 18681 20417 18693 20420
rect 18635 20411 18693 20417
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19081 20380 19109 20488
rect 19702 20476 19708 20488
rect 19760 20476 19766 20528
rect 21192 20525 21220 20556
rect 21177 20519 21235 20525
rect 21177 20516 21189 20519
rect 20260 20488 21189 20516
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20417 19211 20451
rect 19613 20451 19671 20457
rect 19613 20448 19625 20451
rect 19153 20411 19211 20417
rect 19536 20420 19625 20448
rect 18064 20352 19109 20380
rect 19168 20324 19196 20411
rect 19536 20392 19564 20420
rect 19613 20417 19625 20420
rect 19659 20417 19671 20451
rect 19613 20411 19671 20417
rect 20162 20408 20168 20460
rect 20220 20457 20226 20460
rect 20220 20448 20229 20457
rect 20260 20448 20288 20488
rect 21177 20485 21189 20488
rect 21223 20485 21235 20519
rect 21177 20479 21235 20485
rect 21450 20476 21456 20528
rect 21508 20516 21514 20528
rect 21545 20519 21603 20525
rect 21545 20516 21557 20519
rect 21508 20488 21557 20516
rect 21508 20476 21514 20488
rect 21545 20485 21557 20488
rect 21591 20485 21603 20519
rect 22373 20519 22431 20525
rect 22373 20516 22385 20519
rect 21545 20479 21603 20485
rect 22112 20488 22385 20516
rect 20220 20420 20288 20448
rect 20349 20451 20407 20457
rect 20220 20411 20229 20420
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 20438 20448 20444 20460
rect 20395 20420 20444 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 20220 20408 20226 20411
rect 20438 20408 20444 20420
rect 20496 20448 20502 20460
rect 21361 20451 21419 20457
rect 21361 20448 21373 20451
rect 20496 20420 21373 20448
rect 20496 20408 20502 20420
rect 21361 20417 21373 20420
rect 21407 20417 21419 20451
rect 21361 20411 21419 20417
rect 21726 20408 21732 20460
rect 21784 20448 21790 20460
rect 21913 20451 21971 20457
rect 21913 20448 21925 20451
rect 21784 20420 21925 20448
rect 21784 20408 21790 20420
rect 21913 20417 21925 20420
rect 21959 20417 21971 20451
rect 21913 20411 21971 20417
rect 22002 20408 22008 20460
rect 22060 20408 22066 20460
rect 22112 20457 22140 20488
rect 22373 20485 22385 20488
rect 22419 20485 22431 20519
rect 22480 20516 22508 20556
rect 22741 20553 22753 20587
rect 22787 20584 22799 20587
rect 23106 20584 23112 20596
rect 22787 20556 23112 20584
rect 22787 20553 22799 20556
rect 22741 20547 22799 20553
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 23477 20587 23535 20593
rect 23477 20584 23489 20587
rect 23440 20556 23489 20584
rect 23440 20544 23446 20556
rect 23477 20553 23489 20556
rect 23523 20553 23535 20587
rect 23477 20547 23535 20553
rect 23934 20544 23940 20596
rect 23992 20544 23998 20596
rect 24762 20544 24768 20596
rect 24820 20544 24826 20596
rect 25590 20544 25596 20596
rect 25648 20544 25654 20596
rect 25682 20544 25688 20596
rect 25740 20544 25746 20596
rect 27338 20584 27344 20596
rect 26068 20556 27344 20584
rect 23014 20516 23020 20528
rect 22480 20488 23020 20516
rect 22373 20479 22431 20485
rect 23014 20476 23020 20488
rect 23072 20476 23078 20528
rect 24780 20516 24808 20544
rect 24688 20488 24808 20516
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20417 22155 20451
rect 22097 20411 22155 20417
rect 19245 20383 19303 20389
rect 19245 20349 19257 20383
rect 19291 20380 19303 20383
rect 19334 20380 19340 20392
rect 19291 20352 19340 20380
rect 19291 20349 19303 20352
rect 19245 20343 19303 20349
rect 19334 20340 19340 20352
rect 19392 20340 19398 20392
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 19150 20312 19156 20324
rect 17880 20284 19156 20312
rect 17359 20281 17371 20284
rect 17313 20275 17371 20281
rect 19150 20272 19156 20284
rect 19208 20312 19214 20324
rect 19720 20312 19748 20343
rect 19978 20340 19984 20392
rect 20036 20340 20042 20392
rect 20530 20340 20536 20392
rect 20588 20380 20594 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 20588 20352 20637 20380
rect 20588 20340 20594 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 20806 20340 20812 20392
rect 20864 20340 20870 20392
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20349 20959 20383
rect 22020 20380 22048 20408
rect 20901 20343 20959 20349
rect 21928 20352 22048 20380
rect 22112 20380 22140 20411
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 22244 20420 22293 20448
rect 22244 20408 22250 20420
rect 22281 20417 22293 20420
rect 22327 20448 22339 20451
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 22327 20420 22569 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 22557 20417 22569 20420
rect 22603 20417 22615 20451
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 22557 20411 22615 20417
rect 22756 20420 23857 20448
rect 22112 20352 22232 20380
rect 19996 20312 20024 20340
rect 19208 20284 19748 20312
rect 19812 20284 20024 20312
rect 19208 20272 19214 20284
rect 18138 20244 18144 20256
rect 17236 20216 18144 20244
rect 17037 20207 17095 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 19058 20244 19064 20256
rect 18656 20216 19064 20244
rect 18656 20204 18662 20216
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19812 20253 19840 20284
rect 20070 20272 20076 20324
rect 20128 20312 20134 20324
rect 20916 20312 20944 20343
rect 21928 20324 21956 20352
rect 22204 20324 22232 20352
rect 20128 20284 20944 20312
rect 20128 20272 20134 20284
rect 21266 20272 21272 20324
rect 21324 20312 21330 20324
rect 21324 20284 21772 20312
rect 21324 20272 21330 20284
rect 19797 20247 19855 20253
rect 19797 20213 19809 20247
rect 19843 20213 19855 20247
rect 19797 20207 19855 20213
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20898 20244 20904 20256
rect 20680 20216 20904 20244
rect 20680 20204 20686 20216
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 21634 20204 21640 20256
rect 21692 20204 21698 20256
rect 21744 20244 21772 20284
rect 21910 20272 21916 20324
rect 21968 20272 21974 20324
rect 22186 20272 22192 20324
rect 22244 20272 22250 20324
rect 22756 20244 22784 20420
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 24578 20448 24584 20460
rect 23845 20411 23903 20417
rect 24044 20420 24584 20448
rect 22830 20340 22836 20392
rect 22888 20380 22894 20392
rect 24044 20380 24072 20420
rect 24578 20408 24584 20420
rect 24636 20408 24642 20460
rect 22888 20352 24072 20380
rect 24121 20383 24179 20389
rect 22888 20340 22894 20352
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24688 20380 24716 20488
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 25133 20451 25191 20457
rect 25133 20417 25145 20451
rect 25179 20417 25191 20451
rect 25700 20448 25728 20544
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 25700 20420 25789 20448
rect 25133 20411 25191 20417
rect 25777 20417 25789 20420
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 24167 20352 24716 20380
rect 24780 20380 24808 20411
rect 25148 20380 25176 20411
rect 26068 20380 26096 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 27614 20544 27620 20596
rect 27672 20584 27678 20596
rect 28258 20584 28264 20596
rect 27672 20556 28264 20584
rect 27672 20544 27678 20556
rect 27908 20528 27936 20556
rect 28258 20544 28264 20556
rect 28316 20544 28322 20596
rect 28350 20544 28356 20596
rect 28408 20584 28414 20596
rect 29086 20584 29092 20596
rect 28408 20556 29092 20584
rect 28408 20544 28414 20556
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 29362 20544 29368 20596
rect 29420 20584 29426 20596
rect 29917 20587 29975 20593
rect 29917 20584 29929 20587
rect 29420 20556 29929 20584
rect 29420 20544 29426 20556
rect 29917 20553 29929 20556
rect 29963 20553 29975 20587
rect 29917 20547 29975 20553
rect 30208 20556 31984 20584
rect 27890 20516 27896 20528
rect 27830 20488 27896 20516
rect 27890 20476 27896 20488
rect 27948 20476 27954 20528
rect 28166 20516 28172 20528
rect 28000 20488 28172 20516
rect 26142 20408 26148 20460
rect 26200 20408 26206 20460
rect 28000 20392 28028 20488
rect 28166 20476 28172 20488
rect 28224 20476 28230 20528
rect 28445 20519 28503 20525
rect 28445 20485 28457 20519
rect 28491 20516 28503 20519
rect 28718 20516 28724 20528
rect 28491 20488 28724 20516
rect 28491 20485 28503 20488
rect 28445 20479 28503 20485
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 30208 20457 30236 20556
rect 30374 20476 30380 20528
rect 30432 20476 30438 20528
rect 30558 20476 30564 20528
rect 30616 20516 30622 20528
rect 31757 20519 31815 20525
rect 31757 20516 31769 20519
rect 30616 20488 31769 20516
rect 30616 20476 30622 20488
rect 31757 20485 31769 20488
rect 31803 20485 31815 20519
rect 31956 20516 31984 20556
rect 32030 20544 32036 20596
rect 32088 20544 32094 20596
rect 33226 20584 33232 20596
rect 32140 20556 33232 20584
rect 32140 20516 32168 20556
rect 33226 20544 33232 20556
rect 33284 20544 33290 20596
rect 33410 20544 33416 20596
rect 33468 20544 33474 20596
rect 33689 20587 33747 20593
rect 33689 20553 33701 20587
rect 33735 20553 33747 20587
rect 33689 20547 33747 20553
rect 31956 20488 32168 20516
rect 31757 20479 31815 20485
rect 32950 20476 32956 20528
rect 33008 20476 33014 20528
rect 30193 20451 30251 20457
rect 24780 20352 25084 20380
rect 25148 20352 26096 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 24210 20272 24216 20324
rect 24268 20312 24274 20324
rect 25056 20312 25084 20352
rect 26234 20340 26240 20392
rect 26292 20380 26298 20392
rect 26329 20383 26387 20389
rect 26329 20380 26341 20383
rect 26292 20352 26341 20380
rect 26292 20340 26298 20352
rect 26329 20349 26341 20352
rect 26375 20349 26387 20383
rect 26329 20343 26387 20349
rect 26605 20383 26663 20389
rect 26605 20349 26617 20383
rect 26651 20380 26663 20383
rect 27614 20380 27620 20392
rect 26651 20352 27620 20380
rect 26651 20349 26663 20352
rect 26605 20343 26663 20349
rect 27614 20340 27620 20352
rect 27672 20340 27678 20392
rect 27982 20340 27988 20392
rect 28040 20340 28046 20392
rect 28166 20340 28172 20392
rect 28224 20340 28230 20392
rect 28994 20380 29000 20392
rect 28276 20352 29000 20380
rect 25866 20312 25872 20324
rect 24268 20284 24992 20312
rect 25056 20284 25872 20312
rect 24268 20272 24274 20284
rect 21744 20216 22784 20244
rect 23385 20247 23443 20253
rect 23385 20213 23397 20247
rect 23431 20244 23443 20247
rect 24394 20244 24400 20256
rect 23431 20216 24400 20244
rect 23431 20213 23443 20216
rect 23385 20207 23443 20213
rect 24394 20204 24400 20216
rect 24452 20244 24458 20256
rect 24964 20253 24992 20284
rect 25866 20272 25872 20284
rect 25924 20272 25930 20324
rect 25961 20315 26019 20321
rect 25961 20281 25973 20315
rect 26007 20281 26019 20315
rect 28276 20312 28304 20352
rect 28994 20340 29000 20352
rect 29052 20340 29058 20392
rect 29178 20340 29184 20392
rect 29236 20380 29242 20392
rect 29564 20380 29592 20434
rect 30193 20417 30205 20451
rect 30239 20417 30251 20451
rect 30392 20448 30420 20476
rect 30653 20451 30711 20457
rect 30653 20448 30665 20451
rect 30392 20420 30665 20448
rect 30193 20411 30251 20417
rect 30653 20417 30665 20420
rect 30699 20417 30711 20451
rect 30653 20411 30711 20417
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20448 30803 20451
rect 30791 20420 30880 20448
rect 30791 20417 30803 20420
rect 30745 20411 30803 20417
rect 30282 20380 30288 20392
rect 29236 20352 30288 20380
rect 29236 20340 29242 20352
rect 25961 20275 26019 20281
rect 28000 20284 28304 20312
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 24452 20216 24593 20244
rect 24452 20204 24458 20216
rect 24581 20213 24593 20216
rect 24627 20213 24639 20247
rect 24581 20207 24639 20213
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25038 20244 25044 20256
rect 24995 20216 25044 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 25314 20204 25320 20256
rect 25372 20204 25378 20256
rect 25976 20244 26004 20275
rect 28000 20244 28028 20284
rect 25976 20216 28028 20244
rect 28074 20204 28080 20256
rect 28132 20204 28138 20256
rect 28258 20204 28264 20256
rect 28316 20244 28322 20256
rect 29472 20244 29500 20352
rect 30282 20340 30288 20352
rect 30340 20340 30346 20392
rect 30009 20315 30067 20321
rect 30009 20281 30021 20315
rect 30055 20312 30067 20315
rect 30466 20312 30472 20324
rect 30055 20284 30472 20312
rect 30055 20281 30067 20284
rect 30009 20275 30067 20281
rect 30466 20272 30472 20284
rect 30524 20272 30530 20324
rect 30558 20272 30564 20324
rect 30616 20312 30622 20324
rect 30852 20312 30880 20420
rect 31110 20408 31116 20460
rect 31168 20448 31174 20460
rect 31481 20451 31539 20457
rect 31481 20448 31493 20451
rect 31168 20420 31493 20448
rect 31168 20408 31174 20420
rect 31481 20417 31493 20420
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 31662 20408 31668 20460
rect 31720 20408 31726 20460
rect 31846 20408 31852 20460
rect 31904 20408 31910 20460
rect 32125 20451 32183 20457
rect 32125 20417 32137 20451
rect 32171 20448 32183 20451
rect 33045 20451 33103 20457
rect 32171 20420 32628 20448
rect 32171 20417 32183 20420
rect 32125 20411 32183 20417
rect 30929 20383 30987 20389
rect 30929 20349 30941 20383
rect 30975 20380 30987 20383
rect 31018 20380 31024 20392
rect 30975 20352 31024 20380
rect 30975 20349 30987 20352
rect 30929 20343 30987 20349
rect 31018 20340 31024 20352
rect 31076 20340 31082 20392
rect 30616 20284 30880 20312
rect 31036 20312 31064 20340
rect 31386 20312 31392 20324
rect 31036 20284 31392 20312
rect 30616 20272 30622 20284
rect 31386 20272 31392 20284
rect 31444 20272 31450 20324
rect 32306 20272 32312 20324
rect 32364 20272 32370 20324
rect 32600 20321 32628 20420
rect 33045 20417 33057 20451
rect 33091 20448 33103 20451
rect 33410 20448 33416 20460
rect 33091 20420 33416 20448
rect 33091 20417 33103 20420
rect 33045 20411 33103 20417
rect 33410 20408 33416 20420
rect 33468 20408 33474 20460
rect 33597 20451 33655 20457
rect 33597 20417 33609 20451
rect 33643 20448 33655 20451
rect 33704 20448 33732 20547
rect 34054 20544 34060 20596
rect 34112 20544 34118 20596
rect 34149 20587 34207 20593
rect 34149 20553 34161 20587
rect 34195 20584 34207 20587
rect 34514 20584 34520 20596
rect 34195 20556 34520 20584
rect 34195 20553 34207 20556
rect 34149 20547 34207 20553
rect 34514 20544 34520 20556
rect 34572 20544 34578 20596
rect 34885 20587 34943 20593
rect 34885 20553 34897 20587
rect 34931 20584 34943 20587
rect 35158 20584 35164 20596
rect 34931 20556 35164 20584
rect 34931 20553 34943 20556
rect 34885 20547 34943 20553
rect 35158 20544 35164 20556
rect 35216 20544 35222 20596
rect 35713 20587 35771 20593
rect 35713 20553 35725 20587
rect 35759 20584 35771 20587
rect 35894 20584 35900 20596
rect 35759 20556 35900 20584
rect 35759 20553 35771 20556
rect 35713 20547 35771 20553
rect 35894 20544 35900 20556
rect 35952 20544 35958 20596
rect 36446 20544 36452 20596
rect 36504 20584 36510 20596
rect 36633 20587 36691 20593
rect 36633 20584 36645 20587
rect 36504 20556 36645 20584
rect 36504 20544 36510 20556
rect 36633 20553 36645 20556
rect 36679 20553 36691 20587
rect 36633 20547 36691 20553
rect 37093 20587 37151 20593
rect 37093 20553 37105 20587
rect 37139 20584 37151 20587
rect 37274 20584 37280 20596
rect 37139 20556 37280 20584
rect 37139 20553 37151 20556
rect 37093 20547 37151 20553
rect 37274 20544 37280 20556
rect 37332 20584 37338 20596
rect 37734 20584 37740 20596
rect 37332 20556 37740 20584
rect 37332 20544 37338 20556
rect 37734 20544 37740 20556
rect 37792 20544 37798 20596
rect 38562 20584 38568 20596
rect 37844 20556 38568 20584
rect 33962 20476 33968 20528
rect 34020 20516 34026 20528
rect 34020 20488 34744 20516
rect 34020 20476 34026 20488
rect 33643 20420 33732 20448
rect 34716 20448 34744 20488
rect 34974 20476 34980 20528
rect 35032 20476 35038 20528
rect 36081 20519 36139 20525
rect 36081 20485 36093 20519
rect 36127 20516 36139 20519
rect 36814 20516 36820 20528
rect 36127 20488 36820 20516
rect 36127 20485 36139 20488
rect 36081 20479 36139 20485
rect 36814 20476 36820 20488
rect 36872 20516 36878 20528
rect 37844 20525 37872 20556
rect 38562 20544 38568 20556
rect 38620 20544 38626 20596
rect 39301 20587 39359 20593
rect 39301 20553 39313 20587
rect 39347 20584 39359 20587
rect 39666 20584 39672 20596
rect 39347 20556 39672 20584
rect 39347 20553 39359 20556
rect 39301 20547 39359 20553
rect 39666 20544 39672 20556
rect 39724 20544 39730 20596
rect 39758 20544 39764 20596
rect 39816 20584 39822 20596
rect 40770 20584 40776 20596
rect 39816 20556 40776 20584
rect 39816 20544 39822 20556
rect 37001 20519 37059 20525
rect 37001 20516 37013 20519
rect 36872 20488 37013 20516
rect 36872 20476 36878 20488
rect 37001 20485 37013 20488
rect 37047 20485 37059 20519
rect 37001 20479 37059 20485
rect 37829 20519 37887 20525
rect 37829 20485 37841 20519
rect 37875 20485 37887 20519
rect 37829 20479 37887 20485
rect 37918 20476 37924 20528
rect 37976 20516 37982 20528
rect 38102 20516 38108 20528
rect 37976 20488 38108 20516
rect 37976 20476 37982 20488
rect 38102 20476 38108 20488
rect 38160 20516 38166 20528
rect 39945 20519 40003 20525
rect 38160 20488 38318 20516
rect 38160 20476 38166 20488
rect 39945 20485 39957 20519
rect 39991 20516 40003 20519
rect 40034 20516 40040 20528
rect 39991 20488 40040 20516
rect 39991 20485 40003 20488
rect 39945 20479 40003 20485
rect 40034 20476 40040 20488
rect 40092 20476 40098 20528
rect 40144 20516 40172 20556
rect 40770 20544 40776 20556
rect 40828 20544 40834 20596
rect 41417 20587 41475 20593
rect 41417 20553 41429 20587
rect 41463 20584 41475 20587
rect 42245 20587 42303 20593
rect 42245 20584 42257 20587
rect 41463 20556 42257 20584
rect 41463 20553 41475 20556
rect 41417 20547 41475 20553
rect 42245 20553 42257 20556
rect 42291 20584 42303 20587
rect 42334 20584 42340 20596
rect 42291 20556 42340 20584
rect 42291 20553 42303 20556
rect 42245 20547 42303 20553
rect 42334 20544 42340 20556
rect 42392 20544 42398 20596
rect 40144 20488 40434 20516
rect 42058 20476 42064 20528
rect 42116 20516 42122 20528
rect 43073 20519 43131 20525
rect 43073 20516 43085 20519
rect 42116 20488 43085 20516
rect 42116 20476 42122 20488
rect 43073 20485 43085 20488
rect 43119 20516 43131 20519
rect 43438 20516 43444 20528
rect 43119 20488 43444 20516
rect 43119 20485 43131 20488
rect 43073 20479 43131 20485
rect 43438 20476 43444 20488
rect 43496 20516 43502 20528
rect 44545 20519 44603 20525
rect 44545 20516 44557 20519
rect 43496 20488 44557 20516
rect 43496 20476 43502 20488
rect 44545 20485 44557 20488
rect 44591 20516 44603 20519
rect 44913 20519 44971 20525
rect 44913 20516 44925 20519
rect 44591 20488 44925 20516
rect 44591 20485 44603 20488
rect 44545 20479 44603 20485
rect 44913 20485 44925 20488
rect 44959 20485 44971 20519
rect 44913 20479 44971 20485
rect 36173 20451 36231 20457
rect 34716 20420 35756 20448
rect 33643 20417 33655 20420
rect 33597 20411 33655 20417
rect 35728 20392 35756 20420
rect 36173 20417 36185 20451
rect 36219 20448 36231 20451
rect 36906 20448 36912 20460
rect 36219 20420 36912 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 36906 20408 36912 20420
rect 36964 20408 36970 20460
rect 41414 20408 41420 20460
rect 41472 20448 41478 20460
rect 42153 20451 42211 20457
rect 42153 20448 42165 20451
rect 41472 20420 42165 20448
rect 41472 20408 41478 20420
rect 42153 20417 42165 20420
rect 42199 20417 42211 20451
rect 42797 20451 42855 20457
rect 42797 20448 42809 20451
rect 42153 20411 42211 20417
rect 42260 20420 42809 20448
rect 33134 20340 33140 20392
rect 33192 20340 33198 20392
rect 33318 20340 33324 20392
rect 33376 20380 33382 20392
rect 34238 20380 34244 20392
rect 33376 20352 34244 20380
rect 33376 20340 33382 20352
rect 34238 20340 34244 20352
rect 34296 20340 34302 20392
rect 34606 20340 34612 20392
rect 34664 20380 34670 20392
rect 35066 20380 35072 20392
rect 34664 20352 35072 20380
rect 34664 20340 34670 20352
rect 35066 20340 35072 20352
rect 35124 20340 35130 20392
rect 35710 20340 35716 20392
rect 35768 20380 35774 20392
rect 36357 20383 36415 20389
rect 36357 20380 36369 20383
rect 35768 20352 36369 20380
rect 35768 20340 35774 20352
rect 36357 20349 36369 20352
rect 36403 20349 36415 20383
rect 36357 20343 36415 20349
rect 32585 20315 32643 20321
rect 32585 20281 32597 20315
rect 32631 20281 32643 20315
rect 32585 20275 32643 20281
rect 34517 20315 34575 20321
rect 34517 20281 34529 20315
rect 34563 20312 34575 20315
rect 34698 20312 34704 20324
rect 34563 20284 34704 20312
rect 34563 20281 34575 20284
rect 34517 20275 34575 20281
rect 34698 20272 34704 20284
rect 34756 20272 34762 20324
rect 36372 20312 36400 20343
rect 37182 20340 37188 20392
rect 37240 20340 37246 20392
rect 37366 20340 37372 20392
rect 37424 20380 37430 20392
rect 37553 20383 37611 20389
rect 37553 20380 37565 20383
rect 37424 20352 37565 20380
rect 37424 20340 37430 20352
rect 37553 20349 37565 20352
rect 37599 20349 37611 20383
rect 38378 20380 38384 20392
rect 37553 20343 37611 20349
rect 37660 20352 38384 20380
rect 37660 20312 37688 20352
rect 38378 20340 38384 20352
rect 38436 20340 38442 20392
rect 39206 20340 39212 20392
rect 39264 20380 39270 20392
rect 39669 20383 39727 20389
rect 39669 20380 39681 20383
rect 39264 20352 39681 20380
rect 39264 20340 39270 20352
rect 39669 20349 39681 20352
rect 39715 20349 39727 20383
rect 39669 20343 39727 20349
rect 41782 20340 41788 20392
rect 41840 20380 41846 20392
rect 42260 20380 42288 20420
rect 42797 20417 42809 20420
rect 42843 20417 42855 20451
rect 42797 20411 42855 20417
rect 41840 20352 42288 20380
rect 41840 20340 41846 20352
rect 42334 20340 42340 20392
rect 42392 20340 42398 20392
rect 39390 20312 39396 20324
rect 36372 20284 37688 20312
rect 38856 20284 39396 20312
rect 28316 20216 29500 20244
rect 30285 20247 30343 20253
rect 28316 20204 28322 20216
rect 30285 20213 30297 20247
rect 30331 20244 30343 20247
rect 30834 20244 30840 20256
rect 30331 20216 30840 20244
rect 30331 20213 30343 20216
rect 30285 20207 30343 20213
rect 30834 20204 30840 20216
rect 30892 20204 30898 20256
rect 35618 20204 35624 20256
rect 35676 20244 35682 20256
rect 38856 20244 38884 20284
rect 39390 20272 39396 20284
rect 39448 20272 39454 20324
rect 41616 20284 43760 20312
rect 35676 20216 38884 20244
rect 35676 20204 35682 20216
rect 38930 20204 38936 20256
rect 38988 20244 38994 20256
rect 41616 20244 41644 20284
rect 38988 20216 41644 20244
rect 38988 20204 38994 20216
rect 41690 20204 41696 20256
rect 41748 20244 41754 20256
rect 41785 20247 41843 20253
rect 41785 20244 41797 20247
rect 41748 20216 41797 20244
rect 41748 20204 41754 20216
rect 41785 20213 41797 20216
rect 41831 20213 41843 20247
rect 41785 20207 41843 20213
rect 42610 20204 42616 20256
rect 42668 20204 42674 20256
rect 43732 20244 43760 20284
rect 43806 20272 43812 20324
rect 43864 20272 43870 20324
rect 44174 20244 44180 20256
rect 43732 20216 44180 20244
rect 44174 20204 44180 20216
rect 44232 20204 44238 20256
rect 44266 20204 44272 20256
rect 44324 20204 44330 20256
rect 460 20154 45540 20176
rect 460 20102 3570 20154
rect 3622 20102 3634 20154
rect 3686 20102 3698 20154
rect 3750 20102 3762 20154
rect 3814 20102 3826 20154
rect 3878 20102 8570 20154
rect 8622 20102 8634 20154
rect 8686 20102 8698 20154
rect 8750 20102 8762 20154
rect 8814 20102 8826 20154
rect 8878 20102 13570 20154
rect 13622 20102 13634 20154
rect 13686 20102 13698 20154
rect 13750 20102 13762 20154
rect 13814 20102 13826 20154
rect 13878 20102 18570 20154
rect 18622 20102 18634 20154
rect 18686 20102 18698 20154
rect 18750 20102 18762 20154
rect 18814 20102 18826 20154
rect 18878 20102 23570 20154
rect 23622 20102 23634 20154
rect 23686 20102 23698 20154
rect 23750 20102 23762 20154
rect 23814 20102 23826 20154
rect 23878 20102 28570 20154
rect 28622 20102 28634 20154
rect 28686 20102 28698 20154
rect 28750 20102 28762 20154
rect 28814 20102 28826 20154
rect 28878 20102 33570 20154
rect 33622 20102 33634 20154
rect 33686 20102 33698 20154
rect 33750 20102 33762 20154
rect 33814 20102 33826 20154
rect 33878 20102 38570 20154
rect 38622 20102 38634 20154
rect 38686 20102 38698 20154
rect 38750 20102 38762 20154
rect 38814 20102 38826 20154
rect 38878 20102 43570 20154
rect 43622 20102 43634 20154
rect 43686 20102 43698 20154
rect 43750 20102 43762 20154
rect 43814 20102 43826 20154
rect 43878 20102 45540 20154
rect 460 20080 45540 20102
rect 3326 20000 3332 20052
rect 3384 20040 3390 20052
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3384 20012 3985 20040
rect 3384 20000 3390 20012
rect 3973 20009 3985 20012
rect 4019 20040 4031 20043
rect 5166 20040 5172 20052
rect 4019 20012 5172 20040
rect 4019 20009 4031 20012
rect 3973 20003 4031 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6880 20012 6929 20040
rect 6880 20000 6886 20012
rect 6917 20009 6929 20012
rect 6963 20040 6975 20043
rect 7653 20043 7711 20049
rect 7653 20040 7665 20043
rect 6963 20012 7665 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7653 20009 7665 20012
rect 7699 20040 7711 20043
rect 8570 20040 8576 20052
rect 7699 20012 8576 20040
rect 7699 20009 7711 20012
rect 7653 20003 7711 20009
rect 8570 20000 8576 20012
rect 8628 20040 8634 20052
rect 8757 20043 8815 20049
rect 8757 20040 8769 20043
rect 8628 20012 8769 20040
rect 8628 20000 8634 20012
rect 8757 20009 8769 20012
rect 8803 20009 8815 20043
rect 8757 20003 8815 20009
rect 9217 20043 9275 20049
rect 9217 20009 9229 20043
rect 9263 20040 9275 20043
rect 10134 20040 10140 20052
rect 9263 20012 10140 20040
rect 9263 20009 9275 20012
rect 9217 20003 9275 20009
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 11422 20000 11428 20052
rect 11480 20040 11486 20052
rect 12342 20040 12348 20052
rect 11480 20012 12348 20040
rect 11480 20000 11486 20012
rect 12342 20000 12348 20012
rect 12400 20040 12406 20052
rect 17681 20043 17739 20049
rect 12400 20012 17264 20040
rect 12400 20000 12406 20012
rect 12526 19932 12532 19984
rect 12584 19972 12590 19984
rect 12805 19975 12863 19981
rect 12805 19972 12817 19975
rect 12584 19944 12817 19972
rect 12584 19932 12590 19944
rect 12805 19941 12817 19944
rect 12851 19972 12863 19975
rect 14185 19975 14243 19981
rect 14185 19972 14197 19975
rect 12851 19944 14197 19972
rect 12851 19941 12863 19944
rect 12805 19935 12863 19941
rect 14185 19941 14197 19944
rect 14231 19972 14243 19975
rect 17236 19972 17264 20012
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 18046 20040 18052 20052
rect 17727 20012 18052 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18693 20043 18751 20049
rect 18693 20040 18705 20043
rect 18472 20012 18705 20040
rect 18472 20000 18478 20012
rect 18693 20009 18705 20012
rect 18739 20009 18751 20043
rect 18693 20003 18751 20009
rect 19058 20000 19064 20052
rect 19116 20040 19122 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19116 20012 19717 20040
rect 19116 20000 19122 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 21266 20040 21272 20052
rect 19705 20003 19763 20009
rect 19996 20012 21272 20040
rect 19996 19972 20024 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21361 20043 21419 20049
rect 21361 20009 21373 20043
rect 21407 20040 21419 20043
rect 21450 20040 21456 20052
rect 21407 20012 21456 20040
rect 21407 20009 21419 20012
rect 21361 20003 21419 20009
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 21634 20000 21640 20052
rect 21692 20000 21698 20052
rect 22002 20000 22008 20052
rect 22060 20040 22066 20052
rect 22554 20040 22560 20052
rect 22060 20012 22560 20040
rect 22060 20000 22066 20012
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 23753 20043 23811 20049
rect 23753 20040 23765 20043
rect 22664 20012 23765 20040
rect 14231 19944 15148 19972
rect 17236 19944 20024 19972
rect 14231 19941 14243 19944
rect 14185 19935 14243 19941
rect 3970 19864 3976 19916
rect 4028 19904 4034 19916
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 4028 19876 5457 19904
rect 4028 19864 4034 19876
rect 5445 19873 5457 19876
rect 5491 19904 5503 19907
rect 5626 19904 5632 19916
rect 5491 19876 5632 19904
rect 5491 19873 5503 19876
rect 5445 19867 5503 19873
rect 5626 19864 5632 19876
rect 5684 19864 5690 19916
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 9640 19876 11284 19904
rect 9640 19864 9646 19876
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19805 9551 19839
rect 9493 19799 9551 19805
rect 7282 19768 7288 19780
rect 6196 19740 7288 19768
rect 3418 19660 3424 19712
rect 3476 19700 3482 19712
rect 4709 19703 4767 19709
rect 4709 19700 4721 19703
rect 3476 19672 4721 19700
rect 3476 19660 3482 19672
rect 4709 19669 4721 19672
rect 4755 19700 4767 19703
rect 5077 19703 5135 19709
rect 5077 19700 5089 19703
rect 4755 19672 5089 19700
rect 4755 19669 4767 19672
rect 4709 19663 4767 19669
rect 5077 19669 5089 19672
rect 5123 19700 5135 19703
rect 5813 19703 5871 19709
rect 5813 19700 5825 19703
rect 5123 19672 5825 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5813 19669 5825 19672
rect 5859 19700 5871 19703
rect 5902 19700 5908 19712
rect 5859 19672 5908 19700
rect 5859 19669 5871 19672
rect 5813 19663 5871 19669
rect 5902 19660 5908 19672
rect 5960 19700 5966 19712
rect 6196 19709 6224 19740
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 9508 19768 9536 19799
rect 9674 19796 9680 19848
rect 9732 19796 9738 19848
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 11020 19808 11086 19836
rect 11020 19796 11026 19808
rect 9858 19768 9864 19780
rect 9508 19740 9864 19768
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 9953 19771 10011 19777
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 10226 19768 10232 19780
rect 9999 19740 10232 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 11256 19768 11284 19876
rect 11422 19864 11428 19916
rect 11480 19904 11486 19916
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 11480 19876 11621 19904
rect 11480 19864 11486 19876
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 13354 19864 13360 19916
rect 13412 19904 13418 19916
rect 15120 19913 15148 19944
rect 20530 19932 20536 19984
rect 20588 19972 20594 19984
rect 21545 19975 21603 19981
rect 21545 19972 21557 19975
rect 20588 19944 21557 19972
rect 20588 19932 20594 19944
rect 21545 19941 21557 19944
rect 21591 19941 21603 19975
rect 21545 19935 21603 19941
rect 13817 19907 13875 19913
rect 13817 19904 13829 19907
rect 13412 19876 13829 19904
rect 13412 19864 13418 19876
rect 13817 19873 13829 19876
rect 13863 19873 13875 19907
rect 13817 19867 13875 19873
rect 14737 19907 14795 19913
rect 14737 19873 14749 19907
rect 14783 19904 14795 19907
rect 15105 19907 15163 19913
rect 14783 19876 15056 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19836 11759 19839
rect 12158 19836 12164 19848
rect 11747 19808 12164 19836
rect 11747 19805 11759 19808
rect 11701 19799 11759 19805
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 14458 19768 14464 19780
rect 11256 19740 14464 19768
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 6181 19703 6239 19709
rect 6181 19700 6193 19703
rect 5960 19672 6193 19700
rect 5960 19660 5966 19672
rect 6181 19669 6193 19672
rect 6227 19669 6239 19703
rect 6181 19663 6239 19669
rect 6641 19703 6699 19709
rect 6641 19669 6653 19703
rect 6687 19700 6699 19703
rect 6730 19700 6736 19712
rect 6687 19672 6736 19700
rect 6687 19669 6699 19672
rect 6641 19663 6699 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 8113 19703 8171 19709
rect 8113 19669 8125 19703
rect 8159 19700 8171 19703
rect 8386 19700 8392 19712
rect 8159 19672 8392 19700
rect 8159 19669 8171 19672
rect 8113 19663 8171 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 9272 19672 9413 19700
rect 9272 19660 9278 19672
rect 9401 19669 9413 19672
rect 9447 19669 9459 19703
rect 9401 19663 9459 19669
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 11425 19703 11483 19709
rect 11425 19700 11437 19703
rect 10928 19672 11437 19700
rect 10928 19660 10934 19672
rect 11425 19669 11437 19672
rect 11471 19669 11483 19703
rect 11425 19663 11483 19669
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12069 19703 12127 19709
rect 12069 19700 12081 19703
rect 11664 19672 12081 19700
rect 11664 19660 11670 19672
rect 12069 19669 12081 19672
rect 12115 19669 12127 19703
rect 12069 19663 12127 19669
rect 13173 19703 13231 19709
rect 13173 19669 13185 19703
rect 13219 19700 13231 19703
rect 13906 19700 13912 19712
rect 13219 19672 13912 19700
rect 13219 19669 13231 19672
rect 13173 19663 13231 19669
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 14366 19660 14372 19712
rect 14424 19660 14430 19712
rect 14660 19700 14688 19799
rect 14826 19796 14832 19848
rect 14884 19796 14890 19848
rect 15028 19768 15056 19876
rect 15105 19873 15117 19907
rect 15151 19873 15163 19907
rect 15105 19867 15163 19873
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 16022 19904 16028 19916
rect 15519 19876 16028 19904
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 16632 19876 17509 19904
rect 16632 19864 16638 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 17586 19864 17592 19916
rect 17644 19864 17650 19916
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19904 18107 19907
rect 18322 19904 18328 19916
rect 18095 19876 18328 19904
rect 18095 19873 18107 19876
rect 18049 19867 18107 19873
rect 18322 19864 18328 19876
rect 18380 19904 18386 19916
rect 18380 19876 18644 19904
rect 18380 19864 18386 19876
rect 15378 19836 15384 19848
rect 15212 19808 15384 19836
rect 15212 19768 15240 19808
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 16942 19836 16948 19848
rect 16592 19808 16948 19836
rect 15028 19740 15240 19768
rect 15838 19728 15844 19780
rect 15896 19728 15902 19780
rect 15470 19700 15476 19712
rect 14660 19672 15476 19700
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 16592 19700 16620 19808
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17126 19796 17132 19848
rect 17184 19836 17190 19848
rect 17604 19836 17632 19864
rect 17681 19839 17739 19845
rect 17681 19836 17693 19839
rect 17184 19808 17356 19836
rect 17604 19808 17693 19836
rect 17184 19796 17190 19808
rect 17221 19771 17279 19777
rect 17221 19768 17233 19771
rect 16914 19740 17233 19768
rect 15988 19672 16620 19700
rect 15988 19660 15994 19672
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 16914 19709 16942 19740
rect 17221 19737 17233 19740
rect 17267 19737 17279 19771
rect 17221 19731 17279 19737
rect 16899 19703 16957 19709
rect 16899 19700 16911 19703
rect 16816 19672 16911 19700
rect 16816 19660 16822 19672
rect 16899 19669 16911 19672
rect 16945 19669 16957 19703
rect 17328 19700 17356 19808
rect 17681 19805 17693 19808
rect 17727 19805 17739 19839
rect 17681 19799 17739 19805
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 18616 19845 18644 19876
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 18748 19876 19073 19904
rect 18748 19864 18754 19876
rect 19061 19873 19073 19876
rect 19107 19904 19119 19907
rect 19518 19904 19524 19916
rect 19107 19876 19524 19904
rect 19107 19873 19119 19876
rect 19061 19867 19119 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 20622 19904 20628 19916
rect 19904 19876 20628 19904
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17828 19808 17969 19836
rect 17828 19796 17834 19808
rect 17957 19805 17969 19808
rect 18003 19805 18015 19839
rect 18141 19839 18199 19845
rect 17957 19799 18015 19805
rect 18046 19786 18052 19838
rect 18104 19836 18110 19838
rect 18141 19836 18153 19839
rect 18104 19808 18153 19836
rect 18104 19786 18110 19808
rect 18141 19805 18153 19808
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18233 19799 18291 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 18601 19839 18659 19845
rect 18463 19808 18552 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 18248 19768 18276 19799
rect 18322 19768 18328 19780
rect 18248 19740 18328 19768
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 18524 19768 18552 19808
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 19337 19839 19395 19845
rect 19337 19836 19349 19839
rect 18601 19799 18659 19805
rect 18708 19808 19349 19836
rect 18708 19768 18736 19808
rect 19337 19805 19349 19808
rect 19383 19836 19395 19839
rect 19426 19836 19432 19848
rect 19383 19808 19432 19836
rect 19383 19805 19395 19808
rect 19337 19799 19395 19805
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 19904 19845 19932 19876
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 20990 19904 20996 19916
rect 20855 19876 20996 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 19852 19808 19901 19836
rect 19852 19796 19858 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19836 20039 19839
rect 20027 19808 20208 19836
rect 20027 19805 20039 19808
rect 19981 19799 20039 19805
rect 20180 19780 20208 19808
rect 20254 19796 20260 19848
rect 20312 19796 20318 19848
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20395 19808 20668 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 18524 19740 18736 19768
rect 18966 19728 18972 19780
rect 19024 19728 19030 19780
rect 19058 19728 19064 19780
rect 19116 19768 19122 19780
rect 19153 19771 19211 19777
rect 19153 19768 19165 19771
rect 19116 19740 19165 19768
rect 19116 19728 19122 19740
rect 19153 19737 19165 19740
rect 19199 19768 19211 19771
rect 19199 19740 20024 19768
rect 19199 19737 19211 19740
rect 19153 19731 19211 19737
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 17328 19672 17877 19700
rect 16899 19663 16957 19669
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 18417 19703 18475 19709
rect 18417 19700 18429 19703
rect 18196 19672 18429 19700
rect 18196 19660 18202 19672
rect 18417 19669 18429 19672
rect 18463 19700 18475 19703
rect 18984 19700 19012 19728
rect 18463 19672 19012 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 19518 19660 19524 19712
rect 19576 19660 19582 19712
rect 19996 19700 20024 19740
rect 20070 19728 20076 19780
rect 20128 19728 20134 19780
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 20640 19768 20668 19808
rect 20714 19796 20720 19848
rect 20772 19796 20778 19848
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19836 21603 19839
rect 21652 19836 21680 20000
rect 21910 19972 21916 19984
rect 21836 19944 21916 19972
rect 21591 19808 21680 19836
rect 21591 19805 21603 19808
rect 21545 19799 21603 19805
rect 20916 19768 20944 19799
rect 21726 19796 21732 19848
rect 21784 19796 21790 19848
rect 21836 19845 21864 19944
rect 21910 19932 21916 19944
rect 21968 19972 21974 19984
rect 22664 19972 22692 20012
rect 23753 20009 23765 20012
rect 23799 20009 23811 20043
rect 23753 20003 23811 20009
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 27985 20043 28043 20049
rect 27985 20040 27997 20043
rect 27580 20012 27997 20040
rect 27580 20000 27586 20012
rect 27985 20009 27997 20012
rect 28031 20009 28043 20043
rect 33134 20040 33140 20052
rect 27985 20003 28043 20009
rect 30576 20012 31340 20040
rect 21968 19944 22692 19972
rect 23201 19975 23259 19981
rect 21968 19932 21974 19944
rect 23201 19941 23213 19975
rect 23247 19972 23259 19975
rect 24118 19972 24124 19984
rect 23247 19944 24124 19972
rect 23247 19941 23259 19944
rect 23201 19935 23259 19941
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 27614 19932 27620 19984
rect 27672 19972 27678 19984
rect 28629 19975 28687 19981
rect 28629 19972 28641 19975
rect 27672 19944 28641 19972
rect 27672 19932 27678 19944
rect 28629 19941 28641 19944
rect 28675 19941 28687 19975
rect 28629 19935 28687 19941
rect 22278 19864 22284 19916
rect 22336 19864 22342 19916
rect 24302 19864 24308 19916
rect 24360 19864 24366 19916
rect 25406 19864 25412 19916
rect 25464 19864 25470 19916
rect 25958 19864 25964 19916
rect 26016 19904 26022 19916
rect 26234 19904 26240 19916
rect 26016 19876 26240 19904
rect 26016 19864 26022 19876
rect 26234 19864 26240 19876
rect 26292 19904 26298 19916
rect 28166 19904 28172 19916
rect 26292 19876 28172 19904
rect 26292 19864 26298 19876
rect 28166 19864 28172 19876
rect 28224 19904 28230 19916
rect 28905 19907 28963 19913
rect 28905 19904 28917 19907
rect 28224 19876 28917 19904
rect 28224 19864 28230 19876
rect 28905 19873 28917 19876
rect 28951 19873 28963 19907
rect 28905 19867 28963 19873
rect 29181 19907 29239 19913
rect 29181 19873 29193 19907
rect 29227 19904 29239 19907
rect 30576 19904 30604 20012
rect 30650 19932 30656 19984
rect 30708 19972 30714 19984
rect 31312 19981 31340 20012
rect 32600 20012 33140 20040
rect 31297 19975 31355 19981
rect 30708 19944 30972 19972
rect 30708 19932 30714 19944
rect 29227 19876 30604 19904
rect 29227 19873 29239 19876
rect 29181 19867 29239 19873
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19805 21971 19839
rect 21913 19799 21971 19805
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 22296 19836 22324 19864
rect 22143 19808 22324 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 21928 19768 21956 19799
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 24213 19839 24271 19845
rect 24213 19836 24225 19839
rect 23348 19808 24225 19836
rect 23348 19796 23354 19808
rect 24213 19805 24225 19808
rect 24259 19836 24271 19839
rect 25317 19839 25375 19845
rect 25317 19836 25329 19839
rect 24259 19808 25329 19836
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 25317 19805 25329 19808
rect 25363 19805 25375 19839
rect 27890 19836 27896 19848
rect 27646 19808 27896 19836
rect 25317 19799 25375 19805
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 27982 19796 27988 19848
rect 28040 19836 28046 19848
rect 28077 19839 28135 19845
rect 28077 19836 28089 19839
rect 28040 19808 28089 19836
rect 28040 19796 28046 19808
rect 28077 19805 28089 19808
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 22186 19768 22192 19780
rect 20640 19740 20944 19768
rect 21192 19740 21588 19768
rect 21928 19740 22192 19768
rect 20640 19712 20668 19740
rect 20254 19700 20260 19712
rect 19996 19672 20260 19700
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20438 19660 20444 19712
rect 20496 19660 20502 19712
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 21192 19700 21220 19740
rect 20864 19672 21220 19700
rect 21560 19700 21588 19740
rect 22186 19728 22192 19740
rect 22244 19768 22250 19780
rect 23474 19768 23480 19780
rect 22244 19740 23480 19768
rect 22244 19728 22250 19740
rect 23474 19728 23480 19740
rect 23532 19728 23538 19780
rect 23569 19771 23627 19777
rect 23569 19737 23581 19771
rect 23615 19768 23627 19771
rect 23934 19768 23940 19780
rect 23615 19740 23940 19768
rect 23615 19737 23627 19740
rect 23569 19731 23627 19737
rect 23934 19728 23940 19740
rect 23992 19728 23998 19780
rect 25225 19771 25283 19777
rect 25225 19737 25237 19771
rect 25271 19768 25283 19771
rect 25271 19740 26464 19768
rect 25271 19737 25283 19740
rect 25225 19731 25283 19737
rect 22002 19700 22008 19712
rect 21560 19672 22008 19700
rect 20864 19660 20870 19672
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 22370 19660 22376 19712
rect 22428 19660 22434 19712
rect 22833 19703 22891 19709
rect 22833 19669 22845 19703
rect 22879 19700 22891 19703
rect 24026 19700 24032 19712
rect 22879 19672 24032 19700
rect 22879 19669 22891 19672
rect 22833 19663 22891 19669
rect 24026 19660 24032 19672
rect 24084 19700 24090 19712
rect 24121 19703 24179 19709
rect 24121 19700 24133 19703
rect 24084 19672 24133 19700
rect 24084 19660 24090 19672
rect 24121 19669 24133 19672
rect 24167 19669 24179 19703
rect 24121 19663 24179 19669
rect 24854 19660 24860 19712
rect 24912 19660 24918 19712
rect 26436 19700 26464 19740
rect 26510 19728 26516 19780
rect 26568 19728 26574 19780
rect 28092 19768 28120 19799
rect 28166 19768 28172 19780
rect 28092 19740 28172 19768
rect 28166 19728 28172 19740
rect 28224 19728 28230 19780
rect 28258 19728 28264 19780
rect 28316 19728 28322 19780
rect 28353 19771 28411 19777
rect 28353 19737 28365 19771
rect 28399 19737 28411 19771
rect 28353 19731 28411 19737
rect 27798 19700 27804 19712
rect 26436 19672 27804 19700
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 28074 19660 28080 19712
rect 28132 19700 28138 19712
rect 28368 19700 28396 19731
rect 28132 19672 28396 19700
rect 28460 19700 28488 19799
rect 30282 19796 30288 19848
rect 30340 19796 30346 19848
rect 30742 19796 30748 19848
rect 30800 19845 30806 19848
rect 30800 19839 30823 19845
rect 30811 19805 30823 19839
rect 30944 19836 30972 19944
rect 31297 19941 31309 19975
rect 31343 19941 31355 19975
rect 31297 19935 31355 19941
rect 31846 19864 31852 19916
rect 31904 19864 31910 19916
rect 32125 19907 32183 19913
rect 32125 19873 32137 19907
rect 32171 19904 32183 19907
rect 32600 19904 32628 20012
rect 33134 20000 33140 20012
rect 33192 20040 33198 20052
rect 34241 20043 34299 20049
rect 34241 20040 34253 20043
rect 33192 20012 34253 20040
rect 33192 20000 33198 20012
rect 32677 19975 32735 19981
rect 32677 19941 32689 19975
rect 32723 19941 32735 19975
rect 32677 19935 32735 19941
rect 32171 19876 32628 19904
rect 32171 19873 32183 19876
rect 32125 19867 32183 19873
rect 31017 19839 31075 19845
rect 31017 19836 31029 19839
rect 30944 19808 31029 19836
rect 30800 19799 30823 19805
rect 31017 19805 31029 19808
rect 31063 19805 31075 19839
rect 31017 19799 31075 19805
rect 30800 19796 30806 19799
rect 31110 19796 31116 19848
rect 31168 19836 31174 19848
rect 31864 19836 31892 19864
rect 31168 19808 31892 19836
rect 32309 19839 32367 19845
rect 31168 19796 31174 19808
rect 32309 19805 32321 19839
rect 32355 19836 32367 19839
rect 32692 19836 32720 19935
rect 33336 19913 33364 20012
rect 34241 20009 34253 20012
rect 34287 20009 34299 20043
rect 34241 20003 34299 20009
rect 35986 20000 35992 20052
rect 36044 20040 36050 20052
rect 36173 20043 36231 20049
rect 36173 20040 36185 20043
rect 36044 20012 36185 20040
rect 36044 20000 36050 20012
rect 36173 20009 36185 20012
rect 36219 20009 36231 20043
rect 36173 20003 36231 20009
rect 36633 20043 36691 20049
rect 36633 20009 36645 20043
rect 36679 20040 36691 20043
rect 37642 20040 37648 20052
rect 36679 20012 37648 20040
rect 36679 20009 36691 20012
rect 36633 20003 36691 20009
rect 37642 20000 37648 20012
rect 37700 20000 37706 20052
rect 41690 20040 41696 20052
rect 38580 20012 41696 20040
rect 38470 19972 38476 19984
rect 37108 19944 38476 19972
rect 33321 19907 33379 19913
rect 33321 19873 33333 19907
rect 33367 19904 33379 19907
rect 33502 19904 33508 19916
rect 33367 19876 33508 19904
rect 33367 19873 33379 19876
rect 33321 19867 33379 19873
rect 33502 19864 33508 19876
rect 33560 19864 33566 19916
rect 35066 19864 35072 19916
rect 35124 19904 35130 19916
rect 37108 19913 37136 19944
rect 35713 19907 35771 19913
rect 35713 19904 35725 19907
rect 35124 19876 35725 19904
rect 35124 19864 35130 19876
rect 35713 19873 35725 19876
rect 35759 19873 35771 19907
rect 35713 19867 35771 19873
rect 37093 19907 37151 19913
rect 37093 19873 37105 19907
rect 37139 19873 37151 19907
rect 37093 19867 37151 19873
rect 37182 19864 37188 19916
rect 37240 19904 37246 19916
rect 38013 19907 38071 19913
rect 38013 19904 38025 19907
rect 37240 19876 38025 19904
rect 37240 19864 37246 19876
rect 38013 19873 38025 19876
rect 38059 19873 38071 19907
rect 38013 19867 38071 19873
rect 32355 19808 32720 19836
rect 33045 19839 33103 19845
rect 32355 19805 32367 19808
rect 32309 19799 32367 19805
rect 33045 19805 33057 19839
rect 33091 19836 33103 19839
rect 33091 19808 34836 19836
rect 33091 19805 33103 19808
rect 33045 19799 33103 19805
rect 30760 19768 30788 19796
rect 30668 19740 30788 19768
rect 30929 19771 30987 19777
rect 28534 19700 28540 19712
rect 28460 19672 28540 19700
rect 28132 19660 28138 19672
rect 28534 19660 28540 19672
rect 28592 19700 28598 19712
rect 28902 19700 28908 19712
rect 28592 19672 28908 19700
rect 28592 19660 28598 19672
rect 28902 19660 28908 19672
rect 28960 19700 28966 19712
rect 29822 19700 29828 19712
rect 28960 19672 29828 19700
rect 28960 19660 28966 19672
rect 29822 19660 29828 19672
rect 29880 19660 29886 19712
rect 30006 19660 30012 19712
rect 30064 19700 30070 19712
rect 30668 19700 30696 19740
rect 30929 19737 30941 19771
rect 30975 19768 30987 19771
rect 31849 19771 31907 19777
rect 30975 19740 31051 19768
rect 30975 19737 30987 19740
rect 30929 19731 30987 19737
rect 30064 19672 30696 19700
rect 30064 19660 30070 19672
rect 30742 19660 30748 19712
rect 30800 19700 30806 19712
rect 31023 19700 31051 19740
rect 31849 19737 31861 19771
rect 31895 19768 31907 19771
rect 32766 19768 32772 19780
rect 31895 19740 32772 19768
rect 31895 19737 31907 19740
rect 31849 19731 31907 19737
rect 32766 19728 32772 19740
rect 32824 19728 32830 19780
rect 33318 19728 33324 19780
rect 33376 19768 33382 19780
rect 34146 19768 34152 19780
rect 33376 19740 34152 19768
rect 33376 19728 33382 19740
rect 34146 19728 34152 19740
rect 34204 19728 34210 19780
rect 34808 19768 34836 19808
rect 34882 19796 34888 19848
rect 34940 19796 34946 19848
rect 35529 19839 35587 19845
rect 35529 19805 35541 19839
rect 35575 19836 35587 19839
rect 35802 19836 35808 19848
rect 35575 19808 35808 19836
rect 35575 19805 35587 19808
rect 35529 19799 35587 19805
rect 35802 19796 35808 19808
rect 35860 19796 35866 19848
rect 37001 19839 37059 19845
rect 37001 19805 37013 19839
rect 37047 19836 37059 19839
rect 37274 19836 37280 19848
rect 37047 19808 37280 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 37274 19796 37280 19808
rect 37332 19796 37338 19848
rect 37829 19839 37887 19845
rect 37829 19805 37841 19839
rect 37875 19836 37887 19839
rect 38120 19836 38148 19944
rect 38470 19932 38476 19944
rect 38528 19932 38534 19984
rect 37875 19808 38148 19836
rect 37875 19805 37887 19808
rect 37829 19799 37887 19805
rect 38470 19796 38476 19848
rect 38528 19796 38534 19848
rect 38580 19768 38608 20012
rect 41690 20000 41696 20012
rect 41748 20000 41754 20052
rect 44174 20000 44180 20052
rect 44232 20040 44238 20052
rect 44545 20043 44603 20049
rect 44545 20040 44557 20043
rect 44232 20012 44557 20040
rect 44232 20000 44238 20012
rect 44545 20009 44557 20012
rect 44591 20009 44603 20043
rect 44545 20003 44603 20009
rect 44910 20000 44916 20052
rect 44968 20000 44974 20052
rect 39390 19932 39396 19984
rect 39448 19932 39454 19984
rect 39850 19864 39856 19916
rect 39908 19904 39914 19916
rect 40129 19907 40187 19913
rect 40129 19904 40141 19907
rect 39908 19876 40141 19904
rect 39908 19864 39914 19876
rect 40129 19873 40141 19876
rect 40175 19873 40187 19907
rect 41414 19904 41420 19916
rect 40129 19867 40187 19873
rect 40328 19876 41420 19904
rect 38746 19796 38752 19848
rect 38804 19796 38810 19848
rect 40037 19839 40095 19845
rect 40037 19805 40049 19839
rect 40083 19836 40095 19839
rect 40328 19836 40356 19876
rect 41414 19864 41420 19876
rect 41472 19864 41478 19916
rect 42245 19907 42303 19913
rect 42245 19904 42257 19907
rect 42076 19876 42257 19904
rect 42076 19848 42104 19876
rect 42245 19873 42257 19876
rect 42291 19873 42303 19907
rect 42245 19867 42303 19873
rect 42521 19907 42579 19913
rect 42521 19873 42533 19907
rect 42567 19904 42579 19907
rect 42610 19904 42616 19916
rect 42567 19876 42616 19904
rect 42567 19873 42579 19876
rect 42521 19867 42579 19873
rect 42610 19864 42616 19876
rect 42668 19864 42674 19916
rect 40083 19808 40356 19836
rect 40405 19839 40463 19845
rect 40083 19805 40095 19808
rect 40037 19799 40095 19805
rect 40405 19805 40417 19839
rect 40451 19805 40463 19839
rect 40405 19799 40463 19805
rect 34808 19740 38608 19768
rect 39206 19728 39212 19780
rect 39264 19768 39270 19780
rect 40420 19768 40448 19799
rect 42058 19796 42064 19848
rect 42116 19796 42122 19848
rect 39264 19740 40448 19768
rect 40681 19771 40739 19777
rect 39264 19728 39270 19740
rect 40681 19737 40693 19771
rect 40727 19737 40739 19771
rect 40681 19731 40739 19737
rect 30800 19672 31051 19700
rect 30800 19660 30806 19672
rect 31478 19660 31484 19712
rect 31536 19660 31542 19712
rect 31938 19660 31944 19712
rect 31996 19660 32002 19712
rect 32490 19660 32496 19712
rect 32548 19660 32554 19712
rect 33134 19660 33140 19712
rect 33192 19660 33198 19712
rect 33781 19703 33839 19709
rect 33781 19669 33793 19703
rect 33827 19700 33839 19703
rect 34422 19700 34428 19712
rect 33827 19672 34428 19700
rect 33827 19669 33839 19672
rect 33781 19663 33839 19669
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 34698 19660 34704 19712
rect 34756 19660 34762 19712
rect 35158 19660 35164 19712
rect 35216 19660 35222 19712
rect 35621 19703 35679 19709
rect 35621 19669 35633 19703
rect 35667 19700 35679 19703
rect 35802 19700 35808 19712
rect 35667 19672 35808 19700
rect 35667 19669 35679 19672
rect 35621 19663 35679 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 37274 19660 37280 19712
rect 37332 19700 37338 19712
rect 37461 19703 37519 19709
rect 37461 19700 37473 19703
rect 37332 19672 37473 19700
rect 37332 19660 37338 19672
rect 37461 19669 37473 19672
rect 37507 19669 37519 19703
rect 37461 19663 37519 19669
rect 37918 19660 37924 19712
rect 37976 19660 37982 19712
rect 38286 19660 38292 19712
rect 38344 19660 38350 19712
rect 39574 19660 39580 19712
rect 39632 19660 39638 19712
rect 39942 19660 39948 19712
rect 40000 19660 40006 19712
rect 40696 19700 40724 19731
rect 40770 19728 40776 19780
rect 40828 19768 40834 19780
rect 40828 19740 41170 19768
rect 40828 19728 40834 19740
rect 42794 19728 42800 19780
rect 42852 19768 42858 19780
rect 42852 19740 43010 19768
rect 42852 19728 42858 19740
rect 40862 19700 40868 19712
rect 40696 19672 40868 19700
rect 40862 19660 40868 19672
rect 40920 19660 40926 19712
rect 42150 19660 42156 19712
rect 42208 19660 42214 19712
rect 43990 19660 43996 19712
rect 44048 19660 44054 19712
rect 460 19610 45540 19632
rect 460 19558 6070 19610
rect 6122 19558 6134 19610
rect 6186 19558 6198 19610
rect 6250 19558 6262 19610
rect 6314 19558 6326 19610
rect 6378 19558 11070 19610
rect 11122 19558 11134 19610
rect 11186 19558 11198 19610
rect 11250 19558 11262 19610
rect 11314 19558 11326 19610
rect 11378 19558 16070 19610
rect 16122 19558 16134 19610
rect 16186 19558 16198 19610
rect 16250 19558 16262 19610
rect 16314 19558 16326 19610
rect 16378 19558 21070 19610
rect 21122 19558 21134 19610
rect 21186 19558 21198 19610
rect 21250 19558 21262 19610
rect 21314 19558 21326 19610
rect 21378 19558 26070 19610
rect 26122 19558 26134 19610
rect 26186 19558 26198 19610
rect 26250 19558 26262 19610
rect 26314 19558 26326 19610
rect 26378 19558 31070 19610
rect 31122 19558 31134 19610
rect 31186 19558 31198 19610
rect 31250 19558 31262 19610
rect 31314 19558 31326 19610
rect 31378 19558 36070 19610
rect 36122 19558 36134 19610
rect 36186 19558 36198 19610
rect 36250 19558 36262 19610
rect 36314 19558 36326 19610
rect 36378 19558 41070 19610
rect 41122 19558 41134 19610
rect 41186 19558 41198 19610
rect 41250 19558 41262 19610
rect 41314 19558 41326 19610
rect 41378 19558 45540 19610
rect 460 19536 45540 19558
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 8294 19496 8300 19508
rect 7791 19468 8300 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 8386 19456 8392 19508
rect 8444 19456 8450 19508
rect 9214 19456 9220 19508
rect 9272 19456 9278 19508
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 10321 19499 10379 19505
rect 10321 19496 10333 19499
rect 9640 19468 10333 19496
rect 9640 19456 9646 19468
rect 10321 19465 10333 19468
rect 10367 19465 10379 19499
rect 10962 19496 10968 19508
rect 10321 19459 10379 19465
rect 10428 19468 10968 19496
rect 5534 19388 5540 19440
rect 5592 19428 5598 19440
rect 8202 19428 8208 19440
rect 5592 19400 8208 19428
rect 5592 19388 5598 19400
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 6822 19360 6828 19372
rect 6288 19332 6828 19360
rect 5537 19159 5595 19165
rect 5537 19125 5549 19159
rect 5583 19156 5595 19159
rect 5644 19156 5672 19320
rect 5994 19156 6000 19168
rect 5583 19128 6000 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5994 19116 6000 19128
rect 6052 19156 6058 19168
rect 6288 19165 6316 19332
rect 6822 19320 6828 19332
rect 6880 19360 6886 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6880 19332 7021 19360
rect 6880 19320 6886 19332
rect 7009 19329 7021 19332
rect 7055 19360 7067 19363
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 7055 19332 7389 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7558 19320 7564 19372
rect 7616 19320 7622 19372
rect 7742 19320 7748 19372
rect 7800 19320 7806 19372
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 8404 19360 8432 19456
rect 8849 19431 8907 19437
rect 8849 19397 8861 19431
rect 8895 19428 8907 19431
rect 9232 19428 9260 19456
rect 10134 19428 10140 19440
rect 8895 19400 9260 19428
rect 10074 19400 10140 19428
rect 8895 19397 8907 19400
rect 8849 19391 8907 19397
rect 10134 19388 10140 19400
rect 10192 19428 10198 19440
rect 10428 19428 10456 19468
rect 10962 19456 10968 19468
rect 11020 19496 11026 19508
rect 11020 19468 11284 19496
rect 11020 19456 11026 19468
rect 10192 19400 10456 19428
rect 10192 19388 10198 19400
rect 10870 19388 10876 19440
rect 10928 19388 10934 19440
rect 11256 19428 11284 19468
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 12621 19499 12679 19505
rect 12621 19496 12633 19499
rect 12216 19468 12633 19496
rect 12216 19456 12222 19468
rect 12621 19465 12633 19468
rect 12667 19465 12679 19499
rect 14734 19496 14740 19508
rect 12621 19459 12679 19465
rect 12912 19468 14740 19496
rect 11256 19400 11638 19428
rect 8168 19332 8432 19360
rect 8168 19320 8174 19332
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 9858 19320 9864 19372
rect 9916 19320 9922 19372
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19329 10471 19363
rect 10413 19323 10471 19329
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19360 10655 19363
rect 10888 19360 10916 19388
rect 10643 19332 10916 19360
rect 12912 19360 12940 19468
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 14826 19456 14832 19508
rect 14884 19456 14890 19508
rect 15930 19496 15936 19508
rect 15764 19468 15936 19496
rect 13906 19388 13912 19440
rect 13964 19388 13970 19440
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 15473 19431 15531 19437
rect 15068 19400 15286 19428
rect 15068 19388 15074 19400
rect 15258 19394 15286 19400
rect 15473 19397 15485 19431
rect 15519 19428 15531 19431
rect 15764 19428 15792 19468
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 16574 19496 16580 19508
rect 16040 19468 16580 19496
rect 15519 19400 15792 19428
rect 15519 19397 15531 19400
rect 13173 19363 13231 19369
rect 15258 19366 15424 19394
rect 15473 19391 15531 19397
rect 13173 19360 13185 19363
rect 12912 19332 13185 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 13173 19329 13185 19332
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 15290 19363 15424 19366
rect 15290 19329 15302 19363
rect 15336 19342 15424 19363
rect 15336 19329 15348 19342
rect 15290 19323 15348 19329
rect 6730 19252 6736 19304
rect 6788 19252 6794 19304
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 8128 19224 8156 19320
rect 8386 19252 8392 19304
rect 8444 19292 8450 19304
rect 8588 19292 8616 19320
rect 8444 19264 8616 19292
rect 9876 19292 9904 19320
rect 10428 19292 10456 19323
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15657 19363 15715 19369
rect 15657 19360 15669 19363
rect 15620 19332 15669 19360
rect 15620 19320 15626 19332
rect 15657 19329 15669 19332
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 15746 19320 15752 19372
rect 15804 19320 15810 19372
rect 16040 19369 16068 19468
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 17460 19468 18184 19496
rect 17460 19456 17466 19468
rect 16758 19428 16764 19440
rect 16316 19400 16764 19428
rect 16316 19369 16344 19400
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 17034 19428 17040 19440
rect 16868 19400 17040 19428
rect 16025 19363 16083 19369
rect 16025 19329 16037 19363
rect 16071 19329 16083 19363
rect 16025 19323 16083 19329
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 16868 19360 16896 19400
rect 17034 19388 17040 19400
rect 17092 19428 17098 19440
rect 17586 19428 17592 19440
rect 17092 19400 17592 19428
rect 17092 19388 17098 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 17678 19388 17684 19440
rect 17736 19428 17742 19440
rect 18156 19428 18184 19468
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18288 19468 18981 19496
rect 18288 19456 18294 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 19150 19456 19156 19508
rect 19208 19456 19214 19508
rect 19518 19456 19524 19508
rect 19576 19456 19582 19508
rect 20162 19496 20168 19508
rect 19904 19468 20168 19496
rect 18690 19428 18696 19440
rect 17736 19400 18000 19428
rect 18156 19400 18696 19428
rect 17736 19388 17742 19400
rect 16715 19332 16896 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 16942 19320 16948 19372
rect 17000 19320 17006 19372
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 17972 19369 18000 19400
rect 18616 19369 18644 19400
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 19168 19428 19196 19456
rect 18800 19400 19196 19428
rect 18800 19369 18828 19400
rect 17957 19363 18015 19369
rect 17552 19332 17908 19360
rect 17552 19320 17558 19332
rect 10686 19292 10692 19304
rect 9876 19264 10692 19292
rect 8444 19252 8450 19264
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10873 19295 10931 19301
rect 10873 19292 10885 19295
rect 10836 19264 10885 19292
rect 10836 19252 10842 19264
rect 10873 19261 10885 19264
rect 10919 19292 10931 19295
rect 12802 19292 12808 19304
rect 10919 19264 12808 19292
rect 10919 19261 10931 19264
rect 10873 19255 10931 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15106 19295 15164 19301
rect 15106 19261 15118 19295
rect 15152 19261 15164 19295
rect 15106 19255 15164 19261
rect 6696 19196 8156 19224
rect 6696 19184 6702 19196
rect 6273 19159 6331 19165
rect 6273 19156 6285 19159
rect 6052 19128 6285 19156
rect 6052 19116 6058 19128
rect 6273 19125 6285 19128
rect 6319 19125 6331 19159
rect 6273 19119 6331 19125
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10505 19159 10563 19165
rect 10505 19156 10517 19159
rect 10468 19128 10517 19156
rect 10468 19116 10474 19128
rect 10505 19125 10517 19128
rect 10551 19125 10563 19159
rect 10505 19119 10563 19125
rect 11136 19159 11194 19165
rect 11136 19125 11148 19159
rect 11182 19156 11194 19159
rect 11606 19156 11612 19168
rect 11182 19128 11612 19156
rect 11182 19125 11194 19128
rect 11136 19119 11194 19125
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 14599 19159 14657 19165
rect 14599 19125 14611 19159
rect 14645 19156 14657 19159
rect 14826 19156 14832 19168
rect 14645 19128 14832 19156
rect 14645 19125 14657 19128
rect 14599 19119 14657 19125
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 15028 19156 15056 19255
rect 15120 19224 15148 19255
rect 15194 19252 15200 19304
rect 15252 19252 15258 19304
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 16206 19292 16212 19304
rect 15436 19264 16212 19292
rect 15436 19252 15442 19264
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 16960 19292 16988 19320
rect 16439 19264 16988 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17678 19292 17684 19304
rect 17276 19264 17684 19292
rect 17276 19252 17282 19264
rect 17678 19252 17684 19264
rect 17736 19252 17742 19304
rect 17880 19292 17908 19332
rect 17957 19329 17969 19363
rect 18003 19329 18015 19363
rect 17957 19323 18015 19329
rect 18233 19363 18291 19369
rect 18233 19329 18245 19363
rect 18279 19360 18291 19363
rect 18601 19363 18659 19369
rect 18279 19332 18368 19360
rect 18279 19329 18291 19332
rect 18233 19323 18291 19329
rect 18340 19292 18368 19332
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19329 18843 19363
rect 18785 19323 18843 19329
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 19024 19332 19073 19360
rect 19024 19320 19030 19332
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19536 19360 19564 19456
rect 19904 19437 19932 19468
rect 20162 19456 20168 19468
rect 20220 19496 20226 19508
rect 20714 19496 20720 19508
rect 20220 19468 20720 19496
rect 20220 19456 20226 19468
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21637 19499 21695 19505
rect 21637 19496 21649 19499
rect 20864 19468 21649 19496
rect 20864 19456 20870 19468
rect 21637 19465 21649 19468
rect 21683 19465 21695 19499
rect 21637 19459 21695 19465
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 24581 19499 24639 19505
rect 24581 19496 24593 19499
rect 23348 19468 24593 19496
rect 23348 19456 23354 19468
rect 24581 19465 24593 19468
rect 24627 19465 24639 19499
rect 24581 19459 24639 19465
rect 24854 19456 24860 19508
rect 24912 19456 24918 19508
rect 25593 19499 25651 19505
rect 25593 19465 25605 19499
rect 25639 19496 25651 19499
rect 26234 19496 26240 19508
rect 25639 19468 26240 19496
rect 25639 19465 25651 19468
rect 25593 19459 25651 19465
rect 26234 19456 26240 19468
rect 26292 19456 26298 19508
rect 26510 19456 26516 19508
rect 26568 19496 26574 19508
rect 27893 19499 27951 19505
rect 27893 19496 27905 19499
rect 26568 19468 27905 19496
rect 26568 19456 26574 19468
rect 27893 19465 27905 19468
rect 27939 19465 27951 19499
rect 27893 19459 27951 19465
rect 28350 19456 28356 19508
rect 28408 19496 28414 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 28408 19468 28917 19496
rect 28408 19456 28414 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 28905 19459 28963 19465
rect 29914 19456 29920 19508
rect 29972 19496 29978 19508
rect 29972 19468 30420 19496
rect 29972 19456 29978 19468
rect 19889 19431 19947 19437
rect 19889 19428 19901 19431
rect 19291 19332 19564 19360
rect 19628 19400 19901 19428
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 17880 19264 18368 19292
rect 15286 19224 15292 19236
rect 15120 19196 15292 19224
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15396 19224 15424 19252
rect 15473 19227 15531 19233
rect 15473 19224 15485 19227
rect 15396 19196 15485 19224
rect 15473 19193 15485 19196
rect 15519 19193 15531 19227
rect 15473 19187 15531 19193
rect 16853 19227 16911 19233
rect 16853 19193 16865 19227
rect 16899 19193 16911 19227
rect 16853 19187 16911 19193
rect 15746 19156 15752 19168
rect 15028 19128 15752 19156
rect 15746 19116 15752 19128
rect 15804 19156 15810 19168
rect 16666 19156 16672 19168
rect 15804 19128 16672 19156
rect 15804 19116 15810 19128
rect 16666 19116 16672 19128
rect 16724 19156 16730 19168
rect 16868 19156 16896 19187
rect 17954 19184 17960 19236
rect 18012 19224 18018 19236
rect 18049 19227 18107 19233
rect 18049 19224 18061 19227
rect 18012 19196 18061 19224
rect 18012 19184 18018 19196
rect 18049 19193 18061 19196
rect 18095 19193 18107 19227
rect 18340 19224 18368 19264
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 19628 19292 19656 19400
rect 19889 19397 19901 19400
rect 19935 19397 19947 19431
rect 19889 19391 19947 19397
rect 21177 19431 21235 19437
rect 21177 19397 21189 19431
rect 21223 19428 21235 19431
rect 21726 19428 21732 19440
rect 21223 19400 21732 19428
rect 21223 19397 21235 19400
rect 21177 19391 21235 19397
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 24872 19428 24900 19456
rect 28166 19428 28172 19440
rect 24872 19400 25820 19428
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 19794 19320 19800 19372
rect 19852 19320 19858 19372
rect 19978 19320 19984 19372
rect 20036 19320 20042 19372
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 20349 19364 20407 19369
rect 20349 19363 20576 19364
rect 20349 19329 20361 19363
rect 20395 19360 20576 19363
rect 20395 19336 20944 19360
rect 20395 19332 20414 19336
rect 20548 19332 20944 19336
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 19484 19264 19656 19292
rect 19484 19252 19490 19264
rect 19613 19227 19671 19233
rect 19613 19224 19625 19227
rect 18340 19196 19625 19224
rect 18049 19187 18107 19193
rect 19613 19193 19625 19196
rect 19659 19193 19671 19227
rect 19613 19187 19671 19193
rect 17310 19156 17316 19168
rect 16724 19128 17316 19156
rect 16724 19116 16730 19128
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17770 19116 17776 19168
rect 17828 19156 17834 19168
rect 18322 19156 18328 19168
rect 17828 19128 18328 19156
rect 17828 19116 17834 19128
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 18785 19159 18843 19165
rect 18785 19125 18797 19159
rect 18831 19156 18843 19159
rect 19720 19156 19748 19320
rect 19886 19184 19892 19236
rect 19944 19224 19950 19236
rect 20088 19224 20116 19323
rect 20272 19292 20300 19323
rect 20916 19304 20944 19332
rect 21450 19320 21456 19372
rect 21508 19369 21514 19372
rect 21508 19363 21527 19369
rect 21515 19329 21527 19363
rect 21508 19323 21527 19329
rect 21508 19320 21514 19323
rect 22278 19320 22284 19372
rect 22336 19320 22342 19372
rect 25792 19369 25820 19400
rect 27356 19400 28172 19428
rect 25133 19363 25191 19369
rect 20272 19264 20392 19292
rect 19944 19196 20116 19224
rect 20364 19224 20392 19264
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20588 19264 20821 19292
rect 20588 19252 20594 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 20898 19252 20904 19304
rect 20956 19252 20962 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19261 21419 19295
rect 21361 19255 21419 19261
rect 21376 19224 21404 19255
rect 22296 19224 22324 19320
rect 22830 19292 22836 19304
rect 20364 19196 20668 19224
rect 21376 19196 22324 19224
rect 22388 19264 22836 19292
rect 19944 19184 19950 19196
rect 20640 19168 20668 19196
rect 18831 19128 19748 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 20622 19116 20628 19168
rect 20680 19116 20686 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21542 19156 21548 19168
rect 21232 19128 21548 19156
rect 21232 19116 21238 19128
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 21968 19128 22293 19156
rect 21968 19116 21974 19128
rect 22281 19125 22293 19128
rect 22327 19156 22339 19159
rect 22388 19156 22416 19264
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 23106 19252 23112 19304
rect 23164 19252 23170 19304
rect 24228 19292 24256 19346
rect 25133 19329 25145 19363
rect 25179 19360 25191 19363
rect 25777 19363 25835 19369
rect 25179 19332 25728 19360
rect 25179 19329 25191 19332
rect 25133 19323 25191 19329
rect 24394 19292 24400 19304
rect 24228 19264 24400 19292
rect 22327 19128 22416 19156
rect 22327 19125 22339 19128
rect 22281 19119 22339 19125
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 22741 19159 22799 19165
rect 22741 19156 22753 19159
rect 22520 19128 22753 19156
rect 22520 19116 22526 19128
rect 22741 19125 22753 19128
rect 22787 19156 22799 19159
rect 24228 19156 24256 19264
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19261 25283 19295
rect 25225 19255 25283 19261
rect 25130 19184 25136 19236
rect 25188 19224 25194 19236
rect 25240 19224 25268 19255
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 25700 19292 25728 19332
rect 25777 19329 25789 19363
rect 25823 19329 25835 19363
rect 26326 19360 26332 19372
rect 25777 19323 25835 19329
rect 25884 19332 26332 19360
rect 25884 19292 25912 19332
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 27356 19369 27384 19400
rect 28166 19388 28172 19400
rect 28224 19428 28230 19440
rect 28224 19400 29408 19428
rect 28224 19388 28230 19400
rect 27341 19363 27399 19369
rect 27341 19329 27353 19363
rect 27387 19329 27399 19363
rect 27341 19323 27399 19329
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 27525 19363 27583 19369
rect 27525 19360 27537 19363
rect 27488 19332 27537 19360
rect 27488 19320 27494 19332
rect 27525 19329 27537 19332
rect 27571 19329 27583 19363
rect 27525 19323 27583 19329
rect 27614 19320 27620 19372
rect 27672 19320 27678 19372
rect 27709 19363 27767 19369
rect 27709 19329 27721 19363
rect 27755 19329 27767 19363
rect 27709 19323 27767 19329
rect 25700 19264 25912 19292
rect 27724 19292 27752 19323
rect 28074 19320 28080 19372
rect 28132 19320 28138 19372
rect 28534 19320 28540 19372
rect 28592 19320 28598 19372
rect 28721 19363 28779 19369
rect 28721 19329 28733 19363
rect 28767 19360 28779 19363
rect 28902 19360 28908 19372
rect 28767 19332 28908 19360
rect 28767 19329 28779 19332
rect 28721 19323 28779 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29380 19369 29408 19400
rect 29638 19388 29644 19440
rect 29696 19388 29702 19440
rect 29748 19400 30144 19428
rect 29748 19372 29776 19400
rect 29365 19363 29423 19369
rect 29365 19329 29377 19363
rect 29411 19329 29423 19363
rect 29365 19323 29423 19329
rect 28552 19292 28580 19320
rect 27724 19264 28580 19292
rect 29380 19292 29408 19323
rect 29546 19320 29552 19372
rect 29604 19320 29610 19372
rect 29730 19320 29736 19372
rect 29788 19320 29794 19372
rect 30006 19320 30012 19372
rect 30064 19320 30070 19372
rect 29454 19292 29460 19304
rect 29380 19264 29460 19292
rect 29454 19252 29460 19264
rect 29512 19292 29518 19304
rect 30024 19292 30052 19320
rect 29512 19264 30052 19292
rect 30116 19292 30144 19400
rect 30190 19388 30196 19440
rect 30248 19388 30254 19440
rect 30285 19431 30343 19437
rect 30285 19397 30297 19431
rect 30331 19428 30343 19431
rect 30392 19428 30420 19468
rect 30834 19456 30840 19508
rect 30892 19456 30898 19508
rect 31662 19456 31668 19508
rect 31720 19456 31726 19508
rect 31846 19456 31852 19508
rect 31904 19496 31910 19508
rect 32950 19496 32956 19508
rect 31904 19468 32956 19496
rect 31904 19456 31910 19468
rect 32950 19456 32956 19468
rect 33008 19456 33014 19508
rect 33410 19456 33416 19508
rect 33468 19496 33474 19508
rect 33597 19499 33655 19505
rect 33597 19496 33609 19499
rect 33468 19468 33609 19496
rect 33468 19456 33474 19468
rect 33597 19465 33609 19468
rect 33643 19465 33655 19499
rect 33597 19459 33655 19465
rect 34517 19499 34575 19505
rect 34517 19465 34529 19499
rect 34563 19496 34575 19499
rect 34882 19496 34888 19508
rect 34563 19468 34888 19496
rect 34563 19465 34575 19468
rect 34517 19459 34575 19465
rect 30331 19400 30420 19428
rect 30331 19397 30343 19400
rect 30285 19391 30343 19397
rect 30401 19364 30459 19369
rect 30392 19363 30604 19364
rect 30392 19332 30413 19363
rect 30401 19329 30413 19332
rect 30447 19360 30604 19363
rect 30852 19360 30880 19456
rect 32214 19428 32220 19440
rect 31312 19400 32220 19428
rect 31312 19372 31340 19400
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 30447 19336 30880 19360
rect 30447 19329 30459 19336
rect 30401 19323 30459 19329
rect 30576 19332 30880 19336
rect 30576 19292 30604 19332
rect 31294 19320 31300 19372
rect 31352 19320 31358 19372
rect 31386 19320 31392 19372
rect 31444 19360 31450 19372
rect 31481 19363 31539 19369
rect 31481 19360 31493 19363
rect 31444 19332 31493 19360
rect 31444 19320 31450 19332
rect 31481 19329 31493 19332
rect 31527 19329 31539 19363
rect 31481 19323 31539 19329
rect 33226 19320 33232 19372
rect 33284 19320 33290 19372
rect 33612 19360 33640 19459
rect 34882 19456 34888 19468
rect 34940 19456 34946 19508
rect 35710 19456 35716 19508
rect 35768 19456 35774 19508
rect 37274 19496 37280 19508
rect 37200 19468 37280 19496
rect 34606 19388 34612 19440
rect 34664 19388 34670 19440
rect 35728 19428 35756 19456
rect 35728 19400 35940 19428
rect 33965 19363 34023 19369
rect 33965 19360 33977 19363
rect 33612 19332 33977 19360
rect 33965 19329 33977 19332
rect 34011 19329 34023 19363
rect 34624 19360 34652 19388
rect 34885 19363 34943 19369
rect 34885 19360 34897 19363
rect 34624 19332 34897 19360
rect 33965 19323 34023 19329
rect 34885 19329 34897 19332
rect 34931 19329 34943 19363
rect 34885 19323 34943 19329
rect 34977 19363 35035 19369
rect 34977 19329 34989 19363
rect 35023 19360 35035 19363
rect 35713 19363 35771 19369
rect 35713 19360 35725 19363
rect 35023 19332 35725 19360
rect 35023 19329 35035 19332
rect 34977 19323 35035 19329
rect 35636 19329 35725 19332
rect 35759 19329 35771 19363
rect 35636 19323 35771 19329
rect 35636 19306 35756 19323
rect 30116 19264 30604 19292
rect 29512 19252 29518 19264
rect 30834 19252 30840 19304
rect 30892 19292 30898 19304
rect 30929 19295 30987 19301
rect 30929 19292 30941 19295
rect 30892 19264 30941 19292
rect 30892 19252 30898 19264
rect 30929 19261 30941 19264
rect 30975 19261 30987 19295
rect 30929 19255 30987 19261
rect 31021 19295 31079 19301
rect 31021 19261 31033 19295
rect 31067 19261 31079 19295
rect 31021 19255 31079 19261
rect 25188 19196 25268 19224
rect 31036 19224 31064 19255
rect 31110 19252 31116 19304
rect 31168 19252 31174 19304
rect 31205 19295 31263 19301
rect 31205 19261 31217 19295
rect 31251 19292 31263 19295
rect 31251 19264 31754 19292
rect 31251 19261 31263 19264
rect 31205 19255 31263 19261
rect 31570 19224 31576 19236
rect 31036 19196 31576 19224
rect 25188 19184 25194 19196
rect 31570 19184 31576 19196
rect 31628 19184 31634 19236
rect 22787 19128 24256 19156
rect 22787 19125 22799 19128
rect 22741 19119 22799 19125
rect 24762 19116 24768 19168
rect 24820 19116 24826 19168
rect 26145 19159 26203 19165
rect 26145 19125 26157 19159
rect 26191 19156 26203 19159
rect 26418 19156 26424 19168
rect 26191 19128 26424 19156
rect 26191 19125 26203 19128
rect 26145 19119 26203 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 26602 19116 26608 19168
rect 26660 19156 26666 19168
rect 26881 19159 26939 19165
rect 26881 19156 26893 19159
rect 26660 19128 26893 19156
rect 26660 19116 26666 19128
rect 26881 19125 26893 19128
rect 26927 19156 26939 19159
rect 27154 19156 27160 19168
rect 26927 19128 27160 19156
rect 26927 19125 26939 19128
rect 26881 19119 26939 19125
rect 27154 19116 27160 19128
rect 27212 19116 27218 19168
rect 28258 19116 28264 19168
rect 28316 19156 28322 19168
rect 28353 19159 28411 19165
rect 28353 19156 28365 19159
rect 28316 19128 28365 19156
rect 28316 19116 28322 19128
rect 28353 19125 28365 19128
rect 28399 19125 28411 19159
rect 28353 19119 28411 19125
rect 29638 19116 29644 19168
rect 29696 19156 29702 19168
rect 29917 19159 29975 19165
rect 29917 19156 29929 19159
rect 29696 19128 29929 19156
rect 29696 19116 29702 19128
rect 29917 19125 29929 19128
rect 29963 19125 29975 19159
rect 29917 19119 29975 19125
rect 30558 19116 30564 19168
rect 30616 19116 30622 19168
rect 30745 19159 30803 19165
rect 30745 19125 30757 19159
rect 30791 19156 30803 19159
rect 31294 19156 31300 19168
rect 30791 19128 31300 19156
rect 30791 19125 30803 19128
rect 30745 19119 30803 19125
rect 31294 19116 31300 19128
rect 31352 19116 31358 19168
rect 31726 19156 31754 19264
rect 31846 19252 31852 19304
rect 31904 19252 31910 19304
rect 32125 19295 32183 19301
rect 32125 19261 32137 19295
rect 32171 19292 32183 19295
rect 33689 19295 33747 19301
rect 33689 19292 33701 19295
rect 32171 19264 33701 19292
rect 32171 19261 32183 19264
rect 32125 19255 32183 19261
rect 33689 19261 33701 19264
rect 33735 19261 33747 19295
rect 33689 19255 33747 19261
rect 33873 19295 33931 19301
rect 33873 19261 33885 19295
rect 33919 19261 33931 19295
rect 33873 19255 33931 19261
rect 33134 19184 33140 19236
rect 33192 19224 33198 19236
rect 33888 19224 33916 19255
rect 34054 19252 34060 19304
rect 34112 19252 34118 19304
rect 34149 19295 34207 19301
rect 34149 19261 34161 19295
rect 34195 19292 34207 19295
rect 34514 19292 34520 19304
rect 34195 19264 34520 19292
rect 34195 19261 34207 19264
rect 34149 19255 34207 19261
rect 34514 19252 34520 19264
rect 34572 19252 34578 19304
rect 35161 19295 35219 19301
rect 35161 19261 35173 19295
rect 35207 19292 35219 19295
rect 35526 19292 35532 19304
rect 35207 19264 35532 19292
rect 35207 19261 35219 19264
rect 35161 19255 35219 19261
rect 33192 19196 33916 19224
rect 33192 19184 33198 19196
rect 34238 19184 34244 19236
rect 34296 19224 34302 19236
rect 35176 19224 35204 19255
rect 35526 19252 35532 19264
rect 35584 19252 35590 19304
rect 34296 19196 35204 19224
rect 35636 19224 35664 19306
rect 35802 19252 35808 19304
rect 35860 19252 35866 19304
rect 35912 19301 35940 19400
rect 37200 19393 37228 19468
rect 37274 19456 37280 19468
rect 37332 19456 37338 19508
rect 38286 19496 38292 19508
rect 37568 19468 38292 19496
rect 37568 19437 37596 19468
rect 38286 19456 38292 19468
rect 38344 19456 38350 19508
rect 39574 19456 39580 19508
rect 39632 19496 39638 19508
rect 39632 19468 40816 19496
rect 39632 19456 39638 19468
rect 37553 19431 37611 19437
rect 37553 19397 37565 19431
rect 37599 19397 37611 19431
rect 37185 19387 37243 19393
rect 37553 19391 37611 19397
rect 38102 19388 38108 19440
rect 38160 19388 38166 19440
rect 39758 19428 39764 19440
rect 39040 19400 39764 19428
rect 35986 19320 35992 19372
rect 36044 19360 36050 19372
rect 36357 19363 36415 19369
rect 36357 19360 36369 19363
rect 36044 19332 36369 19360
rect 36044 19320 36050 19332
rect 36357 19329 36369 19332
rect 36403 19329 36415 19363
rect 37185 19353 37197 19387
rect 37231 19353 37243 19387
rect 37185 19347 37243 19353
rect 36357 19323 36415 19329
rect 35897 19295 35955 19301
rect 35897 19261 35909 19295
rect 35943 19261 35955 19295
rect 37274 19292 37280 19304
rect 35897 19255 35955 19261
rect 36924 19264 37280 19292
rect 36078 19224 36084 19236
rect 35636 19196 36084 19224
rect 34296 19184 34302 19196
rect 35912 19168 35940 19196
rect 36078 19184 36084 19196
rect 36136 19184 36142 19236
rect 36924 19168 36952 19264
rect 37274 19252 37280 19264
rect 37332 19292 37338 19304
rect 38010 19292 38016 19304
rect 37332 19264 38016 19292
rect 37332 19252 37338 19264
rect 38010 19252 38016 19264
rect 38068 19252 38074 19304
rect 38102 19252 38108 19304
rect 38160 19292 38166 19304
rect 39040 19292 39068 19400
rect 39758 19388 39764 19400
rect 39816 19428 39822 19440
rect 39816 19400 39974 19428
rect 39816 19388 39822 19400
rect 40788 19360 40816 19468
rect 40862 19456 40868 19508
rect 40920 19496 40926 19508
rect 41325 19499 41383 19505
rect 41325 19496 41337 19499
rect 40920 19468 41337 19496
rect 40920 19456 40926 19468
rect 41325 19465 41337 19468
rect 41371 19465 41383 19499
rect 41325 19459 41383 19465
rect 41690 19456 41696 19508
rect 41748 19456 41754 19508
rect 41782 19456 41788 19508
rect 41840 19456 41846 19508
rect 42150 19456 42156 19508
rect 42208 19456 42214 19508
rect 42245 19499 42303 19505
rect 42245 19465 42257 19499
rect 42291 19496 42303 19499
rect 43073 19499 43131 19505
rect 43073 19496 43085 19499
rect 42291 19468 43085 19496
rect 42291 19465 42303 19468
rect 42245 19459 42303 19465
rect 43073 19465 43085 19468
rect 43119 19496 43131 19499
rect 43990 19496 43996 19508
rect 43119 19468 43996 19496
rect 43119 19465 43131 19468
rect 43073 19459 43131 19465
rect 43990 19456 43996 19468
rect 44048 19456 44054 19508
rect 41708 19428 41736 19456
rect 41708 19400 42656 19428
rect 41233 19363 41291 19369
rect 41233 19360 41245 19363
rect 40788 19332 41245 19360
rect 41233 19329 41245 19332
rect 41279 19329 41291 19363
rect 41233 19323 41291 19329
rect 41506 19320 41512 19372
rect 41564 19320 41570 19372
rect 38160 19264 39068 19292
rect 38160 19252 38166 19264
rect 39206 19252 39212 19304
rect 39264 19301 39270 19304
rect 39264 19292 39274 19301
rect 39485 19295 39543 19301
rect 39264 19264 39309 19292
rect 39264 19255 39274 19264
rect 39485 19261 39497 19295
rect 39531 19292 39543 19295
rect 39531 19264 41092 19292
rect 39531 19261 39543 19264
rect 39485 19255 39543 19261
rect 39264 19252 39270 19255
rect 41064 19233 41092 19264
rect 41598 19252 41604 19304
rect 41656 19292 41662 19304
rect 42334 19292 42340 19304
rect 41656 19264 42340 19292
rect 41656 19252 41662 19264
rect 42334 19252 42340 19264
rect 42392 19252 42398 19304
rect 41049 19227 41107 19233
rect 41049 19193 41061 19227
rect 41095 19193 41107 19227
rect 41049 19187 41107 19193
rect 41414 19184 41420 19236
rect 41472 19184 41478 19236
rect 42628 19233 42656 19400
rect 42702 19388 42708 19440
rect 42760 19428 42766 19440
rect 42981 19431 43039 19437
rect 42981 19428 42993 19431
rect 42760 19400 42993 19428
rect 42760 19388 42766 19400
rect 42981 19397 42993 19400
rect 43027 19397 43039 19431
rect 42981 19391 43039 19397
rect 43438 19388 43444 19440
rect 43496 19428 43502 19440
rect 44085 19431 44143 19437
rect 44085 19428 44097 19431
rect 43496 19400 44097 19428
rect 43496 19388 43502 19400
rect 44085 19397 44097 19400
rect 44131 19397 44143 19431
rect 44085 19391 44143 19397
rect 43162 19252 43168 19304
rect 43220 19252 43226 19304
rect 44726 19252 44732 19304
rect 44784 19252 44790 19304
rect 42613 19227 42671 19233
rect 42613 19193 42625 19227
rect 42659 19193 42671 19227
rect 42613 19187 42671 19193
rect 42794 19184 42800 19236
rect 42852 19224 42858 19236
rect 43625 19227 43683 19233
rect 43625 19224 43637 19227
rect 42852 19196 43637 19224
rect 42852 19184 42858 19196
rect 43625 19193 43637 19196
rect 43671 19224 43683 19227
rect 44361 19227 44419 19233
rect 44361 19224 44373 19227
rect 43671 19196 44373 19224
rect 43671 19193 43683 19196
rect 43625 19187 43683 19193
rect 44361 19193 44373 19196
rect 44407 19224 44419 19227
rect 45097 19227 45155 19233
rect 45097 19224 45109 19227
rect 44407 19196 45109 19224
rect 44407 19193 44419 19196
rect 44361 19187 44419 19193
rect 45097 19193 45109 19196
rect 45143 19193 45155 19227
rect 45097 19187 45155 19193
rect 32766 19156 32772 19168
rect 31726 19128 32772 19156
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 35342 19116 35348 19168
rect 35400 19116 35406 19168
rect 35894 19116 35900 19168
rect 35952 19116 35958 19168
rect 36170 19116 36176 19168
rect 36228 19116 36234 19168
rect 36262 19116 36268 19168
rect 36320 19156 36326 19168
rect 36906 19156 36912 19168
rect 36320 19128 36912 19156
rect 36320 19116 36326 19128
rect 36906 19116 36912 19128
rect 36964 19116 36970 19168
rect 37001 19159 37059 19165
rect 37001 19125 37013 19159
rect 37047 19156 37059 19159
rect 37090 19156 37096 19168
rect 37047 19128 37096 19156
rect 37047 19125 37059 19128
rect 37001 19119 37059 19125
rect 37090 19116 37096 19128
rect 37148 19116 37154 19168
rect 39022 19116 39028 19168
rect 39080 19116 39086 19168
rect 40957 19159 41015 19165
rect 40957 19125 40969 19159
rect 41003 19156 41015 19159
rect 41432 19156 41460 19184
rect 41003 19128 41460 19156
rect 41003 19125 41015 19128
rect 40957 19119 41015 19125
rect 460 19066 45540 19088
rect 460 19014 3570 19066
rect 3622 19014 3634 19066
rect 3686 19014 3698 19066
rect 3750 19014 3762 19066
rect 3814 19014 3826 19066
rect 3878 19014 8570 19066
rect 8622 19014 8634 19066
rect 8686 19014 8698 19066
rect 8750 19014 8762 19066
rect 8814 19014 8826 19066
rect 8878 19014 13570 19066
rect 13622 19014 13634 19066
rect 13686 19014 13698 19066
rect 13750 19014 13762 19066
rect 13814 19014 13826 19066
rect 13878 19014 18570 19066
rect 18622 19014 18634 19066
rect 18686 19014 18698 19066
rect 18750 19014 18762 19066
rect 18814 19014 18826 19066
rect 18878 19014 23570 19066
rect 23622 19014 23634 19066
rect 23686 19014 23698 19066
rect 23750 19014 23762 19066
rect 23814 19014 23826 19066
rect 23878 19014 28570 19066
rect 28622 19014 28634 19066
rect 28686 19014 28698 19066
rect 28750 19014 28762 19066
rect 28814 19014 28826 19066
rect 28878 19014 33570 19066
rect 33622 19014 33634 19066
rect 33686 19014 33698 19066
rect 33750 19014 33762 19066
rect 33814 19014 33826 19066
rect 33878 19014 38570 19066
rect 38622 19014 38634 19066
rect 38686 19014 38698 19066
rect 38750 19014 38762 19066
rect 38814 19014 38826 19066
rect 38878 19014 43570 19066
rect 43622 19014 43634 19066
rect 43686 19014 43698 19066
rect 43750 19014 43762 19066
rect 43814 19014 43826 19066
rect 43878 19014 45540 19066
rect 460 18992 45540 19014
rect 5445 18955 5503 18961
rect 5445 18921 5457 18955
rect 5491 18952 5503 18955
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 5491 18924 6469 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 6457 18921 6469 18924
rect 6503 18952 6515 18955
rect 6638 18952 6644 18964
rect 6503 18924 6644 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 7098 18952 7104 18964
rect 6748 18924 7104 18952
rect 5994 18844 6000 18896
rect 6052 18844 6058 18896
rect 4430 18776 4436 18828
rect 4488 18776 4494 18828
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 5442 18748 5448 18760
rect 4571 18720 5448 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18748 5595 18751
rect 5626 18748 5632 18760
rect 5583 18720 5632 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 5626 18708 5632 18720
rect 5684 18708 5690 18760
rect 6748 18757 6776 18924
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 8738 18955 8796 18961
rect 8738 18952 8750 18955
rect 8067 18924 8750 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 8738 18921 8750 18924
rect 8784 18921 8796 18955
rect 8738 18915 8796 18921
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10413 18955 10471 18961
rect 10413 18952 10425 18955
rect 10284 18924 10425 18952
rect 10284 18912 10290 18924
rect 10413 18921 10425 18924
rect 10459 18921 10471 18955
rect 10413 18915 10471 18921
rect 10965 18955 11023 18961
rect 10965 18921 10977 18955
rect 11011 18952 11023 18955
rect 11422 18952 11428 18964
rect 11011 18924 11428 18952
rect 11011 18921 11023 18924
rect 10965 18915 11023 18921
rect 7006 18844 7012 18896
rect 7064 18844 7070 18896
rect 7742 18884 7748 18896
rect 7668 18856 7748 18884
rect 7024 18816 7052 18844
rect 7668 18825 7696 18856
rect 7742 18844 7748 18856
rect 7800 18844 7806 18896
rect 7101 18819 7159 18825
rect 7101 18816 7113 18819
rect 7024 18788 7113 18816
rect 7101 18785 7113 18788
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18785 7711 18819
rect 9122 18816 9128 18828
rect 7653 18779 7711 18785
rect 7760 18788 9128 18816
rect 7760 18757 7788 18788
rect 9122 18776 9128 18788
rect 9180 18816 9186 18828
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 9180 18788 10241 18816
rect 9180 18776 9186 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10980 18816 11008 18915
rect 11422 18912 11428 18924
rect 11480 18952 11486 18964
rect 11882 18952 11888 18964
rect 11480 18924 11888 18952
rect 11480 18912 11486 18924
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 14550 18952 14556 18964
rect 13219 18924 14556 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 14734 18912 14740 18964
rect 14792 18952 14798 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 14792 18924 16681 18952
rect 14792 18912 14798 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 16669 18915 16727 18921
rect 17696 18924 18368 18952
rect 17696 18884 17724 18924
rect 14568 18856 17724 18884
rect 14568 18828 14596 18856
rect 18230 18844 18236 18896
rect 18288 18844 18294 18896
rect 18340 18884 18368 18924
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18472 18924 18613 18952
rect 18472 18912 18478 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 19334 18952 19340 18964
rect 18601 18915 18659 18921
rect 18984 18924 19340 18952
rect 18984 18884 19012 18924
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 20438 18952 20444 18964
rect 19536 18924 20444 18952
rect 19444 18884 19472 18912
rect 18340 18856 19012 18884
rect 19076 18856 19472 18884
rect 13449 18819 13507 18825
rect 13449 18816 13461 18819
rect 10229 18779 10287 18785
rect 10520 18788 11008 18816
rect 13004 18788 13461 18816
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 6549 18751 6607 18757
rect 6549 18748 6561 18751
rect 5767 18720 6561 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 6549 18717 6561 18720
rect 6595 18717 6607 18751
rect 6549 18711 6607 18717
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 6564 18624 6592 18711
rect 7024 18680 7052 18711
rect 8386 18708 8392 18760
rect 8444 18748 8450 18760
rect 8481 18751 8539 18757
rect 8481 18748 8493 18751
rect 8444 18720 8493 18748
rect 8444 18708 8450 18720
rect 8481 18717 8493 18720
rect 8527 18717 8539 18751
rect 10134 18748 10140 18760
rect 9890 18720 10140 18748
rect 8481 18711 8539 18717
rect 7834 18680 7840 18692
rect 7024 18652 7840 18680
rect 7834 18640 7840 18652
rect 7892 18640 7898 18692
rect 4890 18572 4896 18624
rect 4948 18572 4954 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 5629 18615 5687 18621
rect 5629 18612 5641 18615
rect 5592 18584 5641 18612
rect 5592 18572 5598 18584
rect 5629 18581 5641 18584
rect 5675 18581 5687 18615
rect 5629 18575 5687 18581
rect 6546 18572 6552 18624
rect 6604 18572 6610 18624
rect 6733 18615 6791 18621
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 6914 18612 6920 18624
rect 6779 18584 6920 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7374 18572 7380 18624
rect 7432 18572 7438 18624
rect 8496 18612 8524 18711
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10410 18748 10416 18760
rect 10367 18720 10416 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10520 18757 10548 18788
rect 13004 18760 13032 18788
rect 13449 18785 13461 18788
rect 13495 18785 13507 18819
rect 13449 18779 13507 18785
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 14366 18816 14372 18828
rect 13863 18788 14372 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 14550 18776 14556 18828
rect 14608 18776 14614 18828
rect 14826 18776 14832 18828
rect 14884 18816 14890 18828
rect 15194 18816 15200 18828
rect 14884 18788 15200 18816
rect 14884 18776 14890 18788
rect 15194 18776 15200 18788
rect 15252 18816 15258 18828
rect 15562 18816 15568 18828
rect 15252 18788 15568 18816
rect 15252 18776 15258 18788
rect 15562 18776 15568 18788
rect 15620 18816 15626 18828
rect 15620 18788 15700 18816
rect 15620 18776 15626 18788
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 10686 18748 10692 18760
rect 10643 18720 10692 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18748 10839 18751
rect 10870 18748 10876 18760
rect 10827 18720 10876 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18717 11115 18751
rect 11057 18711 11115 18717
rect 11072 18680 11100 18711
rect 12986 18708 12992 18760
rect 13044 18708 13050 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 13127 18720 13584 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 10796 18652 11100 18680
rect 11333 18683 11391 18689
rect 10796 18624 10824 18652
rect 11333 18649 11345 18683
rect 11379 18680 11391 18683
rect 11606 18680 11612 18692
rect 11379 18652 11612 18680
rect 11379 18649 11391 18652
rect 11333 18643 11391 18649
rect 11606 18640 11612 18652
rect 11664 18640 11670 18692
rect 13170 18680 13176 18692
rect 12558 18652 13176 18680
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 8570 18612 8576 18624
rect 8496 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 10778 18572 10784 18624
rect 10836 18572 10842 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 12124 18584 12817 18612
rect 12124 18572 12130 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 13556 18612 13584 18720
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 15344 18720 15393 18748
rect 15344 18708 15350 18720
rect 15381 18717 15393 18720
rect 15427 18717 15439 18751
rect 15672 18748 15700 18788
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 15804 18788 16160 18816
rect 15804 18776 15810 18788
rect 16132 18757 16160 18788
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17000 18788 17618 18816
rect 17000 18776 17006 18788
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18380 18788 19012 18816
rect 18380 18776 18386 18788
rect 15866 18751 15924 18757
rect 15866 18748 15878 18751
rect 15672 18720 15878 18748
rect 15381 18711 15439 18717
rect 15866 18717 15878 18720
rect 15912 18717 15924 18751
rect 15866 18711 15924 18717
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18717 16175 18751
rect 16117 18711 16175 18717
rect 14734 18640 14740 18692
rect 14792 18640 14798 18692
rect 15881 18680 15909 18711
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 16264 18720 16313 18748
rect 16264 18708 16270 18720
rect 16301 18717 16313 18720
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17218 18748 17224 18760
rect 17083 18720 17224 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17494 18748 17500 18760
rect 17451 18720 17500 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17920 18720 17969 18748
rect 17920 18708 17926 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18046 18708 18052 18760
rect 18104 18708 18110 18760
rect 18616 18757 18644 18788
rect 18984 18760 19012 18788
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18785 18751 18843 18757
rect 18785 18717 18797 18751
rect 18831 18717 18843 18751
rect 18785 18711 18843 18717
rect 16393 18683 16451 18689
rect 16393 18680 16405 18683
rect 15881 18652 16405 18680
rect 16393 18649 16405 18652
rect 16439 18649 16451 18683
rect 18064 18680 18092 18708
rect 18800 18680 18828 18711
rect 18966 18708 18972 18760
rect 19024 18708 19030 18760
rect 19076 18757 19104 18856
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19199 18788 19441 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 19536 18757 19564 18924
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 22833 18955 22891 18961
rect 22833 18952 22845 18955
rect 20548 18924 22845 18952
rect 19889 18887 19947 18893
rect 19889 18853 19901 18887
rect 19935 18853 19947 18887
rect 19889 18847 19947 18853
rect 19061 18751 19119 18757
rect 19061 18717 19073 18751
rect 19107 18717 19119 18751
rect 19061 18711 19119 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19904 18748 19932 18847
rect 20162 18844 20168 18896
rect 20220 18884 20226 18896
rect 20548 18884 20576 18924
rect 22833 18921 22845 18924
rect 22879 18921 22891 18955
rect 22833 18915 22891 18921
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 23753 18955 23811 18961
rect 23753 18952 23765 18955
rect 23532 18924 23765 18952
rect 23532 18912 23538 18924
rect 23753 18921 23765 18924
rect 23799 18921 23811 18955
rect 23753 18915 23811 18921
rect 24026 18912 24032 18964
rect 24084 18952 24090 18964
rect 25590 18952 25596 18964
rect 24084 18924 25596 18952
rect 24084 18912 24090 18924
rect 25590 18912 25596 18924
rect 25648 18912 25654 18964
rect 26234 18912 26240 18964
rect 26292 18912 26298 18964
rect 27798 18912 27804 18964
rect 27856 18952 27862 18964
rect 28166 18952 28172 18964
rect 27856 18924 28172 18952
rect 27856 18912 27862 18924
rect 28166 18912 28172 18924
rect 28224 18912 28230 18964
rect 28902 18912 28908 18964
rect 28960 18952 28966 18964
rect 29457 18955 29515 18961
rect 29457 18952 29469 18955
rect 28960 18924 29469 18952
rect 28960 18912 28966 18924
rect 29457 18921 29469 18924
rect 29503 18921 29515 18955
rect 29457 18915 29515 18921
rect 30484 18924 31892 18952
rect 20220 18856 20576 18884
rect 20220 18844 20226 18856
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 21910 18816 21916 18828
rect 20671 18788 21916 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 23477 18819 23535 18825
rect 23477 18785 23489 18819
rect 23523 18816 23535 18819
rect 24026 18816 24032 18828
rect 23523 18788 24032 18816
rect 23523 18785 23535 18788
rect 23477 18779 23535 18785
rect 24026 18776 24032 18788
rect 24084 18816 24090 18828
rect 24302 18816 24308 18828
rect 24084 18788 24308 18816
rect 24084 18776 24090 18788
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 26252 18816 26280 18912
rect 27982 18844 27988 18896
rect 28040 18884 28046 18896
rect 28629 18887 28687 18893
rect 28629 18884 28641 18887
rect 28040 18856 28641 18884
rect 28040 18844 28046 18856
rect 28629 18853 28641 18856
rect 28675 18853 28687 18887
rect 28629 18847 28687 18853
rect 29178 18844 29184 18896
rect 29236 18884 29242 18896
rect 30484 18884 30512 18924
rect 31864 18896 31892 18924
rect 31938 18912 31944 18964
rect 31996 18952 32002 18964
rect 32217 18955 32275 18961
rect 32217 18952 32229 18955
rect 31996 18924 32229 18952
rect 31996 18912 32002 18924
rect 32217 18921 32229 18924
rect 32263 18921 32275 18955
rect 33134 18952 33140 18964
rect 32217 18915 32275 18921
rect 32508 18924 33140 18952
rect 29236 18856 30512 18884
rect 29236 18844 29242 18856
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 24596 18788 26096 18816
rect 26252 18788 26709 18816
rect 19981 18751 20039 18757
rect 19981 18748 19993 18751
rect 19904 18720 19993 18748
rect 19521 18711 19579 18717
rect 19981 18717 19993 18720
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 18064 18652 18828 18680
rect 19260 18680 19288 18711
rect 20254 18708 20260 18760
rect 20312 18708 20318 18760
rect 20346 18708 20352 18760
rect 20404 18708 20410 18760
rect 20548 18720 20660 18748
rect 19886 18680 19892 18692
rect 19260 18652 19892 18680
rect 16393 18643 16451 18649
rect 19886 18640 19892 18652
rect 19944 18640 19950 18692
rect 20162 18640 20168 18692
rect 20220 18640 20226 18692
rect 15010 18612 15016 18624
rect 13556 18584 15016 18612
rect 12805 18575 12863 18581
rect 15010 18572 15016 18584
rect 15068 18612 15074 18624
rect 15243 18615 15301 18621
rect 15243 18612 15255 18615
rect 15068 18584 15255 18612
rect 15068 18572 15074 18584
rect 15243 18581 15255 18584
rect 15289 18581 15301 18615
rect 15243 18575 15301 18581
rect 15654 18572 15660 18624
rect 15712 18572 15718 18624
rect 16022 18572 16028 18624
rect 16080 18572 16086 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 17402 18612 17408 18624
rect 16816 18584 17408 18612
rect 16816 18572 16822 18584
rect 17402 18572 17408 18584
rect 17460 18612 17466 18624
rect 17954 18612 17960 18624
rect 17460 18584 17960 18612
rect 17460 18572 17466 18584
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 20548 18621 20576 18720
rect 20632 18680 20660 18720
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 24118 18708 24124 18760
rect 24176 18748 24182 18760
rect 24486 18748 24492 18760
rect 24176 18720 24492 18748
rect 24176 18708 24182 18720
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 24596 18757 24624 18788
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 25958 18708 25964 18760
rect 26016 18708 26022 18760
rect 26068 18748 26096 18788
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 30009 18819 30067 18825
rect 30009 18816 30021 18819
rect 26697 18779 26755 18785
rect 28276 18788 30021 18816
rect 28276 18760 28304 18788
rect 30009 18785 30021 18788
rect 30055 18816 30067 18819
rect 30374 18816 30380 18828
rect 30055 18788 30380 18816
rect 30055 18785 30067 18788
rect 30009 18779 30067 18785
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 30484 18825 30512 18856
rect 31846 18844 31852 18896
rect 31904 18884 31910 18896
rect 32030 18884 32036 18896
rect 31904 18856 32036 18884
rect 31904 18844 31910 18856
rect 32030 18844 32036 18856
rect 32088 18844 32094 18896
rect 30469 18819 30527 18825
rect 30469 18785 30481 18819
rect 30515 18785 30527 18819
rect 30469 18779 30527 18785
rect 30834 18776 30840 18828
rect 30892 18816 30898 18828
rect 31754 18816 31760 18828
rect 30892 18788 31760 18816
rect 30892 18776 30898 18788
rect 31754 18776 31760 18788
rect 31812 18816 31818 18828
rect 32508 18825 32536 18924
rect 33134 18912 33140 18924
rect 33192 18912 33198 18964
rect 36170 18912 36176 18964
rect 36228 18912 36234 18964
rect 38105 18955 38163 18961
rect 38105 18921 38117 18955
rect 38151 18952 38163 18955
rect 38470 18952 38476 18964
rect 38151 18924 38476 18952
rect 38151 18921 38163 18924
rect 38105 18915 38163 18921
rect 38470 18912 38476 18924
rect 38528 18912 38534 18964
rect 39942 18912 39948 18964
rect 40000 18952 40006 18964
rect 40954 18952 40960 18964
rect 40000 18924 40960 18952
rect 40000 18912 40006 18924
rect 40954 18912 40960 18924
rect 41012 18912 41018 18964
rect 41049 18955 41107 18961
rect 41049 18921 41061 18955
rect 41095 18952 41107 18955
rect 41506 18952 41512 18964
rect 41095 18924 41512 18952
rect 41095 18921 41107 18924
rect 41049 18915 41107 18921
rect 41506 18912 41512 18924
rect 41564 18912 41570 18964
rect 41598 18912 41604 18964
rect 41656 18912 41662 18964
rect 32953 18887 33011 18893
rect 32953 18853 32965 18887
rect 32999 18884 33011 18887
rect 32999 18856 33640 18884
rect 32999 18853 33011 18856
rect 32953 18847 33011 18853
rect 32493 18819 32551 18825
rect 32493 18816 32505 18819
rect 31812 18788 32505 18816
rect 31812 18776 31818 18788
rect 32493 18785 32505 18788
rect 32539 18785 32551 18819
rect 32493 18779 32551 18785
rect 32585 18819 32643 18825
rect 32585 18785 32597 18819
rect 32631 18816 32643 18819
rect 33410 18816 33416 18828
rect 32631 18788 33416 18816
rect 32631 18785 32643 18788
rect 32585 18779 32643 18785
rect 33410 18776 33416 18788
rect 33468 18776 33474 18828
rect 33502 18776 33508 18828
rect 33560 18776 33566 18828
rect 26418 18748 26424 18760
rect 26068 18720 26424 18748
rect 26418 18708 26424 18720
rect 26476 18708 26482 18760
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 28442 18708 28448 18760
rect 28500 18708 28506 18760
rect 29822 18708 29828 18760
rect 29880 18708 29886 18760
rect 29914 18708 29920 18760
rect 29972 18708 29978 18760
rect 32398 18748 32404 18760
rect 31878 18720 32404 18748
rect 32398 18708 32404 18720
rect 32456 18708 32462 18760
rect 32677 18751 32735 18757
rect 32677 18717 32689 18751
rect 32723 18717 32735 18751
rect 32677 18711 32735 18717
rect 32769 18751 32827 18757
rect 32769 18717 32781 18751
rect 32815 18748 32827 18751
rect 32858 18748 32864 18760
rect 32815 18720 32864 18748
rect 32815 18717 32827 18720
rect 32769 18711 32827 18717
rect 20901 18683 20959 18689
rect 20901 18680 20913 18683
rect 20632 18652 20913 18680
rect 20901 18649 20913 18652
rect 20947 18649 20959 18683
rect 22462 18680 22468 18692
rect 22126 18652 22468 18680
rect 20901 18643 20959 18649
rect 22462 18640 22468 18652
rect 22520 18640 22526 18692
rect 23293 18683 23351 18689
rect 23293 18649 23305 18683
rect 23339 18680 23351 18683
rect 23339 18652 24624 18680
rect 23339 18649 23351 18652
rect 23293 18643 23351 18649
rect 20533 18615 20591 18621
rect 20533 18581 20545 18615
rect 20579 18581 20591 18615
rect 20533 18575 20591 18581
rect 21542 18572 21548 18624
rect 21600 18612 21606 18624
rect 22373 18615 22431 18621
rect 22373 18612 22385 18615
rect 21600 18584 22385 18612
rect 21600 18572 21606 18584
rect 22373 18581 22385 18584
rect 22419 18581 22431 18615
rect 22373 18575 22431 18581
rect 22554 18572 22560 18624
rect 22612 18572 22618 18624
rect 23198 18572 23204 18624
rect 23256 18572 23262 18624
rect 24213 18615 24271 18621
rect 24213 18581 24225 18615
rect 24259 18612 24271 18615
rect 24302 18612 24308 18624
rect 24259 18584 24308 18612
rect 24259 18581 24271 18584
rect 24213 18575 24271 18581
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 24596 18612 24624 18652
rect 24854 18640 24860 18692
rect 24912 18640 24918 18692
rect 26436 18680 26464 18708
rect 26786 18680 26792 18692
rect 26436 18652 26792 18680
rect 26786 18640 26792 18652
rect 26844 18640 26850 18692
rect 27154 18640 27160 18692
rect 27212 18640 27218 18692
rect 30742 18640 30748 18692
rect 30800 18640 30806 18692
rect 32490 18640 32496 18692
rect 32548 18680 32554 18692
rect 32692 18680 32720 18711
rect 32858 18708 32864 18720
rect 32916 18708 32922 18760
rect 33612 18748 33640 18856
rect 34698 18776 34704 18828
rect 34756 18776 34762 18828
rect 36188 18816 36216 18912
rect 41616 18884 41644 18912
rect 38672 18856 39344 18884
rect 36541 18819 36599 18825
rect 36541 18816 36553 18819
rect 36188 18788 36553 18816
rect 36541 18785 36553 18788
rect 36587 18785 36599 18819
rect 36541 18779 36599 18785
rect 36998 18776 37004 18828
rect 37056 18816 37062 18828
rect 37274 18816 37280 18828
rect 37056 18788 37280 18816
rect 37056 18776 37062 18788
rect 37274 18776 37280 18788
rect 37332 18776 37338 18828
rect 37550 18776 37556 18828
rect 37608 18816 37614 18828
rect 38378 18816 38384 18828
rect 37608 18788 38384 18816
rect 37608 18776 37614 18788
rect 38378 18776 38384 18788
rect 38436 18816 38442 18828
rect 38672 18825 38700 18856
rect 38657 18819 38715 18825
rect 38657 18816 38669 18819
rect 38436 18788 38669 18816
rect 38436 18776 38442 18788
rect 38657 18785 38669 18788
rect 38703 18785 38715 18819
rect 38657 18779 38715 18785
rect 39022 18776 39028 18828
rect 39080 18776 39086 18828
rect 39206 18776 39212 18828
rect 39264 18776 39270 18828
rect 39316 18816 39344 18856
rect 40512 18856 42472 18884
rect 40512 18816 40540 18856
rect 39316 18788 40540 18816
rect 40954 18776 40960 18828
rect 41012 18816 41018 18828
rect 41601 18819 41659 18825
rect 41601 18816 41613 18819
rect 41012 18788 41613 18816
rect 41012 18776 41018 18788
rect 41601 18785 41613 18788
rect 41647 18785 41659 18819
rect 42150 18816 42156 18828
rect 41601 18779 41659 18785
rect 41800 18788 42156 18816
rect 34057 18751 34115 18757
rect 34057 18748 34069 18751
rect 33612 18720 34069 18748
rect 34057 18717 34069 18720
rect 34103 18717 34115 18751
rect 34057 18711 34115 18717
rect 34425 18751 34483 18757
rect 34425 18717 34437 18751
rect 34471 18717 34483 18751
rect 34425 18711 34483 18717
rect 33321 18683 33379 18689
rect 32548 18652 32812 18680
rect 32548 18640 32554 18652
rect 25130 18612 25136 18624
rect 24596 18584 25136 18612
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 28350 18612 28356 18624
rect 26384 18584 28356 18612
rect 26384 18572 26390 18584
rect 28350 18572 28356 18584
rect 28408 18572 28414 18624
rect 31110 18572 31116 18624
rect 31168 18612 31174 18624
rect 32122 18612 32128 18624
rect 31168 18584 32128 18612
rect 31168 18572 31174 18584
rect 32122 18572 32128 18584
rect 32180 18572 32186 18624
rect 32306 18572 32312 18624
rect 32364 18572 32370 18624
rect 32784 18612 32812 18652
rect 33321 18649 33333 18683
rect 33367 18680 33379 18683
rect 34146 18680 34152 18692
rect 33367 18652 34152 18680
rect 33367 18649 33379 18652
rect 33321 18643 33379 18649
rect 34146 18640 34152 18652
rect 34204 18640 34210 18692
rect 34440 18680 34468 18711
rect 36262 18708 36268 18760
rect 36320 18708 36326 18760
rect 37918 18708 37924 18760
rect 37976 18748 37982 18760
rect 38470 18748 38476 18760
rect 37976 18720 38476 18748
rect 37976 18708 37982 18720
rect 38470 18708 38476 18720
rect 38528 18708 38534 18760
rect 38565 18751 38623 18757
rect 38565 18717 38577 18751
rect 38611 18748 38623 18751
rect 39040 18748 39068 18776
rect 38611 18720 39068 18748
rect 38611 18717 38623 18720
rect 38565 18711 38623 18717
rect 36998 18680 37004 18692
rect 34440 18652 34652 18680
rect 34624 18624 34652 18652
rect 34900 18652 35190 18680
rect 36004 18652 37004 18680
rect 34900 18624 34928 18652
rect 34054 18612 34060 18624
rect 32784 18584 34060 18612
rect 34054 18572 34060 18584
rect 34112 18572 34118 18624
rect 34238 18572 34244 18624
rect 34296 18572 34302 18624
rect 34606 18572 34612 18624
rect 34664 18572 34670 18624
rect 34882 18572 34888 18624
rect 34940 18612 34946 18624
rect 36004 18612 36032 18652
rect 36998 18640 37004 18652
rect 37056 18640 37062 18692
rect 38102 18640 38108 18692
rect 38160 18680 38166 18692
rect 39224 18680 39252 18776
rect 41414 18708 41420 18760
rect 41472 18708 41478 18760
rect 41506 18708 41512 18760
rect 41564 18748 41570 18760
rect 41800 18748 41828 18788
rect 42150 18776 42156 18788
rect 42208 18776 42214 18828
rect 42444 18825 42472 18856
rect 42429 18819 42487 18825
rect 42429 18785 42441 18819
rect 42475 18785 42487 18819
rect 42429 18779 42487 18785
rect 42889 18751 42947 18757
rect 42889 18748 42901 18751
rect 41564 18720 41828 18748
rect 41892 18720 42901 18748
rect 41564 18708 41570 18720
rect 38160 18652 39252 18680
rect 38160 18640 38166 18652
rect 34940 18584 36032 18612
rect 34940 18572 34946 18584
rect 36078 18572 36084 18624
rect 36136 18612 36142 18624
rect 36173 18615 36231 18621
rect 36173 18612 36185 18615
rect 36136 18584 36185 18612
rect 36136 18572 36142 18584
rect 36173 18581 36185 18584
rect 36219 18581 36231 18615
rect 36173 18575 36231 18581
rect 36446 18572 36452 18624
rect 36504 18612 36510 18624
rect 36814 18612 36820 18624
rect 36504 18584 36820 18612
rect 36504 18572 36510 18584
rect 36814 18572 36820 18584
rect 36872 18612 36878 18624
rect 38013 18615 38071 18621
rect 38013 18612 38025 18615
rect 36872 18584 38025 18612
rect 36872 18572 36878 18584
rect 38013 18581 38025 18584
rect 38059 18581 38071 18615
rect 39224 18612 39252 18652
rect 39482 18640 39488 18692
rect 39540 18640 39546 18692
rect 39758 18640 39764 18692
rect 39816 18680 39822 18692
rect 39816 18652 39974 18680
rect 39816 18640 39822 18652
rect 41690 18612 41696 18624
rect 39224 18584 41696 18612
rect 38013 18575 38071 18581
rect 41690 18572 41696 18584
rect 41748 18572 41754 18624
rect 41892 18621 41920 18720
rect 42889 18717 42901 18720
rect 42935 18717 42947 18751
rect 42889 18711 42947 18717
rect 42337 18683 42395 18689
rect 42337 18649 42349 18683
rect 42383 18680 42395 18683
rect 42978 18680 42984 18692
rect 42383 18652 42984 18680
rect 42383 18649 42395 18652
rect 42337 18643 42395 18649
rect 42978 18640 42984 18652
rect 43036 18640 43042 18692
rect 41877 18615 41935 18621
rect 41877 18581 41889 18615
rect 41923 18581 41935 18615
rect 41877 18575 41935 18581
rect 42242 18572 42248 18624
rect 42300 18572 42306 18624
rect 42702 18572 42708 18624
rect 42760 18572 42766 18624
rect 43257 18615 43315 18621
rect 43257 18581 43269 18615
rect 43303 18612 43315 18615
rect 43533 18615 43591 18621
rect 43533 18612 43545 18615
rect 43303 18584 43545 18612
rect 43303 18581 43315 18584
rect 43257 18575 43315 18581
rect 43533 18581 43545 18584
rect 43579 18612 43591 18615
rect 43714 18612 43720 18624
rect 43579 18584 43720 18612
rect 43579 18581 43591 18584
rect 43533 18575 43591 18581
rect 43714 18572 43720 18584
rect 43772 18572 43778 18624
rect 43806 18572 43812 18624
rect 43864 18612 43870 18624
rect 43901 18615 43959 18621
rect 43901 18612 43913 18615
rect 43864 18584 43913 18612
rect 43864 18572 43870 18584
rect 43901 18581 43913 18584
rect 43947 18612 43959 18615
rect 44545 18615 44603 18621
rect 44545 18612 44557 18615
rect 43947 18584 44557 18612
rect 43947 18581 43959 18584
rect 43901 18575 43959 18581
rect 44545 18581 44557 18584
rect 44591 18581 44603 18615
rect 44545 18575 44603 18581
rect 44818 18572 44824 18624
rect 44876 18612 44882 18624
rect 44913 18615 44971 18621
rect 44913 18612 44925 18615
rect 44876 18584 44925 18612
rect 44876 18572 44882 18584
rect 44913 18581 44925 18584
rect 44959 18581 44971 18615
rect 44913 18575 44971 18581
rect 460 18522 45540 18544
rect 460 18470 6070 18522
rect 6122 18470 6134 18522
rect 6186 18470 6198 18522
rect 6250 18470 6262 18522
rect 6314 18470 6326 18522
rect 6378 18470 11070 18522
rect 11122 18470 11134 18522
rect 11186 18470 11198 18522
rect 11250 18470 11262 18522
rect 11314 18470 11326 18522
rect 11378 18470 16070 18522
rect 16122 18470 16134 18522
rect 16186 18470 16198 18522
rect 16250 18470 16262 18522
rect 16314 18470 16326 18522
rect 16378 18470 21070 18522
rect 21122 18470 21134 18522
rect 21186 18470 21198 18522
rect 21250 18470 21262 18522
rect 21314 18470 21326 18522
rect 21378 18470 26070 18522
rect 26122 18470 26134 18522
rect 26186 18470 26198 18522
rect 26250 18470 26262 18522
rect 26314 18470 26326 18522
rect 26378 18470 31070 18522
rect 31122 18470 31134 18522
rect 31186 18470 31198 18522
rect 31250 18470 31262 18522
rect 31314 18470 31326 18522
rect 31378 18470 36070 18522
rect 36122 18470 36134 18522
rect 36186 18470 36198 18522
rect 36250 18470 36262 18522
rect 36314 18470 36326 18522
rect 36378 18470 41070 18522
rect 41122 18470 41134 18522
rect 41186 18470 41198 18522
rect 41250 18470 41262 18522
rect 41314 18470 41326 18522
rect 41378 18470 45540 18522
rect 460 18448 45540 18470
rect 4890 18408 4896 18420
rect 4080 18380 4896 18408
rect 4080 18349 4108 18380
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 5500 18380 5549 18408
rect 5500 18368 5506 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 5537 18371 5595 18377
rect 4065 18343 4123 18349
rect 4065 18309 4077 18343
rect 4111 18309 4123 18343
rect 4065 18303 4123 18309
rect 4614 18300 4620 18352
rect 4672 18300 4678 18352
rect 3786 18232 3792 18284
rect 3844 18232 3850 18284
rect 5552 18068 5580 18371
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 6089 18411 6147 18417
rect 6089 18408 6101 18411
rect 5684 18380 6101 18408
rect 5684 18368 5690 18380
rect 6089 18377 6101 18380
rect 6135 18377 6147 18411
rect 7374 18408 7380 18420
rect 6089 18371 6147 18377
rect 7024 18380 7380 18408
rect 7024 18349 7052 18380
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 7834 18368 7840 18420
rect 7892 18408 7898 18420
rect 8386 18408 8392 18420
rect 7892 18380 8392 18408
rect 7892 18368 7898 18380
rect 8386 18368 8392 18380
rect 8444 18408 8450 18420
rect 8481 18411 8539 18417
rect 8481 18408 8493 18411
rect 8444 18380 8493 18408
rect 8444 18368 8450 18380
rect 8481 18377 8493 18380
rect 8527 18377 8539 18411
rect 8481 18371 8539 18377
rect 11606 18368 11612 18420
rect 11664 18408 11670 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 11664 18380 12449 18408
rect 11664 18368 11670 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 12986 18368 12992 18420
rect 13044 18368 13050 18420
rect 13541 18411 13599 18417
rect 13541 18377 13553 18411
rect 13587 18408 13599 18411
rect 13587 18380 13952 18408
rect 13587 18377 13599 18380
rect 13541 18371 13599 18377
rect 6273 18343 6331 18349
rect 6273 18309 6285 18343
rect 6319 18340 6331 18343
rect 7009 18343 7067 18349
rect 6319 18312 6592 18340
rect 6319 18309 6331 18312
rect 6273 18303 6331 18309
rect 6564 18284 6592 18312
rect 7009 18309 7021 18343
rect 7055 18309 7067 18343
rect 7009 18303 7067 18309
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 8849 18343 8907 18349
rect 8849 18340 8861 18343
rect 8352 18312 8861 18340
rect 8352 18300 8358 18312
rect 8849 18309 8861 18312
rect 8895 18309 8907 18343
rect 10134 18340 10140 18352
rect 10074 18312 10140 18340
rect 8849 18303 8907 18309
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 11793 18343 11851 18349
rect 11793 18309 11805 18343
rect 11839 18340 11851 18343
rect 13004 18340 13032 18368
rect 11839 18312 12388 18340
rect 13004 18312 13860 18340
rect 11839 18309 11851 18312
rect 11793 18303 11851 18309
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5684 18244 5733 18272
rect 5684 18232 5690 18244
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18241 6515 18275
rect 6457 18235 6515 18241
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6196 18204 6224 18235
rect 5868 18176 6224 18204
rect 5868 18164 5874 18176
rect 6472 18136 6500 18235
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 8110 18232 8116 18284
rect 8168 18232 8174 18284
rect 8570 18232 8576 18284
rect 8628 18232 8634 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 7098 18204 7104 18216
rect 6840 18176 7104 18204
rect 6840 18136 6868 18176
rect 7098 18164 7104 18176
rect 7156 18204 7162 18216
rect 8588 18204 8616 18232
rect 10597 18207 10655 18213
rect 10597 18204 10609 18207
rect 7156 18176 8156 18204
rect 8588 18176 10609 18204
rect 7156 18164 7162 18176
rect 6472 18108 6868 18136
rect 8128 18080 8156 18176
rect 10597 18173 10609 18176
rect 10643 18204 10655 18207
rect 10778 18204 10784 18216
rect 10643 18176 10784 18204
rect 10643 18173 10655 18176
rect 10597 18167 10655 18173
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 11532 18204 11560 18235
rect 11882 18232 11888 18284
rect 11940 18232 11946 18284
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12069 18275 12127 18281
rect 12069 18272 12081 18275
rect 12032 18244 12081 18272
rect 12032 18232 12038 18244
rect 12069 18241 12081 18244
rect 12115 18272 12127 18275
rect 12158 18272 12164 18284
rect 12115 18244 12164 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12360 18281 12388 18312
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 13354 18232 13360 18284
rect 13412 18272 13418 18284
rect 13832 18281 13860 18312
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13412 18244 13737 18272
rect 13412 18232 13418 18244
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18241 13875 18275
rect 13924 18272 13952 18380
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 15896 18380 16436 18408
rect 15896 18368 15902 18380
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 13924 18244 14197 18272
rect 13817 18235 13875 18241
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 11606 18204 11612 18216
rect 11532 18176 11612 18204
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18173 11851 18207
rect 12544 18204 12572 18232
rect 11793 18167 11851 18173
rect 12268 18176 12572 18204
rect 5718 18068 5724 18080
rect 5552 18040 5724 18068
rect 5718 18028 5724 18040
rect 5776 18068 5782 18080
rect 5859 18071 5917 18077
rect 5859 18068 5871 18071
rect 5776 18040 5871 18068
rect 5776 18028 5782 18040
rect 5859 18037 5871 18040
rect 5905 18037 5917 18071
rect 5859 18031 5917 18037
rect 5994 18028 6000 18080
rect 6052 18028 6058 18080
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 7006 18068 7012 18080
rect 6687 18040 7012 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 8110 18028 8116 18080
rect 8168 18028 8174 18080
rect 9950 18028 9956 18080
rect 10008 18068 10014 18080
rect 10321 18071 10379 18077
rect 10321 18068 10333 18071
rect 10008 18040 10333 18068
rect 10008 18028 10014 18040
rect 10321 18037 10333 18040
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 11330 18028 11336 18080
rect 11388 18028 11394 18080
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 11609 18071 11667 18077
rect 11609 18068 11621 18071
rect 11572 18040 11621 18068
rect 11572 18028 11578 18040
rect 11609 18037 11621 18040
rect 11655 18037 11667 18071
rect 11808 18068 11836 18167
rect 12268 18145 12296 18176
rect 12253 18139 12311 18145
rect 12253 18105 12265 18139
rect 12299 18105 12311 18139
rect 12253 18099 12311 18105
rect 12066 18068 12072 18080
rect 11808 18040 12072 18068
rect 11609 18031 11667 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 13170 18028 13176 18080
rect 13228 18068 13234 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 13228 18040 13461 18068
rect 13228 18028 13234 18040
rect 13449 18037 13461 18040
rect 13495 18068 13507 18071
rect 14734 18068 14740 18080
rect 13495 18040 14740 18068
rect 13495 18037 13507 18040
rect 13449 18031 13507 18037
rect 14734 18028 14740 18040
rect 14792 18068 14798 18080
rect 14936 18068 14964 18326
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 16209 18343 16267 18349
rect 16209 18340 16221 18343
rect 15988 18312 16221 18340
rect 15988 18300 15994 18312
rect 16209 18309 16221 18312
rect 16255 18309 16267 18343
rect 16408 18340 16436 18380
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 17687 18411 17745 18417
rect 17687 18408 17699 18411
rect 16540 18380 17699 18408
rect 16540 18368 16546 18380
rect 17687 18377 17699 18380
rect 17733 18377 17745 18411
rect 17687 18371 17745 18377
rect 17773 18411 17831 18417
rect 17773 18377 17785 18411
rect 17819 18408 17831 18411
rect 17954 18408 17960 18420
rect 17819 18380 17960 18408
rect 17819 18377 17831 18380
rect 17773 18371 17831 18377
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 19886 18408 19892 18420
rect 19668 18380 19892 18408
rect 19668 18368 19674 18380
rect 19886 18368 19892 18380
rect 19944 18408 19950 18420
rect 20162 18408 20168 18420
rect 19944 18380 20168 18408
rect 19944 18368 19950 18380
rect 20162 18368 20168 18380
rect 20220 18408 20226 18420
rect 20220 18380 20484 18408
rect 20220 18368 20226 18380
rect 16574 18340 16580 18352
rect 16408 18312 16580 18340
rect 16209 18303 16267 18309
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 16666 18300 16672 18352
rect 16724 18300 16730 18352
rect 16758 18300 16764 18352
rect 16816 18300 16822 18352
rect 17126 18340 17132 18352
rect 16914 18312 17132 18340
rect 16668 18297 16726 18300
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 16025 18275 16083 18281
rect 16025 18272 16037 18275
rect 15068 18244 16037 18272
rect 15068 18232 15074 18244
rect 16025 18241 16037 18244
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16298 18232 16304 18284
rect 16356 18232 16362 18284
rect 16393 18275 16451 18281
rect 16393 18241 16405 18275
rect 16439 18272 16451 18275
rect 16482 18272 16488 18284
rect 16439 18244 16488 18272
rect 16439 18241 16451 18244
rect 16393 18235 16451 18241
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16408 18204 16436 18235
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16668 18263 16680 18297
rect 16714 18263 16726 18297
rect 16914 18281 16942 18312
rect 17126 18300 17132 18312
rect 17184 18300 17190 18352
rect 17310 18300 17316 18352
rect 17368 18349 17374 18352
rect 17368 18343 17387 18349
rect 17375 18340 17387 18343
rect 17375 18312 17908 18340
rect 17375 18309 17387 18312
rect 17368 18303 17387 18309
rect 17368 18300 17374 18303
rect 16668 18257 16726 18263
rect 16895 18275 16953 18281
rect 16895 18241 16907 18275
rect 16941 18241 16953 18275
rect 16895 18235 16953 18241
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18272 17095 18275
rect 17494 18272 17500 18284
rect 17083 18244 17500 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 17494 18232 17500 18244
rect 17552 18272 17558 18284
rect 17589 18275 17647 18281
rect 17589 18272 17601 18275
rect 17552 18244 17601 18272
rect 17552 18232 17558 18244
rect 17589 18241 17601 18244
rect 17635 18241 17647 18275
rect 17589 18235 17647 18241
rect 17678 18232 17684 18284
rect 17736 18272 17742 18284
rect 17880 18281 17908 18312
rect 19334 18300 19340 18352
rect 19392 18300 19398 18352
rect 20456 18340 20484 18380
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 20680 18380 21833 18408
rect 20680 18368 20686 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 21821 18371 21879 18377
rect 22462 18368 22468 18420
rect 22520 18368 22526 18420
rect 22554 18368 22560 18420
rect 22612 18368 22618 18420
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 22796 18380 24685 18408
rect 22796 18368 22802 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 24762 18368 24768 18420
rect 24820 18368 24826 18420
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25501 18411 25559 18417
rect 25501 18408 25513 18411
rect 24912 18380 25513 18408
rect 24912 18368 24918 18380
rect 25501 18377 25513 18380
rect 25547 18377 25559 18411
rect 25501 18371 25559 18377
rect 25682 18368 25688 18420
rect 25740 18408 25746 18420
rect 28261 18411 28319 18417
rect 28261 18408 28273 18411
rect 25740 18380 28273 18408
rect 25740 18368 25746 18380
rect 28261 18377 28273 18380
rect 28307 18377 28319 18411
rect 28261 18371 28319 18377
rect 29178 18368 29184 18420
rect 29236 18368 29242 18420
rect 30190 18408 30196 18420
rect 29288 18380 30196 18408
rect 20533 18343 20591 18349
rect 20533 18340 20545 18343
rect 20456 18312 20545 18340
rect 20533 18309 20545 18312
rect 20579 18309 20591 18343
rect 20533 18303 20591 18309
rect 20990 18300 20996 18352
rect 21048 18340 21054 18352
rect 21269 18343 21327 18349
rect 21269 18340 21281 18343
rect 21048 18312 21281 18340
rect 21048 18300 21054 18312
rect 21269 18309 21281 18312
rect 21315 18309 21327 18343
rect 21269 18303 21327 18309
rect 21542 18300 21548 18352
rect 21600 18340 21606 18352
rect 22572 18340 22600 18368
rect 23109 18343 23167 18349
rect 23109 18340 23121 18343
rect 21600 18312 21956 18340
rect 22572 18312 23121 18340
rect 21600 18300 21606 18312
rect 17865 18275 17923 18281
rect 17865 18272 17877 18275
rect 17736 18244 17877 18272
rect 17736 18232 17742 18244
rect 17865 18241 17877 18244
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 17954 18232 17960 18284
rect 18012 18232 18018 18284
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18241 18199 18275
rect 18141 18235 18199 18241
rect 18156 18204 18184 18235
rect 20254 18232 20260 18284
rect 20312 18232 20318 18284
rect 20346 18232 20352 18284
rect 20404 18232 20410 18284
rect 20438 18232 20444 18284
rect 20496 18232 20502 18284
rect 20651 18275 20709 18281
rect 20651 18241 20663 18275
rect 20697 18241 20709 18275
rect 20651 18235 20709 18241
rect 15896 18176 16436 18204
rect 16960 18196 18184 18204
rect 16776 18176 18184 18196
rect 18325 18207 18383 18213
rect 15896 18164 15902 18176
rect 16776 18168 16988 18176
rect 18325 18173 18337 18207
rect 18371 18173 18383 18207
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 16577 18139 16635 18145
rect 16577 18136 16589 18139
rect 15160 18108 16589 18136
rect 15160 18096 15166 18108
rect 16577 18105 16589 18108
rect 16623 18105 16635 18139
rect 16577 18099 16635 18105
rect 14792 18040 14964 18068
rect 15611 18071 15669 18077
rect 14792 18028 14798 18040
rect 15611 18037 15623 18071
rect 15657 18068 15669 18071
rect 16022 18068 16028 18080
rect 15657 18040 16028 18068
rect 15657 18037 15669 18040
rect 15611 18031 15669 18037
rect 16022 18028 16028 18040
rect 16080 18068 16086 18080
rect 16776 18068 16804 18168
rect 18325 18167 18383 18173
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18204 18659 18207
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 18647 18176 20177 18204
rect 18647 18173 18659 18176
rect 18601 18167 18659 18173
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20272 18204 20300 18232
rect 20666 18204 20694 18235
rect 21174 18232 21180 18284
rect 21232 18232 21238 18284
rect 21358 18232 21364 18284
rect 21416 18232 21422 18284
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18241 21511 18275
rect 21560 18272 21588 18300
rect 21928 18281 21956 18312
rect 23109 18309 23121 18312
rect 23155 18309 23167 18343
rect 24780 18340 24808 18368
rect 27341 18343 27399 18349
rect 24780 18312 25728 18340
rect 23109 18303 23167 18309
rect 21628 18275 21686 18281
rect 21628 18272 21640 18275
rect 21560 18244 21640 18272
rect 21453 18235 21511 18241
rect 21628 18241 21640 18244
rect 21674 18241 21686 18275
rect 21753 18275 21811 18281
rect 21753 18272 21765 18275
rect 21628 18235 21686 18241
rect 21752 18241 21765 18272
rect 21799 18241 21811 18275
rect 21752 18235 21811 18241
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18241 21971 18275
rect 21913 18235 21971 18241
rect 20272 18176 20694 18204
rect 20809 18207 20867 18213
rect 20165 18167 20223 18173
rect 20809 18173 20821 18207
rect 20855 18204 20867 18207
rect 21376 18204 21404 18232
rect 20855 18176 21404 18204
rect 21468 18204 21496 18235
rect 21542 18204 21548 18216
rect 21468 18176 21548 18204
rect 20855 18173 20867 18176
rect 20809 18167 20867 18173
rect 17034 18096 17040 18148
rect 17092 18096 17098 18148
rect 17862 18136 17868 18148
rect 17144 18108 17868 18136
rect 17144 18080 17172 18108
rect 17862 18096 17868 18108
rect 17920 18136 17926 18148
rect 18049 18139 18107 18145
rect 18049 18136 18061 18139
rect 17920 18108 18061 18136
rect 17920 18096 17926 18108
rect 18049 18105 18061 18108
rect 18095 18105 18107 18139
rect 18340 18136 18368 18167
rect 18049 18099 18107 18105
rect 18156 18108 18368 18136
rect 20073 18139 20131 18145
rect 18156 18080 18184 18108
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20438 18136 20444 18148
rect 20119 18108 20444 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 20438 18096 20444 18108
rect 20496 18136 20502 18148
rect 20824 18136 20852 18167
rect 21542 18164 21548 18176
rect 21600 18204 21606 18216
rect 21752 18204 21780 18235
rect 22738 18232 22744 18284
rect 22796 18232 22802 18284
rect 22830 18232 22836 18284
rect 22888 18232 22894 18284
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24394 18272 24400 18284
rect 24268 18244 24400 18272
rect 24268 18232 24274 18244
rect 24394 18232 24400 18244
rect 24452 18272 24458 18284
rect 24854 18272 24860 18284
rect 24452 18244 24860 18272
rect 24452 18232 24458 18244
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 24946 18232 24952 18284
rect 25004 18272 25010 18284
rect 25041 18275 25099 18281
rect 25041 18272 25053 18275
rect 25004 18244 25053 18272
rect 25004 18232 25010 18244
rect 25041 18241 25053 18244
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 25590 18232 25596 18284
rect 25648 18232 25654 18284
rect 25700 18281 25728 18312
rect 26620 18312 27108 18340
rect 26620 18281 26648 18312
rect 25685 18275 25743 18281
rect 25685 18241 25697 18275
rect 25731 18241 25743 18275
rect 25685 18235 25743 18241
rect 26605 18275 26663 18281
rect 26605 18241 26617 18275
rect 26651 18241 26663 18275
rect 26605 18235 26663 18241
rect 26881 18275 26939 18281
rect 26881 18241 26893 18275
rect 26927 18272 26939 18275
rect 26970 18272 26976 18284
rect 26927 18244 26976 18272
rect 26927 18241 26939 18244
rect 26881 18235 26939 18241
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 27080 18272 27108 18312
rect 27341 18309 27353 18343
rect 27387 18340 27399 18343
rect 27522 18340 27528 18352
rect 27387 18312 27528 18340
rect 27387 18309 27399 18312
rect 27341 18303 27399 18309
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 27614 18300 27620 18352
rect 27672 18340 27678 18352
rect 28813 18343 28871 18349
rect 28813 18340 28825 18343
rect 27672 18312 28825 18340
rect 27672 18300 27678 18312
rect 28813 18309 28825 18312
rect 28859 18309 28871 18343
rect 29196 18340 29224 18368
rect 29288 18352 29316 18380
rect 28813 18303 28871 18309
rect 29104 18312 29224 18340
rect 27080 18244 27568 18272
rect 23106 18204 23112 18216
rect 21600 18176 21780 18204
rect 22940 18176 23112 18204
rect 21600 18164 21606 18176
rect 20496 18108 20852 18136
rect 22557 18139 22615 18145
rect 20496 18096 20502 18108
rect 22557 18105 22569 18139
rect 22603 18136 22615 18139
rect 22940 18136 22968 18176
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 25148 18204 25176 18232
rect 24627 18176 25176 18204
rect 25225 18207 25283 18213
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25225 18173 25237 18207
rect 25271 18173 25283 18207
rect 25608 18204 25636 18232
rect 27433 18207 27491 18213
rect 27433 18204 27445 18207
rect 25608 18176 27445 18204
rect 25225 18167 25283 18173
rect 27433 18173 27445 18176
rect 27479 18173 27491 18207
rect 27433 18167 27491 18173
rect 25240 18136 25268 18167
rect 22603 18108 22968 18136
rect 24872 18108 25268 18136
rect 22603 18105 22615 18108
rect 22557 18099 22615 18105
rect 24872 18080 24900 18108
rect 25958 18096 25964 18148
rect 26016 18136 26022 18148
rect 26053 18139 26111 18145
rect 26053 18136 26065 18139
rect 26016 18108 26065 18136
rect 26016 18096 26022 18108
rect 26053 18105 26065 18108
rect 26099 18136 26111 18139
rect 26099 18108 26648 18136
rect 26099 18105 26111 18108
rect 26053 18099 26111 18105
rect 26620 18080 26648 18108
rect 26970 18096 26976 18148
rect 27028 18096 27034 18148
rect 27540 18136 27568 18244
rect 27890 18232 27896 18284
rect 27948 18272 27954 18284
rect 29104 18281 29132 18312
rect 29270 18300 29276 18352
rect 29328 18300 29334 18352
rect 29365 18343 29423 18349
rect 29365 18309 29377 18343
rect 29411 18340 29423 18343
rect 29638 18340 29644 18352
rect 29411 18312 29644 18340
rect 29411 18309 29423 18312
rect 29365 18303 29423 18309
rect 29638 18300 29644 18312
rect 29696 18300 29702 18352
rect 29827 18312 29855 18380
rect 30190 18368 30196 18380
rect 30248 18368 30254 18420
rect 30742 18368 30748 18420
rect 30800 18408 30806 18420
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 30800 18380 31493 18408
rect 30800 18368 30806 18380
rect 31481 18377 31493 18380
rect 31527 18377 31539 18411
rect 31481 18371 31539 18377
rect 32306 18368 32312 18420
rect 32364 18408 32370 18420
rect 32364 18380 32628 18408
rect 32364 18368 32370 18380
rect 30834 18300 30840 18352
rect 30892 18340 30898 18352
rect 30929 18343 30987 18349
rect 30929 18340 30941 18343
rect 30892 18312 30941 18340
rect 30892 18300 30898 18312
rect 30929 18309 30941 18312
rect 30975 18309 30987 18343
rect 31145 18343 31203 18349
rect 31145 18340 31157 18343
rect 30929 18303 30987 18309
rect 31023 18312 31157 18340
rect 28169 18275 28227 18281
rect 28169 18272 28181 18275
rect 27948 18244 28181 18272
rect 27948 18232 27954 18244
rect 28169 18241 28181 18244
rect 28215 18272 28227 18275
rect 28629 18275 28687 18281
rect 28629 18272 28641 18275
rect 28215 18244 28641 18272
rect 28215 18241 28227 18244
rect 28169 18235 28227 18241
rect 28629 18241 28641 18244
rect 28675 18241 28687 18275
rect 28629 18235 28687 18241
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18241 29147 18275
rect 31023 18272 31051 18312
rect 31145 18309 31157 18312
rect 31191 18340 31203 18343
rect 32122 18340 32128 18352
rect 31191 18312 31524 18340
rect 31191 18309 31203 18312
rect 31145 18303 31203 18309
rect 31496 18284 31524 18312
rect 31864 18312 32128 18340
rect 29089 18235 29147 18241
rect 30576 18244 31051 18272
rect 27617 18207 27675 18213
rect 27617 18173 27629 18207
rect 27663 18204 27675 18207
rect 28353 18207 28411 18213
rect 28353 18204 28365 18207
rect 27663 18176 28365 18204
rect 27663 18173 27675 18176
rect 27617 18167 27675 18173
rect 28353 18173 28365 18176
rect 28399 18204 28411 18207
rect 28902 18204 28908 18216
rect 28399 18176 28908 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 28902 18164 28908 18176
rect 28960 18164 28966 18216
rect 30006 18164 30012 18216
rect 30064 18204 30070 18216
rect 30576 18204 30604 18244
rect 31478 18232 31484 18284
rect 31536 18232 31542 18284
rect 31662 18232 31668 18284
rect 31720 18232 31726 18284
rect 31754 18232 31760 18284
rect 31812 18232 31818 18284
rect 31864 18281 31892 18312
rect 32122 18300 32128 18312
rect 32180 18340 32186 18352
rect 32490 18340 32496 18352
rect 32180 18312 32496 18340
rect 32180 18300 32186 18312
rect 32490 18300 32496 18312
rect 32548 18300 32554 18352
rect 32600 18349 32628 18380
rect 33410 18368 33416 18420
rect 33468 18408 33474 18420
rect 34057 18411 34115 18417
rect 34057 18408 34069 18411
rect 33468 18380 34069 18408
rect 33468 18368 33474 18380
rect 34057 18377 34069 18380
rect 34103 18377 34115 18411
rect 34057 18371 34115 18377
rect 34514 18368 34520 18420
rect 34572 18368 34578 18420
rect 35802 18368 35808 18420
rect 35860 18408 35866 18420
rect 36449 18411 36507 18417
rect 36449 18408 36461 18411
rect 35860 18380 36461 18408
rect 35860 18368 35866 18380
rect 36449 18377 36461 18380
rect 36495 18377 36507 18411
rect 38749 18411 38807 18417
rect 38749 18408 38761 18411
rect 36449 18371 36507 18377
rect 36556 18380 38761 18408
rect 32585 18343 32643 18349
rect 32585 18309 32597 18343
rect 32631 18309 32643 18343
rect 32585 18303 32643 18309
rect 33226 18300 33232 18352
rect 33284 18300 33290 18352
rect 34149 18343 34207 18349
rect 34149 18309 34161 18343
rect 34195 18309 34207 18343
rect 34149 18303 34207 18309
rect 31849 18275 31907 18281
rect 31849 18241 31861 18275
rect 31895 18241 31907 18275
rect 31849 18235 31907 18241
rect 30064 18176 30604 18204
rect 30837 18207 30895 18213
rect 30064 18164 30070 18176
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 30926 18204 30932 18216
rect 30883 18176 30932 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 30926 18164 30932 18176
rect 30984 18164 30990 18216
rect 31941 18207 31999 18213
rect 31941 18173 31953 18207
rect 31987 18173 31999 18207
rect 31941 18167 31999 18173
rect 27801 18139 27859 18145
rect 27801 18136 27813 18139
rect 27540 18108 27813 18136
rect 27801 18105 27813 18108
rect 27847 18105 27859 18139
rect 27801 18099 27859 18105
rect 31297 18139 31355 18145
rect 31297 18105 31309 18139
rect 31343 18136 31355 18139
rect 31956 18136 31984 18167
rect 32030 18164 32036 18216
rect 32088 18204 32094 18216
rect 32306 18204 32312 18216
rect 32088 18176 32312 18204
rect 32088 18164 32094 18176
rect 32306 18164 32312 18176
rect 32364 18164 32370 18216
rect 32674 18164 32680 18216
rect 32732 18204 32738 18216
rect 34164 18204 34192 18303
rect 34238 18300 34244 18352
rect 34296 18340 34302 18352
rect 34349 18343 34407 18349
rect 34349 18340 34361 18343
rect 34296 18312 34361 18340
rect 34296 18300 34302 18312
rect 34349 18309 34361 18312
rect 34395 18309 34407 18343
rect 34349 18303 34407 18309
rect 34882 18300 34888 18352
rect 34940 18340 34946 18352
rect 34940 18312 35466 18340
rect 34940 18300 34946 18312
rect 34701 18275 34759 18281
rect 34701 18241 34713 18275
rect 34747 18241 34759 18275
rect 34701 18235 34759 18241
rect 32732 18176 34192 18204
rect 32732 18164 32738 18176
rect 34514 18164 34520 18216
rect 34572 18204 34578 18216
rect 34716 18204 34744 18235
rect 34572 18176 34744 18204
rect 34572 18164 34578 18176
rect 34974 18164 34980 18216
rect 35032 18164 35038 18216
rect 31343 18108 31984 18136
rect 31343 18105 31355 18108
rect 31297 18099 31355 18105
rect 34146 18096 34152 18148
rect 34204 18136 34210 18148
rect 34204 18108 34836 18136
rect 34204 18096 34210 18108
rect 16080 18040 16804 18068
rect 16080 18028 16086 18040
rect 17126 18028 17132 18080
rect 17184 18028 17190 18080
rect 17310 18028 17316 18080
rect 17368 18028 17374 18080
rect 17494 18028 17500 18080
rect 17552 18028 17558 18080
rect 18138 18028 18144 18080
rect 18196 18028 18202 18080
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20806 18068 20812 18080
rect 20036 18040 20812 18068
rect 20036 18028 20042 18040
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21545 18071 21603 18077
rect 21545 18068 21557 18071
rect 20956 18040 21557 18068
rect 20956 18028 20962 18040
rect 21545 18037 21557 18040
rect 21591 18037 21603 18071
rect 21545 18031 21603 18037
rect 24854 18028 24860 18080
rect 24912 18028 24918 18080
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25130 18068 25136 18080
rect 25004 18040 25136 18068
rect 25004 18028 25010 18040
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 26418 18028 26424 18080
rect 26476 18028 26482 18080
rect 26602 18028 26608 18080
rect 26660 18028 26666 18080
rect 26697 18071 26755 18077
rect 26697 18037 26709 18071
rect 26743 18068 26755 18071
rect 27154 18068 27160 18080
rect 26743 18040 27160 18068
rect 26743 18037 26755 18040
rect 26697 18031 26755 18037
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 28994 18028 29000 18080
rect 29052 18028 29058 18080
rect 31110 18028 31116 18080
rect 31168 18068 31174 18080
rect 33226 18068 33232 18080
rect 31168 18040 33232 18068
rect 31168 18028 31174 18040
rect 33226 18028 33232 18040
rect 33284 18068 33290 18080
rect 34333 18071 34391 18077
rect 34333 18068 34345 18071
rect 33284 18040 34345 18068
rect 33284 18028 33290 18040
rect 34333 18037 34345 18040
rect 34379 18037 34391 18071
rect 34808 18068 34836 18108
rect 36556 18068 36584 18380
rect 38749 18377 38761 18380
rect 38795 18377 38807 18411
rect 38749 18371 38807 18377
rect 39022 18368 39028 18420
rect 39080 18408 39086 18420
rect 39209 18411 39267 18417
rect 39209 18408 39221 18411
rect 39080 18380 39221 18408
rect 39080 18368 39086 18380
rect 39209 18377 39221 18380
rect 39255 18377 39267 18411
rect 39209 18371 39267 18377
rect 39298 18368 39304 18420
rect 39356 18368 39362 18420
rect 40034 18368 40040 18420
rect 40092 18368 40098 18420
rect 41233 18411 41291 18417
rect 41233 18377 41245 18411
rect 41279 18408 41291 18411
rect 41506 18408 41512 18420
rect 41279 18380 41512 18408
rect 41279 18377 41291 18380
rect 41233 18371 41291 18377
rect 41506 18368 41512 18380
rect 41564 18368 41570 18420
rect 42702 18408 42708 18420
rect 42076 18380 42708 18408
rect 37090 18300 37096 18352
rect 37148 18340 37154 18352
rect 37185 18343 37243 18349
rect 37185 18340 37197 18343
rect 37148 18312 37197 18340
rect 37148 18300 37154 18312
rect 37185 18309 37197 18312
rect 37231 18309 37243 18343
rect 37185 18303 37243 18309
rect 37274 18300 37280 18352
rect 37332 18340 37338 18352
rect 39117 18343 39175 18349
rect 37332 18312 37674 18340
rect 37332 18300 37338 18312
rect 39117 18309 39129 18343
rect 39163 18340 39175 18343
rect 39316 18340 39344 18368
rect 40954 18340 40960 18352
rect 39163 18312 39344 18340
rect 40328 18312 40960 18340
rect 39163 18309 39175 18312
rect 39117 18303 39175 18309
rect 39945 18275 40003 18281
rect 39945 18272 39957 18275
rect 38672 18244 39957 18272
rect 36906 18164 36912 18216
rect 36964 18164 36970 18216
rect 38470 18096 38476 18148
rect 38528 18136 38534 18148
rect 38672 18145 38700 18244
rect 39945 18241 39957 18244
rect 39991 18241 40003 18275
rect 39945 18235 40003 18241
rect 40328 18216 40356 18312
rect 40954 18300 40960 18312
rect 41012 18340 41018 18352
rect 42076 18349 42104 18380
rect 42702 18368 42708 18380
rect 42760 18368 42766 18420
rect 42978 18368 42984 18420
rect 43036 18408 43042 18420
rect 43533 18411 43591 18417
rect 43533 18408 43545 18411
rect 43036 18380 43545 18408
rect 43036 18368 43042 18380
rect 43533 18377 43545 18380
rect 43579 18377 43591 18411
rect 43533 18371 43591 18377
rect 43714 18368 43720 18420
rect 43772 18408 43778 18420
rect 44177 18411 44235 18417
rect 44177 18408 44189 18411
rect 43772 18380 44189 18408
rect 43772 18368 43778 18380
rect 44177 18377 44189 18380
rect 44223 18408 44235 18411
rect 44818 18408 44824 18420
rect 44223 18380 44824 18408
rect 44223 18377 44235 18380
rect 44177 18371 44235 18377
rect 44818 18368 44824 18380
rect 44876 18408 44882 18420
rect 44913 18411 44971 18417
rect 44913 18408 44925 18411
rect 44876 18380 44925 18408
rect 44876 18368 44882 18380
rect 44913 18377 44925 18380
rect 44959 18377 44971 18411
rect 44913 18371 44971 18377
rect 42061 18343 42119 18349
rect 41012 18312 41460 18340
rect 41012 18300 41018 18312
rect 40773 18275 40831 18281
rect 40773 18241 40785 18275
rect 40819 18272 40831 18275
rect 40819 18244 40908 18272
rect 40819 18241 40831 18244
rect 40773 18235 40831 18241
rect 38930 18164 38936 18216
rect 38988 18204 38994 18216
rect 39301 18207 39359 18213
rect 39301 18204 39313 18207
rect 38988 18176 39313 18204
rect 38988 18164 38994 18176
rect 39301 18173 39313 18176
rect 39347 18173 39359 18207
rect 39301 18167 39359 18173
rect 39850 18164 39856 18216
rect 39908 18204 39914 18216
rect 40129 18207 40187 18213
rect 40129 18204 40141 18207
rect 39908 18176 40141 18204
rect 39908 18164 39914 18176
rect 40129 18173 40141 18176
rect 40175 18204 40187 18207
rect 40310 18204 40316 18216
rect 40175 18176 40316 18204
rect 40175 18173 40187 18176
rect 40129 18167 40187 18173
rect 40310 18164 40316 18176
rect 40368 18164 40374 18216
rect 40880 18145 40908 18244
rect 41432 18213 41460 18312
rect 42061 18309 42073 18343
rect 42107 18309 42119 18343
rect 42061 18303 42119 18309
rect 42794 18300 42800 18352
rect 42852 18300 42858 18352
rect 41690 18232 41696 18284
rect 41748 18272 41754 18284
rect 41748 18244 41828 18272
rect 41748 18232 41754 18244
rect 41800 18213 41828 18244
rect 41325 18207 41383 18213
rect 41325 18173 41337 18207
rect 41371 18173 41383 18207
rect 41325 18167 41383 18173
rect 41417 18207 41475 18213
rect 41417 18173 41429 18207
rect 41463 18173 41475 18207
rect 41417 18167 41475 18173
rect 41785 18207 41843 18213
rect 41785 18173 41797 18207
rect 41831 18204 41843 18207
rect 42058 18204 42064 18216
rect 41831 18176 42064 18204
rect 41831 18173 41843 18176
rect 41785 18167 41843 18173
rect 38657 18139 38715 18145
rect 38657 18136 38669 18139
rect 38528 18108 38669 18136
rect 38528 18096 38534 18108
rect 38657 18105 38669 18108
rect 38703 18105 38715 18139
rect 38657 18099 38715 18105
rect 40865 18139 40923 18145
rect 40865 18105 40877 18139
rect 40911 18105 40923 18139
rect 41340 18136 41368 18167
rect 42058 18164 42064 18176
rect 42116 18164 42122 18216
rect 42794 18164 42800 18216
rect 42852 18204 42858 18216
rect 43806 18204 43812 18216
rect 42852 18176 43812 18204
rect 42852 18164 42858 18176
rect 43806 18164 43812 18176
rect 43864 18204 43870 18216
rect 44545 18207 44603 18213
rect 44545 18204 44557 18207
rect 43864 18176 44557 18204
rect 43864 18164 43870 18176
rect 44545 18173 44557 18176
rect 44591 18173 44603 18207
rect 44545 18167 44603 18173
rect 41340 18108 41460 18136
rect 40865 18099 40923 18105
rect 34808 18040 36584 18068
rect 34333 18031 34391 18037
rect 37274 18028 37280 18080
rect 37332 18068 37338 18080
rect 38930 18068 38936 18080
rect 37332 18040 38936 18068
rect 37332 18028 37338 18040
rect 38930 18028 38936 18040
rect 38988 18028 38994 18080
rect 39022 18028 39028 18080
rect 39080 18068 39086 18080
rect 39577 18071 39635 18077
rect 39577 18068 39589 18071
rect 39080 18040 39589 18068
rect 39080 18028 39086 18040
rect 39577 18037 39589 18040
rect 39623 18037 39635 18071
rect 39577 18031 39635 18037
rect 40586 18028 40592 18080
rect 40644 18028 40650 18080
rect 41432 18068 41460 18108
rect 41506 18068 41512 18080
rect 41432 18040 41512 18068
rect 41506 18028 41512 18040
rect 41564 18068 41570 18080
rect 42242 18068 42248 18080
rect 41564 18040 42248 18068
rect 41564 18028 41570 18040
rect 42242 18028 42248 18040
rect 42300 18028 42306 18080
rect 460 17978 45540 18000
rect 460 17926 3570 17978
rect 3622 17926 3634 17978
rect 3686 17926 3698 17978
rect 3750 17926 3762 17978
rect 3814 17926 3826 17978
rect 3878 17926 8570 17978
rect 8622 17926 8634 17978
rect 8686 17926 8698 17978
rect 8750 17926 8762 17978
rect 8814 17926 8826 17978
rect 8878 17926 13570 17978
rect 13622 17926 13634 17978
rect 13686 17926 13698 17978
rect 13750 17926 13762 17978
rect 13814 17926 13826 17978
rect 13878 17926 18570 17978
rect 18622 17926 18634 17978
rect 18686 17926 18698 17978
rect 18750 17926 18762 17978
rect 18814 17926 18826 17978
rect 18878 17926 23570 17978
rect 23622 17926 23634 17978
rect 23686 17926 23698 17978
rect 23750 17926 23762 17978
rect 23814 17926 23826 17978
rect 23878 17926 28570 17978
rect 28622 17926 28634 17978
rect 28686 17926 28698 17978
rect 28750 17926 28762 17978
rect 28814 17926 28826 17978
rect 28878 17926 33570 17978
rect 33622 17926 33634 17978
rect 33686 17926 33698 17978
rect 33750 17926 33762 17978
rect 33814 17926 33826 17978
rect 33878 17926 38570 17978
rect 38622 17926 38634 17978
rect 38686 17926 38698 17978
rect 38750 17926 38762 17978
rect 38814 17926 38826 17978
rect 38878 17926 43570 17978
rect 43622 17926 43634 17978
rect 43686 17926 43698 17978
rect 43750 17926 43762 17978
rect 43814 17926 43826 17978
rect 43878 17926 45540 17978
rect 460 17904 45540 17926
rect 3881 17867 3939 17873
rect 3881 17864 3893 17867
rect 3528 17836 3893 17864
rect 3528 17669 3556 17836
rect 3881 17833 3893 17836
rect 3927 17833 3939 17867
rect 3881 17827 3939 17833
rect 4430 17824 4436 17876
rect 4488 17824 4494 17876
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 6822 17864 6828 17876
rect 6420 17836 6828 17864
rect 6420 17824 6426 17836
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7742 17824 7748 17876
rect 7800 17824 7806 17876
rect 8386 17824 8392 17876
rect 8444 17824 8450 17876
rect 9306 17824 9312 17876
rect 9364 17824 9370 17876
rect 9582 17824 9588 17876
rect 9640 17824 9646 17876
rect 9858 17824 9864 17876
rect 9916 17824 9922 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 12710 17864 12716 17876
rect 10827 17836 12716 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 12986 17824 12992 17876
rect 13044 17864 13050 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 13044 17836 13185 17864
rect 13044 17824 13050 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 15381 17867 15439 17873
rect 15381 17864 15393 17867
rect 13412 17836 15393 17864
rect 13412 17824 13418 17836
rect 15381 17833 15393 17836
rect 15427 17833 15439 17867
rect 15381 17827 15439 17833
rect 16298 17824 16304 17876
rect 16356 17824 16362 17876
rect 17037 17867 17095 17873
rect 17037 17833 17049 17867
rect 17083 17864 17095 17867
rect 17865 17867 17923 17873
rect 17083 17836 17264 17864
rect 17083 17833 17095 17836
rect 17037 17827 17095 17833
rect 4448 17796 4476 17824
rect 3712 17768 4476 17796
rect 7760 17796 7788 17824
rect 8757 17799 8815 17805
rect 8757 17796 8769 17799
rect 7760 17768 8769 17796
rect 3712 17669 3740 17768
rect 8757 17765 8769 17768
rect 8803 17796 8815 17799
rect 9217 17799 9275 17805
rect 9217 17796 9229 17799
rect 8803 17768 9229 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 9217 17765 9229 17768
rect 9263 17765 9275 17799
rect 9217 17759 9275 17765
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 5534 17728 5540 17740
rect 4847 17700 5540 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5534 17688 5540 17700
rect 5592 17688 5598 17740
rect 5920 17700 7788 17728
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17629 3571 17663
rect 3513 17623 3571 17629
rect 3697 17663 3755 17669
rect 3697 17629 3709 17663
rect 3743 17629 3755 17663
rect 3697 17623 3755 17629
rect 3789 17663 3847 17669
rect 3789 17629 3801 17663
rect 3835 17629 3847 17663
rect 3789 17623 3847 17629
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17660 4031 17663
rect 4019 17632 4292 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 3804 17592 3832 17623
rect 4065 17595 4123 17601
rect 4065 17592 4077 17595
rect 3804 17564 4077 17592
rect 4065 17561 4077 17564
rect 4111 17592 4123 17595
rect 4154 17592 4160 17604
rect 4111 17564 4160 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 4154 17552 4160 17564
rect 4212 17552 4218 17604
rect 4264 17601 4292 17632
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4488 17632 4537 17660
rect 4488 17620 4494 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 5920 17646 5948 17700
rect 4525 17623 4583 17629
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 7760 17660 7788 17700
rect 8110 17688 8116 17740
rect 8168 17688 8174 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8527 17700 8892 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8018 17660 8024 17672
rect 7760 17646 8024 17660
rect 7774 17632 8024 17646
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 8128 17660 8156 17688
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 8128 17632 8585 17660
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17561 4307 17595
rect 4249 17555 4307 17561
rect 3418 17484 3424 17536
rect 3476 17484 3482 17536
rect 3697 17527 3755 17533
rect 3697 17493 3709 17527
rect 3743 17524 3755 17527
rect 3970 17524 3976 17536
rect 3743 17496 3976 17524
rect 3743 17493 3755 17496
rect 3697 17487 3755 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4264 17524 4292 17555
rect 6638 17552 6644 17604
rect 6696 17552 6702 17604
rect 8297 17595 8355 17601
rect 8297 17561 8309 17595
rect 8343 17561 8355 17595
rect 8297 17555 8355 17561
rect 5626 17524 5632 17536
rect 4264 17496 5632 17524
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 5868 17496 6285 17524
rect 5868 17484 5874 17496
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6273 17487 6331 17493
rect 6546 17484 6552 17536
rect 6604 17524 6610 17536
rect 8312 17524 8340 17555
rect 8864 17536 8892 17700
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 9232 17660 9260 17759
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 9600 17728 9628 17824
rect 11330 17756 11336 17808
rect 11388 17796 11394 17808
rect 11388 17768 13492 17796
rect 11388 17756 11394 17768
rect 9447 17700 9628 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 11425 17731 11483 17737
rect 11425 17728 11437 17731
rect 10192 17700 11437 17728
rect 10192 17688 10198 17700
rect 11425 17697 11437 17700
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 12250 17728 12256 17740
rect 12207 17700 12256 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 12526 17688 12532 17740
rect 12584 17688 12590 17740
rect 13464 17728 13492 17768
rect 15194 17756 15200 17808
rect 15252 17805 15258 17808
rect 15252 17799 15301 17805
rect 15252 17765 15255 17799
rect 15289 17796 15301 17799
rect 16316 17796 16344 17824
rect 16758 17796 16764 17808
rect 15289 17768 16344 17796
rect 16408 17768 16764 17796
rect 15289 17765 15301 17768
rect 15252 17759 15301 17765
rect 15252 17756 15258 17759
rect 13817 17731 13875 17737
rect 13464 17700 13768 17728
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 9232 17632 9505 17660
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9585 17663 9643 17669
rect 9585 17629 9597 17663
rect 9631 17629 9643 17663
rect 9585 17623 9643 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 12342 17660 12348 17672
rect 11287 17632 12348 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 9140 17592 9168 17620
rect 9600 17592 9628 17623
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 13354 17660 13360 17672
rect 12483 17632 13360 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17629 13507 17663
rect 13740 17660 13768 17700
rect 13817 17697 13829 17731
rect 13863 17728 13875 17731
rect 15102 17728 15108 17740
rect 13863 17700 15108 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15838 17688 15844 17740
rect 15896 17688 15902 17740
rect 16022 17688 16028 17740
rect 16080 17688 16086 17740
rect 16408 17728 16436 17768
rect 16758 17756 16764 17768
rect 16816 17756 16822 17808
rect 16942 17756 16948 17808
rect 17000 17756 17006 17808
rect 17236 17796 17264 17836
rect 17865 17833 17877 17867
rect 17911 17864 17923 17867
rect 17954 17864 17960 17876
rect 17911 17836 17960 17864
rect 17911 17833 17923 17836
rect 17865 17827 17923 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 19061 17867 19119 17873
rect 19061 17833 19073 17867
rect 19107 17864 19119 17867
rect 19610 17864 19616 17876
rect 19107 17836 19616 17864
rect 19107 17833 19119 17836
rect 19061 17827 19119 17833
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 19978 17864 19984 17876
rect 19720 17836 19984 17864
rect 19245 17799 19303 17805
rect 19245 17796 19257 17799
rect 17236 17768 19257 17796
rect 19245 17765 19257 17768
rect 19291 17765 19303 17799
rect 19720 17796 19748 17836
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20073 17867 20131 17873
rect 20073 17833 20085 17867
rect 20119 17864 20131 17867
rect 20346 17864 20352 17876
rect 20119 17836 20352 17864
rect 20119 17833 20131 17836
rect 20073 17827 20131 17833
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20806 17824 20812 17876
rect 20864 17824 20870 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 22005 17867 22063 17873
rect 22005 17864 22017 17867
rect 21968 17836 22017 17864
rect 21968 17824 21974 17836
rect 22005 17833 22017 17836
rect 22051 17864 22063 17867
rect 22370 17864 22376 17876
rect 22051 17836 22376 17864
rect 22051 17833 22063 17836
rect 22005 17827 22063 17833
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22796 17836 22845 17864
rect 22796 17824 22802 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 27522 17824 27528 17876
rect 27580 17864 27586 17876
rect 28261 17867 28319 17873
rect 28261 17864 28273 17867
rect 27580 17836 28273 17864
rect 27580 17824 27586 17836
rect 28261 17833 28273 17836
rect 28307 17833 28319 17867
rect 28261 17827 28319 17833
rect 20717 17799 20775 17805
rect 20717 17796 20729 17799
rect 19245 17759 19303 17765
rect 19352 17768 19748 17796
rect 19812 17768 20729 17796
rect 16316 17700 16436 17728
rect 16485 17731 16543 17737
rect 13906 17660 13912 17672
rect 13740 17632 13912 17660
rect 13449 17623 13507 17629
rect 9140 17564 9628 17592
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 10321 17595 10379 17601
rect 10321 17592 10333 17595
rect 9824 17564 10333 17592
rect 9824 17552 9830 17564
rect 10321 17561 10333 17564
rect 10367 17561 10379 17595
rect 10321 17555 10379 17561
rect 11348 17564 12204 17592
rect 6604 17496 8340 17524
rect 6604 17484 6610 17496
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 9950 17524 9956 17536
rect 8904 17496 9956 17524
rect 8904 17484 8910 17496
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11348 17533 11376 17564
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10836 17496 10885 17524
rect 10836 17484 10842 17496
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 10873 17487 10931 17493
rect 11333 17527 11391 17533
rect 11333 17493 11345 17527
rect 11379 17493 11391 17527
rect 12176 17524 12204 17564
rect 12986 17552 12992 17604
rect 13044 17592 13050 17604
rect 13464 17592 13492 17623
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 16316 17669 16344 17700
rect 16485 17697 16497 17731
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16390 17620 16396 17672
rect 16448 17620 16454 17672
rect 16500 17660 16528 17691
rect 16850 17688 16856 17740
rect 16908 17688 16914 17740
rect 16960 17728 16988 17756
rect 17037 17731 17095 17737
rect 17037 17728 17049 17731
rect 16960 17700 17049 17728
rect 17037 17697 17049 17700
rect 17083 17697 17095 17731
rect 17037 17691 17095 17697
rect 17310 17688 17316 17740
rect 17368 17688 17374 17740
rect 17678 17688 17684 17740
rect 17736 17728 17742 17740
rect 18969 17731 19027 17737
rect 17736 17700 17816 17728
rect 17736 17688 17742 17700
rect 16574 17660 16580 17672
rect 16500 17632 16580 17660
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 16868 17660 16896 17688
rect 16715 17632 17080 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 17052 17604 17080 17632
rect 17126 17620 17132 17672
rect 17184 17620 17190 17672
rect 17328 17660 17356 17688
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17328 17632 17417 17660
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 17494 17620 17500 17672
rect 17552 17620 17558 17672
rect 17586 17620 17592 17672
rect 17644 17620 17650 17672
rect 17788 17669 17816 17700
rect 18969 17697 18981 17731
rect 19015 17728 19027 17731
rect 19352 17728 19380 17768
rect 19702 17728 19708 17740
rect 19015 17700 19380 17728
rect 19444 17700 19708 17728
rect 19015 17697 19027 17700
rect 18969 17691 19027 17697
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 19444 17669 19472 17700
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 19812 17669 19840 17768
rect 20717 17765 20729 17768
rect 20763 17796 20775 17799
rect 20990 17796 20996 17808
rect 20763 17768 20996 17796
rect 20763 17765 20775 17768
rect 20717 17759 20775 17765
rect 20990 17756 20996 17768
rect 21048 17756 21054 17808
rect 23753 17799 23811 17805
rect 23753 17796 23765 17799
rect 22756 17768 23765 17796
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 21174 17728 21180 17740
rect 20303 17700 21180 17728
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 21174 17688 21180 17700
rect 21232 17728 21238 17740
rect 22002 17728 22008 17740
rect 21232 17700 22008 17728
rect 21232 17688 21238 17700
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18196 17632 18337 17660
rect 18196 17620 18202 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 19061 17663 19119 17669
rect 19061 17629 19073 17663
rect 19107 17629 19119 17663
rect 19061 17623 19119 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 20073 17663 20131 17669
rect 20073 17660 20085 17663
rect 19797 17623 19855 17629
rect 19904 17632 20085 17660
rect 15749 17595 15807 17601
rect 13044 17564 13492 17592
rect 14108 17564 14214 17592
rect 13044 17552 13050 17564
rect 12434 17524 12440 17536
rect 12176 17496 12440 17524
rect 11333 17487 11391 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12802 17484 12808 17536
rect 12860 17484 12866 17536
rect 14108 17524 14136 17564
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 15795 17564 16711 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 14274 17524 14280 17536
rect 14108 17496 14280 17524
rect 14274 17484 14280 17496
rect 14332 17524 14338 17536
rect 14734 17524 14740 17536
rect 14332 17496 14740 17524
rect 14332 17484 14338 17496
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16540 17496 16589 17524
rect 16540 17484 16546 17496
rect 16577 17493 16589 17496
rect 16623 17493 16635 17527
rect 16683 17524 16711 17564
rect 16850 17552 16856 17604
rect 16908 17552 16914 17604
rect 17034 17552 17040 17604
rect 17092 17552 17098 17604
rect 17512 17592 17540 17620
rect 17144 17564 17540 17592
rect 17604 17592 17632 17620
rect 18601 17595 18659 17601
rect 18601 17592 18613 17595
rect 17604 17564 18613 17592
rect 17144 17524 17172 17564
rect 18601 17561 18613 17564
rect 18647 17561 18659 17595
rect 19076 17592 19104 17623
rect 19334 17592 19340 17604
rect 19076 17564 19340 17592
rect 18601 17555 18659 17561
rect 19334 17552 19340 17564
rect 19392 17592 19398 17604
rect 19628 17592 19656 17623
rect 19392 17564 19656 17592
rect 19392 17552 19398 17564
rect 16683 17496 17172 17524
rect 16577 17487 16635 17493
rect 17310 17484 17316 17536
rect 17368 17484 17374 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 18874 17524 18880 17536
rect 17635 17496 18880 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 18874 17484 18880 17496
rect 18932 17524 18938 17536
rect 19426 17524 19432 17536
rect 18932 17496 19432 17524
rect 18932 17484 18938 17496
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19518 17484 19524 17536
rect 19576 17484 19582 17536
rect 19904 17524 19932 17632
rect 20073 17629 20085 17632
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17660 20407 17663
rect 20438 17660 20444 17672
rect 20395 17632 20444 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 22756 17669 22784 17768
rect 23753 17765 23765 17768
rect 23799 17765 23811 17799
rect 23753 17759 23811 17765
rect 23290 17688 23296 17740
rect 23348 17688 23354 17740
rect 23382 17688 23388 17740
rect 23440 17728 23446 17740
rect 24305 17731 24363 17737
rect 24305 17728 24317 17731
rect 23440 17700 24317 17728
rect 23440 17688 23446 17700
rect 24305 17697 24317 17700
rect 24351 17728 24363 17731
rect 24854 17728 24860 17740
rect 24351 17700 24860 17728
rect 24351 17697 24363 17700
rect 24305 17691 24363 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17728 25099 17731
rect 25087 17700 26832 17728
rect 25087 17697 25099 17700
rect 25041 17691 25099 17697
rect 26804 17672 26832 17700
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 19978 17552 19984 17604
rect 20036 17592 20042 17604
rect 20622 17592 20628 17604
rect 20036 17564 20628 17592
rect 20036 17552 20042 17564
rect 20622 17552 20628 17564
rect 20680 17592 20686 17604
rect 21284 17592 21312 17623
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 27154 17669 27160 17672
rect 26881 17663 26939 17669
rect 26881 17660 26893 17663
rect 26844 17632 26893 17660
rect 26844 17620 26850 17632
rect 26881 17629 26893 17632
rect 26927 17629 26939 17663
rect 26881 17623 26939 17629
rect 27137 17663 27160 17669
rect 27137 17629 27149 17663
rect 27137 17623 27160 17629
rect 27154 17620 27160 17623
rect 27212 17620 27218 17672
rect 28276 17660 28304 17827
rect 29914 17824 29920 17876
rect 29972 17864 29978 17876
rect 30653 17867 30711 17873
rect 30653 17864 30665 17867
rect 29972 17836 30665 17864
rect 29972 17824 29978 17836
rect 30653 17833 30665 17836
rect 30699 17833 30711 17867
rect 30653 17827 30711 17833
rect 31021 17867 31079 17873
rect 31021 17833 31033 17867
rect 31067 17864 31079 17867
rect 31110 17864 31116 17876
rect 31067 17836 31116 17864
rect 31067 17833 31079 17836
rect 31021 17827 31079 17833
rect 31110 17824 31116 17836
rect 31168 17824 31174 17876
rect 31202 17824 31208 17876
rect 31260 17824 31266 17876
rect 31570 17824 31576 17876
rect 31628 17864 31634 17876
rect 32858 17864 32864 17876
rect 31628 17836 32864 17864
rect 31628 17824 31634 17836
rect 32858 17824 32864 17836
rect 32916 17824 32922 17876
rect 32950 17824 32956 17876
rect 33008 17864 33014 17876
rect 33689 17867 33747 17873
rect 33689 17864 33701 17867
rect 33008 17836 33701 17864
rect 33008 17824 33014 17836
rect 33689 17833 33701 17836
rect 33735 17833 33747 17867
rect 33689 17827 33747 17833
rect 34974 17824 34980 17876
rect 35032 17864 35038 17876
rect 35069 17867 35127 17873
rect 35069 17864 35081 17867
rect 35032 17836 35081 17864
rect 35032 17824 35038 17836
rect 35069 17833 35081 17836
rect 35115 17833 35127 17867
rect 35069 17827 35127 17833
rect 35713 17867 35771 17873
rect 35713 17833 35725 17867
rect 35759 17864 35771 17867
rect 35986 17864 35992 17876
rect 35759 17836 35992 17864
rect 35759 17833 35771 17836
rect 35713 17827 35771 17833
rect 35986 17824 35992 17836
rect 36044 17824 36050 17876
rect 36906 17824 36912 17876
rect 36964 17864 36970 17876
rect 37093 17867 37151 17873
rect 37093 17864 37105 17867
rect 36964 17836 37105 17864
rect 36964 17824 36970 17836
rect 37093 17833 37105 17836
rect 37139 17833 37151 17867
rect 37093 17827 37151 17833
rect 37645 17867 37703 17873
rect 37645 17833 37657 17867
rect 37691 17864 37703 17867
rect 38194 17864 38200 17876
rect 37691 17836 38200 17864
rect 37691 17833 37703 17836
rect 37645 17827 37703 17833
rect 38194 17824 38200 17836
rect 38252 17824 38258 17876
rect 38381 17867 38439 17873
rect 38381 17833 38393 17867
rect 38427 17864 38439 17867
rect 39482 17864 39488 17876
rect 38427 17836 39488 17864
rect 38427 17833 38439 17836
rect 38381 17827 38439 17833
rect 39482 17824 39488 17836
rect 39540 17824 39546 17876
rect 40034 17824 40040 17876
rect 40092 17824 40098 17876
rect 40310 17824 40316 17876
rect 40368 17824 40374 17876
rect 40420 17836 42012 17864
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 28721 17799 28779 17805
rect 28721 17796 28733 17799
rect 28500 17768 28733 17796
rect 28500 17756 28506 17768
rect 28721 17765 28733 17768
rect 28767 17765 28779 17799
rect 28721 17759 28779 17765
rect 30558 17756 30564 17808
rect 30616 17756 30622 17808
rect 31662 17796 31668 17808
rect 31496 17768 31668 17796
rect 28534 17688 28540 17740
rect 28592 17728 28598 17740
rect 28905 17731 28963 17737
rect 28905 17728 28917 17731
rect 28592 17700 28917 17728
rect 28592 17688 28598 17700
rect 28905 17697 28917 17700
rect 28951 17697 28963 17731
rect 28905 17691 28963 17697
rect 29181 17731 29239 17737
rect 29181 17697 29193 17731
rect 29227 17728 29239 17731
rect 30576 17728 30604 17756
rect 31496 17737 31524 17768
rect 31662 17756 31668 17768
rect 31720 17756 31726 17808
rect 31846 17756 31852 17808
rect 31904 17756 31910 17808
rect 40052 17796 40080 17824
rect 40420 17796 40448 17836
rect 33244 17768 39344 17796
rect 40052 17768 40448 17796
rect 41984 17796 42012 17836
rect 42242 17824 42248 17876
rect 42300 17864 42306 17876
rect 42429 17867 42487 17873
rect 42429 17864 42441 17867
rect 42300 17836 42441 17864
rect 42300 17824 42306 17836
rect 42429 17833 42441 17836
rect 42475 17833 42487 17867
rect 42429 17827 42487 17833
rect 44910 17824 44916 17876
rect 44968 17824 44974 17876
rect 44928 17796 44956 17824
rect 41984 17768 44956 17796
rect 29227 17700 30604 17728
rect 31481 17731 31539 17737
rect 29227 17697 29239 17700
rect 29181 17691 29239 17697
rect 31481 17697 31493 17731
rect 31527 17697 31539 17731
rect 31481 17691 31539 17697
rect 31573 17731 31631 17737
rect 31573 17697 31585 17731
rect 31619 17728 31631 17731
rect 31864 17728 31892 17756
rect 31619 17700 31892 17728
rect 31619 17697 31631 17700
rect 31573 17691 31631 17697
rect 32214 17688 32220 17740
rect 32272 17688 32278 17740
rect 32582 17688 32588 17740
rect 32640 17728 32646 17740
rect 33244 17728 33272 17768
rect 32640 17700 33272 17728
rect 32640 17688 32646 17700
rect 33778 17688 33784 17740
rect 33836 17728 33842 17740
rect 34701 17731 34759 17737
rect 34701 17728 34713 17731
rect 33836 17700 34713 17728
rect 33836 17688 33842 17700
rect 34701 17697 34713 17700
rect 34747 17728 34759 17731
rect 35618 17728 35624 17740
rect 34747 17700 35624 17728
rect 34747 17697 34759 17700
rect 34701 17691 34759 17697
rect 35618 17688 35624 17700
rect 35676 17688 35682 17740
rect 36357 17731 36415 17737
rect 36357 17728 36369 17731
rect 35728 17700 36369 17728
rect 28353 17663 28411 17669
rect 28353 17660 28365 17663
rect 28276 17632 28365 17660
rect 28353 17629 28365 17632
rect 28399 17629 28411 17663
rect 28353 17623 28411 17629
rect 28460 17632 28856 17660
rect 20680 17564 21312 17592
rect 24213 17595 24271 17601
rect 20680 17552 20686 17564
rect 24213 17561 24225 17595
rect 24259 17592 24271 17595
rect 24302 17592 24308 17604
rect 24259 17564 24308 17592
rect 24259 17561 24271 17564
rect 24213 17555 24271 17561
rect 24302 17552 24308 17564
rect 24360 17552 24366 17604
rect 25317 17595 25375 17601
rect 25317 17592 25329 17595
rect 24780 17564 25329 17592
rect 20346 17524 20352 17536
rect 19904 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21177 17527 21235 17533
rect 21177 17524 21189 17527
rect 21048 17496 21189 17524
rect 21048 17484 21054 17496
rect 21177 17493 21189 17496
rect 21223 17493 21235 17527
rect 21177 17487 21235 17493
rect 21634 17484 21640 17536
rect 21692 17484 21698 17536
rect 21910 17484 21916 17536
rect 21968 17524 21974 17536
rect 22373 17527 22431 17533
rect 22373 17524 22385 17527
rect 21968 17496 22385 17524
rect 21968 17484 21974 17496
rect 22373 17493 22385 17496
rect 22419 17493 22431 17527
rect 22373 17487 22431 17493
rect 22554 17484 22560 17536
rect 22612 17484 22618 17536
rect 23198 17484 23204 17536
rect 23256 17484 23262 17536
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 24780 17533 24808 17564
rect 25317 17561 25329 17564
rect 25363 17561 25375 17595
rect 26602 17592 26608 17604
rect 26542 17564 26608 17592
rect 25317 17555 25375 17561
rect 26602 17552 26608 17564
rect 26660 17552 26666 17604
rect 28460 17592 28488 17632
rect 26804 17564 28488 17592
rect 28537 17595 28595 17601
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 23532 17496 24133 17524
rect 23532 17484 23538 17496
rect 24121 17493 24133 17496
rect 24167 17493 24179 17527
rect 24121 17487 24179 17493
rect 24765 17527 24823 17533
rect 24765 17493 24777 17527
rect 24811 17493 24823 17527
rect 24765 17487 24823 17493
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 26804 17533 26832 17564
rect 28537 17561 28549 17595
rect 28583 17561 28595 17595
rect 28537 17555 28595 17561
rect 26789 17527 26847 17533
rect 26789 17524 26801 17527
rect 25464 17496 26801 17524
rect 25464 17484 25470 17496
rect 26789 17493 26801 17496
rect 26835 17493 26847 17527
rect 26789 17487 26847 17493
rect 27338 17484 27344 17536
rect 27396 17524 27402 17536
rect 27614 17524 27620 17536
rect 27396 17496 27620 17524
rect 27396 17484 27402 17496
rect 27614 17484 27620 17496
rect 27672 17524 27678 17536
rect 28552 17524 28580 17555
rect 28718 17524 28724 17536
rect 27672 17496 28724 17524
rect 27672 17484 27678 17496
rect 28718 17484 28724 17496
rect 28776 17484 28782 17536
rect 28828 17524 28856 17632
rect 30466 17620 30472 17672
rect 30524 17660 30530 17672
rect 31665 17663 31723 17669
rect 30524 17635 31096 17660
rect 30524 17632 31125 17635
rect 30524 17620 30530 17632
rect 31067 17629 31125 17632
rect 30190 17552 30196 17604
rect 30248 17552 30254 17604
rect 30834 17552 30840 17604
rect 30892 17552 30898 17604
rect 31067 17595 31079 17629
rect 31113 17595 31125 17629
rect 31665 17629 31677 17663
rect 31711 17629 31723 17663
rect 31665 17623 31723 17629
rect 31067 17589 31125 17595
rect 30558 17524 30564 17536
rect 28828 17496 30564 17524
rect 30558 17484 30564 17496
rect 30616 17484 30622 17536
rect 31297 17527 31355 17533
rect 31297 17493 31309 17527
rect 31343 17524 31355 17527
rect 31478 17524 31484 17536
rect 31343 17496 31484 17524
rect 31343 17493 31355 17496
rect 31297 17487 31355 17493
rect 31478 17484 31484 17496
rect 31536 17484 31542 17536
rect 31680 17524 31708 17623
rect 31754 17620 31760 17672
rect 31812 17620 31818 17672
rect 31930 17663 31988 17669
rect 31930 17660 31942 17663
rect 31864 17632 31942 17660
rect 31864 17592 31892 17632
rect 31930 17629 31942 17632
rect 31976 17629 31988 17663
rect 31930 17623 31988 17629
rect 34977 17663 35035 17669
rect 34977 17629 34989 17663
rect 35023 17629 35035 17663
rect 34977 17623 35035 17629
rect 35253 17663 35311 17669
rect 35253 17629 35265 17663
rect 35299 17660 35311 17663
rect 35342 17660 35348 17672
rect 35299 17632 35348 17660
rect 35299 17629 35311 17632
rect 35253 17623 35311 17629
rect 32306 17592 32312 17604
rect 31864 17564 32312 17592
rect 32306 17552 32312 17564
rect 32364 17552 32370 17604
rect 34333 17595 34391 17601
rect 32416 17564 32706 17592
rect 32416 17536 32444 17564
rect 34333 17561 34345 17595
rect 34379 17592 34391 17595
rect 34514 17592 34520 17604
rect 34379 17564 34520 17592
rect 34379 17561 34391 17564
rect 34333 17555 34391 17561
rect 34514 17552 34520 17564
rect 34572 17592 34578 17604
rect 34992 17592 35020 17623
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 35526 17620 35532 17672
rect 35584 17660 35590 17672
rect 35728 17660 35756 17700
rect 36357 17697 36369 17700
rect 36403 17728 36415 17731
rect 37182 17728 37188 17740
rect 36403 17700 37188 17728
rect 36403 17697 36415 17700
rect 36357 17691 36415 17697
rect 37182 17688 37188 17700
rect 37240 17728 37246 17740
rect 38013 17731 38071 17737
rect 38013 17728 38025 17731
rect 37240 17700 38025 17728
rect 37240 17688 37246 17700
rect 38013 17697 38025 17700
rect 38059 17697 38071 17731
rect 39022 17728 39028 17740
rect 38013 17691 38071 17697
rect 38580 17700 39028 17728
rect 36081 17663 36139 17669
rect 36081 17660 36093 17663
rect 35584 17632 35756 17660
rect 36004 17632 36093 17660
rect 35584 17620 35590 17632
rect 36004 17604 36032 17632
rect 36081 17629 36093 17632
rect 36127 17629 36139 17663
rect 36081 17623 36139 17629
rect 36170 17620 36176 17672
rect 36228 17620 36234 17672
rect 37734 17620 37740 17672
rect 37792 17660 37798 17672
rect 38580 17669 38608 17700
rect 39022 17688 39028 17700
rect 39080 17688 39086 17740
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37792 17632 37841 17660
rect 37792 17620 37798 17632
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 38565 17663 38623 17669
rect 38565 17629 38577 17663
rect 38611 17629 38623 17663
rect 38565 17623 38623 17629
rect 38841 17663 38899 17669
rect 38841 17629 38853 17663
rect 38887 17660 38899 17663
rect 39316 17660 39344 17768
rect 39482 17688 39488 17740
rect 39540 17728 39546 17740
rect 39761 17731 39819 17737
rect 39761 17728 39773 17731
rect 39540 17700 39773 17728
rect 39540 17688 39546 17700
rect 39761 17697 39773 17700
rect 39807 17697 39819 17731
rect 39761 17691 39819 17697
rect 40681 17731 40739 17737
rect 40681 17697 40693 17731
rect 40727 17728 40739 17731
rect 41322 17728 41328 17740
rect 40727 17700 41328 17728
rect 40727 17697 40739 17700
rect 40681 17691 40739 17697
rect 41322 17688 41328 17700
rect 41380 17688 41386 17740
rect 42978 17688 42984 17740
rect 43036 17688 43042 17740
rect 43070 17688 43076 17740
rect 43128 17688 43134 17740
rect 38887 17632 39252 17660
rect 39316 17632 40448 17660
rect 38887 17629 38899 17632
rect 38841 17623 38899 17629
rect 35894 17592 35900 17604
rect 34572 17564 34928 17592
rect 34992 17564 35900 17592
rect 34572 17552 34578 17564
rect 32122 17524 32128 17536
rect 31680 17496 32128 17524
rect 32122 17484 32128 17496
rect 32180 17484 32186 17536
rect 32398 17484 32404 17536
rect 32456 17524 32462 17536
rect 33042 17524 33048 17536
rect 32456 17496 33048 17524
rect 32456 17484 32462 17496
rect 33042 17484 33048 17496
rect 33100 17484 33106 17536
rect 34790 17484 34796 17536
rect 34848 17484 34854 17536
rect 34900 17524 34928 17564
rect 35894 17552 35900 17564
rect 35952 17552 35958 17604
rect 35986 17552 35992 17604
rect 36044 17552 36050 17604
rect 36096 17564 36952 17592
rect 35621 17527 35679 17533
rect 35621 17524 35633 17527
rect 34900 17496 35633 17524
rect 35621 17493 35633 17496
rect 35667 17524 35679 17527
rect 36096 17524 36124 17564
rect 36924 17536 36952 17564
rect 37274 17552 37280 17604
rect 37332 17592 37338 17604
rect 37369 17595 37427 17601
rect 37369 17592 37381 17595
rect 37332 17564 37381 17592
rect 37332 17552 37338 17564
rect 37369 17561 37381 17564
rect 37415 17561 37427 17595
rect 37369 17555 37427 17561
rect 35667 17496 36124 17524
rect 35667 17493 35679 17496
rect 35621 17487 35679 17493
rect 36446 17484 36452 17536
rect 36504 17524 36510 17536
rect 36725 17527 36783 17533
rect 36725 17524 36737 17527
rect 36504 17496 36737 17524
rect 36504 17484 36510 17496
rect 36725 17493 36737 17496
rect 36771 17493 36783 17527
rect 36725 17487 36783 17493
rect 36906 17484 36912 17536
rect 36964 17524 36970 17536
rect 37458 17524 37464 17536
rect 36964 17496 37464 17524
rect 36964 17484 36970 17496
rect 37458 17484 37464 17496
rect 37516 17484 37522 17536
rect 38657 17527 38715 17533
rect 38657 17493 38669 17527
rect 38703 17524 38715 17527
rect 39114 17524 39120 17536
rect 38703 17496 39120 17524
rect 38703 17493 38715 17496
rect 38657 17487 38715 17493
rect 39114 17484 39120 17496
rect 39172 17484 39178 17536
rect 39224 17533 39252 17632
rect 39577 17595 39635 17601
rect 39577 17561 39589 17595
rect 39623 17592 39635 17595
rect 39623 17564 40080 17592
rect 39623 17561 39635 17564
rect 39577 17555 39635 17561
rect 40052 17536 40080 17564
rect 40126 17552 40132 17604
rect 40184 17592 40190 17604
rect 40221 17595 40279 17601
rect 40221 17592 40233 17595
rect 40184 17564 40233 17592
rect 40184 17552 40190 17564
rect 40221 17561 40233 17564
rect 40267 17561 40279 17595
rect 40221 17555 40279 17561
rect 39209 17527 39267 17533
rect 39209 17493 39221 17527
rect 39255 17493 39267 17527
rect 39209 17487 39267 17493
rect 39390 17484 39396 17536
rect 39448 17524 39454 17536
rect 39669 17527 39727 17533
rect 39669 17524 39681 17527
rect 39448 17496 39681 17524
rect 39448 17484 39454 17496
rect 39669 17493 39681 17496
rect 39715 17493 39727 17527
rect 39669 17487 39727 17493
rect 40034 17484 40040 17536
rect 40092 17484 40098 17536
rect 40420 17524 40448 17632
rect 40586 17620 40592 17672
rect 40644 17620 40650 17672
rect 42889 17663 42947 17669
rect 42889 17629 42901 17663
rect 42935 17660 42947 17663
rect 43254 17660 43260 17672
rect 42935 17632 43260 17660
rect 42935 17629 42947 17632
rect 42889 17623 42947 17629
rect 43254 17620 43260 17632
rect 43312 17620 43318 17672
rect 40604 17592 40632 17620
rect 40957 17595 41015 17601
rect 40957 17592 40969 17595
rect 40604 17564 40969 17592
rect 40957 17561 40969 17564
rect 41003 17561 41015 17595
rect 40957 17555 41015 17561
rect 41414 17552 41420 17604
rect 41472 17552 41478 17604
rect 42426 17552 42432 17604
rect 42484 17592 42490 17604
rect 42484 17564 44588 17592
rect 42484 17552 42490 17564
rect 42521 17527 42579 17533
rect 42521 17524 42533 17527
rect 40420 17496 42533 17524
rect 42521 17493 42533 17496
rect 42567 17493 42579 17527
rect 42521 17487 42579 17493
rect 43530 17484 43536 17536
rect 43588 17524 43594 17536
rect 43898 17524 43904 17536
rect 43588 17496 43904 17524
rect 43588 17484 43594 17496
rect 43898 17484 43904 17496
rect 43956 17484 43962 17536
rect 44560 17533 44588 17564
rect 44545 17527 44603 17533
rect 44545 17493 44557 17527
rect 44591 17493 44603 17527
rect 44545 17487 44603 17493
rect 44910 17484 44916 17536
rect 44968 17484 44974 17536
rect 460 17434 45540 17456
rect 460 17382 6070 17434
rect 6122 17382 6134 17434
rect 6186 17382 6198 17434
rect 6250 17382 6262 17434
rect 6314 17382 6326 17434
rect 6378 17382 11070 17434
rect 11122 17382 11134 17434
rect 11186 17382 11198 17434
rect 11250 17382 11262 17434
rect 11314 17382 11326 17434
rect 11378 17382 16070 17434
rect 16122 17382 16134 17434
rect 16186 17382 16198 17434
rect 16250 17382 16262 17434
rect 16314 17382 16326 17434
rect 16378 17382 21070 17434
rect 21122 17382 21134 17434
rect 21186 17382 21198 17434
rect 21250 17382 21262 17434
rect 21314 17382 21326 17434
rect 21378 17382 26070 17434
rect 26122 17382 26134 17434
rect 26186 17382 26198 17434
rect 26250 17382 26262 17434
rect 26314 17382 26326 17434
rect 26378 17382 31070 17434
rect 31122 17382 31134 17434
rect 31186 17382 31198 17434
rect 31250 17382 31262 17434
rect 31314 17382 31326 17434
rect 31378 17382 36070 17434
rect 36122 17382 36134 17434
rect 36186 17382 36198 17434
rect 36250 17382 36262 17434
rect 36314 17382 36326 17434
rect 36378 17382 41070 17434
rect 41122 17382 41134 17434
rect 41186 17382 41198 17434
rect 41250 17382 41262 17434
rect 41314 17382 41326 17434
rect 41378 17382 45540 17434
rect 460 17360 45540 17382
rect 5537 17323 5595 17329
rect 5537 17289 5549 17323
rect 5583 17320 5595 17323
rect 5626 17320 5632 17332
rect 5583 17292 5632 17320
rect 5583 17289 5595 17292
rect 5537 17283 5595 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6546 17320 6552 17332
rect 6227 17292 6552 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 6696 17292 7021 17320
rect 6696 17280 6702 17292
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 7009 17283 7067 17289
rect 7558 17280 7564 17332
rect 7616 17320 7622 17332
rect 7653 17323 7711 17329
rect 7653 17320 7665 17323
rect 7616 17292 7665 17320
rect 7616 17280 7622 17292
rect 7653 17289 7665 17292
rect 7699 17289 7711 17323
rect 7653 17283 7711 17289
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 8076 17292 8125 17320
rect 8076 17280 8082 17292
rect 8113 17289 8125 17292
rect 8159 17289 8171 17323
rect 8113 17283 8171 17289
rect 8846 17280 8852 17332
rect 8904 17280 8910 17332
rect 9766 17280 9772 17332
rect 9824 17280 9830 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17289 9919 17323
rect 9861 17283 9919 17289
rect 3697 17255 3755 17261
rect 3697 17221 3709 17255
rect 3743 17252 3755 17255
rect 4522 17252 4528 17264
rect 3743 17224 4528 17252
rect 3743 17221 3755 17224
rect 3697 17215 3755 17221
rect 4522 17212 4528 17224
rect 4580 17212 4586 17264
rect 4614 17212 4620 17264
rect 4672 17212 4678 17264
rect 5644 17252 5672 17280
rect 5644 17224 6040 17252
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5500 17156 5733 17184
rect 5500 17144 5506 17156
rect 5721 17153 5733 17156
rect 5767 17184 5779 17187
rect 5902 17184 5908 17196
rect 5767 17156 5908 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 6012 17193 6040 17224
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 7852 17184 7880 17280
rect 7423 17156 7880 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3789 17119 3847 17125
rect 3789 17116 3801 17119
rect 3384 17088 3801 17116
rect 3384 17076 3390 17088
rect 3789 17085 3801 17088
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 5460 17116 5488 17144
rect 4212 17088 5488 17116
rect 4212 17076 4218 17088
rect 5810 17076 5816 17128
rect 5868 17076 5874 17128
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7116 17116 7144 17147
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7064 17088 7481 17116
rect 7064 17076 7070 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 7469 17079 7527 17085
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 8864 17116 8892 17280
rect 9876 17252 9904 17283
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 12860 17292 13032 17320
rect 12860 17280 12866 17292
rect 13004 17261 13032 17292
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 13412 17292 14473 17320
rect 13412 17280 13418 17292
rect 14461 17289 14473 17292
rect 14507 17320 14519 17323
rect 15039 17323 15097 17329
rect 14507 17292 14964 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 11149 17255 11207 17261
rect 11149 17252 11161 17255
rect 9876 17224 11161 17252
rect 11149 17221 11161 17224
rect 11195 17221 11207 17255
rect 11149 17215 11207 17221
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17221 13047 17255
rect 12989 17215 13047 17221
rect 14826 17212 14832 17264
rect 14884 17212 14890 17264
rect 14936 17252 14964 17292
rect 15039 17289 15051 17323
rect 15085 17320 15097 17323
rect 15194 17320 15200 17332
rect 15085 17292 15200 17320
rect 15085 17289 15097 17292
rect 15039 17283 15097 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16577 17323 16635 17329
rect 15795 17292 16528 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 16500 17252 16528 17292
rect 16577 17289 16589 17323
rect 16623 17320 16635 17323
rect 16666 17320 16672 17332
rect 16623 17292 16672 17320
rect 16623 17289 16635 17292
rect 16577 17283 16635 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17092 17292 18736 17320
rect 17092 17280 17098 17292
rect 18708 17261 18736 17292
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19518 17320 19524 17332
rect 19076 17292 19524 17320
rect 18693 17255 18751 17261
rect 14936 17224 15884 17252
rect 16500 17224 18644 17252
rect 15856 17196 15884 17224
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17184 9091 17187
rect 9674 17184 9680 17196
rect 9079 17156 9680 17184
rect 9079 17153 9091 17156
rect 9033 17147 9091 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 7699 17088 8892 17116
rect 9048 17088 9137 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 9048 16992 9076 17088
rect 9125 17085 9137 17088
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 9950 17116 9956 17128
rect 9355 17088 9956 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10060 17116 10088 17147
rect 10318 17144 10324 17196
rect 10376 17144 10382 17196
rect 10686 17144 10692 17196
rect 10744 17144 10750 17196
rect 10778 17144 10784 17196
rect 10836 17144 10842 17196
rect 10870 17144 10876 17196
rect 10928 17144 10934 17196
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 14274 17184 14280 17196
rect 14122 17156 14280 17184
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 10796 17116 10824 17144
rect 10060 17088 10824 17116
rect 10888 17116 10916 17144
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 10888 17088 12725 17116
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 15304 17116 15332 17147
rect 15562 17144 15568 17196
rect 15620 17193 15626 17196
rect 15620 17184 15629 17193
rect 15620 17156 15665 17184
rect 15620 17147 15629 17156
rect 15620 17144 15626 17147
rect 15838 17144 15844 17196
rect 15896 17144 15902 17196
rect 16393 17187 16451 17193
rect 16393 17153 16405 17187
rect 16439 17184 16451 17187
rect 16574 17184 16580 17196
rect 16439 17156 16580 17184
rect 16439 17153 16451 17156
rect 16393 17147 16451 17153
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 16942 17184 16948 17196
rect 16899 17156 16948 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17236 17193 17264 17224
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 17267 17156 17301 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 16298 17116 16304 17128
rect 15304 17088 16304 17116
rect 12713 17079 12771 17085
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16408 17088 16681 17116
rect 16408 17060 16436 17088
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 15197 17051 15255 17057
rect 15197 17017 15209 17051
rect 15243 17048 15255 17051
rect 15286 17048 15292 17060
rect 15243 17020 15292 17048
rect 15243 17017 15255 17020
rect 15197 17011 15255 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 15562 17008 15568 17060
rect 15620 17048 15626 17060
rect 15620 17020 16252 17048
rect 15620 17008 15626 17020
rect 5718 16940 5724 16992
rect 5776 16940 5782 16992
rect 6822 16940 6828 16992
rect 6880 16940 6886 16992
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 8168 16952 8493 16980
rect 8168 16940 8174 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 8481 16943 8539 16949
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 8665 16983 8723 16989
rect 8665 16980 8677 16983
rect 8628 16952 8677 16980
rect 8628 16940 8634 16952
rect 8665 16949 8677 16952
rect 8711 16949 8723 16983
rect 8665 16943 8723 16949
rect 9030 16940 9036 16992
rect 9088 16940 9094 16992
rect 10042 16940 10048 16992
rect 10100 16980 10106 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 10100 16952 10149 16980
rect 10100 16940 10106 16952
rect 10137 16949 10149 16952
rect 10183 16949 10195 16983
rect 10137 16943 10195 16949
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10778 16980 10784 16992
rect 10551 16952 10784 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12621 16983 12679 16989
rect 12621 16980 12633 16983
rect 12492 16952 12633 16980
rect 12492 16940 12498 16952
rect 12621 16949 12633 16952
rect 12667 16949 12679 16983
rect 12621 16943 12679 16949
rect 15010 16940 15016 16992
rect 15068 16940 15074 16992
rect 15381 16983 15439 16989
rect 15381 16949 15393 16983
rect 15427 16980 15439 16983
rect 15470 16980 15476 16992
rect 15427 16952 15476 16980
rect 15427 16949 15439 16952
rect 15381 16943 15439 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 15988 16952 16129 16980
rect 15988 16940 15994 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16224 16980 16252 17020
rect 16390 17008 16396 17060
rect 16448 17008 16454 17060
rect 16684 17048 16712 17079
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 17144 17116 17172 17147
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 17862 17184 17868 17196
rect 17727 17156 17868 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 18288 17156 18337 17184
rect 18288 17144 18294 17156
rect 18325 17153 18337 17156
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17153 18567 17187
rect 18509 17147 18567 17153
rect 17880 17116 17908 17144
rect 18524 17116 18552 17147
rect 17144 17088 17724 17116
rect 17880 17088 18552 17116
rect 18616 17116 18644 17224
rect 18693 17221 18705 17255
rect 18739 17221 18751 17255
rect 18693 17215 18751 17221
rect 18892 17184 18920 17280
rect 19076 17261 19104 17292
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 19978 17320 19984 17332
rect 19812 17292 19984 17320
rect 19061 17255 19119 17261
rect 19061 17221 19073 17255
rect 19107 17221 19119 17255
rect 19061 17215 19119 17221
rect 19153 17255 19211 17261
rect 19153 17221 19165 17255
rect 19199 17252 19211 17255
rect 19426 17252 19432 17264
rect 19199 17224 19432 17252
rect 19199 17221 19211 17224
rect 19153 17215 19211 17221
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 19812 17261 19840 17292
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 20438 17280 20444 17332
rect 20496 17280 20502 17332
rect 20622 17280 20628 17332
rect 20680 17280 20686 17332
rect 22370 17280 22376 17332
rect 22428 17280 22434 17332
rect 22554 17280 22560 17332
rect 22612 17320 22618 17332
rect 22612 17292 22876 17320
rect 22612 17280 22618 17292
rect 19797 17255 19855 17261
rect 19797 17221 19809 17255
rect 19843 17221 19855 17255
rect 20272 17252 20300 17280
rect 19797 17215 19855 17221
rect 18969 17187 19027 17193
rect 18969 17184 18981 17187
rect 18892 17156 18981 17184
rect 18969 17153 18981 17156
rect 19015 17153 19027 17187
rect 19271 17187 19329 17193
rect 19271 17184 19283 17187
rect 18969 17147 19027 17153
rect 19076 17156 19283 17184
rect 19076 17116 19104 17156
rect 19271 17153 19283 17156
rect 19317 17184 19329 17187
rect 19317 17156 19564 17184
rect 19317 17153 19329 17156
rect 19271 17147 19329 17153
rect 18616 17088 19104 17116
rect 19429 17119 19487 17125
rect 17126 17048 17132 17060
rect 16684 17020 17132 17048
rect 17126 17008 17132 17020
rect 17184 17008 17190 17060
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 17236 17020 17509 17048
rect 17236 16980 17264 17020
rect 17497 17017 17509 17020
rect 17543 17017 17555 17051
rect 17497 17011 17555 17017
rect 17696 16992 17724 17088
rect 19429 17085 19441 17119
rect 19475 17085 19487 17119
rect 19536 17116 19564 17156
rect 19702 17144 19708 17196
rect 19760 17144 19766 17196
rect 19886 17178 19892 17230
rect 19944 17178 19950 17230
rect 20042 17224 20300 17252
rect 20042 17193 20070 17224
rect 20027 17187 20085 17193
rect 19890 17153 19902 17178
rect 19936 17153 19948 17178
rect 19890 17147 19948 17153
rect 20027 17153 20039 17187
rect 20073 17153 20085 17187
rect 20027 17147 20085 17153
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 20042 17116 20070 17147
rect 19536 17088 20070 17116
rect 19429 17079 19487 17085
rect 18414 17008 18420 17060
rect 18472 17048 18478 17060
rect 18785 17051 18843 17057
rect 18785 17048 18797 17051
rect 18472 17020 18797 17048
rect 18472 17008 18478 17020
rect 18785 17017 18797 17020
rect 18831 17017 18843 17051
rect 18785 17011 18843 17017
rect 19334 17008 19340 17060
rect 19392 17048 19398 17060
rect 19444 17048 19472 17079
rect 20162 17076 20168 17128
rect 20220 17076 20226 17128
rect 20272 17116 20300 17147
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 20990 17184 20996 17196
rect 20404 17156 20996 17184
rect 20404 17144 20410 17156
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 22388 17184 22416 17280
rect 22848 17261 22876 17292
rect 24302 17280 24308 17332
rect 24360 17280 24366 17332
rect 24946 17280 24952 17332
rect 25004 17320 25010 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 25004 17292 25053 17320
rect 25004 17280 25010 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 25406 17280 25412 17332
rect 25464 17280 25470 17332
rect 27890 17280 27896 17332
rect 27948 17280 27954 17332
rect 28000 17292 28580 17320
rect 22833 17255 22891 17261
rect 22833 17221 22845 17255
rect 22879 17221 22891 17255
rect 24210 17252 24216 17264
rect 24058 17224 24216 17252
rect 22833 17215 22891 17221
rect 24210 17212 24216 17224
rect 24268 17212 24274 17264
rect 24320 17252 24348 17280
rect 25501 17255 25559 17261
rect 25501 17252 25513 17255
rect 24320 17224 25513 17252
rect 25501 17221 25513 17224
rect 25547 17221 25559 17255
rect 25501 17215 25559 17221
rect 26418 17212 26424 17264
rect 26476 17252 26482 17264
rect 26758 17255 26816 17261
rect 26758 17252 26770 17255
rect 26476 17224 26770 17252
rect 26476 17212 26482 17224
rect 26758 17221 26770 17224
rect 26804 17221 26816 17255
rect 26758 17215 26816 17221
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 22388 17156 22569 17184
rect 22557 17153 22569 17156
rect 22603 17153 22615 17187
rect 22557 17147 22615 17153
rect 24394 17144 24400 17196
rect 24452 17144 24458 17196
rect 24946 17144 24952 17196
rect 25004 17144 25010 17196
rect 28000 17193 28028 17292
rect 28552 17264 28580 17292
rect 28994 17280 29000 17332
rect 29052 17280 29058 17332
rect 29457 17323 29515 17329
rect 29457 17289 29469 17323
rect 29503 17320 29515 17323
rect 29546 17320 29552 17332
rect 29503 17292 29552 17320
rect 29503 17289 29515 17292
rect 29457 17283 29515 17289
rect 29546 17280 29552 17292
rect 29604 17320 29610 17332
rect 30374 17320 30380 17332
rect 29604 17292 30380 17320
rect 29604 17280 29610 17292
rect 30374 17280 30380 17292
rect 30432 17280 30438 17332
rect 30466 17280 30472 17332
rect 30524 17320 30530 17332
rect 30834 17320 30840 17332
rect 30524 17292 30840 17320
rect 30524 17280 30530 17292
rect 30834 17280 30840 17292
rect 30892 17320 30898 17332
rect 31297 17323 31355 17329
rect 30892 17292 30972 17320
rect 30892 17280 30898 17292
rect 28350 17212 28356 17264
rect 28408 17252 28414 17264
rect 28408 17224 28488 17252
rect 28408 17212 28414 17224
rect 28258 17193 28264 17196
rect 27985 17187 28043 17193
rect 27985 17184 27997 17187
rect 27586 17156 27997 17184
rect 20272 17088 20392 17116
rect 20364 17060 20392 17088
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 20625 17119 20683 17125
rect 20625 17116 20637 17119
rect 20588 17088 20637 17116
rect 20588 17076 20594 17088
rect 20625 17085 20637 17088
rect 20671 17085 20683 17119
rect 20625 17079 20683 17085
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25593 17119 25651 17125
rect 25593 17116 25605 17119
rect 25280 17088 25605 17116
rect 25280 17076 25286 17088
rect 25593 17085 25605 17088
rect 25639 17085 25651 17119
rect 25593 17079 25651 17085
rect 26145 17119 26203 17125
rect 26145 17085 26157 17119
rect 26191 17116 26203 17119
rect 26513 17119 26571 17125
rect 26513 17116 26525 17119
rect 26191 17088 26525 17116
rect 26191 17085 26203 17088
rect 26145 17079 26203 17085
rect 26513 17085 26525 17088
rect 26559 17085 26571 17119
rect 26513 17079 26571 17085
rect 19392 17020 19472 17048
rect 19392 17008 19398 17020
rect 20346 17008 20352 17060
rect 20404 17008 20410 17060
rect 20898 17008 20904 17060
rect 20956 17008 20962 17060
rect 22005 17051 22063 17057
rect 22005 17048 22017 17051
rect 21652 17020 22017 17048
rect 21652 16992 21680 17020
rect 22005 17017 22017 17020
rect 22051 17048 22063 17051
rect 22278 17048 22284 17060
rect 22051 17020 22284 17048
rect 22051 17017 22063 17020
rect 22005 17011 22063 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 16224 16952 17264 16980
rect 16117 16943 16175 16949
rect 17402 16940 17408 16992
rect 17460 16940 17466 16992
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16980 18291 16983
rect 18322 16980 18328 16992
rect 18279 16952 18328 16980
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 19518 16940 19524 16992
rect 19576 16940 19582 16992
rect 21634 16940 21640 16992
rect 21692 16940 21698 16992
rect 21729 16983 21787 16989
rect 21729 16949 21741 16983
rect 21775 16980 21787 16983
rect 22370 16980 22376 16992
rect 21775 16952 22376 16980
rect 21775 16949 21787 16952
rect 21729 16943 21787 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23934 16940 23940 16992
rect 23992 16980 23998 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 23992 16952 24593 16980
rect 23992 16940 23998 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 24762 16940 24768 16992
rect 24820 16940 24826 16992
rect 26528 16980 26556 17079
rect 26786 16980 26792 16992
rect 26528 16952 26792 16980
rect 26786 16940 26792 16952
rect 26844 16980 26850 16992
rect 27586 16980 27614 17156
rect 27985 17153 27997 17156
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28252 17147 28264 17193
rect 28258 17144 28264 17147
rect 28316 17144 28322 17196
rect 28460 17184 28488 17224
rect 28534 17212 28540 17264
rect 28592 17212 28598 17264
rect 29012 17252 29040 17280
rect 30944 17261 30972 17292
rect 31297 17289 31309 17323
rect 31343 17320 31355 17323
rect 31754 17320 31760 17332
rect 31343 17292 31760 17320
rect 31343 17289 31355 17292
rect 31297 17283 31355 17289
rect 31754 17280 31760 17292
rect 31812 17280 31818 17332
rect 31849 17323 31907 17329
rect 31849 17289 31861 17323
rect 31895 17289 31907 17323
rect 31849 17283 31907 17289
rect 30929 17255 30987 17261
rect 29012 17224 29960 17252
rect 28460 17156 29040 17184
rect 29012 17116 29040 17156
rect 29270 17144 29276 17196
rect 29328 17184 29334 17196
rect 29932 17193 29960 17224
rect 30116 17224 30880 17252
rect 30116 17193 30144 17224
rect 29687 17187 29745 17193
rect 29687 17184 29699 17187
rect 29328 17156 29699 17184
rect 29328 17144 29334 17156
rect 29687 17153 29699 17156
rect 29733 17153 29745 17187
rect 29687 17147 29745 17153
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17153 29883 17187
rect 29825 17147 29883 17153
rect 29922 17187 29980 17193
rect 29922 17153 29934 17187
rect 29968 17153 29980 17187
rect 29922 17147 29980 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17153 30159 17187
rect 30101 17147 30159 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 29837 17116 29865 17147
rect 29012 17088 29865 17116
rect 29288 17020 29868 17048
rect 29288 16992 29316 17020
rect 26844 16952 27614 16980
rect 26844 16940 26850 16952
rect 28718 16940 28724 16992
rect 28776 16980 28782 16992
rect 28994 16980 29000 16992
rect 28776 16952 29000 16980
rect 28776 16940 28782 16952
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 29270 16940 29276 16992
rect 29328 16940 29334 16992
rect 29362 16940 29368 16992
rect 29420 16940 29426 16992
rect 29840 16980 29868 17020
rect 29914 17008 29920 17060
rect 29972 17048 29978 17060
rect 30193 17051 30251 17057
rect 30193 17048 30205 17051
rect 29972 17020 30205 17048
rect 29972 17008 29978 17020
rect 30193 17017 30205 17020
rect 30239 17017 30251 17051
rect 30193 17011 30251 17017
rect 30484 16980 30512 17147
rect 30558 17144 30564 17196
rect 30616 17144 30622 17196
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 30852 17193 30880 17224
rect 30929 17221 30941 17255
rect 30975 17221 30987 17255
rect 30929 17215 30987 17221
rect 31129 17255 31187 17261
rect 31129 17221 31141 17255
rect 31175 17221 31187 17255
rect 31129 17215 31187 17221
rect 31573 17255 31631 17261
rect 31573 17221 31585 17255
rect 31619 17252 31631 17255
rect 31864 17252 31892 17283
rect 32030 17280 32036 17332
rect 32088 17320 32094 17332
rect 32306 17320 32312 17332
rect 32088 17292 32312 17320
rect 32088 17280 32094 17292
rect 32306 17280 32312 17292
rect 32364 17320 32370 17332
rect 32364 17292 32812 17320
rect 32364 17280 32370 17292
rect 31619 17224 31892 17252
rect 32217 17255 32275 17261
rect 31619 17221 31631 17224
rect 31573 17215 31631 17221
rect 32217 17221 32229 17255
rect 32263 17252 32275 17255
rect 32582 17252 32588 17264
rect 32263 17224 32588 17252
rect 32263 17221 32275 17224
rect 32217 17215 32275 17221
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 30852 17116 30880 17147
rect 30576 17088 30880 17116
rect 30944 17116 30972 17215
rect 31018 17144 31024 17196
rect 31076 17184 31082 17196
rect 31144 17184 31172 17215
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 32674 17212 32680 17264
rect 32732 17212 32738 17264
rect 32784 17252 32812 17292
rect 32858 17280 32864 17332
rect 32916 17329 32922 17332
rect 32916 17323 32935 17329
rect 32923 17289 32935 17323
rect 32916 17283 32935 17289
rect 32916 17280 32922 17283
rect 33134 17280 33140 17332
rect 33192 17320 33198 17332
rect 33778 17320 33784 17332
rect 33192 17292 33784 17320
rect 33192 17280 33198 17292
rect 33778 17280 33784 17292
rect 33836 17280 33842 17332
rect 34514 17280 34520 17332
rect 34572 17280 34578 17332
rect 34790 17320 34796 17332
rect 34716 17292 34796 17320
rect 34532 17252 34560 17280
rect 34716 17261 34744 17292
rect 34790 17280 34796 17292
rect 34848 17280 34854 17332
rect 34882 17280 34888 17332
rect 34940 17280 34946 17332
rect 39022 17280 39028 17332
rect 39080 17320 39086 17332
rect 41233 17323 41291 17329
rect 39080 17292 41092 17320
rect 39080 17280 39086 17292
rect 32784 17224 34100 17252
rect 31076 17156 31172 17184
rect 31076 17144 31082 17156
rect 31754 17144 31760 17196
rect 31812 17144 31818 17196
rect 31846 17144 31852 17196
rect 31904 17144 31910 17196
rect 31864 17116 31892 17144
rect 32306 17116 32312 17128
rect 30944 17088 31800 17116
rect 31864 17088 32312 17116
rect 30576 17060 30604 17088
rect 30558 17008 30564 17060
rect 30616 17008 30622 17060
rect 31772 17048 31800 17088
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 32490 17076 32496 17128
rect 32548 17076 32554 17128
rect 32692 17048 32720 17212
rect 34072 17196 34100 17224
rect 34440 17224 34560 17252
rect 34701 17255 34759 17261
rect 32766 17144 32772 17196
rect 32824 17144 32830 17196
rect 34054 17144 34060 17196
rect 34112 17184 34118 17196
rect 34440 17193 34468 17224
rect 34701 17221 34713 17255
rect 34747 17221 34759 17255
rect 34900 17252 34928 17280
rect 34900 17224 35190 17252
rect 34701 17215 34759 17221
rect 38194 17212 38200 17264
rect 38252 17212 38258 17264
rect 38930 17212 38936 17264
rect 38988 17212 38994 17264
rect 40034 17212 40040 17264
rect 40092 17252 40098 17264
rect 41064 17252 41092 17292
rect 41233 17289 41245 17323
rect 41279 17320 41291 17323
rect 41506 17320 41512 17332
rect 41279 17292 41512 17320
rect 41279 17289 41291 17292
rect 41233 17283 41291 17289
rect 41506 17280 41512 17292
rect 41564 17280 41570 17332
rect 42794 17280 42800 17332
rect 42852 17320 42858 17332
rect 43162 17320 43168 17332
rect 42852 17292 43168 17320
rect 42852 17280 42858 17292
rect 43162 17280 43168 17292
rect 43220 17320 43226 17332
rect 43898 17320 43904 17332
rect 43220 17292 43904 17320
rect 43220 17280 43226 17292
rect 43898 17280 43904 17292
rect 43956 17320 43962 17332
rect 44269 17323 44327 17329
rect 44269 17320 44281 17323
rect 43956 17292 44281 17320
rect 43956 17280 43962 17292
rect 44269 17289 44281 17292
rect 44315 17320 44327 17323
rect 45005 17323 45063 17329
rect 45005 17320 45017 17323
rect 44315 17292 45017 17320
rect 44315 17289 44327 17292
rect 44269 17283 44327 17289
rect 45005 17289 45017 17292
rect 45051 17289 45063 17323
rect 45005 17283 45063 17289
rect 42426 17252 42432 17264
rect 40092 17224 41000 17252
rect 41064 17224 42432 17252
rect 40092 17212 40098 17224
rect 40972 17196 41000 17224
rect 42426 17212 42432 17224
rect 42484 17212 42490 17264
rect 34149 17187 34207 17193
rect 34149 17184 34161 17187
rect 34112 17156 34161 17184
rect 34112 17144 34118 17156
rect 34149 17153 34161 17156
rect 34195 17184 34207 17187
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34195 17156 34437 17184
rect 34195 17153 34207 17156
rect 34149 17147 34207 17153
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34425 17147 34483 17153
rect 36814 17144 36820 17196
rect 36872 17144 36878 17196
rect 37458 17144 37464 17196
rect 37516 17184 37522 17196
rect 37921 17187 37979 17193
rect 37921 17184 37933 17187
rect 37516 17156 37933 17184
rect 37516 17144 37522 17156
rect 37921 17153 37933 17156
rect 37967 17153 37979 17187
rect 37921 17147 37979 17153
rect 39574 17144 39580 17196
rect 39632 17184 39638 17196
rect 39945 17187 40003 17193
rect 39945 17184 39957 17187
rect 39632 17156 39957 17184
rect 39632 17144 39638 17156
rect 39945 17153 39957 17156
rect 39991 17153 40003 17187
rect 39945 17147 40003 17153
rect 40126 17144 40132 17196
rect 40184 17144 40190 17196
rect 40773 17187 40831 17193
rect 40773 17153 40785 17187
rect 40819 17184 40831 17187
rect 40819 17156 40908 17184
rect 40819 17153 40831 17156
rect 40773 17147 40831 17153
rect 31772 17020 32720 17048
rect 32784 17048 32812 17144
rect 37292 17088 39896 17116
rect 37292 17060 37320 17088
rect 33045 17051 33103 17057
rect 33045 17048 33057 17051
rect 32784 17020 33057 17048
rect 33045 17017 33057 17020
rect 33091 17017 33103 17051
rect 33045 17011 33103 17017
rect 37274 17008 37280 17060
rect 37332 17008 37338 17060
rect 39758 17008 39764 17060
rect 39816 17008 39822 17060
rect 39868 17048 39896 17088
rect 40880 17057 40908 17156
rect 40954 17144 40960 17196
rect 41012 17144 41018 17196
rect 41325 17187 41383 17193
rect 41325 17153 41337 17187
rect 41371 17184 41383 17187
rect 41598 17184 41604 17196
rect 41371 17156 41604 17184
rect 41371 17153 41383 17156
rect 41325 17147 41383 17153
rect 41598 17144 41604 17156
rect 41656 17184 41662 17196
rect 42153 17187 42211 17193
rect 42153 17184 42165 17187
rect 41656 17156 42165 17184
rect 41656 17144 41662 17156
rect 42153 17153 42165 17156
rect 42199 17153 42211 17187
rect 42153 17147 42211 17153
rect 42245 17187 42303 17193
rect 42245 17153 42257 17187
rect 42291 17184 42303 17187
rect 43346 17184 43352 17196
rect 42291 17156 43352 17184
rect 42291 17153 42303 17156
rect 42245 17147 42303 17153
rect 43346 17144 43352 17156
rect 43404 17144 43410 17196
rect 44910 17144 44916 17196
rect 44968 17144 44974 17196
rect 41046 17076 41052 17128
rect 41104 17116 41110 17128
rect 41417 17119 41475 17125
rect 41417 17116 41429 17119
rect 41104 17088 41429 17116
rect 41104 17076 41110 17088
rect 41417 17085 41429 17088
rect 41463 17116 41475 17119
rect 41506 17116 41512 17128
rect 41463 17088 41512 17116
rect 41463 17085 41475 17088
rect 41417 17079 41475 17085
rect 41506 17076 41512 17088
rect 41564 17076 41570 17128
rect 41874 17076 41880 17128
rect 41932 17116 41938 17128
rect 42337 17119 42395 17125
rect 42337 17116 42349 17119
rect 41932 17088 42349 17116
rect 41932 17076 41938 17088
rect 42337 17085 42349 17088
rect 42383 17085 42395 17119
rect 42337 17079 42395 17085
rect 40865 17051 40923 17057
rect 39868 17020 40816 17048
rect 29840 16952 30512 16980
rect 31110 16940 31116 16992
rect 31168 16980 31174 16992
rect 32861 16983 32919 16989
rect 32861 16980 32873 16983
rect 31168 16952 32873 16980
rect 31168 16940 31174 16952
rect 32861 16949 32873 16952
rect 32907 16980 32919 16983
rect 33226 16980 33232 16992
rect 32907 16952 33232 16980
rect 32907 16949 32919 16952
rect 32861 16943 32919 16949
rect 33226 16940 33232 16952
rect 33284 16940 33290 16992
rect 33413 16983 33471 16989
rect 33413 16949 33425 16983
rect 33459 16980 33471 16983
rect 34514 16980 34520 16992
rect 33459 16952 34520 16980
rect 33459 16949 33471 16952
rect 33413 16943 33471 16949
rect 34514 16940 34520 16952
rect 34572 16940 34578 16992
rect 36170 16940 36176 16992
rect 36228 16940 36234 16992
rect 36630 16940 36636 16992
rect 36688 16940 36694 16992
rect 37182 16940 37188 16992
rect 37240 16940 37246 16992
rect 37458 16940 37464 16992
rect 37516 16940 37522 16992
rect 38930 16940 38936 16992
rect 38988 16980 38994 16992
rect 39574 16980 39580 16992
rect 38988 16952 39580 16980
rect 38988 16940 38994 16952
rect 39574 16940 39580 16952
rect 39632 16980 39638 16992
rect 39669 16983 39727 16989
rect 39669 16980 39681 16983
rect 39632 16952 39681 16980
rect 39632 16940 39638 16952
rect 39669 16949 39681 16952
rect 39715 16949 39727 16983
rect 39669 16943 39727 16949
rect 39850 16940 39856 16992
rect 39908 16980 39914 16992
rect 40313 16983 40371 16989
rect 40313 16980 40325 16983
rect 39908 16952 40325 16980
rect 39908 16940 39914 16952
rect 40313 16949 40325 16952
rect 40359 16949 40371 16983
rect 40313 16943 40371 16949
rect 40586 16940 40592 16992
rect 40644 16940 40650 16992
rect 40788 16980 40816 17020
rect 40865 17017 40877 17051
rect 40911 17017 40923 17051
rect 44928 17048 44956 17144
rect 40865 17011 40923 17017
rect 41386 17020 44956 17048
rect 41386 16980 41414 17020
rect 40788 16952 41414 16980
rect 41782 16940 41788 16992
rect 41840 16940 41846 16992
rect 42794 16940 42800 16992
rect 42852 16980 42858 16992
rect 43165 16983 43223 16989
rect 43165 16980 43177 16983
rect 42852 16952 43177 16980
rect 42852 16940 42858 16952
rect 43165 16949 43177 16952
rect 43211 16980 43223 16983
rect 43530 16980 43536 16992
rect 43211 16952 43536 16980
rect 43211 16949 43223 16952
rect 43165 16943 43223 16949
rect 43530 16940 43536 16952
rect 43588 16980 43594 16992
rect 44634 16980 44640 16992
rect 43588 16952 44640 16980
rect 43588 16940 43594 16952
rect 44634 16940 44640 16952
rect 44692 16940 44698 16992
rect 460 16890 45540 16912
rect 460 16838 3570 16890
rect 3622 16838 3634 16890
rect 3686 16838 3698 16890
rect 3750 16838 3762 16890
rect 3814 16838 3826 16890
rect 3878 16838 8570 16890
rect 8622 16838 8634 16890
rect 8686 16838 8698 16890
rect 8750 16838 8762 16890
rect 8814 16838 8826 16890
rect 8878 16838 13570 16890
rect 13622 16838 13634 16890
rect 13686 16838 13698 16890
rect 13750 16838 13762 16890
rect 13814 16838 13826 16890
rect 13878 16838 18570 16890
rect 18622 16838 18634 16890
rect 18686 16838 18698 16890
rect 18750 16838 18762 16890
rect 18814 16838 18826 16890
rect 18878 16838 23570 16890
rect 23622 16838 23634 16890
rect 23686 16838 23698 16890
rect 23750 16838 23762 16890
rect 23814 16838 23826 16890
rect 23878 16838 28570 16890
rect 28622 16838 28634 16890
rect 28686 16838 28698 16890
rect 28750 16838 28762 16890
rect 28814 16838 28826 16890
rect 28878 16838 33570 16890
rect 33622 16838 33634 16890
rect 33686 16838 33698 16890
rect 33750 16838 33762 16890
rect 33814 16838 33826 16890
rect 33878 16838 38570 16890
rect 38622 16838 38634 16890
rect 38686 16838 38698 16890
rect 38750 16838 38762 16890
rect 38814 16838 38826 16890
rect 38878 16838 43570 16890
rect 43622 16838 43634 16890
rect 43686 16838 43698 16890
rect 43750 16838 43762 16890
rect 43814 16838 43826 16890
rect 43878 16838 45540 16890
rect 460 16816 45540 16838
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 8018 16776 8024 16788
rect 7432 16748 8024 16776
rect 7432 16736 7438 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9950 16776 9956 16788
rect 9784 16748 9956 16776
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4672 16612 4721 16640
rect 4672 16600 4678 16612
rect 4709 16609 4721 16612
rect 4755 16640 4767 16643
rect 4755 16612 6224 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 4430 16572 4436 16584
rect 4264 16544 4436 16572
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 4264 16445 4292 16544
rect 4430 16532 4436 16544
rect 4488 16572 4494 16584
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 4488 16544 4813 16572
rect 4488 16532 4494 16544
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 6196 16572 6224 16612
rect 6638 16572 6644 16584
rect 6196 16558 6644 16572
rect 6210 16544 6644 16558
rect 4801 16535 4859 16541
rect 6638 16532 6644 16544
rect 6696 16572 6702 16584
rect 7392 16572 7420 16736
rect 9674 16708 9680 16720
rect 9324 16680 9680 16708
rect 9324 16649 9352 16680
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9784 16640 9812 16748
rect 9950 16736 9956 16748
rect 10008 16776 10014 16788
rect 10134 16776 10140 16788
rect 10008 16748 10140 16776
rect 10008 16736 10014 16748
rect 10134 16736 10140 16748
rect 10192 16776 10198 16788
rect 10410 16776 10416 16788
rect 10192 16748 10416 16776
rect 10192 16736 10198 16748
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 10744 16748 12357 16776
rect 10744 16736 10750 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 12986 16736 12992 16788
rect 13044 16776 13050 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13044 16748 14105 16776
rect 13044 16736 13050 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14660 16748 15976 16776
rect 10980 16680 12112 16708
rect 9539 16612 9812 16640
rect 9953 16643 10011 16649
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 10042 16640 10048 16652
rect 9999 16612 10048 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10980 16640 11008 16680
rect 11882 16640 11888 16652
rect 10468 16612 11008 16640
rect 11072 16612 11888 16640
rect 10468 16600 10474 16612
rect 6696 16544 7420 16572
rect 6696 16532 6702 16544
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 8803 16544 8892 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 5074 16464 5080 16516
rect 5132 16464 5138 16516
rect 3513 16439 3571 16445
rect 3513 16436 3525 16439
rect 3384 16408 3525 16436
rect 3384 16396 3390 16408
rect 3513 16405 3525 16408
rect 3559 16436 3571 16439
rect 3881 16439 3939 16445
rect 3881 16436 3893 16439
rect 3559 16408 3893 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 3881 16405 3893 16408
rect 3927 16436 3939 16439
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 3927 16408 4261 16436
rect 3927 16405 3939 16408
rect 3881 16399 3939 16405
rect 4249 16405 4261 16408
rect 4295 16405 4307 16439
rect 4249 16399 4307 16405
rect 6546 16396 6552 16448
rect 6604 16396 6610 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6880 16408 7021 16436
rect 6880 16396 6886 16408
rect 7009 16405 7021 16408
rect 7055 16436 7067 16439
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7055 16408 7665 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7653 16405 7665 16408
rect 7699 16436 7711 16439
rect 8110 16436 8116 16448
rect 7699 16408 8116 16436
rect 7699 16405 7711 16408
rect 7653 16399 7711 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8294 16396 8300 16448
rect 8352 16396 8358 16448
rect 8570 16396 8576 16448
rect 8628 16396 8634 16448
rect 8864 16445 8892 16544
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 9640 16544 9689 16572
rect 9640 16532 9646 16544
rect 9677 16541 9689 16544
rect 9723 16541 9735 16575
rect 11072 16558 11100 16612
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12084 16649 12112 16680
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12115 16612 12909 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 14108 16640 14136 16739
rect 14550 16640 14556 16652
rect 14108 16612 14556 16640
rect 12897 16603 12955 16609
rect 9677 16535 9735 16541
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 11992 16572 12020 16603
rect 14550 16600 14556 16612
rect 14608 16640 14614 16652
rect 14660 16649 14688 16748
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 14608 16612 14657 16640
rect 14608 16600 14614 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15286 16640 15292 16652
rect 14967 16612 15292 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15948 16640 15976 16748
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 17034 16776 17040 16788
rect 16540 16748 17040 16776
rect 16540 16736 16546 16748
rect 17034 16736 17040 16748
rect 17092 16736 17098 16788
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 20162 16776 20168 16788
rect 19668 16748 20168 16776
rect 19668 16736 19674 16748
rect 20162 16736 20168 16748
rect 20220 16776 20226 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 20220 16748 20361 16776
rect 20220 16736 20226 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 20349 16739 20407 16745
rect 20364 16708 20392 16739
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21048 16748 21189 16776
rect 21048 16736 21054 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 23198 16776 23204 16788
rect 21177 16739 21235 16745
rect 22066 16748 23204 16776
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 20364 16680 21097 16708
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 15948 16612 16497 16640
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 17402 16640 17408 16652
rect 16899 16612 17408 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 17678 16600 17684 16652
rect 17736 16640 17742 16652
rect 18279 16643 18337 16649
rect 18279 16640 18291 16643
rect 17736 16612 18291 16640
rect 17736 16600 17742 16612
rect 18279 16609 18291 16612
rect 18325 16609 18337 16643
rect 18279 16603 18337 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16640 18935 16643
rect 19518 16640 19524 16652
rect 18923 16612 19524 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 12158 16572 12164 16584
rect 11480 16544 12164 16572
rect 11480 16532 11486 16544
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18196 16544 18613 16572
rect 18196 16532 18202 16544
rect 18601 16541 18613 16544
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16572 20775 16575
rect 20806 16572 20812 16584
rect 20763 16544 20812 16572
rect 20763 16541 20775 16544
rect 20717 16535 20775 16541
rect 11606 16504 11612 16516
rect 9232 16476 10364 16504
rect 9232 16448 9260 16476
rect 8849 16439 8907 16445
rect 8849 16405 8861 16439
rect 8895 16405 8907 16439
rect 8849 16399 8907 16405
rect 9214 16396 9220 16448
rect 9272 16396 9278 16448
rect 10336 16436 10364 16476
rect 11440 16476 11612 16504
rect 11440 16445 11468 16476
rect 11606 16464 11612 16476
rect 11664 16464 11670 16516
rect 12805 16507 12863 16513
rect 12805 16504 12817 16507
rect 11900 16476 12817 16504
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 10336 16408 11437 16436
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11425 16399 11483 16405
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 11900 16445 11928 16476
rect 12805 16473 12817 16476
rect 12851 16473 12863 16507
rect 19334 16504 19340 16516
rect 16146 16476 16252 16504
rect 17894 16476 17954 16504
rect 12805 16467 12863 16473
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11848 16408 11897 16436
rect 11848 16396 11854 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 12713 16439 12771 16445
rect 12713 16436 12725 16439
rect 12492 16408 12725 16436
rect 12492 16396 12498 16408
rect 12713 16405 12725 16408
rect 12759 16405 12771 16439
rect 12820 16436 12848 16467
rect 13354 16436 13360 16448
rect 12820 16408 13360 16436
rect 12713 16399 12771 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 14274 16436 14280 16448
rect 13863 16408 14280 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 14274 16396 14280 16408
rect 14332 16436 14338 16448
rect 14553 16439 14611 16445
rect 14553 16436 14565 16439
rect 14332 16408 14565 16436
rect 14332 16396 14338 16408
rect 14553 16405 14565 16408
rect 14599 16436 14611 16439
rect 16224 16436 16252 16476
rect 17926 16436 17954 16476
rect 18524 16476 19340 16504
rect 18524 16448 18552 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20346 16504 20352 16516
rect 20180 16476 20352 16504
rect 20180 16448 20208 16476
rect 20346 16464 20352 16476
rect 20404 16504 20410 16516
rect 20441 16507 20499 16513
rect 20441 16504 20453 16507
rect 20404 16476 20453 16504
rect 20404 16464 20410 16476
rect 20441 16473 20453 16476
rect 20487 16473 20499 16507
rect 20441 16467 20499 16473
rect 18322 16436 18328 16448
rect 14599 16408 18328 16436
rect 14599 16405 14611 16408
rect 14553 16399 14611 16405
rect 18322 16396 18328 16408
rect 18380 16436 18386 16448
rect 18506 16436 18512 16448
rect 18380 16408 18512 16436
rect 18380 16396 18386 16408
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 20162 16396 20168 16448
rect 20220 16396 20226 16448
rect 20640 16436 20668 16535
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 20898 16532 20904 16584
rect 20956 16532 20962 16584
rect 21008 16581 21036 16680
rect 21085 16677 21097 16680
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 22066 16640 22094 16748
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 24581 16779 24639 16785
rect 24581 16745 24593 16779
rect 24627 16776 24639 16779
rect 24946 16776 24952 16788
rect 24627 16748 24952 16776
rect 24627 16745 24639 16748
rect 24581 16739 24639 16745
rect 24946 16736 24952 16748
rect 25004 16736 25010 16788
rect 28258 16736 28264 16788
rect 28316 16776 28322 16788
rect 28537 16779 28595 16785
rect 28537 16776 28549 16779
rect 28316 16748 28549 16776
rect 28316 16736 28322 16748
rect 28537 16745 28549 16748
rect 28583 16745 28595 16779
rect 28537 16739 28595 16745
rect 30101 16779 30159 16785
rect 30101 16745 30113 16779
rect 30147 16776 30159 16779
rect 30650 16776 30656 16788
rect 30147 16748 30656 16776
rect 30147 16745 30159 16748
rect 30101 16739 30159 16745
rect 30650 16736 30656 16748
rect 30708 16736 30714 16788
rect 31110 16776 31116 16788
rect 30760 16748 31116 16776
rect 28905 16711 28963 16717
rect 28905 16708 28917 16711
rect 22480 16680 25084 16708
rect 22480 16649 22508 16680
rect 21284 16612 22094 16640
rect 22465 16643 22523 16649
rect 21284 16584 21312 16612
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21266 16532 21272 16584
rect 21324 16532 21330 16584
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16572 21419 16575
rect 21450 16572 21456 16584
rect 21407 16544 21456 16572
rect 21407 16541 21419 16544
rect 21361 16535 21419 16541
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 21560 16581 21588 16612
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22649 16643 22707 16649
rect 22649 16609 22661 16643
rect 22695 16640 22707 16643
rect 23201 16643 23259 16649
rect 23201 16640 23213 16643
rect 22695 16612 23213 16640
rect 22695 16609 22707 16612
rect 22649 16603 22707 16609
rect 23201 16609 23213 16612
rect 23247 16640 23259 16643
rect 24394 16640 24400 16652
rect 23247 16612 24400 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 22278 16532 22284 16584
rect 22336 16572 22342 16584
rect 22664 16572 22692 16603
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 25056 16649 25084 16680
rect 28736 16680 28917 16708
rect 25041 16643 25099 16649
rect 25041 16609 25053 16643
rect 25087 16640 25099 16643
rect 25130 16640 25136 16652
rect 25087 16612 25136 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 25222 16600 25228 16652
rect 25280 16640 25286 16652
rect 25961 16643 26019 16649
rect 25961 16640 25973 16643
rect 25280 16612 25973 16640
rect 25280 16600 25286 16612
rect 25961 16609 25973 16612
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 26602 16640 26608 16652
rect 26476 16612 26608 16640
rect 26476 16600 26482 16612
rect 26602 16600 26608 16612
rect 26660 16640 26666 16652
rect 27157 16643 27215 16649
rect 27157 16640 27169 16643
rect 26660 16612 27169 16640
rect 26660 16600 26666 16612
rect 27157 16609 27169 16612
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 27338 16600 27344 16652
rect 27396 16600 27402 16652
rect 22336 16544 22692 16572
rect 22925 16575 22983 16581
rect 22336 16532 22342 16544
rect 22925 16541 22937 16575
rect 22971 16572 22983 16575
rect 24026 16572 24032 16584
rect 22971 16544 24032 16572
rect 22971 16541 22983 16544
rect 22925 16535 22983 16541
rect 24026 16532 24032 16544
rect 24084 16532 24090 16584
rect 25777 16575 25835 16581
rect 25777 16541 25789 16575
rect 25823 16572 25835 16575
rect 26970 16572 26976 16584
rect 25823 16544 26976 16572
rect 25823 16541 25835 16544
rect 25777 16535 25835 16541
rect 26970 16532 26976 16544
rect 27028 16532 27034 16584
rect 27356 16572 27384 16600
rect 27356 16544 27568 16572
rect 21726 16464 21732 16516
rect 21784 16504 21790 16516
rect 27540 16513 27568 16544
rect 27890 16532 27896 16584
rect 27948 16572 27954 16584
rect 28077 16575 28135 16581
rect 28077 16572 28089 16575
rect 27948 16544 28089 16572
rect 27948 16532 27954 16544
rect 28077 16541 28089 16544
rect 28123 16541 28135 16575
rect 28077 16535 28135 16541
rect 28166 16532 28172 16584
rect 28224 16532 28230 16584
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16572 28319 16575
rect 28350 16572 28356 16584
rect 28307 16544 28356 16572
rect 28307 16541 28319 16544
rect 28261 16535 28319 16541
rect 28350 16532 28356 16544
rect 28408 16532 28414 16584
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16572 28503 16575
rect 28626 16572 28632 16584
rect 28491 16544 28632 16572
rect 28491 16541 28503 16544
rect 28445 16535 28503 16541
rect 28626 16532 28632 16544
rect 28684 16532 28690 16584
rect 28736 16581 28764 16680
rect 28905 16677 28917 16680
rect 28951 16677 28963 16711
rect 28905 16671 28963 16677
rect 28994 16668 29000 16720
rect 29052 16708 29058 16720
rect 29052 16680 29960 16708
rect 29052 16668 29058 16680
rect 29457 16643 29515 16649
rect 29457 16640 29469 16643
rect 28920 16612 29469 16640
rect 28721 16575 28779 16581
rect 28721 16541 28733 16575
rect 28767 16541 28779 16575
rect 28721 16535 28779 16541
rect 28920 16516 28948 16612
rect 29457 16609 29469 16612
rect 29503 16609 29515 16643
rect 29457 16603 29515 16609
rect 29932 16584 29960 16680
rect 30650 16600 30656 16652
rect 30708 16640 30714 16652
rect 30760 16640 30788 16748
rect 31110 16736 31116 16748
rect 31168 16736 31174 16788
rect 31662 16736 31668 16788
rect 31720 16776 31726 16788
rect 32214 16776 32220 16788
rect 31720 16748 32220 16776
rect 31720 16736 31726 16748
rect 32214 16736 32220 16748
rect 32272 16736 32278 16788
rect 32306 16736 32312 16788
rect 32364 16776 32370 16788
rect 32585 16779 32643 16785
rect 32585 16776 32597 16779
rect 32364 16748 32597 16776
rect 32364 16736 32370 16748
rect 32585 16745 32597 16748
rect 32631 16745 32643 16779
rect 32585 16739 32643 16745
rect 35894 16736 35900 16788
rect 35952 16736 35958 16788
rect 36725 16779 36783 16785
rect 36725 16745 36737 16779
rect 36771 16776 36783 16779
rect 36814 16776 36820 16788
rect 36771 16748 36820 16776
rect 36771 16745 36783 16748
rect 36725 16739 36783 16745
rect 36814 16736 36820 16748
rect 36872 16736 36878 16788
rect 37182 16736 37188 16788
rect 37240 16776 37246 16788
rect 37737 16779 37795 16785
rect 37240 16748 37596 16776
rect 37240 16736 37246 16748
rect 32122 16668 32128 16720
rect 32180 16708 32186 16720
rect 33318 16708 33324 16720
rect 32180 16680 33324 16708
rect 32180 16668 32186 16680
rect 33318 16668 33324 16680
rect 33376 16668 33382 16720
rect 33689 16711 33747 16717
rect 33689 16677 33701 16711
rect 33735 16677 33747 16711
rect 33689 16671 33747 16677
rect 30708 16612 30788 16640
rect 31113 16643 31171 16649
rect 30708 16600 30714 16612
rect 31113 16609 31125 16643
rect 31159 16640 31171 16643
rect 31478 16640 31484 16652
rect 31159 16612 31484 16640
rect 31159 16609 31171 16612
rect 31113 16603 31171 16609
rect 31478 16600 31484 16612
rect 31536 16600 31542 16652
rect 32306 16600 32312 16652
rect 32364 16600 32370 16652
rect 32490 16600 32496 16652
rect 32548 16640 32554 16652
rect 33229 16643 33287 16649
rect 33229 16640 33241 16643
rect 32548 16612 33241 16640
rect 32548 16600 32554 16612
rect 33229 16609 33241 16612
rect 33275 16640 33287 16643
rect 33410 16640 33416 16652
rect 33275 16612 33416 16640
rect 33275 16609 33287 16612
rect 33229 16603 33287 16609
rect 33410 16600 33416 16612
rect 33468 16600 33474 16652
rect 29273 16575 29331 16581
rect 29273 16541 29285 16575
rect 29319 16572 29331 16575
rect 29362 16572 29368 16584
rect 29319 16544 29368 16572
rect 29319 16541 29331 16544
rect 29273 16535 29331 16541
rect 29362 16532 29368 16544
rect 29420 16572 29426 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29420 16544 29745 16572
rect 29420 16532 29426 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 29914 16532 29920 16584
rect 29972 16532 29978 16584
rect 30558 16572 30564 16584
rect 30024 16544 30564 16572
rect 21913 16507 21971 16513
rect 21913 16504 21925 16507
rect 21784 16476 21925 16504
rect 21784 16464 21790 16476
rect 21913 16473 21925 16476
rect 21959 16473 21971 16507
rect 24213 16507 24271 16513
rect 24213 16504 24225 16507
rect 21913 16467 21971 16473
rect 23308 16476 24225 16504
rect 23308 16448 23336 16476
rect 24213 16473 24225 16476
rect 24259 16504 24271 16507
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 24259 16476 25881 16504
rect 24259 16473 24271 16476
rect 24213 16467 24271 16473
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 27341 16507 27399 16513
rect 27341 16473 27353 16507
rect 27387 16473 27399 16507
rect 27341 16467 27399 16473
rect 27525 16507 27583 16513
rect 27525 16473 27537 16507
rect 27571 16473 27583 16507
rect 27525 16467 27583 16473
rect 21266 16436 21272 16448
rect 20640 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 22002 16396 22008 16448
rect 22060 16396 22066 16448
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 23014 16436 23020 16448
rect 22428 16408 23020 16436
rect 22428 16396 22434 16408
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23750 16396 23756 16448
rect 23808 16396 23814 16448
rect 24118 16396 24124 16448
rect 24176 16396 24182 16448
rect 24946 16396 24952 16448
rect 25004 16396 25010 16448
rect 25406 16396 25412 16448
rect 25464 16396 25470 16448
rect 25498 16396 25504 16448
rect 25556 16436 25562 16448
rect 26421 16439 26479 16445
rect 26421 16436 26433 16439
rect 25556 16408 26433 16436
rect 25556 16396 25562 16408
rect 26421 16405 26433 16408
rect 26467 16405 26479 16439
rect 26421 16399 26479 16405
rect 26878 16396 26884 16448
rect 26936 16396 26942 16448
rect 27356 16436 27384 16467
rect 28902 16464 28908 16516
rect 28960 16464 28966 16516
rect 29104 16476 29500 16504
rect 27614 16436 27620 16448
rect 27356 16408 27620 16436
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 27706 16396 27712 16448
rect 27764 16396 27770 16448
rect 27801 16439 27859 16445
rect 27801 16405 27813 16439
rect 27847 16436 27859 16439
rect 29104 16436 29132 16476
rect 27847 16408 29132 16436
rect 27847 16405 27859 16408
rect 27801 16399 27859 16405
rect 29178 16396 29184 16448
rect 29236 16436 29242 16448
rect 29365 16439 29423 16445
rect 29365 16436 29377 16439
rect 29236 16408 29377 16436
rect 29236 16396 29242 16408
rect 29365 16405 29377 16408
rect 29411 16405 29423 16439
rect 29472 16436 29500 16476
rect 29546 16464 29552 16516
rect 29604 16504 29610 16516
rect 30024 16504 30052 16544
rect 30558 16532 30564 16544
rect 30616 16532 30622 16584
rect 30837 16575 30895 16581
rect 30837 16541 30849 16575
rect 30883 16541 30895 16575
rect 32324 16572 32352 16600
rect 33505 16575 33563 16581
rect 33505 16572 33517 16575
rect 32246 16544 32352 16572
rect 32692 16544 33517 16572
rect 30837 16535 30895 16541
rect 29604 16476 30052 16504
rect 30469 16507 30527 16513
rect 29604 16464 29610 16476
rect 30469 16473 30481 16507
rect 30515 16504 30527 16507
rect 30852 16504 30880 16535
rect 30515 16476 30972 16504
rect 30515 16473 30527 16476
rect 30469 16467 30527 16473
rect 30944 16448 30972 16476
rect 30282 16436 30288 16448
rect 29472 16408 30288 16436
rect 29365 16399 29423 16405
rect 30282 16396 30288 16408
rect 30340 16436 30346 16448
rect 30834 16436 30840 16448
rect 30340 16408 30840 16436
rect 30340 16396 30346 16408
rect 30834 16396 30840 16408
rect 30892 16396 30898 16448
rect 30926 16396 30932 16448
rect 30984 16396 30990 16448
rect 32692 16445 32720 16544
rect 33505 16541 33517 16544
rect 33551 16541 33563 16575
rect 33505 16535 33563 16541
rect 33704 16516 33732 16671
rect 34333 16643 34391 16649
rect 34333 16609 34345 16643
rect 34379 16640 34391 16643
rect 35986 16640 35992 16652
rect 34379 16612 35992 16640
rect 34379 16609 34391 16612
rect 34333 16603 34391 16609
rect 35986 16600 35992 16612
rect 36044 16600 36050 16652
rect 36449 16643 36507 16649
rect 36449 16609 36461 16643
rect 36495 16640 36507 16643
rect 37182 16640 37188 16652
rect 36495 16612 37188 16640
rect 36495 16609 36507 16612
rect 36449 16603 36507 16609
rect 34054 16532 34060 16584
rect 34112 16532 34118 16584
rect 35802 16532 35808 16584
rect 35860 16572 35866 16584
rect 36464 16572 36492 16603
rect 37182 16600 37188 16612
rect 37240 16640 37246 16652
rect 37277 16643 37335 16649
rect 37277 16640 37289 16643
rect 37240 16612 37289 16640
rect 37240 16600 37246 16612
rect 37277 16609 37289 16612
rect 37323 16609 37335 16643
rect 37568 16640 37596 16748
rect 37737 16745 37749 16779
rect 37783 16776 37795 16779
rect 38194 16776 38200 16788
rect 37783 16748 38200 16776
rect 37783 16745 37795 16748
rect 37737 16739 37795 16745
rect 38194 16736 38200 16748
rect 38252 16736 38258 16788
rect 39114 16736 39120 16788
rect 39172 16736 39178 16788
rect 39942 16776 39948 16788
rect 39224 16748 39948 16776
rect 38764 16680 39068 16708
rect 38764 16649 38792 16680
rect 39040 16652 39068 16680
rect 38749 16643 38807 16649
rect 37568 16612 38608 16640
rect 37277 16603 37335 16609
rect 35860 16544 36492 16572
rect 37921 16575 37979 16581
rect 35860 16532 35866 16544
rect 37921 16541 37933 16575
rect 37967 16541 37979 16575
rect 37921 16535 37979 16541
rect 38197 16575 38255 16581
rect 38197 16541 38209 16575
rect 38243 16572 38255 16575
rect 38286 16572 38292 16584
rect 38243 16544 38292 16572
rect 38243 16541 38255 16544
rect 38197 16535 38255 16541
rect 33137 16507 33195 16513
rect 33137 16504 33149 16507
rect 32968 16476 33149 16504
rect 32968 16448 32996 16476
rect 33137 16473 33149 16476
rect 33183 16473 33195 16507
rect 33137 16467 33195 16473
rect 33686 16464 33692 16516
rect 33744 16464 33750 16516
rect 34790 16464 34796 16516
rect 34848 16464 34854 16516
rect 36357 16507 36415 16513
rect 36357 16473 36369 16507
rect 36403 16504 36415 16507
rect 36446 16504 36452 16516
rect 36403 16476 36452 16504
rect 36403 16473 36415 16476
rect 36357 16467 36415 16473
rect 36446 16464 36452 16476
rect 36504 16464 36510 16516
rect 37093 16507 37151 16513
rect 37093 16473 37105 16507
rect 37139 16504 37151 16507
rect 37936 16504 37964 16535
rect 38286 16532 38292 16544
rect 38344 16532 38350 16584
rect 37139 16476 37872 16504
rect 37936 16476 38332 16504
rect 37139 16473 37151 16476
rect 37093 16467 37151 16473
rect 32677 16439 32735 16445
rect 32677 16405 32689 16439
rect 32723 16405 32735 16439
rect 32677 16399 32735 16405
rect 32950 16396 32956 16448
rect 33008 16396 33014 16448
rect 33042 16396 33048 16448
rect 33100 16396 33106 16448
rect 35710 16396 35716 16448
rect 35768 16436 35774 16448
rect 35805 16439 35863 16445
rect 35805 16436 35817 16439
rect 35768 16408 35817 16436
rect 35768 16396 35774 16408
rect 35805 16405 35817 16408
rect 35851 16405 35863 16439
rect 35805 16399 35863 16405
rect 35894 16396 35900 16448
rect 35952 16436 35958 16448
rect 36170 16436 36176 16448
rect 35952 16408 36176 16436
rect 35952 16396 35958 16408
rect 36170 16396 36176 16408
rect 36228 16436 36234 16448
rect 36265 16439 36323 16445
rect 36265 16436 36277 16439
rect 36228 16408 36277 16436
rect 36228 16396 36234 16408
rect 36265 16405 36277 16408
rect 36311 16405 36323 16439
rect 36265 16399 36323 16405
rect 36906 16396 36912 16448
rect 36964 16436 36970 16448
rect 37185 16439 37243 16445
rect 37185 16436 37197 16439
rect 36964 16408 37197 16436
rect 36964 16396 36970 16408
rect 37185 16405 37197 16408
rect 37231 16405 37243 16439
rect 37844 16436 37872 16476
rect 37918 16436 37924 16448
rect 37844 16408 37924 16436
rect 37185 16399 37243 16405
rect 37918 16396 37924 16408
rect 37976 16396 37982 16448
rect 38010 16396 38016 16448
rect 38068 16396 38074 16448
rect 38304 16445 38332 16476
rect 38289 16439 38347 16445
rect 38289 16405 38301 16439
rect 38335 16405 38347 16439
rect 38580 16436 38608 16612
rect 38749 16609 38761 16643
rect 38795 16609 38807 16643
rect 38749 16603 38807 16609
rect 38838 16600 38844 16652
rect 38896 16600 38902 16652
rect 39022 16600 39028 16652
rect 39080 16600 39086 16652
rect 39132 16640 39160 16736
rect 39224 16720 39252 16748
rect 39942 16736 39948 16748
rect 40000 16736 40006 16788
rect 40586 16736 40592 16788
rect 40644 16736 40650 16788
rect 40954 16736 40960 16788
rect 41012 16736 41018 16788
rect 43070 16736 43076 16788
rect 43128 16736 43134 16788
rect 43898 16736 43904 16788
rect 43956 16736 43962 16788
rect 44634 16736 44640 16788
rect 44692 16776 44698 16788
rect 44913 16779 44971 16785
rect 44913 16776 44925 16779
rect 44692 16748 44925 16776
rect 44692 16736 44698 16748
rect 44913 16745 44925 16748
rect 44959 16745 44971 16779
rect 44913 16739 44971 16745
rect 39206 16668 39212 16720
rect 39264 16668 39270 16720
rect 39485 16643 39543 16649
rect 39485 16640 39497 16643
rect 39132 16612 39497 16640
rect 39485 16609 39497 16612
rect 39531 16609 39543 16643
rect 40604 16640 40632 16736
rect 43088 16708 43116 16736
rect 43088 16680 43484 16708
rect 41325 16643 41383 16649
rect 41325 16640 41337 16643
rect 40604 16612 41337 16640
rect 39485 16603 39543 16609
rect 41325 16609 41337 16612
rect 41371 16609 41383 16643
rect 43088 16640 43116 16680
rect 41325 16603 41383 16609
rect 42812 16612 43116 16640
rect 38657 16575 38715 16581
rect 38657 16541 38669 16575
rect 38703 16572 38715 16575
rect 38930 16572 38936 16584
rect 38703 16544 38936 16572
rect 38703 16541 38715 16544
rect 38657 16535 38715 16541
rect 38930 16532 38936 16544
rect 38988 16532 38994 16584
rect 39114 16532 39120 16584
rect 39172 16572 39178 16584
rect 39209 16575 39267 16581
rect 39209 16572 39221 16575
rect 39172 16544 39221 16572
rect 39172 16532 39178 16544
rect 39209 16541 39221 16544
rect 39255 16541 39267 16575
rect 39209 16535 39267 16541
rect 40954 16532 40960 16584
rect 41012 16572 41018 16584
rect 41049 16575 41107 16581
rect 41049 16572 41061 16575
rect 41012 16544 41061 16572
rect 41012 16532 41018 16544
rect 41049 16541 41061 16544
rect 41095 16541 41107 16575
rect 41049 16535 41107 16541
rect 38838 16464 38844 16516
rect 38896 16504 38902 16516
rect 39482 16504 39488 16516
rect 38896 16476 39488 16504
rect 38896 16464 38902 16476
rect 39482 16464 39488 16476
rect 39540 16464 39546 16516
rect 39942 16464 39948 16516
rect 40000 16464 40006 16516
rect 41322 16504 41328 16516
rect 40710 16476 41328 16504
rect 41322 16464 41328 16476
rect 41380 16504 41386 16516
rect 41380 16476 41814 16504
rect 41380 16464 41386 16476
rect 42702 16464 42708 16516
rect 42760 16504 42766 16516
rect 42812 16504 42840 16612
rect 43346 16600 43352 16652
rect 43404 16600 43410 16652
rect 43456 16649 43484 16680
rect 43441 16643 43499 16649
rect 43441 16609 43453 16643
rect 43487 16609 43499 16643
rect 43441 16603 43499 16609
rect 44174 16600 44180 16652
rect 44232 16640 44238 16652
rect 44545 16643 44603 16649
rect 44545 16640 44557 16643
rect 44232 16612 44557 16640
rect 44232 16600 44238 16612
rect 44545 16609 44557 16612
rect 44591 16609 44603 16643
rect 44545 16603 44603 16609
rect 43257 16575 43315 16581
rect 43257 16541 43269 16575
rect 43303 16572 43315 16575
rect 44358 16572 44364 16584
rect 43303 16544 44364 16572
rect 43303 16541 43315 16544
rect 43257 16535 43315 16541
rect 44358 16532 44364 16544
rect 44416 16532 44422 16584
rect 42760 16476 42840 16504
rect 42760 16464 42766 16476
rect 40770 16436 40776 16448
rect 38580 16408 40776 16436
rect 38289 16399 38347 16405
rect 40770 16396 40776 16408
rect 40828 16396 40834 16448
rect 41598 16396 41604 16448
rect 41656 16436 41662 16448
rect 42797 16439 42855 16445
rect 42797 16436 42809 16439
rect 41656 16408 42809 16436
rect 41656 16396 41662 16408
rect 42797 16405 42809 16408
rect 42843 16405 42855 16439
rect 42797 16399 42855 16405
rect 42886 16396 42892 16448
rect 42944 16396 42950 16448
rect 460 16346 45540 16368
rect 460 16294 6070 16346
rect 6122 16294 6134 16346
rect 6186 16294 6198 16346
rect 6250 16294 6262 16346
rect 6314 16294 6326 16346
rect 6378 16294 11070 16346
rect 11122 16294 11134 16346
rect 11186 16294 11198 16346
rect 11250 16294 11262 16346
rect 11314 16294 11326 16346
rect 11378 16294 16070 16346
rect 16122 16294 16134 16346
rect 16186 16294 16198 16346
rect 16250 16294 16262 16346
rect 16314 16294 16326 16346
rect 16378 16294 21070 16346
rect 21122 16294 21134 16346
rect 21186 16294 21198 16346
rect 21250 16294 21262 16346
rect 21314 16294 21326 16346
rect 21378 16294 26070 16346
rect 26122 16294 26134 16346
rect 26186 16294 26198 16346
rect 26250 16294 26262 16346
rect 26314 16294 26326 16346
rect 26378 16294 31070 16346
rect 31122 16294 31134 16346
rect 31186 16294 31198 16346
rect 31250 16294 31262 16346
rect 31314 16294 31326 16346
rect 31378 16294 36070 16346
rect 36122 16294 36134 16346
rect 36186 16294 36198 16346
rect 36250 16294 36262 16346
rect 36314 16294 36326 16346
rect 36378 16294 41070 16346
rect 41122 16294 41134 16346
rect 41186 16294 41198 16346
rect 41250 16294 41262 16346
rect 41314 16294 41326 16346
rect 41378 16294 45540 16346
rect 460 16272 45540 16294
rect 4338 16192 4344 16244
rect 4396 16232 4402 16244
rect 4614 16232 4620 16244
rect 4396 16204 4620 16232
rect 4396 16192 4402 16204
rect 4614 16192 4620 16204
rect 4672 16232 4678 16244
rect 4709 16235 4767 16241
rect 4709 16232 4721 16235
rect 4672 16204 4721 16232
rect 4672 16192 4678 16204
rect 4709 16201 4721 16204
rect 4755 16201 4767 16235
rect 4709 16195 4767 16201
rect 5074 16192 5080 16244
rect 5132 16232 5138 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 5132 16204 5365 16232
rect 5132 16192 5138 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 5500 16204 6101 16232
rect 5500 16192 5506 16204
rect 6089 16201 6101 16204
rect 6135 16201 6147 16235
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6089 16195 6147 16201
rect 6196 16204 6561 16232
rect 6196 16164 6224 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6549 16195 6607 16201
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 7374 16232 7380 16244
rect 7147 16204 7380 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7374 16192 7380 16204
rect 7432 16232 7438 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7432 16204 7757 16232
rect 7432 16192 7438 16204
rect 5276 16136 6224 16164
rect 5276 16105 5304 16136
rect 6274 16121 6332 16127
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5442 16056 5448 16108
rect 5500 16056 5506 16108
rect 6274 16106 6286 16121
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5644 16068 5733 16096
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3384 16000 3617 16028
rect 3384 15988 3390 16000
rect 3605 15997 3617 16000
rect 3651 16028 3663 16031
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 3651 16000 4353 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 4341 15997 4353 16000
rect 4387 16028 4399 16031
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4387 16000 5089 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 5644 15960 5672 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 6104 16096 6286 16106
rect 5721 16059 5779 16065
rect 5828 16087 6286 16096
rect 6320 16087 6332 16121
rect 5828 16081 6332 16087
rect 6365 16099 6423 16105
rect 5828 16078 6317 16081
rect 5828 16068 6132 16078
rect 5828 16040 5856 16068
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 5810 15988 5816 16040
rect 5868 15988 5874 16040
rect 6380 16028 6408 16059
rect 6289 16000 6408 16028
rect 6289 15960 6317 16000
rect 6546 15988 6552 16040
rect 6604 15988 6610 16040
rect 7668 16028 7696 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 8570 16192 8576 16244
rect 8628 16192 8634 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 9953 16235 10011 16241
rect 9272 16204 9904 16232
rect 9272 16192 9278 16204
rect 8110 16164 8116 16176
rect 7944 16136 8116 16164
rect 7944 16105 7972 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 8205 16167 8263 16173
rect 8205 16133 8217 16167
rect 8251 16164 8263 16167
rect 8588 16164 8616 16192
rect 8251 16136 8616 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 9324 16028 9352 16082
rect 7668 16000 9352 16028
rect 9876 16028 9904 16204
rect 9953 16201 9965 16235
rect 9999 16232 10011 16235
rect 10318 16232 10324 16244
rect 9999 16204 10324 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 13556 16204 14320 16232
rect 11422 16164 11428 16176
rect 10336 16136 11428 16164
rect 10336 16105 10364 16136
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 13556 16164 13584 16204
rect 12820 16136 13584 16164
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 12820 16096 12848 16136
rect 14292 16108 14320 16204
rect 15286 16192 15292 16244
rect 15344 16192 15350 16244
rect 16390 16192 16396 16244
rect 16448 16192 16454 16244
rect 16850 16192 16856 16244
rect 16908 16232 16914 16244
rect 17037 16235 17095 16241
rect 17037 16232 17049 16235
rect 16908 16204 17049 16232
rect 16908 16192 16914 16204
rect 17037 16201 17049 16204
rect 17083 16201 17095 16235
rect 17037 16195 17095 16201
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17276 16204 17509 16232
rect 17276 16192 17282 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17586 16192 17592 16244
rect 17644 16232 17650 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 17644 16204 18061 16232
rect 17644 16192 17650 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 19702 16192 19708 16244
rect 19760 16232 19766 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 19760 16204 20637 16232
rect 19760 16192 19766 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 20625 16195 20683 16201
rect 21542 16192 21548 16244
rect 21600 16192 21606 16244
rect 24026 16192 24032 16244
rect 24084 16232 24090 16244
rect 24121 16235 24179 16241
rect 24121 16232 24133 16235
rect 24084 16204 24133 16232
rect 24084 16192 24090 16204
rect 24121 16201 24133 16204
rect 24167 16201 24179 16235
rect 24121 16195 24179 16201
rect 26881 16235 26939 16241
rect 26881 16201 26893 16235
rect 26927 16201 26939 16235
rect 26881 16195 26939 16201
rect 16408 16164 16436 16192
rect 16408 16136 16712 16164
rect 12308 16068 12848 16096
rect 12308 16056 12314 16068
rect 12894 16056 12900 16108
rect 12952 16056 12958 16108
rect 14274 16056 14280 16108
rect 14332 16056 14338 16108
rect 15470 16056 15476 16108
rect 15528 16056 15534 16108
rect 15562 16056 15568 16108
rect 15620 16056 15626 16108
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 15930 16096 15936 16108
rect 15795 16068 15936 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 16114 16056 16120 16108
rect 16172 16056 16178 16108
rect 16298 16056 16304 16108
rect 16356 16056 16362 16108
rect 16393 16099 16451 16105
rect 16393 16065 16405 16099
rect 16439 16096 16451 16099
rect 16574 16096 16580 16108
rect 16439 16068 16580 16096
rect 16439 16065 16451 16068
rect 16393 16059 16451 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 16684 16105 16712 16136
rect 16942 16124 16948 16176
rect 17000 16164 17006 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 17000 16136 17141 16164
rect 17000 16124 17006 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 17328 16136 17724 16164
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16850 16056 16856 16108
rect 16908 16056 16914 16108
rect 17328 16105 17356 16136
rect 17696 16108 17724 16136
rect 18414 16124 18420 16176
rect 18472 16124 18478 16176
rect 18506 16124 18512 16176
rect 18564 16164 18570 16176
rect 18564 16136 18906 16164
rect 18564 16124 18570 16136
rect 20254 16124 20260 16176
rect 20312 16124 20318 16176
rect 21361 16167 21419 16173
rect 21361 16133 21373 16167
rect 21407 16164 21419 16167
rect 21726 16164 21732 16176
rect 21407 16136 21732 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 24210 16164 24216 16176
rect 23874 16136 24216 16164
rect 24210 16124 24216 16136
rect 24268 16124 24274 16176
rect 24489 16167 24547 16173
rect 24489 16133 24501 16167
rect 24535 16164 24547 16167
rect 24762 16164 24768 16176
rect 24535 16136 24768 16164
rect 24535 16133 24547 16136
rect 24489 16127 24547 16133
rect 24762 16124 24768 16136
rect 24820 16124 24826 16176
rect 26896 16164 26924 16195
rect 27614 16192 27620 16244
rect 27672 16232 27678 16244
rect 28537 16235 28595 16241
rect 28537 16232 28549 16235
rect 27672 16204 28549 16232
rect 27672 16192 27678 16204
rect 28537 16201 28549 16204
rect 28583 16201 28595 16235
rect 28537 16195 28595 16201
rect 28718 16192 28724 16244
rect 28776 16232 28782 16244
rect 29546 16232 29552 16244
rect 28776 16204 29552 16232
rect 28776 16192 28782 16204
rect 29546 16192 29552 16204
rect 29604 16192 29610 16244
rect 30098 16192 30104 16244
rect 30156 16232 30162 16244
rect 31205 16235 31263 16241
rect 31205 16232 31217 16235
rect 30156 16204 31217 16232
rect 30156 16192 30162 16204
rect 31205 16201 31217 16204
rect 31251 16201 31263 16235
rect 31205 16195 31263 16201
rect 32030 16192 32036 16244
rect 32088 16192 32094 16244
rect 33042 16192 33048 16244
rect 33100 16232 33106 16244
rect 33100 16204 35940 16232
rect 33100 16192 33106 16204
rect 27402 16167 27460 16173
rect 27402 16164 27414 16167
rect 26896 16136 27414 16164
rect 27402 16133 27414 16136
rect 27448 16133 27460 16167
rect 27402 16127 27460 16133
rect 27724 16136 28856 16164
rect 27724 16108 27752 16136
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 9876 16000 10425 16028
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 6564 15960 6592 15988
rect 10520 15960 10548 15991
rect 5500 15932 6317 15960
rect 6380 15932 6592 15960
rect 10152 15932 10548 15960
rect 5500 15920 5506 15932
rect 3329 15895 3387 15901
rect 3329 15861 3341 15895
rect 3375 15892 3387 15895
rect 3418 15892 3424 15904
rect 3375 15864 3424 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 3418 15852 3424 15864
rect 3476 15892 3482 15904
rect 4062 15892 4068 15904
rect 3476 15864 4068 15892
rect 3476 15852 3482 15864
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 5905 15895 5963 15901
rect 5905 15861 5917 15895
rect 5951 15892 5963 15895
rect 6380 15892 6408 15932
rect 10152 15904 10180 15932
rect 5951 15864 6408 15892
rect 5951 15861 5963 15864
rect 5905 15855 5963 15861
rect 9674 15852 9680 15904
rect 9732 15852 9738 15904
rect 10134 15852 10140 15904
rect 10192 15852 10198 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10888 15892 10916 15991
rect 11146 15988 11152 16040
rect 11204 15988 11210 16040
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 14182 16028 14188 16040
rect 13219 16000 14188 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14792 16000 14933 16028
rect 14792 15988 14798 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 16028 15715 16031
rect 16482 16028 16488 16040
rect 15703 16000 16488 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 16592 16028 16620 16056
rect 17328 16028 17356 16059
rect 17586 16056 17592 16108
rect 17644 16056 17650 16108
rect 17678 16056 17684 16108
rect 17736 16056 17742 16108
rect 17770 16056 17776 16108
rect 17828 16056 17834 16108
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16096 20131 16099
rect 20162 16096 20168 16108
rect 20119 16068 20168 16096
rect 20119 16065 20131 16068
rect 20073 16059 20131 16065
rect 17880 16028 17908 16059
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 16592 16000 17356 16028
rect 17696 16000 17908 16028
rect 12710 15920 12716 15972
rect 12768 15920 12774 15972
rect 16117 15963 16175 15969
rect 16117 15929 16129 15963
rect 16163 15960 16175 15963
rect 16666 15960 16672 15972
rect 16163 15932 16672 15960
rect 16163 15929 16175 15932
rect 16117 15923 16175 15929
rect 16666 15920 16672 15932
rect 16724 15920 16730 15972
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 17586 15960 17592 15972
rect 16816 15932 17592 15960
rect 16816 15920 16822 15932
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 10468 15864 10916 15892
rect 10468 15852 10474 15864
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12618 15892 12624 15904
rect 12216 15864 12624 15892
rect 12216 15852 12222 15864
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 12728 15892 12756 15920
rect 14274 15892 14280 15904
rect 12728 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 16853 15895 16911 15901
rect 16853 15861 16865 15895
rect 16899 15892 16911 15895
rect 16942 15892 16948 15904
rect 16899 15864 16948 15892
rect 16899 15861 16911 15864
rect 16853 15855 16911 15861
rect 16942 15852 16948 15864
rect 17000 15892 17006 15904
rect 17696 15892 17724 16000
rect 18138 15988 18144 16040
rect 18196 15988 18202 16040
rect 20364 16028 20392 16059
rect 20438 16056 20444 16108
rect 20496 16056 20502 16108
rect 20806 16056 20812 16108
rect 20864 16096 20870 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20864 16068 21281 16096
rect 20864 16056 20870 16068
rect 21269 16065 21281 16068
rect 21315 16096 21327 16099
rect 21315 16068 21864 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 19904 16000 20392 16028
rect 19904 15972 19932 16000
rect 19886 15920 19892 15972
rect 19944 15920 19950 15972
rect 21082 15960 21088 15972
rect 19996 15932 21088 15960
rect 17000 15864 17724 15892
rect 17000 15852 17006 15864
rect 18230 15852 18236 15904
rect 18288 15892 18294 15904
rect 19996 15892 20024 15932
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 21836 15960 21864 16068
rect 21910 16056 21916 16108
rect 21968 16056 21974 16108
rect 26326 16096 26332 16108
rect 25622 16068 26332 16096
rect 26326 16056 26332 16068
rect 26384 16056 26390 16108
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 27706 16056 27712 16108
rect 27764 16056 27770 16108
rect 28258 16056 28264 16108
rect 28316 16096 28322 16108
rect 28629 16099 28687 16105
rect 28629 16096 28641 16099
rect 28316 16068 28641 16096
rect 28316 16056 28322 16068
rect 28629 16065 28641 16068
rect 28675 16096 28687 16099
rect 28718 16096 28724 16108
rect 28675 16068 28724 16096
rect 28675 16065 28687 16068
rect 28629 16059 28687 16065
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 28828 16105 28856 16136
rect 30190 16124 30196 16176
rect 30248 16124 30254 16176
rect 32048 16164 32076 16192
rect 31496 16136 32076 16164
rect 28813 16099 28871 16105
rect 28813 16065 28825 16099
rect 28859 16065 28871 16099
rect 28813 16059 28871 16065
rect 28905 16099 28963 16105
rect 28905 16065 28917 16099
rect 28951 16065 28963 16099
rect 29270 16096 29276 16108
rect 29013 16095 29276 16096
rect 28905 16059 28963 16065
rect 28998 16089 29276 16095
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 16028 22063 16031
rect 22094 16028 22100 16040
rect 22051 16000 22100 16028
rect 22051 15997 22063 16000
rect 22005 15991 22063 15997
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 22189 16031 22247 16037
rect 22189 15997 22201 16031
rect 22235 16028 22247 16031
rect 22278 16028 22284 16040
rect 22235 16000 22284 16028
rect 22235 15997 22247 16000
rect 22189 15991 22247 15997
rect 22204 15960 22232 15991
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 15997 22431 16031
rect 22373 15991 22431 15997
rect 21836 15932 22232 15960
rect 18288 15864 20024 15892
rect 18288 15852 18294 15864
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20864 15864 20913 15892
rect 20864 15852 20870 15864
rect 20901 15861 20913 15864
rect 20947 15892 20959 15895
rect 21910 15892 21916 15904
rect 20947 15864 21916 15892
rect 20947 15861 20959 15864
rect 20901 15855 20959 15861
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22388 15892 22416 15991
rect 22646 15988 22652 16040
rect 22704 15988 22710 16040
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 16028 24271 16031
rect 24854 16028 24860 16040
rect 24259 16000 24860 16028
rect 24259 15997 24271 16000
rect 24213 15991 24271 15997
rect 22462 15892 22468 15904
rect 22388 15864 22468 15892
rect 22462 15852 22468 15864
rect 22520 15892 22526 15904
rect 24228 15892 24256 15991
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 24946 15988 24952 16040
rect 25004 16028 25010 16040
rect 25004 16000 26004 16028
rect 25004 15988 25010 16000
rect 25976 15969 26004 16000
rect 26878 15988 26884 16040
rect 26936 16028 26942 16040
rect 27157 16031 27215 16037
rect 27157 16028 27169 16031
rect 26936 16000 27169 16028
rect 26936 15988 26942 16000
rect 27157 15997 27169 16000
rect 27203 15997 27215 16031
rect 27157 15991 27215 15997
rect 25961 15963 26019 15969
rect 25961 15929 25973 15963
rect 26007 15929 26019 15963
rect 25961 15923 26019 15929
rect 22520 15864 24256 15892
rect 25976 15892 26004 15923
rect 26510 15920 26516 15972
rect 26568 15920 26574 15972
rect 28920 15892 28948 16059
rect 28998 16055 29010 16089
rect 29044 16068 29276 16089
rect 29044 16055 29056 16068
rect 29270 16056 29276 16068
rect 29328 16056 29334 16108
rect 31496 16105 31524 16136
rect 32306 16124 32312 16176
rect 32364 16124 32370 16176
rect 34054 16164 34060 16176
rect 33520 16136 34060 16164
rect 33520 16105 33548 16136
rect 34054 16124 34060 16136
rect 34112 16124 34118 16176
rect 35805 16167 35863 16173
rect 35805 16164 35817 16167
rect 35544 16136 35817 16164
rect 31481 16099 31539 16105
rect 31481 16065 31493 16099
rect 31527 16065 31539 16099
rect 31481 16059 31539 16065
rect 33505 16099 33563 16105
rect 33505 16065 33517 16099
rect 33551 16065 33563 16099
rect 33505 16059 33563 16065
rect 28998 16049 29056 16055
rect 25976 15864 28948 15892
rect 29013 15892 29041 16049
rect 29086 15988 29092 16040
rect 29144 15988 29150 16040
rect 29457 16031 29515 16037
rect 29457 15997 29469 16031
rect 29503 16028 29515 16031
rect 29503 16000 29592 16028
rect 29503 15997 29515 16000
rect 29457 15991 29515 15997
rect 29104 15960 29132 15988
rect 29273 15963 29331 15969
rect 29273 15960 29285 15963
rect 29104 15932 29285 15960
rect 29273 15929 29285 15932
rect 29319 15929 29331 15963
rect 29273 15923 29331 15929
rect 29086 15892 29092 15904
rect 29013 15864 29092 15892
rect 22520 15852 22526 15864
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 29564 15892 29592 16000
rect 29730 15988 29736 16040
rect 29788 15988 29794 16040
rect 30926 15988 30932 16040
rect 30984 16028 30990 16040
rect 31496 16028 31524 16059
rect 34790 16056 34796 16108
rect 34848 16096 34854 16108
rect 35544 16096 35572 16136
rect 35805 16133 35817 16136
rect 35851 16133 35863 16167
rect 35912 16164 35940 16204
rect 35986 16192 35992 16244
rect 36044 16232 36050 16244
rect 36173 16235 36231 16241
rect 36173 16232 36185 16235
rect 36044 16204 36185 16232
rect 36044 16192 36050 16204
rect 36173 16201 36185 16204
rect 36219 16201 36231 16235
rect 36173 16195 36231 16201
rect 36556 16204 40080 16232
rect 36556 16164 36584 16204
rect 35912 16136 36584 16164
rect 35805 16127 35863 16133
rect 36630 16124 36636 16176
rect 36688 16164 36694 16176
rect 36909 16167 36967 16173
rect 36909 16164 36921 16167
rect 36688 16136 36921 16164
rect 36688 16124 36694 16136
rect 36909 16133 36921 16136
rect 36955 16133 36967 16167
rect 39206 16164 39212 16176
rect 38134 16136 39212 16164
rect 36909 16127 36967 16133
rect 39206 16124 39212 16136
rect 39264 16124 39270 16176
rect 40052 16164 40080 16204
rect 40126 16192 40132 16244
rect 40184 16232 40190 16244
rect 40678 16232 40684 16244
rect 40184 16204 40684 16232
rect 40184 16192 40190 16204
rect 40678 16192 40684 16204
rect 40736 16192 40742 16244
rect 42886 16232 42892 16244
rect 40788 16204 42892 16232
rect 40788 16164 40816 16204
rect 42886 16192 42892 16204
rect 42944 16192 42950 16244
rect 43346 16192 43352 16244
rect 43404 16232 43410 16244
rect 43533 16235 43591 16241
rect 43533 16232 43545 16235
rect 43404 16204 43545 16232
rect 43404 16192 43410 16204
rect 43533 16201 43545 16204
rect 43579 16201 43591 16235
rect 43533 16195 43591 16201
rect 42061 16167 42119 16173
rect 42061 16164 42073 16167
rect 40052 16136 40816 16164
rect 41432 16136 42073 16164
rect 34848 16068 34914 16096
rect 35268 16068 35572 16096
rect 34848 16056 34854 16068
rect 35268 16040 35296 16068
rect 35710 16056 35716 16108
rect 35768 16056 35774 16108
rect 36357 16099 36415 16105
rect 36357 16065 36369 16099
rect 36403 16065 36415 16099
rect 36357 16059 36415 16065
rect 30984 16000 31524 16028
rect 31757 16031 31815 16037
rect 30984 15988 30990 16000
rect 31757 15997 31769 16031
rect 31803 16028 31815 16031
rect 32766 16028 32772 16040
rect 31803 16000 32772 16028
rect 31803 15997 31815 16000
rect 31757 15991 31815 15997
rect 32766 15988 32772 16000
rect 32824 15988 32830 16040
rect 33410 15988 33416 16040
rect 33468 16028 33474 16040
rect 33781 16031 33839 16037
rect 33781 16028 33793 16031
rect 33468 16000 33793 16028
rect 33468 15988 33474 16000
rect 33781 15997 33793 16000
rect 33827 15997 33839 16031
rect 33781 15991 33839 15997
rect 35250 15988 35256 16040
rect 35308 15988 35314 16040
rect 35434 15988 35440 16040
rect 35492 16028 35498 16040
rect 35802 16028 35808 16040
rect 35492 16000 35808 16028
rect 35492 15988 35498 16000
rect 35802 15988 35808 16000
rect 35860 16028 35866 16040
rect 35897 16031 35955 16037
rect 35897 16028 35909 16031
rect 35860 16000 35909 16028
rect 35860 15988 35866 16000
rect 35897 15997 35909 16000
rect 35943 15997 35955 16031
rect 35897 15991 35955 15997
rect 30944 15892 30972 15988
rect 35345 15963 35403 15969
rect 35345 15929 35357 15963
rect 35391 15960 35403 15963
rect 36372 15960 36400 16059
rect 37918 16056 37924 16108
rect 37976 16056 37982 16108
rect 40770 16056 40776 16108
rect 40828 16056 40834 16108
rect 41325 16099 41383 16105
rect 41325 16065 41337 16099
rect 41371 16065 41383 16099
rect 41325 16059 41383 16065
rect 36630 15988 36636 16040
rect 36688 16028 36694 16040
rect 37458 16028 37464 16040
rect 36688 16000 37464 16028
rect 36688 15988 36694 16000
rect 37458 15988 37464 16000
rect 37516 15988 37522 16040
rect 37936 16028 37964 16056
rect 38381 16031 38439 16037
rect 38381 16028 38393 16031
rect 37936 16000 38393 16028
rect 38381 15997 38393 16000
rect 38427 15997 38439 16031
rect 38381 15991 38439 15997
rect 38470 15988 38476 16040
rect 38528 15988 38534 16040
rect 38749 16031 38807 16037
rect 38749 16028 38761 16031
rect 38580 16000 38761 16028
rect 35391 15932 36400 15960
rect 35391 15929 35403 15932
rect 35345 15923 35403 15929
rect 38010 15920 38016 15972
rect 38068 15960 38074 15972
rect 38580 15960 38608 16000
rect 38749 15997 38761 16000
rect 38795 15997 38807 16031
rect 38749 15991 38807 15997
rect 39482 15988 39488 16040
rect 39540 16028 39546 16040
rect 40865 16031 40923 16037
rect 40865 16028 40877 16031
rect 39540 16000 40877 16028
rect 39540 15988 39546 16000
rect 40865 15997 40877 16000
rect 40911 15997 40923 16031
rect 40865 15991 40923 15997
rect 38068 15932 38608 15960
rect 40313 15963 40371 15969
rect 38068 15920 38074 15932
rect 40313 15929 40325 15963
rect 40359 15960 40371 15963
rect 41340 15960 41368 16059
rect 41432 15969 41460 16136
rect 42061 16133 42073 16136
rect 42107 16133 42119 16167
rect 42061 16127 42119 16133
rect 41598 16056 41604 16108
rect 41656 16056 41662 16108
rect 43162 16056 43168 16108
rect 43220 16096 43226 16108
rect 43220 16068 43944 16096
rect 43220 16056 43226 16068
rect 41782 15988 41788 16040
rect 41840 15988 41846 16040
rect 40359 15932 41368 15960
rect 41417 15963 41475 15969
rect 40359 15929 40371 15932
rect 40313 15923 40371 15929
rect 41417 15929 41429 15963
rect 41463 15929 41475 15963
rect 41417 15923 41475 15929
rect 43916 15960 43944 16068
rect 44545 15963 44603 15969
rect 44545 15960 44557 15963
rect 43916 15932 44557 15960
rect 43916 15904 43944 15932
rect 44545 15929 44557 15932
rect 44591 15960 44603 15963
rect 44913 15963 44971 15969
rect 44913 15960 44925 15963
rect 44591 15932 44925 15960
rect 44591 15929 44603 15932
rect 44545 15923 44603 15929
rect 44913 15929 44925 15932
rect 44959 15929 44971 15963
rect 44913 15923 44971 15929
rect 29564 15864 30972 15892
rect 32950 15852 32956 15904
rect 33008 15892 33014 15904
rect 33229 15895 33287 15901
rect 33229 15892 33241 15895
rect 33008 15864 33241 15892
rect 33008 15852 33014 15864
rect 33229 15861 33241 15864
rect 33275 15861 33287 15895
rect 33229 15855 33287 15861
rect 35066 15852 35072 15904
rect 35124 15892 35130 15904
rect 35253 15895 35311 15901
rect 35253 15892 35265 15895
rect 35124 15864 35265 15892
rect 35124 15852 35130 15864
rect 35253 15861 35265 15864
rect 35299 15861 35311 15895
rect 35253 15855 35311 15861
rect 38194 15852 38200 15904
rect 38252 15892 38258 15904
rect 39758 15892 39764 15904
rect 38252 15864 39764 15892
rect 38252 15852 38258 15864
rect 39758 15852 39764 15864
rect 39816 15892 39822 15904
rect 40221 15895 40279 15901
rect 40221 15892 40233 15895
rect 39816 15864 40233 15892
rect 39816 15852 39822 15864
rect 40221 15861 40233 15864
rect 40267 15861 40279 15895
rect 40221 15855 40279 15861
rect 40494 15852 40500 15904
rect 40552 15892 40558 15904
rect 41141 15895 41199 15901
rect 41141 15892 41153 15895
rect 40552 15864 41153 15892
rect 40552 15852 40558 15864
rect 41141 15861 41153 15864
rect 41187 15861 41199 15895
rect 41141 15855 41199 15861
rect 43898 15852 43904 15904
rect 43956 15852 43962 15904
rect 44269 15895 44327 15901
rect 44269 15861 44281 15895
rect 44315 15892 44327 15895
rect 44358 15892 44364 15904
rect 44315 15864 44364 15892
rect 44315 15861 44327 15864
rect 44269 15855 44327 15861
rect 44358 15852 44364 15864
rect 44416 15852 44422 15904
rect 460 15802 45540 15824
rect 460 15750 3570 15802
rect 3622 15750 3634 15802
rect 3686 15750 3698 15802
rect 3750 15750 3762 15802
rect 3814 15750 3826 15802
rect 3878 15750 8570 15802
rect 8622 15750 8634 15802
rect 8686 15750 8698 15802
rect 8750 15750 8762 15802
rect 8814 15750 8826 15802
rect 8878 15750 13570 15802
rect 13622 15750 13634 15802
rect 13686 15750 13698 15802
rect 13750 15750 13762 15802
rect 13814 15750 13826 15802
rect 13878 15750 18570 15802
rect 18622 15750 18634 15802
rect 18686 15750 18698 15802
rect 18750 15750 18762 15802
rect 18814 15750 18826 15802
rect 18878 15750 23570 15802
rect 23622 15750 23634 15802
rect 23686 15750 23698 15802
rect 23750 15750 23762 15802
rect 23814 15750 23826 15802
rect 23878 15750 28570 15802
rect 28622 15750 28634 15802
rect 28686 15750 28698 15802
rect 28750 15750 28762 15802
rect 28814 15750 28826 15802
rect 28878 15750 33570 15802
rect 33622 15750 33634 15802
rect 33686 15750 33698 15802
rect 33750 15750 33762 15802
rect 33814 15750 33826 15802
rect 33878 15750 38570 15802
rect 38622 15750 38634 15802
rect 38686 15750 38698 15802
rect 38750 15750 38762 15802
rect 38814 15750 38826 15802
rect 38878 15750 43570 15802
rect 43622 15750 43634 15802
rect 43686 15750 43698 15802
rect 43750 15750 43762 15802
rect 43814 15750 43826 15802
rect 43878 15750 45540 15802
rect 460 15728 45540 15750
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4338 15688 4344 15700
rect 4019 15660 4344 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 5810 15688 5816 15700
rect 4448 15660 5816 15688
rect 4448 15484 4476 15660
rect 5810 15648 5816 15660
rect 5868 15688 5874 15700
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 5868 15660 6837 15688
rect 5868 15648 5874 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 10134 15688 10140 15700
rect 6825 15651 6883 15657
rect 8036 15660 10140 15688
rect 7377 15623 7435 15629
rect 7377 15589 7389 15623
rect 7423 15589 7435 15623
rect 7377 15583 7435 15589
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4580 15524 4721 15552
rect 4580 15512 4586 15524
rect 4709 15521 4721 15524
rect 4755 15552 4767 15555
rect 5442 15552 5448 15564
rect 4755 15524 5448 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4448 15456 4629 15484
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4617 15447 4675 15453
rect 4908 15456 5089 15484
rect 4908 15416 4936 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 6638 15484 6644 15496
rect 6486 15456 6644 15484
rect 5077 15447 5135 15453
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7285 15487 7343 15493
rect 7285 15453 7297 15487
rect 7331 15484 7343 15487
rect 7392 15484 7420 15583
rect 8036 15564 8064 15660
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 11514 15688 11520 15700
rect 10520 15660 11520 15688
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 10410 15620 10416 15632
rect 9640 15592 10416 15620
rect 9640 15580 9646 15592
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 9600 15552 9628 15580
rect 8312 15524 9628 15552
rect 7331 15456 7420 15484
rect 7745 15487 7803 15493
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 7745 15453 7757 15487
rect 7791 15484 7803 15487
rect 8110 15484 8116 15496
rect 7791 15456 8116 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8312 15493 8340 15524
rect 9766 15512 9772 15564
rect 9824 15512 9830 15564
rect 8297 15487 8355 15493
rect 8297 15484 8309 15487
rect 8260 15456 8309 15484
rect 8260 15444 8266 15456
rect 8297 15453 8309 15456
rect 8343 15453 8355 15487
rect 9784 15484 9812 15512
rect 9706 15456 9812 15484
rect 8297 15447 8355 15453
rect 5353 15419 5411 15425
rect 5353 15416 5365 15419
rect 4264 15388 4936 15416
rect 5000 15388 5365 15416
rect 3418 15308 3424 15360
rect 3476 15348 3482 15360
rect 4264 15357 4292 15388
rect 5000 15357 5028 15388
rect 5353 15385 5365 15388
rect 5399 15385 5411 15419
rect 8573 15419 8631 15425
rect 8573 15416 8585 15419
rect 5353 15379 5411 15385
rect 7116 15388 8585 15416
rect 7116 15357 7144 15388
rect 8573 15385 8585 15388
rect 8619 15385 8631 15419
rect 10428 15416 10456 15580
rect 10520 15493 10548 15660
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 12676 15660 13584 15688
rect 12676 15648 12682 15660
rect 13556 15629 13584 15660
rect 14182 15648 14188 15700
rect 14240 15648 14246 15700
rect 14550 15648 14556 15700
rect 14608 15648 14614 15700
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 17034 15688 17040 15700
rect 16816 15660 17040 15688
rect 16816 15648 16822 15660
rect 17034 15648 17040 15660
rect 17092 15688 17098 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 17092 15660 17233 15688
rect 17092 15648 17098 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 17328 15660 17816 15688
rect 13449 15623 13507 15629
rect 13449 15620 13461 15623
rect 13188 15592 13461 15620
rect 13188 15561 13216 15592
rect 13449 15589 13461 15592
rect 13495 15589 13507 15623
rect 13449 15583 13507 15589
rect 13541 15623 13599 15629
rect 13541 15589 13553 15623
rect 13587 15589 13599 15623
rect 14568 15620 14596 15648
rect 16669 15623 16727 15629
rect 14568 15592 14964 15620
rect 13541 15583 13599 15589
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 13171 15555 13229 15561
rect 12759 15524 13032 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15453 10655 15487
rect 12250 15484 12256 15496
rect 12006 15456 12256 15484
rect 10597 15447 10655 15453
rect 10612 15416 10640 15447
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 10428 15388 10640 15416
rect 8573 15379 8631 15385
rect 10778 15376 10784 15428
rect 10836 15416 10842 15428
rect 10873 15419 10931 15425
rect 10873 15416 10885 15419
rect 10836 15388 10885 15416
rect 10836 15376 10842 15388
rect 10873 15385 10885 15388
rect 10919 15385 10931 15419
rect 10873 15379 10931 15385
rect 11146 15376 11152 15428
rect 11204 15376 11210 15428
rect 12544 15416 12572 15447
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 13004 15484 13032 15524
rect 13171 15521 13183 15555
rect 13217 15521 13229 15555
rect 13909 15555 13967 15561
rect 13909 15552 13921 15555
rect 13171 15515 13229 15521
rect 13280 15524 13921 15552
rect 13280 15486 13308 15524
rect 13909 15521 13921 15524
rect 13955 15521 13967 15555
rect 14734 15552 14740 15564
rect 13909 15515 13967 15521
rect 14016 15524 14740 15552
rect 13096 15484 13308 15486
rect 13004 15458 13308 15484
rect 13004 15456 13124 15458
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13412 15456 13461 15484
rect 13412 15444 13418 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 14016 15484 14044 15524
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 14936 15561 14964 15592
rect 16669 15589 16681 15623
rect 16715 15620 16727 15623
rect 16850 15620 16856 15632
rect 16715 15592 16856 15620
rect 16715 15589 16727 15592
rect 16669 15583 16727 15589
rect 16850 15580 16856 15592
rect 16908 15620 16914 15632
rect 17328 15620 17356 15660
rect 16908 15592 17356 15620
rect 17405 15623 17463 15629
rect 16908 15580 16914 15592
rect 17405 15589 17417 15623
rect 17451 15589 17463 15623
rect 17405 15583 17463 15589
rect 14921 15555 14979 15561
rect 14921 15521 14933 15555
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15552 15255 15555
rect 15243 15524 16988 15552
rect 15243 15521 15255 15524
rect 15197 15515 15255 15521
rect 13863 15456 14044 15484
rect 14093 15487 14151 15493
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 13924 15428 13952 15456
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 12544 15388 13216 15416
rect 3513 15351 3571 15357
rect 3513 15348 3525 15351
rect 3476 15320 3525 15348
rect 3476 15308 3482 15320
rect 3513 15317 3525 15320
rect 3559 15348 3571 15351
rect 4249 15351 4307 15357
rect 4249 15348 4261 15351
rect 3559 15320 4261 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 4249 15317 4261 15320
rect 4295 15317 4307 15351
rect 4249 15311 4307 15317
rect 4985 15351 5043 15357
rect 4985 15317 4997 15351
rect 5031 15317 5043 15351
rect 4985 15311 5043 15317
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15317 7159 15351
rect 7101 15311 7159 15317
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 9950 15348 9956 15360
rect 7883 15320 9956 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 9950 15308 9956 15320
rect 10008 15348 10014 15360
rect 10045 15351 10103 15357
rect 10045 15348 10057 15351
rect 10008 15320 10057 15348
rect 10008 15308 10014 15320
rect 10045 15317 10057 15320
rect 10091 15317 10103 15351
rect 10045 15311 10103 15317
rect 10321 15351 10379 15357
rect 10321 15317 10333 15351
rect 10367 15348 10379 15351
rect 11164 15348 11192 15376
rect 10367 15320 11192 15348
rect 10367 15317 10379 15320
rect 10321 15311 10379 15317
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 12345 15351 12403 15357
rect 12345 15348 12357 15351
rect 11848 15320 12357 15348
rect 11848 15308 11854 15320
rect 12345 15317 12357 15320
rect 12391 15317 12403 15351
rect 12345 15311 12403 15317
rect 12986 15308 12992 15360
rect 13044 15308 13050 15360
rect 13078 15308 13084 15360
rect 13136 15308 13142 15360
rect 13188 15348 13216 15388
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 13725 15419 13783 15425
rect 13725 15416 13737 15419
rect 13320 15388 13737 15416
rect 13320 15376 13326 15388
rect 13725 15385 13737 15388
rect 13771 15385 13783 15419
rect 13725 15379 13783 15385
rect 13906 15376 13912 15428
rect 13964 15376 13970 15428
rect 14108 15348 14136 15447
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 14826 15444 14832 15496
rect 14884 15444 14890 15496
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 15654 15416 15660 15428
rect 14976 15388 15660 15416
rect 14976 15376 14982 15388
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 16960 15416 16988 15524
rect 17420 15484 17448 15583
rect 17788 15496 17816 15660
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19484 15660 19809 15688
rect 19484 15648 19490 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 19797 15651 19855 15657
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20898 15688 20904 15700
rect 20395 15660 20904 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 21082 15648 21088 15700
rect 21140 15648 21146 15700
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 21637 15691 21695 15697
rect 21637 15688 21649 15691
rect 21508 15660 21649 15688
rect 21508 15648 21514 15660
rect 21637 15657 21649 15660
rect 21683 15657 21695 15691
rect 21637 15651 21695 15657
rect 21910 15648 21916 15700
rect 21968 15688 21974 15700
rect 22554 15688 22560 15700
rect 21968 15660 22560 15688
rect 21968 15648 21974 15660
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23014 15648 23020 15700
rect 23072 15688 23078 15700
rect 25498 15688 25504 15700
rect 23072 15660 25504 15688
rect 23072 15648 23078 15660
rect 25498 15648 25504 15660
rect 25556 15688 25562 15700
rect 25556 15660 27108 15688
rect 25556 15648 25562 15660
rect 19337 15623 19395 15629
rect 19337 15589 19349 15623
rect 19383 15620 19395 15623
rect 20806 15620 20812 15632
rect 19383 15592 20812 15620
rect 19383 15589 19395 15592
rect 19337 15583 19395 15589
rect 20806 15580 20812 15592
rect 20864 15580 20870 15632
rect 22833 15623 22891 15629
rect 21008 15592 22508 15620
rect 21008 15561 21036 15592
rect 22480 15564 22508 15592
rect 22833 15589 22845 15623
rect 22879 15620 22891 15623
rect 23658 15620 23664 15632
rect 22879 15592 23664 15620
rect 22879 15589 22891 15592
rect 22833 15583 22891 15589
rect 23658 15580 23664 15592
rect 23716 15580 23722 15632
rect 26970 15580 26976 15632
rect 27028 15580 27034 15632
rect 27080 15620 27108 15660
rect 27154 15648 27160 15700
rect 27212 15688 27218 15700
rect 27709 15691 27767 15697
rect 27709 15688 27721 15691
rect 27212 15660 27721 15688
rect 27212 15648 27218 15660
rect 27709 15657 27721 15660
rect 27755 15657 27767 15691
rect 28902 15688 28908 15700
rect 27709 15651 27767 15657
rect 28276 15660 28908 15688
rect 28166 15620 28172 15632
rect 27080 15592 28172 15620
rect 28166 15580 28172 15592
rect 28224 15580 28230 15632
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15552 20223 15555
rect 20993 15555 21051 15561
rect 20211 15524 20852 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17420 15456 17693 15484
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17828 15456 17877 15484
rect 17828 15444 17834 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 19886 15484 19892 15496
rect 19659 15456 19892 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15484 20315 15487
rect 20349 15487 20407 15493
rect 20349 15484 20361 15487
rect 20303 15456 20361 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 20349 15453 20361 15456
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 20533 15487 20591 15493
rect 20533 15453 20545 15487
rect 20579 15484 20591 15487
rect 20714 15484 20720 15496
rect 20579 15456 20720 15484
rect 20579 15453 20591 15456
rect 20533 15447 20591 15453
rect 17497 15419 17555 15425
rect 17497 15416 17509 15419
rect 16960 15388 17509 15416
rect 17497 15385 17509 15388
rect 17543 15385 17555 15419
rect 17497 15379 17555 15385
rect 19429 15419 19487 15425
rect 19429 15385 19441 15419
rect 19475 15385 19487 15419
rect 20088 15416 20116 15447
rect 20162 15416 20168 15428
rect 20088 15388 20168 15416
rect 19429 15379 19487 15385
rect 13188 15320 14136 15348
rect 14645 15351 14703 15357
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 15378 15348 15384 15360
rect 14691 15320 15384 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 17218 15348 17224 15360
rect 16540 15320 17224 15348
rect 16540 15308 16546 15320
rect 17218 15308 17224 15320
rect 17276 15308 17282 15360
rect 18325 15351 18383 15357
rect 18325 15317 18337 15351
rect 18371 15348 18383 15351
rect 18414 15348 18420 15360
rect 18371 15320 18420 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 18414 15308 18420 15320
rect 18472 15308 18478 15360
rect 18782 15308 18788 15360
rect 18840 15348 18846 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 18840 15320 18889 15348
rect 18840 15308 18846 15320
rect 18877 15317 18889 15320
rect 18923 15317 18935 15351
rect 19444 15348 19472 15379
rect 20162 15376 20168 15388
rect 20220 15376 20226 15428
rect 20364 15416 20392 15447
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 20824 15493 20852 15524
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 22278 15552 22284 15564
rect 20993 15515 21051 15521
rect 21284 15524 22284 15552
rect 21284 15493 21312 15524
rect 22278 15512 22284 15524
rect 22336 15552 22342 15564
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 22336 15524 22385 15552
rect 22336 15512 22342 15524
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 22373 15515 22431 15521
rect 22462 15512 22468 15564
rect 22520 15512 22526 15564
rect 23290 15512 23296 15564
rect 23348 15512 23354 15564
rect 23382 15512 23388 15564
rect 23440 15512 23446 15564
rect 25501 15555 25559 15561
rect 25501 15552 25513 15555
rect 23676 15524 25513 15552
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15453 20867 15487
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 20809 15447 20867 15453
rect 20916 15456 21281 15484
rect 20916 15416 20944 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 22152 15456 23213 15484
rect 22152 15444 22158 15456
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 23308 15484 23336 15512
rect 23676 15484 23704 15524
rect 25501 15521 25513 15524
rect 25547 15521 25559 15555
rect 25501 15515 25559 15521
rect 25869 15555 25927 15561
rect 25869 15521 25881 15555
rect 25915 15552 25927 15555
rect 26602 15552 26608 15564
rect 25915 15524 26608 15552
rect 25915 15521 25927 15524
rect 25869 15515 25927 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 26988 15552 27016 15580
rect 26988 15524 27476 15552
rect 23308 15456 23704 15484
rect 23753 15487 23811 15493
rect 23201 15447 23259 15453
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 20364 15388 20944 15416
rect 20990 15376 20996 15428
rect 21048 15416 21054 15428
rect 21177 15419 21235 15425
rect 21177 15416 21189 15419
rect 21048 15388 21189 15416
rect 21048 15376 21054 15388
rect 21177 15385 21189 15388
rect 21223 15385 21235 15419
rect 21177 15379 21235 15385
rect 21453 15419 21511 15425
rect 21453 15385 21465 15419
rect 21499 15416 21511 15419
rect 22002 15416 22008 15428
rect 21499 15388 22008 15416
rect 21499 15385 21511 15388
rect 21453 15379 21511 15385
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 22189 15419 22247 15425
rect 22189 15385 22201 15419
rect 22235 15416 22247 15419
rect 22370 15416 22376 15428
rect 22235 15388 22376 15416
rect 22235 15385 22247 15388
rect 22189 15379 22247 15385
rect 22370 15376 22376 15388
rect 22428 15376 22434 15428
rect 20438 15348 20444 15360
rect 19444 15320 20444 15348
rect 18877 15311 18935 15317
rect 20438 15308 20444 15320
rect 20496 15348 20502 15360
rect 21821 15351 21879 15357
rect 21821 15348 21833 15351
rect 20496 15320 21833 15348
rect 20496 15308 20502 15320
rect 21821 15317 21833 15320
rect 21867 15317 21879 15351
rect 21821 15311 21879 15317
rect 22281 15351 22339 15357
rect 22281 15317 22293 15351
rect 22327 15348 22339 15351
rect 23474 15348 23480 15360
rect 22327 15320 23480 15348
rect 22327 15317 22339 15320
rect 22281 15311 22339 15317
rect 23474 15308 23480 15320
rect 23532 15308 23538 15360
rect 23768 15348 23796 15447
rect 25314 15444 25320 15496
rect 25372 15484 25378 15496
rect 25593 15487 25651 15493
rect 25593 15484 25605 15487
rect 25372 15456 25605 15484
rect 25372 15444 25378 15456
rect 25593 15453 25605 15456
rect 25639 15453 25651 15487
rect 25593 15447 25651 15453
rect 24026 15376 24032 15428
rect 24084 15376 24090 15428
rect 26326 15416 26332 15428
rect 25254 15388 26332 15416
rect 26326 15376 26332 15388
rect 26384 15376 26390 15428
rect 26418 15376 26424 15428
rect 26476 15376 26482 15428
rect 27448 15416 27476 15524
rect 27614 15512 27620 15564
rect 27672 15512 27678 15564
rect 27798 15512 27804 15564
rect 27856 15552 27862 15564
rect 28276 15561 28304 15660
rect 28902 15648 28908 15660
rect 28960 15648 28966 15700
rect 29380 15660 29684 15688
rect 28537 15623 28595 15629
rect 28537 15589 28549 15623
rect 28583 15620 28595 15623
rect 28994 15620 29000 15632
rect 28583 15592 29000 15620
rect 28583 15589 28595 15592
rect 28537 15583 28595 15589
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 28261 15555 28319 15561
rect 28261 15552 28273 15555
rect 27856 15524 28273 15552
rect 27856 15512 27862 15524
rect 28261 15521 28273 15524
rect 28307 15521 28319 15555
rect 28261 15515 28319 15521
rect 28828 15524 29316 15552
rect 27632 15484 27660 15512
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 27632 15456 28089 15484
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 28166 15444 28172 15496
rect 28224 15444 28230 15496
rect 28442 15444 28448 15496
rect 28500 15484 28506 15496
rect 28721 15487 28779 15493
rect 28721 15484 28733 15487
rect 28500 15456 28733 15484
rect 28500 15444 28506 15456
rect 28721 15453 28733 15456
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 28828 15416 28856 15524
rect 29086 15444 29092 15496
rect 29144 15484 29150 15496
rect 29288 15493 29316 15524
rect 29380 15493 29408 15660
rect 29656 15552 29684 15660
rect 29730 15648 29736 15700
rect 29788 15688 29794 15700
rect 30193 15691 30251 15697
rect 30193 15688 30205 15691
rect 29788 15660 30205 15688
rect 29788 15648 29794 15660
rect 30193 15657 30205 15660
rect 30239 15657 30251 15691
rect 30193 15651 30251 15657
rect 30650 15648 30656 15700
rect 30708 15648 30714 15700
rect 30837 15691 30895 15697
rect 30837 15657 30849 15691
rect 30883 15688 30895 15691
rect 33134 15688 33140 15700
rect 30883 15660 33140 15688
rect 30883 15657 30895 15660
rect 30837 15651 30895 15657
rect 33134 15648 33140 15660
rect 33192 15648 33198 15700
rect 33410 15648 33416 15700
rect 33468 15688 33474 15700
rect 33689 15691 33747 15697
rect 33689 15688 33701 15691
rect 33468 15660 33701 15688
rect 33468 15648 33474 15660
rect 33689 15657 33701 15660
rect 33735 15657 33747 15691
rect 33689 15651 33747 15657
rect 37918 15648 37924 15700
rect 37976 15648 37982 15700
rect 38286 15648 38292 15700
rect 38344 15648 38350 15700
rect 40494 15648 40500 15700
rect 40552 15648 40558 15700
rect 40678 15648 40684 15700
rect 40736 15688 40742 15700
rect 40957 15691 41015 15697
rect 40957 15688 40969 15691
rect 40736 15660 40969 15688
rect 40736 15648 40742 15660
rect 40957 15657 40969 15660
rect 41003 15657 41015 15691
rect 40957 15651 41015 15657
rect 32214 15580 32220 15632
rect 32272 15620 32278 15632
rect 32858 15620 32864 15632
rect 32272 15592 32864 15620
rect 32272 15580 32278 15592
rect 32858 15580 32864 15592
rect 32916 15620 32922 15632
rect 38930 15620 38936 15632
rect 32916 15592 32996 15620
rect 32916 15580 32922 15592
rect 30650 15552 30656 15564
rect 29656 15524 30656 15552
rect 30650 15512 30656 15524
rect 30708 15512 30714 15564
rect 30926 15512 30932 15564
rect 30984 15512 30990 15564
rect 32968 15561 32996 15592
rect 37246 15592 38936 15620
rect 37246 15564 37274 15592
rect 31205 15555 31263 15561
rect 31205 15521 31217 15555
rect 31251 15552 31263 15555
rect 32769 15555 32827 15561
rect 32769 15552 32781 15555
rect 31251 15524 32781 15552
rect 31251 15521 31263 15524
rect 31205 15515 31263 15521
rect 32769 15521 32781 15524
rect 32815 15521 32827 15555
rect 32769 15515 32827 15521
rect 32953 15555 33011 15561
rect 32953 15521 32965 15555
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 33137 15555 33195 15561
rect 33137 15521 33149 15555
rect 33183 15552 33195 15555
rect 35342 15552 35348 15564
rect 33183 15524 33364 15552
rect 33183 15521 33195 15524
rect 33137 15515 33195 15521
rect 33336 15496 33364 15524
rect 33612 15524 35348 15552
rect 29181 15487 29239 15493
rect 29181 15484 29193 15487
rect 29144 15456 29193 15484
rect 29144 15444 29150 15456
rect 29181 15453 29193 15456
rect 29227 15453 29239 15487
rect 29181 15447 29239 15453
rect 29273 15487 29331 15493
rect 29273 15453 29285 15487
rect 29319 15453 29331 15487
rect 29273 15447 29331 15453
rect 29365 15487 29423 15493
rect 29365 15453 29377 15487
rect 29411 15453 29423 15487
rect 29365 15447 29423 15453
rect 29546 15444 29552 15496
rect 29604 15444 29610 15496
rect 29638 15444 29644 15496
rect 29696 15444 29702 15496
rect 29730 15444 29736 15496
rect 29788 15484 29794 15496
rect 30009 15487 30067 15493
rect 30009 15484 30021 15487
rect 29788 15456 30021 15484
rect 29788 15444 29794 15456
rect 30009 15453 30021 15456
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30098 15444 30104 15496
rect 30156 15444 30162 15496
rect 32306 15444 32312 15496
rect 32364 15444 32370 15496
rect 33045 15487 33103 15493
rect 33045 15453 33057 15487
rect 33091 15453 33103 15487
rect 33045 15447 33103 15453
rect 33229 15487 33287 15493
rect 33229 15453 33241 15487
rect 33275 15453 33287 15487
rect 33229 15447 33287 15453
rect 27448 15388 28856 15416
rect 28905 15419 28963 15425
rect 28905 15385 28917 15419
rect 28951 15416 28963 15419
rect 29825 15419 29883 15425
rect 29825 15416 29837 15419
rect 28951 15388 29837 15416
rect 28951 15385 28963 15388
rect 28905 15379 28963 15385
rect 29825 15385 29837 15388
rect 29871 15385 29883 15419
rect 29825 15379 29883 15385
rect 29917 15419 29975 15425
rect 29917 15385 29929 15419
rect 29963 15416 29975 15419
rect 30116 15416 30144 15444
rect 29963 15388 30144 15416
rect 29963 15385 29975 15388
rect 29917 15379 29975 15385
rect 24854 15348 24860 15360
rect 23768 15320 24860 15348
rect 24854 15308 24860 15320
rect 24912 15348 24918 15360
rect 25314 15348 25320 15360
rect 24912 15320 25320 15348
rect 24912 15308 24918 15320
rect 25314 15308 25320 15320
rect 25372 15308 25378 15360
rect 25498 15308 25504 15360
rect 25556 15348 25562 15360
rect 25774 15348 25780 15360
rect 25556 15320 25780 15348
rect 25556 15308 25562 15320
rect 25774 15308 25780 15320
rect 25832 15308 25838 15360
rect 26510 15308 26516 15360
rect 26568 15348 26574 15360
rect 27154 15348 27160 15360
rect 26568 15320 27160 15348
rect 26568 15308 26574 15320
rect 27154 15308 27160 15320
rect 27212 15348 27218 15360
rect 27341 15351 27399 15357
rect 27341 15348 27353 15351
rect 27212 15320 27353 15348
rect 27212 15308 27218 15320
rect 27341 15317 27353 15320
rect 27387 15317 27399 15351
rect 27341 15311 27399 15317
rect 28810 15308 28816 15360
rect 28868 15348 28874 15360
rect 29730 15348 29736 15360
rect 28868 15320 29736 15348
rect 28868 15308 28874 15320
rect 29730 15308 29736 15320
rect 29788 15308 29794 15360
rect 29840 15348 29868 15379
rect 30190 15376 30196 15428
rect 30248 15376 30254 15428
rect 30466 15376 30472 15428
rect 30524 15376 30530 15428
rect 33060 15416 33088 15447
rect 32692 15388 33088 15416
rect 30208 15348 30236 15376
rect 29840 15320 30236 15348
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 30679 15351 30737 15357
rect 30679 15348 30691 15351
rect 30432 15320 30691 15348
rect 30432 15308 30438 15320
rect 30679 15317 30691 15320
rect 30725 15348 30737 15351
rect 31846 15348 31852 15360
rect 30725 15320 31852 15348
rect 30725 15317 30737 15320
rect 30679 15311 30737 15317
rect 31846 15308 31852 15320
rect 31904 15308 31910 15360
rect 32582 15308 32588 15360
rect 32640 15348 32646 15360
rect 32692 15357 32720 15388
rect 32677 15351 32735 15357
rect 32677 15348 32689 15351
rect 32640 15320 32689 15348
rect 32640 15308 32646 15320
rect 32677 15317 32689 15320
rect 32723 15317 32735 15351
rect 32677 15311 32735 15317
rect 32766 15308 32772 15360
rect 32824 15348 32830 15360
rect 33244 15348 33272 15447
rect 33318 15444 33324 15496
rect 33376 15444 33382 15496
rect 33612 15493 33640 15524
rect 35342 15512 35348 15524
rect 35400 15512 35406 15564
rect 35897 15555 35955 15561
rect 35897 15521 35909 15555
rect 35943 15552 35955 15555
rect 36630 15552 36636 15564
rect 35943 15524 36636 15552
rect 35943 15521 35955 15524
rect 35897 15515 35955 15521
rect 36630 15512 36636 15524
rect 36688 15512 36694 15564
rect 37182 15512 37188 15564
rect 37240 15524 37274 15564
rect 38856 15561 38884 15592
rect 38930 15580 38936 15592
rect 38988 15580 38994 15632
rect 38841 15555 38899 15561
rect 37240 15512 37246 15524
rect 38841 15521 38853 15555
rect 38887 15521 38899 15555
rect 38841 15515 38899 15521
rect 39485 15555 39543 15561
rect 39485 15521 39497 15555
rect 39531 15552 39543 15555
rect 40512 15552 40540 15648
rect 40770 15580 40776 15632
rect 40828 15620 40834 15632
rect 42242 15620 42248 15632
rect 40828 15592 42248 15620
rect 40828 15580 40834 15592
rect 42242 15580 42248 15592
rect 42300 15580 42306 15632
rect 39531 15524 40540 15552
rect 39531 15521 39543 15524
rect 39485 15515 39543 15521
rect 41414 15512 41420 15564
rect 41472 15552 41478 15564
rect 41877 15555 41935 15561
rect 41877 15552 41889 15555
rect 41472 15524 41889 15552
rect 41472 15512 41478 15524
rect 41877 15521 41889 15524
rect 41923 15552 41935 15555
rect 42058 15552 42064 15564
rect 41923 15524 42064 15552
rect 41923 15521 41935 15524
rect 41877 15515 41935 15521
rect 42058 15512 42064 15524
rect 42116 15512 42122 15564
rect 42702 15512 42708 15564
rect 42760 15512 42766 15564
rect 33597 15487 33655 15493
rect 33597 15453 33609 15487
rect 33643 15453 33655 15487
rect 33597 15447 33655 15453
rect 33870 15444 33876 15496
rect 33928 15444 33934 15496
rect 34054 15444 34060 15496
rect 34112 15444 34118 15496
rect 38194 15444 38200 15496
rect 38252 15484 38258 15496
rect 38657 15487 38715 15493
rect 38657 15484 38669 15487
rect 38252 15456 38669 15484
rect 38252 15444 38258 15456
rect 38657 15453 38669 15456
rect 38703 15453 38715 15487
rect 38657 15447 38715 15453
rect 38746 15444 38752 15496
rect 38804 15484 38810 15496
rect 39114 15484 39120 15496
rect 38804 15456 39120 15484
rect 38804 15444 38810 15456
rect 39114 15444 39120 15456
rect 39172 15484 39178 15496
rect 39209 15487 39267 15493
rect 39209 15484 39221 15487
rect 39172 15456 39221 15484
rect 39172 15444 39178 15456
rect 39209 15453 39221 15456
rect 39255 15453 39267 15487
rect 39209 15447 39267 15453
rect 41233 15487 41291 15493
rect 41233 15453 41245 15487
rect 41279 15484 41291 15487
rect 41279 15456 41368 15484
rect 41279 15453 41291 15456
rect 41233 15447 41291 15453
rect 34333 15419 34391 15425
rect 34333 15416 34345 15419
rect 33428 15388 34345 15416
rect 33428 15357 33456 15388
rect 34333 15385 34345 15388
rect 34379 15385 34391 15419
rect 36173 15419 36231 15425
rect 34333 15379 34391 15385
rect 34716 15388 34822 15416
rect 34716 15360 34744 15388
rect 36173 15385 36185 15419
rect 36219 15416 36231 15419
rect 36446 15416 36452 15428
rect 36219 15388 36452 15416
rect 36219 15385 36231 15388
rect 36173 15379 36231 15385
rect 36446 15376 36452 15388
rect 36504 15376 36510 15428
rect 37550 15416 37556 15428
rect 37398 15388 37556 15416
rect 37550 15376 37556 15388
rect 37608 15376 37614 15428
rect 37737 15419 37795 15425
rect 37737 15416 37749 15419
rect 37660 15388 37749 15416
rect 37660 15360 37688 15388
rect 37737 15385 37749 15388
rect 37783 15385 37795 15419
rect 37737 15379 37795 15385
rect 37953 15419 38011 15425
rect 37953 15385 37965 15419
rect 37999 15416 38011 15419
rect 37999 15388 39896 15416
rect 37999 15385 38011 15388
rect 37953 15379 38011 15385
rect 39868 15360 39896 15388
rect 40034 15376 40040 15428
rect 40092 15376 40098 15428
rect 32824 15320 33272 15348
rect 33413 15351 33471 15357
rect 32824 15308 32830 15320
rect 33413 15317 33425 15351
rect 33459 15317 33471 15351
rect 33413 15311 33471 15317
rect 34698 15308 34704 15360
rect 34756 15308 34762 15360
rect 35802 15308 35808 15360
rect 35860 15308 35866 15360
rect 37642 15308 37648 15360
rect 37700 15308 37706 15360
rect 38102 15308 38108 15360
rect 38160 15308 38166 15360
rect 38749 15351 38807 15357
rect 38749 15317 38761 15351
rect 38795 15348 38807 15351
rect 39114 15348 39120 15360
rect 38795 15320 39120 15348
rect 38795 15317 38807 15320
rect 38749 15311 38807 15317
rect 39114 15308 39120 15320
rect 39172 15308 39178 15360
rect 39850 15308 39856 15360
rect 39908 15308 39914 15360
rect 41046 15308 41052 15360
rect 41104 15308 41110 15360
rect 41340 15357 41368 15456
rect 41690 15444 41696 15496
rect 41748 15444 41754 15496
rect 42794 15444 42800 15496
rect 42852 15484 42858 15496
rect 43165 15487 43223 15493
rect 43165 15484 43177 15487
rect 42852 15456 43177 15484
rect 42852 15444 42858 15456
rect 43165 15453 43177 15456
rect 43211 15453 43223 15487
rect 43165 15447 43223 15453
rect 43438 15444 43444 15496
rect 43496 15484 43502 15496
rect 44913 15487 44971 15493
rect 44913 15484 44925 15487
rect 43496 15456 44925 15484
rect 43496 15444 43502 15456
rect 44913 15453 44925 15456
rect 44959 15453 44971 15487
rect 44913 15447 44971 15453
rect 45002 15444 45008 15496
rect 45060 15444 45066 15496
rect 41785 15419 41843 15425
rect 41785 15416 41797 15419
rect 41524 15388 41797 15416
rect 41524 15360 41552 15388
rect 41785 15385 41797 15388
rect 41831 15385 41843 15419
rect 41785 15379 41843 15385
rect 42521 15419 42579 15425
rect 42521 15385 42533 15419
rect 42567 15416 42579 15419
rect 45020 15416 45048 15444
rect 42567 15388 45048 15416
rect 42567 15385 42579 15388
rect 42521 15379 42579 15385
rect 41325 15351 41383 15357
rect 41325 15317 41337 15351
rect 41371 15317 41383 15351
rect 41325 15311 41383 15317
rect 41506 15308 41512 15360
rect 41564 15308 41570 15360
rect 41598 15308 41604 15360
rect 41656 15348 41662 15360
rect 42153 15351 42211 15357
rect 42153 15348 42165 15351
rect 41656 15320 42165 15348
rect 41656 15308 41662 15320
rect 42153 15317 42165 15320
rect 42199 15317 42211 15351
rect 42153 15311 42211 15317
rect 42610 15308 42616 15360
rect 42668 15308 42674 15360
rect 42978 15308 42984 15360
rect 43036 15308 43042 15360
rect 43070 15308 43076 15360
rect 43128 15348 43134 15360
rect 43441 15351 43499 15357
rect 43441 15348 43453 15351
rect 43128 15320 43453 15348
rect 43128 15308 43134 15320
rect 43441 15317 43453 15320
rect 43487 15317 43499 15351
rect 43441 15311 43499 15317
rect 43898 15308 43904 15360
rect 43956 15308 43962 15360
rect 44358 15308 44364 15360
rect 44416 15348 44422 15360
rect 44545 15351 44603 15357
rect 44545 15348 44557 15351
rect 44416 15320 44557 15348
rect 44416 15308 44422 15320
rect 44545 15317 44557 15320
rect 44591 15317 44603 15351
rect 44545 15311 44603 15317
rect 460 15258 45540 15280
rect 460 15206 6070 15258
rect 6122 15206 6134 15258
rect 6186 15206 6198 15258
rect 6250 15206 6262 15258
rect 6314 15206 6326 15258
rect 6378 15206 11070 15258
rect 11122 15206 11134 15258
rect 11186 15206 11198 15258
rect 11250 15206 11262 15258
rect 11314 15206 11326 15258
rect 11378 15206 16070 15258
rect 16122 15206 16134 15258
rect 16186 15206 16198 15258
rect 16250 15206 16262 15258
rect 16314 15206 16326 15258
rect 16378 15206 21070 15258
rect 21122 15206 21134 15258
rect 21186 15206 21198 15258
rect 21250 15206 21262 15258
rect 21314 15206 21326 15258
rect 21378 15206 26070 15258
rect 26122 15206 26134 15258
rect 26186 15206 26198 15258
rect 26250 15206 26262 15258
rect 26314 15206 26326 15258
rect 26378 15206 31070 15258
rect 31122 15206 31134 15258
rect 31186 15206 31198 15258
rect 31250 15206 31262 15258
rect 31314 15206 31326 15258
rect 31378 15206 36070 15258
rect 36122 15206 36134 15258
rect 36186 15206 36198 15258
rect 36250 15206 36262 15258
rect 36314 15206 36326 15258
rect 36378 15206 41070 15258
rect 41122 15206 41134 15258
rect 41186 15206 41198 15258
rect 41250 15206 41262 15258
rect 41314 15206 41326 15258
rect 41378 15206 45540 15258
rect 460 15184 45540 15206
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 4338 15144 4344 15156
rect 4019 15116 4344 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 4663 15116 6040 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 6012 15085 6040 15116
rect 9766 15104 9772 15156
rect 9824 15104 9830 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10318 15144 10324 15156
rect 10008 15116 10324 15144
rect 10008 15104 10014 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 11606 15144 11612 15156
rect 11256 15116 11612 15144
rect 5997 15079 6055 15085
rect 5997 15045 6009 15079
rect 6043 15045 6055 15079
rect 5997 15039 6055 15045
rect 6638 15036 6644 15088
rect 6696 15036 6702 15088
rect 8021 15079 8079 15085
rect 8021 15045 8033 15079
rect 8067 15076 8079 15079
rect 8294 15076 8300 15088
rect 8067 15048 8300 15076
rect 8067 15045 8079 15048
rect 8021 15039 8079 15045
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 9784 15076 9812 15104
rect 10597 15079 10655 15085
rect 10597 15076 10609 15079
rect 9246 15048 10609 15076
rect 10597 15045 10609 15048
rect 10643 15045 10655 15079
rect 10597 15039 10655 15045
rect 934 14968 940 15020
rect 992 14968 998 15020
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4448 14872 4476 14971
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 4580 14980 4629 15008
rect 4580 14968 4586 14980
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 4755 14980 4844 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 4816 14952 4844 14980
rect 4890 14968 4896 15020
rect 4948 15006 4954 15020
rect 11256 15017 11284 15116
rect 11606 15104 11612 15116
rect 11664 15144 11670 15156
rect 13262 15144 13268 15156
rect 11664 15116 13268 15144
rect 11664 15104 11670 15116
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 14277 15147 14335 15153
rect 14277 15113 14289 15147
rect 14323 15144 14335 15147
rect 14550 15144 14556 15156
rect 14323 15116 14556 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 14826 15104 14832 15156
rect 14884 15144 14890 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 14884 15116 15117 15144
rect 14884 15104 14890 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 15105 15107 15163 15113
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 15519 15116 17325 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 18230 15104 18236 15156
rect 18288 15104 18294 15156
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 20671 15116 22600 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 16850 15076 16856 15088
rect 12860 15048 13952 15076
rect 12860 15036 12866 15048
rect 5077 15011 5135 15017
rect 5077 15006 5089 15011
rect 4948 14978 5089 15006
rect 4948 14968 4954 14978
rect 5077 14977 5089 14978
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 11241 15011 11299 15017
rect 5307 14980 5672 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 5644 14952 5672 14980
rect 9508 14980 10272 15008
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5031 14932 5120 14940
rect 5031 14912 5304 14932
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5092 14904 5304 14912
rect 4893 14875 4951 14881
rect 4893 14872 4905 14875
rect 4448 14844 4905 14872
rect 4893 14841 4905 14844
rect 4939 14841 4951 14875
rect 4893 14835 4951 14841
rect 5276 14872 5304 14904
rect 5626 14900 5632 14952
rect 5684 14900 5690 14952
rect 5718 14900 5724 14952
rect 5776 14900 5782 14952
rect 7742 14900 7748 14952
rect 7800 14900 7806 14952
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 9030 14940 9036 14952
rect 8168 14912 9036 14940
rect 8168 14900 8174 14912
rect 9030 14900 9036 14912
rect 9088 14940 9094 14952
rect 9508 14949 9536 14980
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 9088 14912 9505 14940
rect 9088 14900 9094 14912
rect 9493 14909 9505 14912
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 5276 14844 5580 14872
rect 750 14764 756 14816
rect 808 14764 814 14816
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 5276 14813 5304 14844
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 4672 14776 4813 14804
rect 4672 14764 4678 14776
rect 4801 14773 4813 14776
rect 4847 14773 4859 14807
rect 4801 14767 4859 14773
rect 5261 14807 5319 14813
rect 5261 14773 5273 14807
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5442 14764 5448 14816
rect 5500 14764 5506 14816
rect 5552 14804 5580 14844
rect 10060 14816 10088 14903
rect 10134 14900 10140 14952
rect 10192 14900 10198 14952
rect 10244 14940 10272 14980
rect 11241 14977 11253 15011
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 11422 14968 11428 15020
rect 11480 14968 11486 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 11931 14980 12449 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 13078 14968 13084 15020
rect 13136 14968 13142 15020
rect 13170 14968 13176 15020
rect 13228 14968 13234 15020
rect 13924 15017 13952 15048
rect 16132 15048 16528 15076
rect 13909 15011 13967 15017
rect 13909 14977 13921 15011
rect 13955 15008 13967 15011
rect 14090 15008 14096 15020
rect 13955 14980 14096 15008
rect 13955 14977 13967 14980
rect 13909 14971 13967 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 16132 15017 16160 15048
rect 16500 15020 16528 15048
rect 16592 15048 16856 15076
rect 16117 15011 16175 15017
rect 14240 14980 15884 15008
rect 14240 14968 14246 14980
rect 12161 14943 12219 14949
rect 10244 14912 11928 14940
rect 11900 14816 11928 14912
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12342 14940 12348 14952
rect 12207 14912 12348 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 15580 14872 15608 14903
rect 15746 14900 15752 14952
rect 15804 14900 15810 14952
rect 15856 14940 15884 14980
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16206 14968 16212 15020
rect 16264 14968 16270 15020
rect 16482 14968 16488 15020
rect 16540 14968 16546 15020
rect 16592 15017 16620 15048
rect 16850 15036 16856 15048
rect 16908 15076 16914 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16908 15048 16957 15076
rect 16908 15036 16914 15048
rect 16945 15045 16957 15048
rect 16991 15045 17003 15079
rect 16945 15039 17003 15045
rect 17126 15036 17132 15088
rect 17184 15085 17190 15088
rect 17184 15079 17203 15085
rect 17191 15045 17203 15079
rect 17494 15076 17500 15088
rect 17184 15039 17203 15045
rect 17236 15048 17500 15076
rect 17184 15036 17190 15039
rect 16577 15011 16635 15017
rect 16577 14977 16589 15011
rect 16623 14977 16635 15011
rect 17236 15008 17264 15048
rect 17494 15036 17500 15048
rect 17552 15036 17558 15088
rect 16577 14971 16635 14977
rect 16776 14980 17264 15008
rect 17405 15011 17463 15017
rect 16224 14940 16252 14968
rect 15856 14912 16252 14940
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16776 14940 16804 14980
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 18248 15008 18276 15104
rect 22572 15085 22600 15116
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22704 15116 22937 15144
rect 22704 15104 22710 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 23382 15144 23388 15156
rect 22925 15107 22983 15113
rect 23032 15116 23388 15144
rect 22557 15079 22615 15085
rect 20548 15048 21588 15076
rect 17451 14980 18276 15008
rect 19797 15011 19855 15017
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 19978 15008 19984 15020
rect 19843 14980 19984 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20548 15017 20576 15048
rect 21560 15020 21588 15048
rect 22557 15045 22569 15079
rect 22603 15045 22615 15079
rect 22557 15039 22615 15045
rect 22741 15079 22799 15085
rect 22741 15045 22753 15079
rect 22787 15076 22799 15079
rect 23032 15076 23060 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15113 23535 15147
rect 23477 15107 23535 15113
rect 23492 15076 23520 15107
rect 23658 15104 23664 15156
rect 23716 15104 23722 15156
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 23934 15144 23940 15156
rect 23891 15116 23940 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 24305 15147 24363 15153
rect 24305 15144 24317 15147
rect 24084 15116 24317 15144
rect 24084 15104 24090 15116
rect 24305 15113 24317 15116
rect 24351 15113 24363 15147
rect 24305 15107 24363 15113
rect 24394 15104 24400 15156
rect 24452 15144 24458 15156
rect 25222 15144 25228 15156
rect 24452 15116 25228 15144
rect 24452 15104 24458 15116
rect 25222 15104 25228 15116
rect 25280 15104 25286 15156
rect 25406 15104 25412 15156
rect 25464 15104 25470 15156
rect 25501 15147 25559 15153
rect 25501 15113 25513 15147
rect 25547 15144 25559 15147
rect 26510 15144 26516 15156
rect 25547 15116 26516 15144
rect 25547 15113 25559 15116
rect 25501 15107 25559 15113
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 26602 15104 26608 15156
rect 26660 15104 26666 15156
rect 26786 15144 26792 15156
rect 26712 15116 26792 15144
rect 22787 15048 23060 15076
rect 23124 15048 23520 15076
rect 23676 15076 23704 15104
rect 25424 15076 25452 15104
rect 23676 15048 24532 15076
rect 22787 15045 22799 15048
rect 22741 15039 22799 15045
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20128 14980 20361 15008
rect 20128 14968 20134 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 20714 14968 20720 15020
rect 20772 14968 20778 15020
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 16347 14912 16804 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16850 14900 16856 14952
rect 16908 14900 16914 14952
rect 17954 14900 17960 14952
rect 18012 14900 18018 14952
rect 16761 14875 16819 14881
rect 16761 14872 16773 14875
rect 15580 14844 16773 14872
rect 16761 14841 16773 14844
rect 16807 14872 16819 14875
rect 17972 14872 18000 14900
rect 16807 14844 18000 14872
rect 16807 14841 16819 14844
rect 16761 14835 16819 14841
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 18601 14875 18659 14881
rect 18601 14872 18613 14875
rect 18472 14844 18613 14872
rect 18472 14832 18478 14844
rect 18601 14841 18613 14844
rect 18647 14872 18659 14875
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 18647 14844 18981 14872
rect 18647 14841 18659 14844
rect 18601 14835 18659 14841
rect 18969 14841 18981 14844
rect 19015 14872 19027 14875
rect 19705 14875 19763 14881
rect 19705 14872 19717 14875
rect 19015 14844 19717 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 19705 14841 19717 14844
rect 19751 14872 19763 14875
rect 20732 14872 20760 14968
rect 20824 14940 20852 14971
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20956 14980 21005 15008
rect 20956 14968 20962 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 21450 15008 21456 15020
rect 21315 14980 21456 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 21542 14968 21548 15020
rect 21600 14968 21606 15020
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22186 15008 22192 15020
rect 22143 14980 22192 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22186 14968 22192 14980
rect 22244 15008 22250 15020
rect 23124 15017 23152 15048
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22244 14980 22385 15008
rect 22244 14968 22250 14980
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 21174 14940 21180 14952
rect 20824 14912 21180 14940
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 21361 14875 21419 14881
rect 21361 14872 21373 14875
rect 19751 14844 20484 14872
rect 20732 14844 21373 14872
rect 19751 14841 19763 14844
rect 19705 14835 19763 14841
rect 20456 14816 20484 14844
rect 21361 14841 21373 14844
rect 21407 14872 21419 14875
rect 21910 14872 21916 14884
rect 21407 14844 21916 14872
rect 21407 14841 21419 14844
rect 21361 14835 21419 14841
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 22296 14872 22324 14903
rect 22554 14900 22560 14952
rect 22612 14940 22618 14952
rect 23216 14940 23244 14971
rect 23382 14968 23388 15020
rect 23440 14968 23446 15020
rect 24394 15008 24400 15020
rect 23492 14980 24400 15008
rect 22612 14912 23244 14940
rect 22612 14900 22618 14912
rect 22462 14872 22468 14884
rect 22296 14844 22468 14872
rect 22462 14832 22468 14844
rect 22520 14872 22526 14884
rect 23492 14872 23520 14980
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 24504 15017 24532 15048
rect 25056 15048 25452 15076
rect 25056 15017 25084 15048
rect 25774 15036 25780 15088
rect 25832 15076 25838 15088
rect 26712 15076 26740 15116
rect 26786 15104 26792 15116
rect 26844 15104 26850 15156
rect 27154 15104 27160 15156
rect 27212 15104 27218 15156
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 29362 15144 29368 15156
rect 27663 15116 29368 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 29362 15104 29368 15116
rect 29420 15144 29426 15156
rect 30006 15144 30012 15156
rect 29420 15116 30012 15144
rect 29420 15104 29426 15116
rect 30006 15104 30012 15116
rect 30064 15104 30070 15156
rect 30466 15104 30472 15156
rect 30524 15104 30530 15156
rect 30650 15104 30656 15156
rect 30708 15104 30714 15156
rect 31849 15147 31907 15153
rect 31849 15144 31861 15147
rect 31726 15116 31861 15144
rect 25832 15048 26188 15076
rect 25832 15036 25838 15048
rect 26160 15017 26188 15048
rect 26620 15048 26740 15076
rect 27172 15076 27200 15104
rect 30193 15079 30251 15085
rect 30193 15076 30205 15079
rect 27172 15048 28028 15076
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 14977 25099 15011
rect 26145 15011 26203 15017
rect 25041 14971 25099 14977
rect 25148 14980 25820 15008
rect 23937 14943 23995 14949
rect 23937 14909 23949 14943
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 24029 14943 24087 14949
rect 24029 14909 24041 14943
rect 24075 14940 24087 14943
rect 24210 14940 24216 14952
rect 24075 14912 24216 14940
rect 24075 14909 24087 14912
rect 24029 14903 24087 14909
rect 22520 14844 23520 14872
rect 23952 14872 23980 14903
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 24118 14872 24124 14884
rect 23952 14844 24124 14872
rect 22520 14832 22526 14844
rect 24118 14832 24124 14844
rect 24176 14872 24182 14884
rect 24780 14872 24808 14900
rect 25148 14881 25176 14980
rect 25406 14900 25412 14952
rect 25464 14940 25470 14952
rect 25593 14943 25651 14949
rect 25593 14940 25605 14943
rect 25464 14912 25605 14940
rect 25464 14900 25470 14912
rect 25593 14909 25605 14912
rect 25639 14909 25651 14943
rect 25593 14903 25651 14909
rect 25682 14900 25688 14952
rect 25740 14900 25746 14952
rect 25133 14875 25191 14881
rect 24176 14844 24532 14872
rect 24780 14844 25084 14872
rect 24176 14832 24182 14844
rect 24504 14816 24532 14844
rect 7469 14807 7527 14813
rect 7469 14804 7481 14807
rect 5552 14776 7481 14804
rect 7469 14773 7481 14776
rect 7515 14773 7527 14807
rect 7469 14767 7527 14773
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 9585 14807 9643 14813
rect 9585 14804 9597 14807
rect 8260 14776 9597 14804
rect 8260 14764 8266 14776
rect 9585 14773 9597 14776
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 11882 14764 11888 14816
rect 11940 14764 11946 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 13320 14776 13645 14804
rect 13320 14764 13326 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 14366 14764 14372 14816
rect 14424 14804 14430 14816
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 14424 14776 14565 14804
rect 14424 14764 14430 14776
rect 14553 14773 14565 14776
rect 14599 14804 14611 14807
rect 14918 14804 14924 14816
rect 14599 14776 14924 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16666 14804 16672 14816
rect 15896 14776 16672 14804
rect 15896 14764 15902 14776
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 17129 14807 17187 14813
rect 17129 14804 17141 14807
rect 17092 14776 17141 14804
rect 17092 14764 17098 14776
rect 17129 14773 17141 14776
rect 17175 14773 17187 14807
rect 17129 14767 17187 14773
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 18138 14804 18144 14816
rect 17644 14776 18144 14804
rect 17644 14764 17650 14776
rect 18138 14764 18144 14776
rect 18196 14804 18202 14816
rect 18782 14804 18788 14816
rect 18196 14776 18788 14804
rect 18196 14764 18202 14776
rect 18782 14764 18788 14776
rect 18840 14804 18846 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 18840 14776 19349 14804
rect 18840 14764 18846 14776
rect 19337 14773 19349 14776
rect 19383 14804 19395 14807
rect 19426 14804 19432 14816
rect 19383 14776 19432 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19886 14764 19892 14816
rect 19944 14804 19950 14816
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19944 14776 19993 14804
rect 19944 14764 19950 14776
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 19981 14767 20039 14773
rect 20162 14764 20168 14816
rect 20220 14764 20226 14816
rect 20438 14764 20444 14816
rect 20496 14764 20502 14816
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 20990 14804 20996 14816
rect 20855 14776 20996 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 22830 14764 22836 14816
rect 22888 14804 22894 14816
rect 23293 14807 23351 14813
rect 23293 14804 23305 14807
rect 22888 14776 23305 14804
rect 22888 14764 22894 14776
rect 23293 14773 23305 14776
rect 23339 14804 23351 14807
rect 23934 14804 23940 14816
rect 23339 14776 23940 14804
rect 23339 14773 23351 14776
rect 23293 14767 23351 14773
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 24486 14764 24492 14816
rect 24544 14764 24550 14816
rect 24854 14764 24860 14816
rect 24912 14764 24918 14816
rect 25056 14804 25084 14844
rect 25133 14841 25145 14875
rect 25179 14841 25191 14875
rect 25792 14872 25820 14980
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26234 14968 26240 15020
rect 26292 15008 26298 15020
rect 26513 15011 26571 15017
rect 26513 15008 26525 15011
rect 26292 14980 26525 15008
rect 26292 14968 26298 14980
rect 26513 14977 26525 14980
rect 26559 14977 26571 15011
rect 26513 14971 26571 14977
rect 26620 14952 26648 15048
rect 26789 15011 26847 15017
rect 26789 15008 26801 15011
rect 26712 14980 26801 15008
rect 26602 14900 26608 14952
rect 26660 14900 26666 14952
rect 26712 14872 26740 14980
rect 26789 14977 26801 14980
rect 26835 14977 26847 15011
rect 26789 14971 26847 14977
rect 27062 14968 27068 15020
rect 27120 14968 27126 15020
rect 27154 14968 27160 15020
rect 27212 14968 27218 15020
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 27890 14968 27896 15020
rect 27948 14968 27954 15020
rect 28000 15017 28028 15048
rect 28092 15048 30205 15076
rect 28092 15017 28120 15048
rect 30193 15045 30205 15048
rect 30239 15045 30251 15079
rect 30193 15039 30251 15045
rect 30282 15036 30288 15088
rect 30340 15036 30346 15088
rect 30484 15076 30512 15104
rect 30929 15079 30987 15085
rect 30929 15076 30941 15079
rect 30484 15048 30941 15076
rect 30929 15045 30941 15048
rect 30975 15076 30987 15079
rect 31018 15076 31024 15088
rect 30975 15048 31024 15076
rect 30975 15045 30987 15048
rect 30929 15039 30987 15045
rect 31018 15036 31024 15048
rect 31076 15036 31082 15088
rect 31573 15079 31631 15085
rect 31159 15045 31217 15051
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 28258 14968 28264 15020
rect 28316 14968 28322 15020
rect 28620 15011 28678 15017
rect 28620 14977 28632 15011
rect 28666 15008 28678 15011
rect 29638 15008 29644 15020
rect 28666 14980 29644 15008
rect 28666 14977 28678 14980
rect 28620 14971 28678 14977
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 29825 15011 29883 15017
rect 29825 15008 29837 15011
rect 29748 14980 29837 15008
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 28350 14940 28356 14952
rect 26936 14912 28356 14940
rect 26936 14900 26942 14912
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 25792 14844 26740 14872
rect 25133 14835 25191 14841
rect 25406 14804 25412 14816
rect 25056 14776 25412 14804
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 25958 14764 25964 14816
rect 26016 14764 26022 14816
rect 26329 14807 26387 14813
rect 26329 14773 26341 14807
rect 26375 14804 26387 14807
rect 26418 14804 26424 14816
rect 26375 14776 26424 14804
rect 26375 14773 26387 14776
rect 26329 14767 26387 14773
rect 26418 14764 26424 14776
rect 26476 14764 26482 14816
rect 26878 14764 26884 14816
rect 26936 14764 26942 14816
rect 27522 14764 27528 14816
rect 27580 14764 27586 14816
rect 28166 14764 28172 14816
rect 28224 14804 28230 14816
rect 29748 14813 29776 14980
rect 29825 14977 29837 14980
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 29914 14968 29920 15020
rect 29972 15008 29978 15020
rect 30009 15011 30067 15017
rect 30009 15008 30021 15011
rect 29972 14980 30021 15008
rect 29972 14968 29978 14980
rect 30009 14977 30021 14980
rect 30055 15008 30067 15011
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 30055 14980 30481 15008
rect 30055 14977 30067 14980
rect 30009 14971 30067 14977
rect 30469 14977 30481 14980
rect 30515 14977 30527 15011
rect 31159 15011 31171 15045
rect 31205 15011 31217 15045
rect 31573 15045 31585 15079
rect 31619 15076 31631 15079
rect 31726 15076 31754 15116
rect 31849 15113 31861 15116
rect 31895 15113 31907 15147
rect 31849 15107 31907 15113
rect 32674 15104 32680 15156
rect 32732 15104 32738 15156
rect 33870 15104 33876 15156
rect 33928 15144 33934 15156
rect 34333 15147 34391 15153
rect 34333 15144 34345 15147
rect 33928 15116 34345 15144
rect 33928 15104 33934 15116
rect 34333 15113 34345 15116
rect 34379 15113 34391 15147
rect 34333 15107 34391 15113
rect 34701 15147 34759 15153
rect 34701 15113 34713 15147
rect 34747 15144 34759 15147
rect 35066 15144 35072 15156
rect 34747 15116 35072 15144
rect 34747 15113 34759 15116
rect 34701 15107 34759 15113
rect 35066 15104 35072 15116
rect 35124 15104 35130 15156
rect 35161 15147 35219 15153
rect 35161 15113 35173 15147
rect 35207 15144 35219 15147
rect 35342 15144 35348 15156
rect 35207 15116 35348 15144
rect 35207 15113 35219 15116
rect 35161 15107 35219 15113
rect 35342 15104 35348 15116
rect 35400 15104 35406 15156
rect 35529 15147 35587 15153
rect 35529 15113 35541 15147
rect 35575 15144 35587 15147
rect 35802 15144 35808 15156
rect 35575 15116 35808 15144
rect 35575 15113 35587 15116
rect 35529 15107 35587 15113
rect 35802 15104 35808 15116
rect 35860 15104 35866 15156
rect 36265 15147 36323 15153
rect 36265 15113 36277 15147
rect 36311 15144 36323 15147
rect 36446 15144 36452 15156
rect 36311 15116 36452 15144
rect 36311 15113 36323 15116
rect 36265 15107 36323 15113
rect 36446 15104 36452 15116
rect 36504 15104 36510 15156
rect 37001 15147 37059 15153
rect 37001 15113 37013 15147
rect 37047 15144 37059 15147
rect 37642 15144 37648 15156
rect 37047 15116 37648 15144
rect 37047 15113 37059 15116
rect 37001 15107 37059 15113
rect 37642 15104 37648 15116
rect 37700 15104 37706 15156
rect 38654 15104 38660 15156
rect 38712 15144 38718 15156
rect 40954 15144 40960 15156
rect 38712 15116 39896 15144
rect 38712 15104 38718 15116
rect 31619 15048 31754 15076
rect 31619 15045 31631 15048
rect 31573 15039 31631 15045
rect 32214 15036 32220 15088
rect 32272 15036 32278 15088
rect 32309 15079 32367 15085
rect 32309 15045 32321 15079
rect 32355 15076 32367 15079
rect 32582 15076 32588 15088
rect 32355 15048 32588 15076
rect 32355 15045 32367 15048
rect 32309 15039 32367 15045
rect 32582 15036 32588 15048
rect 32640 15036 32646 15088
rect 33597 15079 33655 15085
rect 33597 15045 33609 15079
rect 33643 15076 33655 15079
rect 34054 15076 34060 15088
rect 33643 15048 34060 15076
rect 33643 15045 33655 15048
rect 33597 15039 33655 15045
rect 34054 15036 34060 15048
rect 34112 15036 34118 15088
rect 34241 15079 34299 15085
rect 34241 15045 34253 15079
rect 34287 15076 34299 15079
rect 35434 15076 35440 15088
rect 34287 15048 35440 15076
rect 34287 15045 34299 15048
rect 34241 15039 34299 15045
rect 35434 15036 35440 15048
rect 35492 15036 35498 15088
rect 37093 15079 37151 15085
rect 37093 15076 37105 15079
rect 35636 15048 37105 15076
rect 31159 15008 31217 15011
rect 32030 15008 32036 15020
rect 30469 14971 30527 14977
rect 30576 14980 32036 15008
rect 30190 14900 30196 14952
rect 30248 14940 30254 14952
rect 30576 14940 30604 14980
rect 32030 14968 32036 14980
rect 32088 14968 32094 15020
rect 32858 15008 32864 15020
rect 32140 14980 32864 15008
rect 30248 14912 30604 14940
rect 30248 14900 30254 14912
rect 30650 14900 30656 14952
rect 30708 14940 30714 14952
rect 32140 14940 32168 14980
rect 32858 14968 32864 14980
rect 32916 14968 32922 15020
rect 32950 14968 32956 15020
rect 33008 14968 33014 15020
rect 33134 14968 33140 15020
rect 33192 14968 33198 15020
rect 33226 14968 33232 15020
rect 33284 15008 33290 15020
rect 35636 15017 35664 15048
rect 37093 15045 37105 15048
rect 37139 15045 37151 15079
rect 37093 15039 37151 15045
rect 33873 15011 33931 15017
rect 33873 15008 33885 15011
rect 33284 14980 33885 15008
rect 33284 14968 33290 14980
rect 33873 14977 33885 14980
rect 33919 14977 33931 15011
rect 35621 15011 35679 15017
rect 35621 15008 35633 15011
rect 33873 14971 33931 14977
rect 34348 14980 35633 15008
rect 30708 14912 32168 14940
rect 30708 14900 30714 14912
rect 32490 14900 32496 14952
rect 32548 14940 32554 14952
rect 32674 14940 32680 14952
rect 32548 14912 32680 14940
rect 32548 14900 32554 14912
rect 32674 14900 32680 14912
rect 32732 14900 32738 14952
rect 33045 14943 33103 14949
rect 33045 14909 33057 14943
rect 33091 14940 33103 14943
rect 33318 14940 33324 14952
rect 33091 14912 33324 14940
rect 33091 14909 33103 14912
rect 33045 14903 33103 14909
rect 33318 14900 33324 14912
rect 33376 14940 33382 14952
rect 34146 14940 34152 14952
rect 33376 14912 34152 14940
rect 33376 14900 33382 14912
rect 34146 14900 34152 14912
rect 34204 14900 34210 14952
rect 31754 14832 31760 14884
rect 31812 14832 31818 14884
rect 32582 14832 32588 14884
rect 32640 14872 32646 14884
rect 34348 14872 34376 14980
rect 35621 14977 35633 14980
rect 35667 14977 35679 15011
rect 35621 14971 35679 14977
rect 36449 15011 36507 15017
rect 36449 14977 36461 15011
rect 36495 15008 36507 15011
rect 37108 15008 37136 15039
rect 37550 15036 37556 15088
rect 37608 15076 37614 15088
rect 38194 15076 38200 15088
rect 37608 15048 38200 15076
rect 37608 15036 37614 15048
rect 38194 15036 38200 15048
rect 38252 15076 38258 15088
rect 38381 15079 38439 15085
rect 38381 15076 38393 15079
rect 38252 15048 38393 15076
rect 38252 15036 38258 15048
rect 38381 15045 38393 15048
rect 38427 15045 38439 15079
rect 39390 15076 39396 15088
rect 38381 15039 38439 15045
rect 39224 15048 39396 15076
rect 39224 15020 39252 15048
rect 39390 15036 39396 15048
rect 39448 15036 39454 15088
rect 37734 15008 37740 15020
rect 36495 14980 36676 15008
rect 37108 14980 37740 15008
rect 36495 14977 36507 14980
rect 36449 14971 36507 14977
rect 34793 14943 34851 14949
rect 34793 14909 34805 14943
rect 34839 14909 34851 14943
rect 34793 14903 34851 14909
rect 34977 14943 35035 14949
rect 34977 14909 34989 14943
rect 35023 14940 35035 14943
rect 35066 14940 35072 14952
rect 35023 14912 35072 14940
rect 35023 14909 35035 14912
rect 34977 14903 35035 14909
rect 32640 14844 34376 14872
rect 32640 14832 32646 14844
rect 29733 14807 29791 14813
rect 29733 14804 29745 14807
rect 28224 14776 29745 14804
rect 28224 14764 28230 14776
rect 29733 14773 29745 14776
rect 29779 14773 29791 14807
rect 29733 14767 29791 14773
rect 30558 14764 30564 14816
rect 30616 14804 30622 14816
rect 31113 14807 31171 14813
rect 31113 14804 31125 14807
rect 30616 14776 31125 14804
rect 30616 14764 30622 14776
rect 31113 14773 31125 14776
rect 31159 14804 31171 14807
rect 31202 14804 31208 14816
rect 31159 14776 31208 14804
rect 31159 14773 31171 14776
rect 31113 14767 31171 14773
rect 31202 14764 31208 14776
rect 31260 14764 31266 14816
rect 31297 14807 31355 14813
rect 31297 14773 31309 14807
rect 31343 14804 31355 14807
rect 32766 14804 32772 14816
rect 31343 14776 32772 14804
rect 31343 14773 31355 14776
rect 31297 14767 31355 14773
rect 32766 14764 32772 14776
rect 32824 14764 32830 14816
rect 33042 14764 33048 14816
rect 33100 14804 33106 14816
rect 34808 14804 34836 14903
rect 35066 14900 35072 14912
rect 35124 14940 35130 14952
rect 35713 14943 35771 14949
rect 35713 14940 35725 14943
rect 35124 14912 35725 14940
rect 35124 14900 35130 14912
rect 35713 14909 35725 14912
rect 35759 14909 35771 14943
rect 35713 14903 35771 14909
rect 36648 14881 36676 14980
rect 37734 14968 37740 14980
rect 37792 14968 37798 15020
rect 39206 14968 39212 15020
rect 39264 14968 39270 15020
rect 39301 15011 39359 15017
rect 39301 14977 39313 15011
rect 39347 15008 39359 15011
rect 39666 15008 39672 15020
rect 39347 14980 39672 15008
rect 39347 14977 39359 14980
rect 39301 14971 39359 14977
rect 39666 14968 39672 14980
rect 39724 14968 39730 15020
rect 39868 15017 39896 15116
rect 40144 15116 40960 15144
rect 40144 15085 40172 15116
rect 40954 15104 40960 15116
rect 41012 15104 41018 15156
rect 42978 15144 42984 15156
rect 42076 15116 42984 15144
rect 40129 15079 40187 15085
rect 40129 15045 40141 15079
rect 40175 15045 40187 15079
rect 40129 15039 40187 15045
rect 40218 15036 40224 15088
rect 40276 15076 40282 15088
rect 40276 15048 40618 15076
rect 40276 15036 40282 15048
rect 41598 15036 41604 15088
rect 41656 15036 41662 15088
rect 42076 15085 42104 15116
rect 42978 15104 42984 15116
rect 43036 15104 43042 15156
rect 42061 15079 42119 15085
rect 42061 15045 42073 15079
rect 42107 15045 42119 15079
rect 42061 15039 42119 15045
rect 39853 15011 39911 15017
rect 39853 14977 39865 15011
rect 39899 14977 39911 15011
rect 39853 14971 39911 14977
rect 37182 14900 37188 14952
rect 37240 14900 37246 14952
rect 39022 14900 39028 14952
rect 39080 14940 39086 14952
rect 39485 14943 39543 14949
rect 39485 14940 39497 14943
rect 39080 14912 39497 14940
rect 39080 14900 39086 14912
rect 39485 14909 39497 14912
rect 39531 14909 39543 14943
rect 41616 14940 41644 15036
rect 43194 14980 43944 15008
rect 39485 14903 39543 14909
rect 39592 14912 41644 14940
rect 36633 14875 36691 14881
rect 36633 14841 36645 14875
rect 36679 14841 36691 14875
rect 36633 14835 36691 14841
rect 36814 14832 36820 14884
rect 36872 14872 36878 14884
rect 39592 14872 39620 14912
rect 41782 14900 41788 14952
rect 41840 14900 41846 14952
rect 36872 14844 39620 14872
rect 36872 14832 36878 14844
rect 41230 14832 41236 14884
rect 41288 14872 41294 14884
rect 41800 14872 41828 14900
rect 41288 14844 41828 14872
rect 41288 14832 41294 14844
rect 43916 14816 43944 14980
rect 45186 14968 45192 15020
rect 45244 14968 45250 15020
rect 36906 14804 36912 14816
rect 33100 14776 36912 14804
rect 33100 14764 33106 14776
rect 36906 14764 36912 14776
rect 36964 14764 36970 14816
rect 37274 14764 37280 14816
rect 37332 14804 37338 14816
rect 37645 14807 37703 14813
rect 37645 14804 37657 14807
rect 37332 14776 37657 14804
rect 37332 14764 37338 14776
rect 37645 14773 37657 14776
rect 37691 14804 37703 14807
rect 38013 14807 38071 14813
rect 38013 14804 38025 14807
rect 37691 14776 38025 14804
rect 37691 14773 37703 14776
rect 37645 14767 37703 14773
rect 38013 14773 38025 14776
rect 38059 14804 38071 14807
rect 38654 14804 38660 14816
rect 38059 14776 38660 14804
rect 38059 14773 38071 14776
rect 38013 14767 38071 14773
rect 38654 14764 38660 14776
rect 38712 14804 38718 14816
rect 38749 14807 38807 14813
rect 38749 14804 38761 14807
rect 38712 14776 38761 14804
rect 38712 14764 38718 14776
rect 38749 14773 38761 14776
rect 38795 14773 38807 14807
rect 38749 14767 38807 14773
rect 38930 14764 38936 14816
rect 38988 14764 38994 14816
rect 39206 14764 39212 14816
rect 39264 14804 39270 14816
rect 40770 14804 40776 14816
rect 39264 14776 40776 14804
rect 39264 14764 39270 14776
rect 40770 14764 40776 14776
rect 40828 14764 40834 14816
rect 41138 14764 41144 14816
rect 41196 14804 41202 14816
rect 41414 14804 41420 14816
rect 41196 14776 41420 14804
rect 41196 14764 41202 14776
rect 41414 14764 41420 14776
rect 41472 14764 41478 14816
rect 41506 14764 41512 14816
rect 41564 14804 41570 14816
rect 41601 14807 41659 14813
rect 41601 14804 41613 14807
rect 41564 14776 41613 14804
rect 41564 14764 41570 14776
rect 41601 14773 41613 14776
rect 41647 14773 41659 14807
rect 41601 14767 41659 14773
rect 42610 14764 42616 14816
rect 42668 14804 42674 14816
rect 43533 14807 43591 14813
rect 43533 14804 43545 14807
rect 42668 14776 43545 14804
rect 42668 14764 42674 14776
rect 43533 14773 43545 14776
rect 43579 14773 43591 14807
rect 43533 14767 43591 14773
rect 43898 14764 43904 14816
rect 43956 14804 43962 14816
rect 44177 14807 44235 14813
rect 44177 14804 44189 14807
rect 43956 14776 44189 14804
rect 43956 14764 43962 14776
rect 44177 14773 44189 14776
rect 44223 14773 44235 14807
rect 44177 14767 44235 14773
rect 44358 14764 44364 14816
rect 44416 14804 44422 14816
rect 44545 14807 44603 14813
rect 44545 14804 44557 14807
rect 44416 14776 44557 14804
rect 44416 14764 44422 14776
rect 44545 14773 44557 14776
rect 44591 14773 44603 14807
rect 44545 14767 44603 14773
rect 45002 14764 45008 14816
rect 45060 14764 45066 14816
rect 460 14714 45540 14736
rect 460 14662 3570 14714
rect 3622 14662 3634 14714
rect 3686 14662 3698 14714
rect 3750 14662 3762 14714
rect 3814 14662 3826 14714
rect 3878 14662 8570 14714
rect 8622 14662 8634 14714
rect 8686 14662 8698 14714
rect 8750 14662 8762 14714
rect 8814 14662 8826 14714
rect 8878 14662 13570 14714
rect 13622 14662 13634 14714
rect 13686 14662 13698 14714
rect 13750 14662 13762 14714
rect 13814 14662 13826 14714
rect 13878 14662 18570 14714
rect 18622 14662 18634 14714
rect 18686 14662 18698 14714
rect 18750 14662 18762 14714
rect 18814 14662 18826 14714
rect 18878 14662 23570 14714
rect 23622 14662 23634 14714
rect 23686 14662 23698 14714
rect 23750 14662 23762 14714
rect 23814 14662 23826 14714
rect 23878 14662 28570 14714
rect 28622 14662 28634 14714
rect 28686 14662 28698 14714
rect 28750 14662 28762 14714
rect 28814 14662 28826 14714
rect 28878 14662 33570 14714
rect 33622 14662 33634 14714
rect 33686 14662 33698 14714
rect 33750 14662 33762 14714
rect 33814 14662 33826 14714
rect 33878 14662 38570 14714
rect 38622 14662 38634 14714
rect 38686 14662 38698 14714
rect 38750 14662 38762 14714
rect 38814 14662 38826 14714
rect 38878 14662 43570 14714
rect 43622 14662 43634 14714
rect 43686 14662 43698 14714
rect 43750 14662 43762 14714
rect 43814 14662 43826 14714
rect 43878 14662 45540 14714
rect 460 14640 45540 14662
rect 4249 14603 4307 14609
rect 4249 14569 4261 14603
rect 4295 14600 4307 14603
rect 4338 14600 4344 14612
rect 4295 14572 4344 14600
rect 4295 14569 4307 14572
rect 4249 14563 4307 14569
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5626 14600 5632 14612
rect 4856 14572 5632 14600
rect 4856 14560 4862 14572
rect 5626 14560 5632 14572
rect 5684 14600 5690 14612
rect 6733 14603 6791 14609
rect 6733 14600 6745 14603
rect 5684 14572 6745 14600
rect 5684 14560 5690 14572
rect 6733 14569 6745 14572
rect 6779 14569 6791 14603
rect 6733 14563 6791 14569
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 12161 14603 12219 14609
rect 9732 14572 11928 14600
rect 9732 14560 9738 14572
rect 4816 14532 4844 14560
rect 4540 14504 4844 14532
rect 4540 14405 4568 14504
rect 6638 14492 6644 14544
rect 6696 14532 6702 14544
rect 7101 14535 7159 14541
rect 7101 14532 7113 14535
rect 6696 14504 7113 14532
rect 6696 14492 6702 14504
rect 7101 14501 7113 14504
rect 7147 14501 7159 14535
rect 7101 14495 7159 14501
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14532 7619 14535
rect 7742 14532 7748 14544
rect 7607 14504 7748 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 7742 14492 7748 14504
rect 7800 14532 7806 14544
rect 7800 14504 8340 14532
rect 7800 14492 7806 14504
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4890 14464 4896 14476
rect 4672 14436 4896 14464
rect 4672 14424 4678 14436
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 5718 14464 5724 14476
rect 5000 14436 5724 14464
rect 5000 14405 5028 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 6656 14396 6684 14492
rect 8202 14464 8208 14476
rect 7852 14436 8208 14464
rect 7852 14405 7880 14436
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8312 14408 8340 14504
rect 10060 14504 11836 14532
rect 10060 14476 10088 14504
rect 9766 14464 9772 14476
rect 9692 14436 9772 14464
rect 6394 14368 6684 14396
rect 7837 14399 7895 14405
rect 4985 14359 5043 14365
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 5000 14328 5028 14359
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 8294 14356 8300 14408
rect 8352 14356 8358 14408
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9692 14396 9720 14436
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10042 14424 10048 14476
rect 10100 14424 10106 14476
rect 11808 14473 11836 14504
rect 11333 14467 11391 14473
rect 11333 14464 11345 14467
rect 10244 14436 11345 14464
rect 9640 14382 9720 14396
rect 9640 14368 9706 14382
rect 9640 14356 9646 14368
rect 3804 14300 5028 14328
rect 5261 14331 5319 14337
rect 3804 14272 3832 14300
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 8573 14331 8631 14337
rect 8573 14328 8585 14331
rect 5261 14291 5319 14297
rect 7668 14300 8585 14328
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5276 14260 5304 14291
rect 7668 14269 7696 14300
rect 8573 14297 8585 14300
rect 8619 14297 8631 14331
rect 8573 14291 8631 14297
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10244 14337 10272 14436
rect 11333 14433 11345 14436
rect 11379 14464 11391 14467
rect 11793 14467 11851 14473
rect 11379 14436 11652 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 10318 14356 10324 14408
rect 10376 14396 10382 14408
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 10376 14368 11529 14396
rect 10376 14356 10382 14368
rect 11517 14365 11529 14368
rect 11563 14365 11575 14399
rect 11624 14396 11652 14436
rect 11793 14433 11805 14467
rect 11839 14433 11851 14467
rect 11900 14464 11928 14572
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 13078 14600 13084 14612
rect 12207 14572 13084 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13596 14572 15148 14600
rect 13596 14560 13602 14572
rect 15120 14544 15148 14572
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 15804 14572 16865 14600
rect 15804 14560 15810 14572
rect 16853 14569 16865 14572
rect 16899 14600 16911 14603
rect 16942 14600 16948 14612
rect 16899 14572 16948 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 18414 14600 18420 14612
rect 17828 14572 18420 14600
rect 17828 14560 17834 14572
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 18690 14560 18696 14612
rect 18748 14600 18754 14612
rect 19242 14600 19248 14612
rect 18748 14572 19248 14600
rect 18748 14560 18754 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19521 14603 19579 14609
rect 19521 14569 19533 14603
rect 19567 14600 19579 14603
rect 19797 14603 19855 14609
rect 19567 14572 19748 14600
rect 19567 14569 19579 14572
rect 19521 14563 19579 14569
rect 13449 14535 13507 14541
rect 13449 14501 13461 14535
rect 13495 14532 13507 14535
rect 13495 14504 14964 14532
rect 13495 14501 13507 14504
rect 13449 14495 13507 14501
rect 12002 14467 12060 14473
rect 12002 14464 12014 14467
rect 11900 14436 12014 14464
rect 11793 14427 11851 14433
rect 12002 14433 12014 14436
rect 12048 14433 12060 14467
rect 12002 14427 12060 14433
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 12400 14436 13185 14464
rect 12400 14424 12406 14436
rect 13173 14433 13185 14436
rect 13219 14464 13231 14467
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13219 14436 14105 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 14093 14433 14105 14436
rect 14139 14464 14151 14467
rect 14826 14464 14832 14476
rect 14139 14436 14832 14464
rect 14139 14433 14151 14436
rect 14093 14427 14151 14433
rect 14826 14424 14832 14436
rect 14884 14424 14890 14476
rect 12360 14396 12388 14424
rect 11624 14368 12388 14396
rect 12437 14399 12495 14405
rect 11517 14359 11575 14365
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 14461 14399 14519 14405
rect 12483 14368 14412 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 9916 14300 10241 14328
rect 9916 14288 9922 14300
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 10229 14291 10287 14297
rect 11057 14331 11115 14337
rect 11057 14297 11069 14331
rect 11103 14328 11115 14331
rect 11103 14300 11560 14328
rect 11103 14297 11115 14300
rect 11057 14291 11115 14297
rect 11532 14272 11560 14300
rect 11882 14288 11888 14340
rect 11940 14288 11946 14340
rect 13817 14331 13875 14337
rect 13817 14297 13829 14331
rect 13863 14328 13875 14331
rect 13998 14328 14004 14340
rect 13863 14300 14004 14328
rect 13863 14297 13875 14300
rect 13817 14291 13875 14297
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 14384 14328 14412 14368
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14936 14396 14964 14504
rect 15102 14492 15108 14544
rect 15160 14492 15166 14544
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 18325 14535 18383 14541
rect 16448 14504 16896 14532
rect 16448 14492 16454 14504
rect 16868 14476 16896 14504
rect 18325 14501 18337 14535
rect 18371 14532 18383 14535
rect 19610 14532 19616 14544
rect 18371 14504 19616 14532
rect 18371 14501 18383 14504
rect 18325 14495 18383 14501
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 19720 14532 19748 14572
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 20070 14600 20076 14612
rect 19843 14572 20076 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 21266 14600 21272 14612
rect 20496 14572 21272 14600
rect 20496 14560 20502 14572
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 21542 14560 21548 14612
rect 21600 14600 21606 14612
rect 21683 14603 21741 14609
rect 21683 14600 21695 14603
rect 21600 14572 21695 14600
rect 21600 14560 21606 14572
rect 21683 14569 21695 14572
rect 21729 14569 21741 14603
rect 21683 14563 21741 14569
rect 23198 14560 23204 14612
rect 23256 14600 23262 14612
rect 23256 14572 24164 14600
rect 23256 14560 23262 14572
rect 19886 14532 19892 14544
rect 19720 14504 19892 14532
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 21450 14492 21456 14544
rect 21508 14532 21514 14544
rect 22738 14532 22744 14544
rect 21508 14504 22744 14532
rect 21508 14492 21514 14504
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 23308 14541 23336 14572
rect 23293 14535 23351 14541
rect 23293 14501 23305 14535
rect 23339 14501 23351 14535
rect 23293 14495 23351 14501
rect 23750 14492 23756 14544
rect 23808 14492 23814 14544
rect 23934 14492 23940 14544
rect 23992 14492 23998 14544
rect 24136 14532 24164 14572
rect 24578 14560 24584 14612
rect 24636 14560 24642 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 24912 14572 25360 14600
rect 24912 14560 24918 14572
rect 25222 14532 25228 14544
rect 24136 14504 25084 14532
rect 15378 14424 15384 14476
rect 15436 14424 15442 14476
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 19521 14467 19579 14473
rect 18800 14436 19104 14464
rect 18800 14408 18828 14436
rect 19076 14408 19104 14436
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 22186 14464 22192 14476
rect 19567 14436 22192 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 22186 14424 22192 14436
rect 22244 14424 22250 14476
rect 23952 14464 23980 14492
rect 25056 14473 25084 14504
rect 25148 14504 25228 14532
rect 25148 14473 25176 14504
rect 25222 14492 25228 14504
rect 25280 14492 25286 14544
rect 25332 14532 25360 14572
rect 27062 14560 27068 14612
rect 27120 14600 27126 14612
rect 27249 14603 27307 14609
rect 27249 14600 27261 14603
rect 27120 14572 27261 14600
rect 27120 14560 27126 14572
rect 27249 14569 27261 14572
rect 27295 14569 27307 14603
rect 27249 14563 27307 14569
rect 28258 14560 28264 14612
rect 28316 14560 28322 14612
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 29086 14600 29092 14612
rect 28408 14572 29092 14600
rect 28408 14560 28414 14572
rect 25332 14504 25544 14532
rect 25041 14467 25099 14473
rect 22664 14436 23428 14464
rect 23952 14436 24072 14464
rect 22664 14408 22692 14436
rect 14507 14368 14964 14396
rect 15105 14399 15163 14405
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 14734 14328 14740 14340
rect 14384 14300 14740 14328
rect 14734 14288 14740 14300
rect 14792 14288 14798 14340
rect 15120 14328 15148 14359
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17736 14368 18153 14396
rect 17736 14356 17742 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 18230 14356 18236 14408
rect 18288 14396 18294 14408
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 18288 14368 18429 14396
rect 18288 14356 18294 14368
rect 18417 14365 18429 14368
rect 18463 14396 18475 14399
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18463 14368 18613 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 18601 14365 18613 14368
rect 18647 14396 18659 14399
rect 18690 14396 18696 14408
rect 18647 14368 18696 14396
rect 18647 14365 18659 14368
rect 18601 14359 18659 14365
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 18782 14356 18788 14408
rect 18840 14356 18846 14408
rect 18966 14356 18972 14408
rect 19024 14356 19030 14408
rect 19058 14356 19064 14408
rect 19116 14356 19122 14408
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19300 14368 19625 14396
rect 19300 14356 19306 14368
rect 19613 14365 19625 14368
rect 19659 14396 19671 14399
rect 19702 14396 19708 14408
rect 19659 14368 19708 14396
rect 19659 14365 19671 14368
rect 19613 14359 19671 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 14936 14300 15148 14328
rect 4939 14232 5304 14260
rect 7653 14263 7711 14269
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 7653 14229 7665 14263
rect 7699 14229 7711 14263
rect 7653 14223 7711 14229
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8386 14260 8392 14272
rect 7975 14232 8392 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 10042 14220 10048 14272
rect 10100 14220 10106 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10321 14263 10379 14269
rect 10321 14260 10333 14263
rect 10192 14232 10333 14260
rect 10192 14220 10198 14232
rect 10321 14229 10333 14232
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 10686 14220 10692 14272
rect 10744 14220 10750 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11422 14260 11428 14272
rect 11195 14232 11428 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 12250 14220 12256 14272
rect 12308 14220 12314 14272
rect 12526 14220 12532 14272
rect 12584 14220 12590 14272
rect 12894 14220 12900 14272
rect 12952 14220 12958 14272
rect 12989 14263 13047 14269
rect 12989 14229 13001 14263
rect 13035 14260 13047 14263
rect 13538 14260 13544 14272
rect 13035 14232 13544 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 13906 14220 13912 14272
rect 13964 14220 13970 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14277 14263 14335 14269
rect 14277 14260 14289 14263
rect 14240 14232 14289 14260
rect 14240 14220 14246 14232
rect 14277 14229 14289 14232
rect 14323 14229 14335 14263
rect 14277 14223 14335 14229
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 14936 14269 14964 14300
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15712 14300 15870 14328
rect 15712 14288 15718 14300
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14608 14232 14933 14260
rect 14608 14220 14614 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 15764 14260 15792 14300
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 17862 14328 17868 14340
rect 16908 14300 17868 14328
rect 16908 14288 16914 14300
rect 17862 14288 17868 14300
rect 17920 14328 17926 14340
rect 18877 14331 18935 14337
rect 18877 14328 18889 14331
rect 17920 14300 18889 14328
rect 17920 14288 17926 14300
rect 18877 14297 18889 14300
rect 18923 14328 18935 14331
rect 18923 14300 19288 14328
rect 18923 14297 18935 14300
rect 18877 14291 18935 14297
rect 17405 14263 17463 14269
rect 17405 14260 17417 14263
rect 15764 14232 17417 14260
rect 14921 14223 14979 14229
rect 17405 14229 17417 14232
rect 17451 14260 17463 14263
rect 17770 14260 17776 14272
rect 17451 14232 17776 14260
rect 17451 14229 17463 14232
rect 17405 14223 17463 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 17957 14263 18015 14269
rect 17957 14229 17969 14263
rect 18003 14260 18015 14263
rect 18322 14260 18328 14272
rect 18003 14232 18328 14260
rect 18003 14229 18015 14232
rect 17957 14223 18015 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18748 14232 19165 14260
rect 18748 14220 18754 14232
rect 19153 14229 19165 14232
rect 19199 14229 19211 14263
rect 19260 14260 19288 14300
rect 19334 14288 19340 14340
rect 19392 14288 19398 14340
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19904 14328 19932 14359
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 20220 14368 20269 14396
rect 20220 14356 20226 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 21174 14356 21180 14408
rect 21232 14396 21238 14408
rect 21232 14368 21404 14396
rect 21232 14356 21238 14368
rect 19484 14300 20024 14328
rect 19484 14288 19490 14300
rect 19886 14260 19892 14272
rect 19260 14232 19892 14260
rect 19153 14223 19211 14229
rect 19886 14220 19892 14232
rect 19944 14220 19950 14272
rect 19996 14260 20024 14300
rect 21266 14288 21272 14340
rect 21324 14288 21330 14340
rect 21376 14328 21404 14368
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21821 14399 21879 14405
rect 21821 14396 21833 14399
rect 21508 14368 21833 14396
rect 21508 14356 21514 14368
rect 21821 14365 21833 14368
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 21910 14356 21916 14408
rect 21968 14396 21974 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 21968 14368 22569 14396
rect 21968 14356 21974 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14396 22799 14399
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22787 14368 22845 14396
rect 22787 14365 22799 14368
rect 22741 14359 22799 14365
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 22922 14356 22928 14408
rect 22980 14396 22986 14408
rect 23400 14405 23428 14436
rect 23017 14399 23075 14405
rect 23017 14396 23029 14399
rect 22980 14368 23029 14396
rect 22980 14356 22986 14368
rect 23017 14365 23029 14368
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 23385 14399 23443 14405
rect 23385 14365 23397 14399
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 23934 14356 23940 14408
rect 23992 14356 23998 14408
rect 24044 14405 24072 14436
rect 25041 14433 25053 14467
rect 25087 14433 25099 14467
rect 25041 14427 25099 14433
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14433 25191 14467
rect 25516 14464 25544 14504
rect 26712 14504 27844 14532
rect 26712 14476 26740 14504
rect 27816 14476 27844 14504
rect 25685 14467 25743 14473
rect 25685 14464 25697 14467
rect 25516 14436 25697 14464
rect 25133 14427 25191 14433
rect 25685 14433 25697 14436
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 26694 14424 26700 14476
rect 26752 14424 26758 14476
rect 27154 14424 27160 14476
rect 27212 14424 27218 14476
rect 27798 14424 27804 14476
rect 27856 14424 27862 14476
rect 28276 14464 28304 14560
rect 28920 14473 28948 14572
rect 29086 14560 29092 14572
rect 29144 14560 29150 14612
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 29328 14572 30604 14600
rect 29328 14560 29334 14572
rect 28905 14467 28963 14473
rect 28276 14436 28396 14464
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14365 24087 14399
rect 24029 14359 24087 14365
rect 24210 14356 24216 14408
rect 24268 14356 24274 14408
rect 24305 14399 24363 14405
rect 24305 14365 24317 14399
rect 24351 14365 24363 14399
rect 24305 14359 24363 14365
rect 22373 14331 22431 14337
rect 22373 14328 22385 14331
rect 21376 14300 22385 14328
rect 21928 14272 21956 14300
rect 22373 14297 22385 14300
rect 22419 14297 22431 14331
rect 22373 14291 22431 14297
rect 20346 14260 20352 14272
rect 19996 14232 20352 14260
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 21910 14220 21916 14272
rect 21968 14220 21974 14272
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22278 14260 22284 14272
rect 22060 14232 22284 14260
rect 22060 14220 22066 14232
rect 22278 14220 22284 14232
rect 22336 14260 22342 14272
rect 23290 14260 23296 14272
rect 22336 14232 23296 14260
rect 22336 14220 22342 14232
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 24026 14220 24032 14272
rect 24084 14260 24090 14272
rect 24320 14260 24348 14359
rect 25406 14356 25412 14408
rect 25464 14356 25470 14408
rect 26786 14356 26792 14408
rect 26844 14356 26850 14408
rect 26970 14356 26976 14408
rect 27028 14356 27034 14408
rect 27172 14396 27200 14424
rect 27617 14399 27675 14405
rect 27617 14396 27629 14399
rect 27172 14368 27629 14396
rect 27617 14365 27629 14368
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 28258 14356 28264 14408
rect 28316 14356 28322 14408
rect 28368 14405 28396 14436
rect 28905 14433 28917 14467
rect 28951 14433 28963 14467
rect 28905 14427 28963 14433
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28994 14356 29000 14408
rect 29052 14396 29058 14408
rect 29161 14399 29219 14405
rect 29161 14396 29173 14399
rect 29052 14368 29173 14396
rect 29052 14356 29058 14368
rect 29161 14365 29173 14368
rect 29207 14365 29219 14399
rect 30576 14396 30604 14572
rect 30742 14560 30748 14612
rect 30800 14600 30806 14612
rect 30800 14572 31248 14600
rect 30800 14560 30806 14572
rect 30760 14532 30788 14560
rect 31110 14532 31116 14544
rect 30760 14504 30880 14532
rect 30650 14424 30656 14476
rect 30708 14464 30714 14476
rect 30852 14473 30880 14504
rect 30944 14504 31116 14532
rect 30944 14473 30972 14504
rect 31110 14492 31116 14504
rect 31168 14492 31174 14544
rect 31220 14532 31248 14572
rect 31294 14560 31300 14612
rect 31352 14600 31358 14612
rect 31389 14603 31447 14609
rect 31389 14600 31401 14603
rect 31352 14572 31401 14600
rect 31352 14560 31358 14572
rect 31389 14569 31401 14572
rect 31435 14600 31447 14603
rect 31662 14600 31668 14612
rect 31435 14572 31668 14600
rect 31435 14569 31447 14572
rect 31389 14563 31447 14569
rect 31662 14560 31668 14572
rect 31720 14560 31726 14612
rect 32122 14560 32128 14612
rect 32180 14600 32186 14612
rect 32217 14603 32275 14609
rect 32217 14600 32229 14603
rect 32180 14572 32229 14600
rect 32180 14560 32186 14572
rect 32217 14569 32229 14572
rect 32263 14600 32275 14603
rect 32490 14600 32496 14612
rect 32263 14572 32496 14600
rect 32263 14569 32275 14572
rect 32217 14563 32275 14569
rect 32490 14560 32496 14572
rect 32548 14600 32554 14612
rect 32585 14603 32643 14609
rect 32585 14600 32597 14603
rect 32548 14572 32597 14600
rect 32548 14560 32554 14572
rect 32585 14569 32597 14572
rect 32631 14569 32643 14603
rect 32585 14563 32643 14569
rect 35618 14560 35624 14612
rect 35676 14600 35682 14612
rect 36630 14600 36636 14612
rect 35676 14572 36636 14600
rect 35676 14560 35682 14572
rect 36630 14560 36636 14572
rect 36688 14600 36694 14612
rect 37090 14600 37096 14612
rect 36688 14572 37096 14600
rect 36688 14560 36694 14572
rect 37090 14560 37096 14572
rect 37148 14560 37154 14612
rect 38289 14603 38347 14609
rect 38289 14569 38301 14603
rect 38335 14600 38347 14603
rect 40126 14600 40132 14612
rect 38335 14572 40132 14600
rect 38335 14569 38347 14572
rect 38289 14563 38347 14569
rect 40126 14560 40132 14572
rect 40184 14560 40190 14612
rect 41693 14603 41751 14609
rect 41693 14569 41705 14603
rect 41739 14600 41751 14603
rect 42794 14600 42800 14612
rect 41739 14572 42800 14600
rect 41739 14569 41751 14572
rect 41693 14563 41751 14569
rect 42794 14560 42800 14572
rect 42852 14560 42858 14612
rect 43901 14603 43959 14609
rect 43901 14569 43913 14603
rect 43947 14600 43959 14603
rect 44266 14600 44272 14612
rect 43947 14572 44272 14600
rect 43947 14569 43959 14572
rect 43901 14563 43959 14569
rect 31478 14532 31484 14544
rect 31220 14504 31484 14532
rect 31478 14492 31484 14504
rect 31536 14492 31542 14544
rect 31573 14535 31631 14541
rect 31573 14501 31585 14535
rect 31619 14501 31631 14535
rect 31573 14495 31631 14501
rect 30745 14467 30803 14473
rect 30745 14464 30757 14467
rect 30708 14436 30757 14464
rect 30708 14424 30714 14436
rect 30745 14433 30757 14436
rect 30791 14433 30803 14467
rect 30745 14427 30803 14433
rect 30837 14467 30895 14473
rect 30837 14433 30849 14467
rect 30883 14433 30895 14467
rect 30837 14427 30895 14433
rect 30929 14467 30987 14473
rect 30929 14433 30941 14467
rect 30975 14433 30987 14467
rect 30929 14427 30987 14433
rect 31021 14467 31079 14473
rect 31021 14433 31033 14467
rect 31067 14464 31079 14467
rect 31588 14464 31616 14495
rect 32950 14492 32956 14544
rect 33008 14492 33014 14544
rect 33318 14492 33324 14544
rect 33376 14492 33382 14544
rect 33502 14492 33508 14544
rect 33560 14492 33566 14544
rect 33597 14535 33655 14541
rect 33597 14501 33609 14535
rect 33643 14532 33655 14535
rect 34330 14532 34336 14544
rect 33643 14504 34336 14532
rect 33643 14501 33655 14504
rect 33597 14495 33655 14501
rect 34330 14492 34336 14504
rect 34388 14492 34394 14544
rect 35526 14532 35532 14544
rect 35176 14504 35532 14532
rect 33520 14464 33548 14492
rect 34609 14467 34667 14473
rect 34609 14464 34621 14467
rect 31067 14436 31616 14464
rect 31864 14436 33088 14464
rect 33520 14436 34621 14464
rect 31067 14433 31079 14436
rect 31021 14427 31079 14433
rect 30576 14392 31754 14396
rect 31864 14392 31892 14436
rect 30576 14368 31892 14392
rect 29161 14359 29219 14365
rect 31726 14364 31892 14368
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14396 31999 14399
rect 32950 14396 32956 14408
rect 31987 14368 32956 14396
rect 31987 14365 31999 14368
rect 31941 14359 31999 14365
rect 32950 14356 32956 14368
rect 33008 14356 33014 14408
rect 33060 14396 33088 14436
rect 34609 14433 34621 14436
rect 34655 14433 34667 14467
rect 35176 14464 35204 14504
rect 35526 14492 35532 14504
rect 35584 14532 35590 14544
rect 35989 14535 36047 14541
rect 35584 14504 35940 14532
rect 35584 14492 35590 14504
rect 34609 14427 34667 14433
rect 34808 14436 35204 14464
rect 35345 14467 35403 14473
rect 33505 14399 33563 14405
rect 33060 14368 33456 14396
rect 24949 14331 25007 14337
rect 24949 14297 24961 14331
rect 24995 14328 25007 14331
rect 24995 14300 26096 14328
rect 24995 14297 25007 14300
rect 24949 14291 25007 14297
rect 24084 14232 24348 14260
rect 24084 14220 24090 14232
rect 25222 14220 25228 14272
rect 25280 14260 25286 14272
rect 25682 14260 25688 14272
rect 25280 14232 25688 14260
rect 25280 14220 25286 14232
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 26068 14260 26096 14300
rect 26602 14260 26608 14272
rect 26068 14232 26608 14260
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 26988 14260 27016 14356
rect 27430 14288 27436 14340
rect 27488 14328 27494 14340
rect 30834 14328 30840 14340
rect 27488 14300 30840 14328
rect 27488 14288 27494 14300
rect 27724 14269 27752 14300
rect 30834 14288 30840 14300
rect 30892 14288 30898 14340
rect 31018 14288 31024 14340
rect 31076 14328 31082 14340
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 31076 14300 31217 14328
rect 31076 14288 31082 14300
rect 31205 14297 31217 14300
rect 31251 14328 31263 14331
rect 32122 14328 32128 14340
rect 31251 14300 32128 14328
rect 31251 14297 31263 14300
rect 31205 14291 31263 14297
rect 32122 14288 32128 14300
rect 32180 14288 32186 14340
rect 33428 14328 33456 14368
rect 33505 14365 33517 14399
rect 33551 14396 33563 14399
rect 33686 14396 33692 14408
rect 33551 14368 33692 14396
rect 33551 14365 33563 14368
rect 33505 14359 33563 14365
rect 33686 14356 33692 14368
rect 33744 14356 33750 14408
rect 33778 14356 33784 14408
rect 33836 14356 33842 14408
rect 34517 14399 34575 14405
rect 34517 14396 34529 14399
rect 33888 14368 34529 14396
rect 33888 14328 33916 14368
rect 34517 14365 34529 14368
rect 34563 14396 34575 14399
rect 34808 14396 34836 14436
rect 35345 14433 35357 14467
rect 35391 14433 35403 14467
rect 35345 14427 35403 14433
rect 34563 14368 34836 14396
rect 34563 14365 34575 14368
rect 34517 14359 34575 14365
rect 34882 14356 34888 14408
rect 34940 14356 34946 14408
rect 35158 14356 35164 14408
rect 35216 14396 35222 14408
rect 35360 14396 35388 14427
rect 35710 14424 35716 14476
rect 35768 14424 35774 14476
rect 35802 14424 35808 14476
rect 35860 14424 35866 14476
rect 35912 14464 35940 14504
rect 35989 14501 36001 14535
rect 36035 14532 36047 14535
rect 37001 14535 37059 14541
rect 37001 14532 37013 14535
rect 36035 14504 37013 14532
rect 36035 14501 36047 14504
rect 35989 14495 36047 14501
rect 37001 14501 37013 14504
rect 37047 14501 37059 14535
rect 37001 14495 37059 14501
rect 37200 14504 39344 14532
rect 36538 14464 36544 14476
rect 35912 14436 36544 14464
rect 36538 14424 36544 14436
rect 36596 14424 36602 14476
rect 35216 14368 35388 14396
rect 35621 14399 35679 14405
rect 35216 14356 35222 14368
rect 35621 14365 35633 14399
rect 35667 14396 35679 14399
rect 35820 14396 35848 14424
rect 35667 14368 35848 14396
rect 35667 14365 35679 14368
rect 35621 14359 35679 14365
rect 35986 14356 35992 14408
rect 36044 14396 36050 14408
rect 37200 14405 37228 14504
rect 38933 14467 38991 14473
rect 38933 14433 38945 14467
rect 38979 14464 38991 14467
rect 39022 14464 39028 14476
rect 38979 14436 39028 14464
rect 38979 14433 38991 14436
rect 38933 14427 38991 14433
rect 39022 14424 39028 14436
rect 39080 14424 39086 14476
rect 39316 14464 39344 14504
rect 41414 14492 41420 14544
rect 41472 14532 41478 14544
rect 43916 14532 43944 14563
rect 44266 14560 44272 14572
rect 44324 14560 44330 14612
rect 41472 14504 43944 14532
rect 41472 14492 41478 14504
rect 39850 14464 39856 14476
rect 39316 14436 39856 14464
rect 39850 14424 39856 14436
rect 39908 14424 39914 14476
rect 40034 14424 40040 14476
rect 40092 14464 40098 14476
rect 40954 14464 40960 14476
rect 40092 14436 40960 14464
rect 40092 14424 40098 14436
rect 40954 14424 40960 14436
rect 41012 14424 41018 14476
rect 41874 14424 41880 14476
rect 41932 14464 41938 14476
rect 42245 14467 42303 14473
rect 42245 14464 42257 14467
rect 41932 14436 42257 14464
rect 41932 14424 41938 14436
rect 42245 14433 42257 14436
rect 42291 14433 42303 14467
rect 42245 14427 42303 14433
rect 36265 14399 36323 14405
rect 36265 14396 36277 14399
rect 36044 14368 36277 14396
rect 36044 14356 36050 14368
rect 36265 14365 36277 14368
rect 36311 14365 36323 14399
rect 36265 14359 36323 14365
rect 37185 14399 37243 14405
rect 37185 14365 37197 14399
rect 37231 14365 37243 14399
rect 37185 14359 37243 14365
rect 38010 14356 38016 14408
rect 38068 14356 38074 14408
rect 38102 14356 38108 14408
rect 38160 14356 38166 14408
rect 38470 14356 38476 14408
rect 38528 14396 38534 14408
rect 38838 14396 38844 14408
rect 38528 14368 38844 14396
rect 38528 14356 38534 14368
rect 38838 14356 38844 14368
rect 38896 14396 38902 14408
rect 39209 14399 39267 14405
rect 39209 14396 39221 14399
rect 38896 14368 39221 14396
rect 38896 14356 38902 14368
rect 39209 14365 39221 14368
rect 39255 14365 39267 14399
rect 39209 14359 39267 14365
rect 42153 14399 42211 14405
rect 42153 14365 42165 14399
rect 42199 14396 42211 14399
rect 42610 14396 42616 14408
rect 42199 14368 42616 14396
rect 42199 14365 42211 14368
rect 42153 14359 42211 14365
rect 42610 14356 42616 14368
rect 42668 14356 42674 14408
rect 33428 14300 33916 14328
rect 34425 14331 34483 14337
rect 34425 14297 34437 14331
rect 34471 14328 34483 14331
rect 34974 14328 34980 14340
rect 34471 14300 34980 14328
rect 34471 14297 34483 14300
rect 34425 14291 34483 14297
rect 34974 14288 34980 14300
rect 35032 14288 35038 14340
rect 35802 14288 35808 14340
rect 35860 14337 35866 14340
rect 35860 14331 35888 14337
rect 35876 14297 35888 14331
rect 35860 14291 35888 14297
rect 37277 14331 37335 14337
rect 37277 14297 37289 14331
rect 37323 14328 37335 14331
rect 38120 14328 38148 14356
rect 37323 14300 38148 14328
rect 38657 14331 38715 14337
rect 37323 14297 37335 14300
rect 37277 14291 37335 14297
rect 38657 14297 38669 14331
rect 38703 14328 38715 14331
rect 38703 14300 39436 14328
rect 38703 14297 38715 14300
rect 38657 14291 38715 14297
rect 35860 14288 35866 14291
rect 27157 14263 27215 14269
rect 27157 14260 27169 14263
rect 26988 14232 27169 14260
rect 27157 14229 27169 14232
rect 27203 14229 27215 14263
rect 27157 14223 27215 14229
rect 27709 14263 27767 14269
rect 27709 14229 27721 14263
rect 27755 14229 27767 14263
rect 27709 14223 27767 14229
rect 28074 14220 28080 14272
rect 28132 14220 28138 14272
rect 28537 14263 28595 14269
rect 28537 14229 28549 14263
rect 28583 14260 28595 14263
rect 28902 14260 28908 14272
rect 28583 14232 28908 14260
rect 28583 14229 28595 14232
rect 28537 14223 28595 14229
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 30282 14260 30288 14272
rect 29052 14232 30288 14260
rect 29052 14220 29058 14232
rect 30282 14220 30288 14232
rect 30340 14220 30346 14272
rect 30558 14220 30564 14272
rect 30616 14220 30622 14272
rect 30926 14220 30932 14272
rect 30984 14260 30990 14272
rect 31405 14263 31463 14269
rect 31405 14260 31417 14263
rect 30984 14232 31417 14260
rect 30984 14220 30990 14232
rect 31405 14229 31417 14232
rect 31451 14260 31463 14263
rect 32398 14260 32404 14272
rect 31451 14232 32404 14260
rect 31451 14229 31463 14232
rect 31405 14223 31463 14229
rect 32398 14220 32404 14232
rect 32456 14220 32462 14272
rect 33962 14220 33968 14272
rect 34020 14260 34026 14272
rect 34057 14263 34115 14269
rect 34057 14260 34069 14263
rect 34020 14232 34069 14260
rect 34020 14220 34026 14232
rect 34057 14229 34069 14232
rect 34103 14229 34115 14263
rect 34057 14223 34115 14229
rect 35066 14220 35072 14272
rect 35124 14260 35130 14272
rect 35710 14260 35716 14272
rect 35124 14232 35716 14260
rect 35124 14220 35130 14232
rect 35710 14220 35716 14232
rect 35768 14220 35774 14272
rect 36081 14263 36139 14269
rect 36081 14229 36093 14263
rect 36127 14260 36139 14263
rect 36446 14260 36452 14272
rect 36127 14232 36452 14260
rect 36127 14229 36139 14232
rect 36081 14223 36139 14229
rect 36446 14220 36452 14232
rect 36504 14220 36510 14272
rect 37366 14220 37372 14272
rect 37424 14220 37430 14272
rect 37550 14220 37556 14272
rect 37608 14220 37614 14272
rect 37826 14220 37832 14272
rect 37884 14220 37890 14272
rect 38749 14263 38807 14269
rect 38749 14229 38761 14263
rect 38795 14260 38807 14263
rect 39114 14260 39120 14272
rect 38795 14232 39120 14260
rect 38795 14229 38807 14232
rect 38749 14223 38807 14229
rect 39114 14220 39120 14232
rect 39172 14220 39178 14272
rect 39408 14260 39436 14300
rect 39482 14288 39488 14340
rect 39540 14288 39546 14340
rect 40218 14288 40224 14340
rect 40276 14288 40282 14340
rect 44174 14328 44180 14340
rect 42812 14300 44180 14328
rect 42812 14272 42840 14300
rect 44174 14288 44180 14300
rect 44232 14288 44238 14340
rect 39758 14260 39764 14272
rect 39408 14232 39764 14260
rect 39758 14220 39764 14232
rect 39816 14220 39822 14272
rect 40862 14220 40868 14272
rect 40920 14260 40926 14272
rect 41230 14260 41236 14272
rect 40920 14232 41236 14260
rect 40920 14220 40926 14232
rect 41230 14220 41236 14232
rect 41288 14220 41294 14272
rect 41506 14220 41512 14272
rect 41564 14260 41570 14272
rect 42061 14263 42119 14269
rect 42061 14260 42073 14263
rect 41564 14232 42073 14260
rect 41564 14220 41570 14232
rect 42061 14229 42073 14232
rect 42107 14229 42119 14263
rect 42061 14223 42119 14229
rect 42794 14220 42800 14272
rect 42852 14220 42858 14272
rect 43070 14220 43076 14272
rect 43128 14220 43134 14272
rect 43438 14220 43444 14272
rect 43496 14220 43502 14272
rect 44358 14220 44364 14272
rect 44416 14260 44422 14272
rect 44545 14263 44603 14269
rect 44545 14260 44557 14263
rect 44416 14232 44557 14260
rect 44416 14220 44422 14232
rect 44545 14229 44557 14232
rect 44591 14229 44603 14263
rect 44545 14223 44603 14229
rect 44726 14220 44732 14272
rect 44784 14260 44790 14272
rect 44913 14263 44971 14269
rect 44913 14260 44925 14263
rect 44784 14232 44925 14260
rect 44784 14220 44790 14232
rect 44913 14229 44925 14232
rect 44959 14229 44971 14263
rect 44913 14223 44971 14229
rect 460 14170 45540 14192
rect 460 14118 6070 14170
rect 6122 14118 6134 14170
rect 6186 14118 6198 14170
rect 6250 14118 6262 14170
rect 6314 14118 6326 14170
rect 6378 14118 11070 14170
rect 11122 14118 11134 14170
rect 11186 14118 11198 14170
rect 11250 14118 11262 14170
rect 11314 14118 11326 14170
rect 11378 14118 16070 14170
rect 16122 14118 16134 14170
rect 16186 14118 16198 14170
rect 16250 14118 16262 14170
rect 16314 14118 16326 14170
rect 16378 14118 21070 14170
rect 21122 14118 21134 14170
rect 21186 14118 21198 14170
rect 21250 14118 21262 14170
rect 21314 14118 21326 14170
rect 21378 14118 26070 14170
rect 26122 14118 26134 14170
rect 26186 14118 26198 14170
rect 26250 14118 26262 14170
rect 26314 14118 26326 14170
rect 26378 14118 31070 14170
rect 31122 14118 31134 14170
rect 31186 14118 31198 14170
rect 31250 14118 31262 14170
rect 31314 14118 31326 14170
rect 31378 14118 36070 14170
rect 36122 14118 36134 14170
rect 36186 14118 36198 14170
rect 36250 14118 36262 14170
rect 36314 14118 36326 14170
rect 36378 14118 41070 14170
rect 41122 14118 41134 14170
rect 41186 14118 41198 14170
rect 41250 14118 41262 14170
rect 41314 14118 41326 14170
rect 41378 14118 45540 14170
rect 460 14096 45540 14118
rect 3513 14059 3571 14065
rect 1872 14028 3464 14056
rect 1872 13988 1900 14028
rect 1780 13960 1900 13988
rect 1780 13929 1808 13960
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 3174 13892 3280 13920
rect 1765 13883 1823 13889
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1872 13824 2053 13852
rect 750 13744 756 13796
rect 808 13784 814 13796
rect 1872 13784 1900 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 808 13756 1900 13784
rect 808 13744 814 13756
rect 3252 13716 3280 13892
rect 3436 13864 3464 14028
rect 3513 14025 3525 14059
rect 3559 14056 3571 14059
rect 3559 14028 4108 14056
rect 3559 14025 3571 14028
rect 3513 14019 3571 14025
rect 4080 13997 4108 14028
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 6917 14059 6975 14065
rect 6917 14056 6929 14059
rect 6696 14028 6929 14056
rect 6696 14016 6702 14028
rect 6917 14025 6929 14028
rect 6963 14056 6975 14059
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6963 14028 7205 14056
rect 6963 14025 6975 14028
rect 6917 14019 6975 14025
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14056 7435 14059
rect 8110 14056 8116 14068
rect 7423 14028 8116 14056
rect 7423 14025 7435 14028
rect 7377 14019 7435 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 10042 14056 10048 14068
rect 8312 14028 10048 14056
rect 4065 13991 4123 13997
rect 4065 13957 4077 13991
rect 4111 13957 4123 13991
rect 4065 13951 4123 13957
rect 4338 13948 4344 14000
rect 4396 13988 4402 14000
rect 7745 13991 7803 13997
rect 4396 13960 4554 13988
rect 4396 13948 4402 13960
rect 7745 13957 7757 13991
rect 7791 13988 7803 13991
rect 8312 13988 8340 14028
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 12805 14059 12863 14065
rect 11716 14028 12756 14056
rect 7791 13960 8340 13988
rect 7791 13957 7803 13960
rect 7745 13951 7803 13957
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 8444 13960 8493 13988
rect 8444 13948 8450 13960
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 7883 13892 8156 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3786 13852 3792 13864
rect 3476 13824 3792 13852
rect 3476 13812 3482 13824
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 8018 13812 8024 13864
rect 8076 13812 8082 13864
rect 8128 13852 8156 13892
rect 8202 13880 8208 13932
rect 8260 13880 8266 13932
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 10134 13920 10140 13932
rect 9640 13892 10140 13920
rect 9640 13880 9646 13892
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10226 13880 10232 13932
rect 10284 13880 10290 13932
rect 10704 13929 10732 14016
rect 11716 13988 11744 14028
rect 12728 13988 12756 14028
rect 12805 14025 12817 14059
rect 12851 14056 12863 14059
rect 13354 14056 13360 14068
rect 12851 14028 13360 14056
rect 12851 14025 12863 14028
rect 12805 14019 12863 14025
rect 13354 14016 13360 14028
rect 13412 14056 13418 14068
rect 13538 14056 13544 14068
rect 13412 14028 13544 14056
rect 13412 14016 13418 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 13998 14016 14004 14068
rect 14056 14056 14062 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14056 14028 15209 14056
rect 14056 14016 14062 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 18414 14056 18420 14068
rect 15197 14019 15255 14025
rect 17880 14028 18420 14056
rect 13630 13988 13636 14000
rect 10980 13960 11822 13988
rect 12728 13960 13636 13988
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 9766 13852 9772 13864
rect 8128 13824 9772 13852
rect 9766 13812 9772 13824
rect 9824 13852 9830 13864
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9824 13824 9965 13852
rect 9824 13812 9830 13824
rect 9953 13821 9965 13824
rect 9999 13821 10011 13855
rect 10152 13852 10180 13880
rect 10980 13852 11008 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 14734 13948 14740 14000
rect 14792 13948 14798 14000
rect 15102 13948 15108 14000
rect 15160 13948 15166 14000
rect 17880 13997 17908 14028
rect 18414 14016 18420 14028
rect 18472 14056 18478 14068
rect 18782 14056 18788 14068
rect 18472 14028 18788 14056
rect 18472 14016 18478 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 20036 14028 20085 14056
rect 20036 14016 20042 14028
rect 20073 14025 20085 14028
rect 20119 14056 20131 14059
rect 20365 14059 20423 14065
rect 20365 14056 20377 14059
rect 20119 14028 20377 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20365 14025 20377 14028
rect 20411 14025 20423 14059
rect 20365 14019 20423 14025
rect 20533 14059 20591 14065
rect 20533 14025 20545 14059
rect 20579 14056 20591 14059
rect 21637 14059 21695 14065
rect 20579 14028 21404 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 17865 13991 17923 13997
rect 17865 13957 17877 13991
rect 17911 13957 17923 13991
rect 17865 13951 17923 13957
rect 17957 13991 18015 13997
rect 17957 13957 17969 13991
rect 18003 13988 18015 13991
rect 18230 13988 18236 14000
rect 18003 13960 18236 13988
rect 18003 13957 18015 13960
rect 17957 13951 18015 13957
rect 18230 13948 18236 13960
rect 18288 13948 18294 14000
rect 18601 13991 18659 13997
rect 18601 13957 18613 13991
rect 18647 13988 18659 13991
rect 18690 13988 18696 14000
rect 18647 13960 18696 13988
rect 18647 13957 18659 13960
rect 18601 13951 18659 13957
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 19150 13948 19156 14000
rect 19208 13948 19214 14000
rect 20165 13991 20223 13997
rect 20165 13957 20177 13991
rect 20211 13988 20223 13991
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 20211 13960 20637 13988
rect 20211 13957 20223 13960
rect 20165 13951 20223 13957
rect 10152 13824 11008 13852
rect 11057 13855 11115 13861
rect 9953 13815 10011 13821
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11330 13852 11336 13864
rect 11103 13824 11336 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 11330 13812 11336 13824
rect 11388 13852 11394 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 11388 13824 12909 13852
rect 11388 13812 11394 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 13964 13824 14657 13852
rect 13964 13812 13970 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14752 13793 14780 13948
rect 15746 13880 15752 13932
rect 15804 13880 15810 13932
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17310 13920 17316 13932
rect 16807 13892 17316 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18138 13920 18144 13932
rect 18095 13892 18144 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 14884 13824 15301 13852
rect 14884 13812 14890 13824
rect 15289 13821 15301 13824
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 16574 13812 16580 13864
rect 16632 13812 16638 13864
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16724 13824 16865 13852
rect 16724 13812 16730 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 16942 13812 16948 13864
rect 17000 13812 17006 13864
rect 17034 13812 17040 13864
rect 17092 13812 17098 13864
rect 17696 13852 17724 13883
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 18248 13892 18337 13920
rect 17954 13852 17960 13864
rect 17696 13824 17960 13852
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 18248 13852 18276 13892
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 18325 13883 18383 13889
rect 20548 13864 20576 13960
rect 20625 13957 20637 13960
rect 20671 13957 20683 13991
rect 20825 13991 20883 13997
rect 20825 13988 20837 13991
rect 20625 13951 20683 13957
rect 20732 13960 20837 13988
rect 20732 13920 20760 13960
rect 20825 13957 20837 13960
rect 20871 13957 20883 13991
rect 20825 13951 20883 13957
rect 20990 13948 20996 14000
rect 21048 13948 21054 14000
rect 21376 13997 21404 14028
rect 21637 14025 21649 14059
rect 21683 14056 21695 14059
rect 24118 14056 24124 14068
rect 21683 14028 24124 14056
rect 21683 14025 21695 14028
rect 21637 14019 21695 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 24670 14016 24676 14068
rect 24728 14056 24734 14068
rect 26053 14059 26111 14065
rect 24728 14028 25360 14056
rect 24728 14016 24734 14028
rect 21361 13991 21419 13997
rect 21361 13957 21373 13991
rect 21407 13957 21419 13991
rect 21361 13951 21419 13957
rect 22557 13991 22615 13997
rect 22557 13957 22569 13991
rect 22603 13988 22615 13991
rect 22603 13960 23244 13988
rect 22603 13957 22615 13960
rect 22557 13951 22615 13957
rect 20640 13892 20760 13920
rect 21008 13920 21036 13948
rect 23216 13932 23244 13960
rect 23750 13948 23756 14000
rect 23808 13988 23814 14000
rect 25332 13997 25360 14028
rect 26053 14025 26065 14059
rect 26099 14056 26111 14059
rect 26694 14056 26700 14068
rect 26099 14028 26700 14056
rect 26099 14025 26111 14028
rect 26053 14019 26111 14025
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 26878 14016 26884 14068
rect 26936 14016 26942 14068
rect 27154 14016 27160 14068
rect 27212 14056 27218 14068
rect 27709 14059 27767 14065
rect 27709 14056 27721 14059
rect 27212 14028 27721 14056
rect 27212 14016 27218 14028
rect 27709 14025 27721 14028
rect 27755 14025 27767 14059
rect 27709 14019 27767 14025
rect 27801 14059 27859 14065
rect 27801 14025 27813 14059
rect 27847 14025 27859 14059
rect 27801 14019 27859 14025
rect 25225 13991 25283 13997
rect 25225 13988 25237 13991
rect 23808 13960 25237 13988
rect 23808 13948 23814 13960
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21008 13892 22017 13920
rect 18064 13824 18276 13852
rect 14737 13787 14795 13793
rect 14737 13753 14749 13787
rect 14783 13753 14795 13787
rect 18064 13784 18092 13824
rect 20530 13812 20536 13864
rect 20588 13812 20594 13864
rect 14737 13747 14795 13753
rect 17604 13756 18092 13784
rect 17604 13728 17632 13756
rect 19702 13744 19708 13796
rect 19760 13784 19766 13796
rect 20640 13784 20668 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 22152 13892 22201 13920
rect 22152 13880 22158 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 21542 13852 21548 13864
rect 21008 13824 21548 13852
rect 21008 13793 21036 13824
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 22204 13852 22232 13883
rect 22462 13880 22468 13932
rect 22520 13880 22526 13932
rect 22646 13880 22652 13932
rect 22704 13880 22710 13932
rect 23106 13880 23112 13932
rect 23164 13880 23170 13932
rect 23198 13880 23204 13932
rect 23256 13880 23262 13932
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 22480 13852 22508 13880
rect 22922 13852 22928 13864
rect 22204 13824 22416 13852
rect 22480 13824 22928 13852
rect 19760 13756 20668 13784
rect 20993 13787 21051 13793
rect 19760 13744 19766 13756
rect 20993 13753 21005 13787
rect 21039 13753 21051 13787
rect 20993 13747 21051 13753
rect 22186 13744 22192 13796
rect 22244 13744 22250 13796
rect 4246 13716 4252 13728
rect 3252 13688 4252 13716
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 5534 13676 5540 13728
rect 5592 13676 5598 13728
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6236 13688 6469 13716
rect 6236 13676 6242 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6457 13679 6515 13685
rect 10042 13676 10048 13728
rect 10100 13676 10106 13728
rect 10502 13676 10508 13728
rect 10560 13676 10566 13728
rect 11320 13719 11378 13725
rect 11320 13685 11332 13719
rect 11366 13716 11378 13719
rect 12434 13716 12440 13728
rect 11366 13688 12440 13716
rect 11366 13685 11378 13688
rect 11320 13679 11378 13685
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 13160 13719 13218 13725
rect 13160 13685 13172 13719
rect 13206 13716 13218 13719
rect 14182 13716 14188 13728
rect 13206 13688 14188 13716
rect 13206 13685 13218 13688
rect 13160 13679 13218 13685
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 15562 13676 15568 13728
rect 15620 13676 15626 13728
rect 16482 13676 16488 13728
rect 16540 13716 16546 13728
rect 17497 13719 17555 13725
rect 17497 13716 17509 13719
rect 16540 13688 17509 13716
rect 16540 13676 16546 13688
rect 17497 13685 17509 13688
rect 17543 13716 17555 13719
rect 17586 13716 17592 13728
rect 17543 13688 17592 13716
rect 17543 13685 17555 13688
rect 17497 13679 17555 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18230 13676 18236 13728
rect 18288 13676 18294 13728
rect 20349 13719 20407 13725
rect 20349 13685 20361 13719
rect 20395 13716 20407 13719
rect 20438 13716 20444 13728
rect 20395 13688 20444 13716
rect 20395 13685 20407 13688
rect 20349 13679 20407 13685
rect 20438 13676 20444 13688
rect 20496 13716 20502 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20496 13688 20821 13716
rect 20496 13676 20502 13688
rect 20809 13685 20821 13688
rect 20855 13685 20867 13719
rect 22388 13716 22416 13824
rect 22922 13812 22928 13824
rect 22980 13852 22986 13864
rect 23400 13852 23428 13883
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23845 13923 23903 13929
rect 23845 13920 23857 13923
rect 23532 13892 23857 13920
rect 23532 13880 23538 13892
rect 23845 13889 23857 13892
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24228 13929 24256 13960
rect 25225 13957 25237 13960
rect 25271 13957 25283 13991
rect 25225 13951 25283 13957
rect 25317 13991 25375 13997
rect 25317 13957 25329 13991
rect 25363 13957 25375 13991
rect 25317 13951 25375 13957
rect 26596 13991 26654 13997
rect 26596 13957 26608 13991
rect 26642 13988 26654 13991
rect 26896 13988 26924 14016
rect 26642 13960 26924 13988
rect 27816 13988 27844 14019
rect 28166 14016 28172 14068
rect 28224 14016 28230 14068
rect 28261 14059 28319 14065
rect 28261 14025 28273 14059
rect 28307 14056 28319 14059
rect 28350 14056 28356 14068
rect 28307 14028 28356 14056
rect 28307 14025 28319 14028
rect 28261 14019 28319 14025
rect 28350 14016 28356 14028
rect 28408 14016 28414 14068
rect 28442 14016 28448 14068
rect 28500 14056 28506 14068
rect 28629 14059 28687 14065
rect 28629 14056 28641 14059
rect 28500 14028 28641 14056
rect 28500 14016 28506 14028
rect 28629 14025 28641 14028
rect 28675 14025 28687 14059
rect 28629 14019 28687 14025
rect 28994 14016 29000 14068
rect 29052 14016 29058 14068
rect 29089 14059 29147 14065
rect 29089 14025 29101 14059
rect 29135 14056 29147 14059
rect 29135 14028 29960 14056
rect 29135 14025 29147 14028
rect 29089 14019 29147 14025
rect 29932 14000 29960 14028
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 31573 14059 31631 14065
rect 31573 14056 31585 14059
rect 30524 14028 31585 14056
rect 30524 14016 30530 14028
rect 31573 14025 31585 14028
rect 31619 14025 31631 14059
rect 32582 14056 32588 14068
rect 31573 14019 31631 14025
rect 31864 14028 32588 14056
rect 29730 13988 29736 14000
rect 27816 13960 29736 13988
rect 26642 13957 26654 13960
rect 26596 13951 26654 13957
rect 29730 13948 29736 13960
rect 29788 13948 29794 14000
rect 29914 13948 29920 14000
rect 29972 13948 29978 14000
rect 31386 13988 31392 14000
rect 31050 13960 31392 13988
rect 31386 13948 31392 13960
rect 31444 13948 31450 14000
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13889 24271 13923
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 24213 13883 24271 13889
rect 24320 13892 24869 13920
rect 22980 13824 23428 13852
rect 23952 13852 23980 13880
rect 24320 13852 24348 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25501 13923 25559 13929
rect 25501 13889 25513 13923
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 25777 13923 25835 13929
rect 25777 13889 25789 13923
rect 25823 13920 25835 13923
rect 27062 13920 27068 13932
rect 25823 13892 27068 13920
rect 25823 13889 25835 13892
rect 25777 13883 25835 13889
rect 23952 13824 24348 13852
rect 22980 13812 22986 13824
rect 24670 13812 24676 13864
rect 24728 13812 24734 13864
rect 25516 13852 25544 13883
rect 24780 13824 25544 13852
rect 24118 13744 24124 13796
rect 24176 13784 24182 13796
rect 24780 13784 24808 13824
rect 24176 13756 24808 13784
rect 24176 13744 24182 13756
rect 24946 13744 24952 13796
rect 25004 13784 25010 13796
rect 25608 13784 25636 13883
rect 27062 13880 27068 13892
rect 27120 13880 27126 13932
rect 28442 13880 28448 13932
rect 28500 13920 28506 13932
rect 28994 13920 29000 13932
rect 28500 13892 29000 13920
rect 28500 13880 28506 13892
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 29086 13880 29092 13932
rect 29144 13920 29150 13932
rect 29549 13923 29607 13929
rect 29549 13920 29561 13923
rect 29144 13892 29561 13920
rect 29144 13880 29150 13892
rect 29549 13889 29561 13892
rect 29595 13889 29607 13923
rect 29549 13883 29607 13889
rect 30834 13880 30840 13932
rect 30892 13880 30898 13932
rect 31478 13880 31484 13932
rect 31536 13880 31542 13932
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 25004 13756 25636 13784
rect 25004 13744 25010 13756
rect 24489 13719 24547 13725
rect 24489 13716 24501 13719
rect 22388 13688 24501 13716
rect 20809 13679 20867 13685
rect 24489 13685 24501 13688
rect 24535 13716 24547 13719
rect 24762 13716 24768 13728
rect 24535 13688 24768 13716
rect 24535 13685 24547 13688
rect 24489 13679 24547 13685
rect 24762 13676 24768 13688
rect 24820 13676 24826 13728
rect 25130 13676 25136 13728
rect 25188 13676 25194 13728
rect 25314 13676 25320 13728
rect 25372 13676 25378 13728
rect 25406 13676 25412 13728
rect 25464 13716 25470 13728
rect 26344 13716 26372 13815
rect 27798 13812 27804 13864
rect 27856 13852 27862 13864
rect 28353 13855 28411 13861
rect 28353 13852 28365 13855
rect 27856 13824 28365 13852
rect 27856 13812 27862 13824
rect 28353 13821 28365 13824
rect 28399 13852 28411 13855
rect 29181 13855 29239 13861
rect 29181 13852 29193 13855
rect 28399 13824 29193 13852
rect 28399 13821 28411 13824
rect 28353 13815 28411 13821
rect 29181 13821 29193 13824
rect 29227 13821 29239 13855
rect 29181 13815 29239 13821
rect 27338 13744 27344 13796
rect 27396 13744 27402 13796
rect 28166 13744 28172 13796
rect 28224 13784 28230 13796
rect 28810 13784 28816 13796
rect 28224 13756 28816 13784
rect 28224 13744 28230 13756
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 30852 13784 30880 13880
rect 31297 13855 31355 13861
rect 31297 13821 31309 13855
rect 31343 13852 31355 13855
rect 31496 13852 31524 13880
rect 31343 13824 31524 13852
rect 31864 13852 31892 14028
rect 32582 14016 32588 14028
rect 32640 14016 32646 14068
rect 32677 14059 32735 14065
rect 32677 14025 32689 14059
rect 32723 14056 32735 14059
rect 32858 14056 32864 14068
rect 32723 14028 32864 14056
rect 32723 14025 32735 14028
rect 32677 14019 32735 14025
rect 32858 14016 32864 14028
rect 32916 14016 32922 14068
rect 33318 14056 33324 14068
rect 33152 14028 33324 14056
rect 32490 13948 32496 14000
rect 32548 13988 32554 14000
rect 33152 13997 33180 14028
rect 33318 14016 33324 14028
rect 33376 14016 33382 14068
rect 33778 14016 33784 14068
rect 33836 14056 33842 14068
rect 34701 14059 34759 14065
rect 34701 14056 34713 14059
rect 33836 14028 34713 14056
rect 33836 14016 33842 14028
rect 34701 14025 34713 14028
rect 34747 14025 34759 14059
rect 34701 14019 34759 14025
rect 35713 14059 35771 14065
rect 35713 14025 35725 14059
rect 35759 14056 35771 14059
rect 35986 14056 35992 14068
rect 35759 14028 35992 14056
rect 35759 14025 35771 14028
rect 35713 14019 35771 14025
rect 35986 14016 35992 14028
rect 36044 14016 36050 14068
rect 36173 14059 36231 14065
rect 36173 14025 36185 14059
rect 36219 14056 36231 14059
rect 36538 14056 36544 14068
rect 36219 14028 36544 14056
rect 36219 14025 36231 14028
rect 36173 14019 36231 14025
rect 36538 14016 36544 14028
rect 36596 14016 36602 14068
rect 36906 14016 36912 14068
rect 36964 14056 36970 14068
rect 38470 14056 38476 14068
rect 36964 14028 38476 14056
rect 36964 14016 36970 14028
rect 38470 14016 38476 14028
rect 38528 14016 38534 14068
rect 39482 14016 39488 14068
rect 39540 14056 39546 14068
rect 41141 14059 41199 14065
rect 41141 14056 41153 14059
rect 39540 14028 41153 14056
rect 39540 14016 39546 14028
rect 41141 14025 41153 14028
rect 41187 14025 41199 14059
rect 41141 14019 41199 14025
rect 41785 14059 41843 14065
rect 41785 14025 41797 14059
rect 41831 14025 41843 14059
rect 41785 14019 41843 14025
rect 33137 13991 33195 13997
rect 32548 13960 32904 13988
rect 32548 13948 32554 13960
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13920 31999 13923
rect 32582 13920 32588 13932
rect 31987 13892 32588 13920
rect 31987 13889 31999 13892
rect 31941 13883 31999 13889
rect 32582 13880 32588 13892
rect 32640 13880 32646 13932
rect 32876 13861 32904 13960
rect 33137 13957 33149 13991
rect 33183 13957 33195 13991
rect 33137 13951 33195 13957
rect 33410 13948 33416 14000
rect 33468 13988 33474 14000
rect 36081 13991 36139 13997
rect 33468 13960 33626 13988
rect 33468 13948 33474 13960
rect 36081 13957 36093 13991
rect 36127 13988 36139 13991
rect 37737 13991 37795 13997
rect 36127 13960 37228 13988
rect 36127 13957 36139 13960
rect 36081 13951 36139 13957
rect 37200 13932 37228 13960
rect 37737 13957 37749 13991
rect 37783 13988 37795 13991
rect 37826 13988 37832 14000
rect 37783 13960 37832 13988
rect 37783 13957 37795 13960
rect 37737 13951 37795 13957
rect 37826 13948 37832 13960
rect 37884 13948 37890 14000
rect 38194 13948 38200 14000
rect 38252 13948 38258 14000
rect 40218 13948 40224 14000
rect 40276 13948 40282 14000
rect 35066 13880 35072 13932
rect 35124 13880 35130 13932
rect 35176 13892 36492 13920
rect 32033 13855 32091 13861
rect 32033 13852 32045 13855
rect 31864 13824 32045 13852
rect 31343 13821 31355 13824
rect 31297 13815 31355 13821
rect 31864 13784 31892 13824
rect 32033 13821 32045 13824
rect 32079 13821 32091 13855
rect 32033 13815 32091 13821
rect 32125 13855 32183 13861
rect 32125 13821 32137 13855
rect 32171 13821 32183 13855
rect 32125 13815 32183 13821
rect 32861 13855 32919 13861
rect 32861 13821 32873 13855
rect 32907 13821 32919 13855
rect 32861 13815 32919 13821
rect 30852 13756 31892 13784
rect 31938 13744 31944 13796
rect 31996 13784 32002 13796
rect 32140 13784 32168 13815
rect 34422 13812 34428 13864
rect 34480 13852 34486 13864
rect 34790 13852 34796 13864
rect 34480 13824 34796 13852
rect 34480 13812 34486 13824
rect 34790 13812 34796 13824
rect 34848 13852 34854 13864
rect 35176 13861 35204 13892
rect 35161 13855 35219 13861
rect 35161 13852 35173 13855
rect 34848 13824 35173 13852
rect 34848 13812 34854 13824
rect 35161 13821 35173 13824
rect 35207 13821 35219 13855
rect 35161 13815 35219 13821
rect 35253 13855 35311 13861
rect 35253 13821 35265 13855
rect 35299 13821 35311 13855
rect 35253 13815 35311 13821
rect 35268 13784 35296 13815
rect 35710 13812 35716 13864
rect 35768 13852 35774 13864
rect 36354 13852 36360 13864
rect 35768 13824 36360 13852
rect 35768 13812 35774 13824
rect 36354 13812 36360 13824
rect 36412 13812 36418 13864
rect 31996 13756 32996 13784
rect 31996 13744 32002 13756
rect 27356 13716 27384 13744
rect 25464 13688 27384 13716
rect 29812 13719 29870 13725
rect 25464 13676 25470 13688
rect 29812 13685 29824 13719
rect 29858 13716 29870 13719
rect 30558 13716 30564 13728
rect 29858 13688 30564 13716
rect 29858 13685 29870 13688
rect 29812 13679 29870 13685
rect 30558 13676 30564 13688
rect 30616 13676 30622 13728
rect 32968 13716 32996 13756
rect 34532 13756 35296 13784
rect 36464 13784 36492 13892
rect 36538 13880 36544 13932
rect 36596 13920 36602 13932
rect 36725 13923 36783 13929
rect 36725 13920 36737 13923
rect 36596 13892 36737 13920
rect 36596 13880 36602 13892
rect 36725 13889 36737 13892
rect 36771 13889 36783 13923
rect 36725 13883 36783 13889
rect 37182 13880 37188 13932
rect 37240 13880 37246 13932
rect 37274 13880 37280 13932
rect 37332 13920 37338 13932
rect 37461 13923 37519 13929
rect 37461 13920 37473 13923
rect 37332 13892 37473 13920
rect 37332 13880 37338 13892
rect 37461 13889 37473 13892
rect 37507 13889 37519 13923
rect 37461 13883 37519 13889
rect 40954 13880 40960 13932
rect 41012 13920 41018 13932
rect 41325 13923 41383 13929
rect 41012 13892 41184 13920
rect 41012 13880 41018 13892
rect 37090 13812 37096 13864
rect 37148 13812 37154 13864
rect 39206 13852 39212 13864
rect 37200 13824 39212 13852
rect 37200 13784 37228 13824
rect 39206 13812 39212 13824
rect 39264 13812 39270 13864
rect 39301 13855 39359 13861
rect 39301 13821 39313 13855
rect 39347 13821 39359 13855
rect 39301 13815 39359 13821
rect 36464 13756 37228 13784
rect 33226 13716 33232 13728
rect 32968 13688 33232 13716
rect 33226 13676 33232 13688
rect 33284 13716 33290 13728
rect 33502 13716 33508 13728
rect 33284 13688 33508 13716
rect 33284 13676 33290 13688
rect 33502 13676 33508 13688
rect 33560 13716 33566 13728
rect 34422 13716 34428 13728
rect 33560 13688 34428 13716
rect 33560 13676 33566 13688
rect 34422 13676 34428 13688
rect 34480 13716 34486 13728
rect 34532 13716 34560 13756
rect 38838 13744 38844 13796
rect 38896 13784 38902 13796
rect 39316 13784 39344 13815
rect 39574 13812 39580 13864
rect 39632 13812 39638 13864
rect 39666 13812 39672 13864
rect 39724 13852 39730 13864
rect 41049 13855 41107 13861
rect 41049 13852 41061 13855
rect 39724 13824 41061 13852
rect 39724 13812 39730 13824
rect 41049 13821 41061 13824
rect 41095 13821 41107 13855
rect 41156 13852 41184 13892
rect 41325 13889 41337 13923
rect 41371 13920 41383 13923
rect 41800 13920 41828 14019
rect 42242 14016 42248 14068
rect 42300 14016 42306 14068
rect 41371 13892 41828 13920
rect 42153 13923 42211 13929
rect 41371 13889 41383 13892
rect 41325 13883 41383 13889
rect 42153 13889 42165 13923
rect 42199 13889 42211 13923
rect 42153 13883 42211 13889
rect 42168 13852 42196 13883
rect 41156 13824 42196 13852
rect 42337 13855 42395 13861
rect 41049 13815 41107 13821
rect 42337 13821 42349 13855
rect 42383 13821 42395 13855
rect 42337 13815 42395 13821
rect 38896 13756 39344 13784
rect 38896 13744 38902 13756
rect 34480 13688 34560 13716
rect 34480 13676 34486 13688
rect 34606 13676 34612 13728
rect 34664 13676 34670 13728
rect 37185 13719 37243 13725
rect 37185 13685 37197 13719
rect 37231 13716 37243 13719
rect 37274 13716 37280 13728
rect 37231 13688 37280 13716
rect 37231 13685 37243 13688
rect 37185 13679 37243 13685
rect 37274 13676 37280 13688
rect 37332 13676 37338 13728
rect 37369 13719 37427 13725
rect 37369 13685 37381 13719
rect 37415 13716 37427 13719
rect 37550 13716 37556 13728
rect 37415 13688 37556 13716
rect 37415 13685 37427 13688
rect 37369 13679 37427 13685
rect 37550 13676 37556 13688
rect 37608 13676 37614 13728
rect 39206 13676 39212 13728
rect 39264 13676 39270 13728
rect 39298 13676 39304 13728
rect 39356 13716 39362 13728
rect 42352 13716 42380 13815
rect 42794 13812 42800 13864
rect 42852 13812 42858 13864
rect 43346 13744 43352 13796
rect 43404 13784 43410 13796
rect 43533 13787 43591 13793
rect 43533 13784 43545 13787
rect 43404 13756 43545 13784
rect 43404 13744 43410 13756
rect 43533 13753 43545 13756
rect 43579 13784 43591 13787
rect 43898 13784 43904 13796
rect 43579 13756 43904 13784
rect 43579 13753 43591 13756
rect 43533 13747 43591 13753
rect 43898 13744 43904 13756
rect 43956 13784 43962 13796
rect 44726 13784 44732 13796
rect 43956 13756 44732 13784
rect 43956 13744 43962 13756
rect 44726 13744 44732 13756
rect 44784 13744 44790 13796
rect 39356 13688 42380 13716
rect 39356 13676 39362 13688
rect 43070 13676 43076 13728
rect 43128 13716 43134 13728
rect 43165 13719 43223 13725
rect 43165 13716 43177 13719
rect 43128 13688 43177 13716
rect 43128 13676 43134 13688
rect 43165 13685 43177 13688
rect 43211 13716 43223 13719
rect 44269 13719 44327 13725
rect 44269 13716 44281 13719
rect 43211 13688 44281 13716
rect 43211 13685 43223 13688
rect 43165 13679 43223 13685
rect 44269 13685 44281 13688
rect 44315 13716 44327 13719
rect 44358 13716 44364 13728
rect 44315 13688 44364 13716
rect 44315 13685 44327 13688
rect 44269 13679 44327 13685
rect 44358 13676 44364 13688
rect 44416 13676 44422 13728
rect 44542 13676 44548 13728
rect 44600 13716 44606 13728
rect 45097 13719 45155 13725
rect 45097 13716 45109 13719
rect 44600 13688 45109 13716
rect 44600 13676 44606 13688
rect 45097 13685 45109 13688
rect 45143 13685 45155 13719
rect 45097 13679 45155 13685
rect 460 13626 45540 13648
rect 460 13574 3570 13626
rect 3622 13574 3634 13626
rect 3686 13574 3698 13626
rect 3750 13574 3762 13626
rect 3814 13574 3826 13626
rect 3878 13574 8570 13626
rect 8622 13574 8634 13626
rect 8686 13574 8698 13626
rect 8750 13574 8762 13626
rect 8814 13574 8826 13626
rect 8878 13574 13570 13626
rect 13622 13574 13634 13626
rect 13686 13574 13698 13626
rect 13750 13574 13762 13626
rect 13814 13574 13826 13626
rect 13878 13574 18570 13626
rect 18622 13574 18634 13626
rect 18686 13574 18698 13626
rect 18750 13574 18762 13626
rect 18814 13574 18826 13626
rect 18878 13574 23570 13626
rect 23622 13574 23634 13626
rect 23686 13574 23698 13626
rect 23750 13574 23762 13626
rect 23814 13574 23826 13626
rect 23878 13574 28570 13626
rect 28622 13574 28634 13626
rect 28686 13574 28698 13626
rect 28750 13574 28762 13626
rect 28814 13574 28826 13626
rect 28878 13574 33570 13626
rect 33622 13574 33634 13626
rect 33686 13574 33698 13626
rect 33750 13574 33762 13626
rect 33814 13574 33826 13626
rect 33878 13574 38570 13626
rect 38622 13574 38634 13626
rect 38686 13574 38698 13626
rect 38750 13574 38762 13626
rect 38814 13574 38826 13626
rect 38878 13574 43570 13626
rect 43622 13574 43634 13626
rect 43686 13574 43698 13626
rect 43750 13574 43762 13626
rect 43814 13574 43826 13626
rect 43878 13574 45540 13626
rect 460 13552 45540 13574
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4246 13512 4252 13524
rect 3927 13484 4252 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4246 13472 4252 13484
rect 4304 13512 4310 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 4304 13484 4721 13512
rect 4304 13472 4310 13484
rect 4709 13481 4721 13484
rect 4755 13512 4767 13515
rect 5537 13515 5595 13521
rect 5537 13512 5549 13515
rect 4755 13484 5549 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 5537 13481 5549 13484
rect 5583 13481 5595 13515
rect 5537 13475 5595 13481
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 7006 13512 7012 13524
rect 5684 13484 7012 13512
rect 5684 13472 5690 13484
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 10226 13512 10232 13524
rect 8803 13484 10232 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11333 13515 11391 13521
rect 11333 13481 11345 13515
rect 11379 13512 11391 13515
rect 11422 13512 11428 13524
rect 11379 13484 11428 13512
rect 11379 13481 11391 13484
rect 11333 13475 11391 13481
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12308 13484 12848 13512
rect 12308 13472 12314 13484
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 5721 13447 5779 13453
rect 5721 13444 5733 13447
rect 5316 13416 5733 13444
rect 5316 13404 5322 13416
rect 5721 13413 5733 13416
rect 5767 13413 5779 13447
rect 5721 13407 5779 13413
rect 9582 13404 9588 13456
rect 9640 13404 9646 13456
rect 12820 13444 12848 13484
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 12952 13484 13185 13512
rect 12952 13472 12958 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 16485 13515 16543 13521
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 17034 13512 17040 13524
rect 16531 13484 17040 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 18012 13484 18429 13512
rect 18012 13472 18018 13484
rect 18417 13481 18429 13484
rect 18463 13512 18475 13515
rect 18690 13512 18696 13524
rect 18463 13484 18696 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 18690 13472 18696 13484
rect 18748 13472 18754 13524
rect 19337 13515 19395 13521
rect 18800 13484 19104 13512
rect 12820 13416 13492 13444
rect 5905 13379 5963 13385
rect 5092 13348 5856 13376
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 5092 13181 5120 13348
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 5828 13308 5856 13348
rect 5905 13345 5917 13379
rect 5951 13376 5963 13379
rect 6914 13376 6920 13388
rect 5951 13348 6920 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13376 9459 13379
rect 9600 13376 9628 13404
rect 9447 13348 9628 13376
rect 9861 13379 9919 13385
rect 9447 13345 9459 13348
rect 9401 13339 9459 13345
rect 9861 13345 9873 13379
rect 9907 13376 9919 13379
rect 10502 13376 10508 13388
rect 9907 13348 10508 13376
rect 9907 13345 9919 13348
rect 9861 13339 9919 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 13464 13376 13492 13416
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 18800 13444 18828 13484
rect 15712 13416 16436 13444
rect 15712 13404 15718 13416
rect 13725 13379 13783 13385
rect 13725 13376 13737 13379
rect 13464 13348 13737 13376
rect 13725 13345 13737 13348
rect 13771 13345 13783 13379
rect 13725 13339 13783 13345
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14332 13348 15976 13376
rect 14332 13336 14338 13348
rect 6178 13308 6184 13320
rect 5828 13280 6184 13308
rect 6178 13268 6184 13280
rect 6236 13308 6242 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6236 13280 6285 13308
rect 6236 13268 6242 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 9490 13308 9496 13320
rect 8711 13280 9496 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9582 13268 9588 13320
rect 9640 13268 9646 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 11388 13280 11437 13308
rect 11388 13268 11394 13280
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 5552 13240 5580 13268
rect 6549 13243 6607 13249
rect 6549 13240 6561 13243
rect 5552 13212 6561 13240
rect 6549 13209 6561 13212
rect 6595 13209 6607 13243
rect 6549 13203 6607 13209
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 9950 13240 9956 13252
rect 6696 13212 7038 13240
rect 8036 13212 9956 13240
rect 6696 13200 6702 13212
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 3476 13144 4353 13172
rect 3476 13132 3482 13144
rect 4341 13141 4353 13144
rect 4387 13172 4399 13175
rect 5077 13175 5135 13181
rect 5077 13172 5089 13175
rect 4387 13144 5089 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 5077 13141 5089 13144
rect 5123 13141 5135 13175
rect 5077 13135 5135 13141
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 8036 13181 8064 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 11440 13240 11468 13271
rect 10192 13212 10350 13240
rect 11440 13212 11652 13240
rect 10192 13200 10198 13212
rect 11624 13184 11652 13212
rect 11698 13200 11704 13252
rect 11756 13200 11762 13252
rect 12158 13200 12164 13252
rect 12216 13200 12222 13252
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8478 13132 8484 13184
rect 8536 13132 8542 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 11514 13172 11520 13184
rect 9263 13144 11520 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 11606 13132 11612 13184
rect 11664 13172 11670 13184
rect 13464 13172 13492 13271
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15948 13317 15976 13348
rect 16022 13336 16028 13388
rect 16080 13336 16086 13388
rect 16408 13317 16436 13416
rect 18064 13416 18828 13444
rect 19076 13444 19104 13484
rect 19337 13481 19349 13515
rect 19383 13481 19395 13515
rect 19337 13475 19395 13481
rect 19153 13447 19211 13453
rect 19153 13444 19165 13447
rect 19076 13416 19165 13444
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13376 17003 13379
rect 18064 13376 18092 13416
rect 19153 13413 19165 13416
rect 19199 13413 19211 13447
rect 19352 13444 19380 13475
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 19484 13484 19717 13512
rect 19484 13472 19490 13484
rect 19705 13481 19717 13484
rect 19751 13481 19763 13515
rect 19705 13475 19763 13481
rect 19978 13472 19984 13524
rect 20036 13472 20042 13524
rect 20152 13515 20210 13521
rect 20152 13481 20164 13515
rect 20198 13512 20210 13515
rect 20898 13512 20904 13524
rect 20198 13484 20904 13512
rect 20198 13481 20210 13484
rect 20152 13475 20210 13481
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21910 13472 21916 13524
rect 21968 13512 21974 13524
rect 22833 13515 22891 13521
rect 21968 13484 22784 13512
rect 21968 13472 21974 13484
rect 19996 13444 20024 13472
rect 22278 13444 22284 13456
rect 19352 13416 20024 13444
rect 22020 13416 22284 13444
rect 19153 13407 19211 13413
rect 16991 13348 18092 13376
rect 16991 13345 17003 13348
rect 16945 13339 17003 13345
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 21910 13376 21916 13388
rect 18564 13348 18828 13376
rect 18564 13336 18570 13348
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16540 13280 16681 13308
rect 16540 13268 16546 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 18690 13308 18696 13320
rect 18647 13280 18696 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 18800 13317 18828 13348
rect 18892 13348 19564 13376
rect 18892 13320 18920 13348
rect 19536 13320 19564 13348
rect 19720 13348 21916 13376
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18874 13268 18880 13320
rect 18932 13268 18938 13320
rect 18966 13268 18972 13320
rect 19024 13268 19030 13320
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 13998 13200 14004 13252
rect 14056 13200 14062 13252
rect 14366 13200 14372 13252
rect 14424 13200 14430 13252
rect 19150 13240 19156 13252
rect 18170 13212 19156 13240
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 19242 13200 19248 13252
rect 19300 13200 19306 13252
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 19444 13240 19472 13271
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19576 13280 19621 13308
rect 19576 13268 19582 13280
rect 19720 13240 19748 13348
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22020 13317 22048 13416
rect 22278 13404 22284 13416
rect 22336 13444 22342 13456
rect 22554 13444 22560 13456
rect 22336 13416 22560 13444
rect 22336 13404 22342 13416
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13376 22155 13379
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22143 13348 22661 13376
rect 22143 13345 22155 13348
rect 22097 13339 22155 13345
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22756 13376 22784 13484
rect 22833 13481 22845 13515
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 22848 13444 22876 13475
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23293 13515 23351 13521
rect 23293 13512 23305 13515
rect 23164 13484 23305 13512
rect 23164 13472 23170 13484
rect 23293 13481 23305 13484
rect 23339 13481 23351 13515
rect 24026 13512 24032 13524
rect 23293 13475 23351 13481
rect 23400 13484 24032 13512
rect 23400 13444 23428 13484
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24305 13515 24363 13521
rect 24305 13481 24317 13515
rect 24351 13512 24363 13515
rect 24394 13512 24400 13524
rect 24351 13484 24400 13512
rect 24351 13481 24363 13484
rect 24305 13475 24363 13481
rect 24394 13472 24400 13484
rect 24452 13512 24458 13524
rect 25498 13512 25504 13524
rect 24452 13484 25504 13512
rect 24452 13472 24458 13484
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 26602 13472 26608 13524
rect 26660 13472 26666 13524
rect 26878 13472 26884 13524
rect 26936 13472 26942 13524
rect 27062 13472 27068 13524
rect 27120 13472 27126 13524
rect 27154 13472 27160 13524
rect 27212 13512 27218 13524
rect 28442 13512 28448 13524
rect 27212 13484 28448 13512
rect 27212 13472 27218 13484
rect 28442 13472 28448 13484
rect 28500 13512 28506 13524
rect 28718 13512 28724 13524
rect 28500 13484 28724 13512
rect 28500 13472 28506 13484
rect 28718 13472 28724 13484
rect 28776 13472 28782 13524
rect 29638 13472 29644 13524
rect 29696 13472 29702 13524
rect 29822 13472 29828 13524
rect 29880 13512 29886 13524
rect 30101 13515 30159 13521
rect 30101 13512 30113 13515
rect 29880 13484 30113 13512
rect 29880 13472 29886 13484
rect 30101 13481 30113 13484
rect 30147 13481 30159 13515
rect 30101 13475 30159 13481
rect 31478 13472 31484 13524
rect 31536 13512 31542 13524
rect 32214 13512 32220 13524
rect 31536 13484 32220 13512
rect 31536 13472 31542 13484
rect 32214 13472 32220 13484
rect 32272 13472 32278 13524
rect 32582 13472 32588 13524
rect 32640 13472 32646 13524
rect 34514 13472 34520 13524
rect 34572 13512 34578 13524
rect 34572 13484 35572 13512
rect 34572 13472 34578 13484
rect 24489 13447 24547 13453
rect 24489 13444 24501 13447
rect 22848 13416 23428 13444
rect 23860 13416 24501 13444
rect 23860 13376 23888 13416
rect 24489 13413 24501 13416
rect 24535 13444 24547 13447
rect 24670 13444 24676 13456
rect 24535 13416 24676 13444
rect 24535 13413 24547 13416
rect 24489 13407 24547 13413
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 28350 13404 28356 13456
rect 28408 13444 28414 13456
rect 28408 13416 30420 13444
rect 28408 13404 28414 13416
rect 24578 13376 24584 13388
rect 22756 13348 23888 13376
rect 23952 13348 24584 13376
rect 22649 13339 22707 13345
rect 22186 13317 22192 13320
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 22005 13311 22063 13317
rect 22005 13277 22017 13311
rect 22051 13277 22063 13311
rect 22183 13308 22192 13317
rect 22147 13280 22192 13308
rect 22005 13271 22063 13277
rect 22183 13271 22192 13280
rect 19392 13212 19748 13240
rect 19392 13200 19398 13212
rect 11664 13144 13492 13172
rect 14016 13172 14044 13200
rect 15197 13175 15255 13181
rect 15197 13172 15209 13175
rect 14016 13144 15209 13172
rect 11664 13132 11670 13144
rect 15197 13141 15209 13144
rect 15243 13141 15255 13175
rect 15197 13135 15255 13141
rect 18414 13132 18420 13184
rect 18472 13172 18478 13184
rect 18690 13172 18696 13184
rect 18472 13144 18696 13172
rect 18472 13132 18478 13144
rect 18690 13132 18696 13144
rect 18748 13172 18754 13184
rect 19794 13172 19800 13184
rect 18748 13144 19800 13172
rect 18748 13132 18754 13144
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 19904 13172 19932 13271
rect 22186 13268 22192 13271
rect 22244 13268 22250 13320
rect 22303 13311 22361 13317
rect 22303 13277 22315 13311
rect 22349 13308 22361 13311
rect 22830 13308 22836 13320
rect 22349 13280 22836 13308
rect 22349 13277 22361 13280
rect 22303 13271 22361 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23492 13317 23520 13348
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 23842 13268 23848 13320
rect 23900 13268 23906 13320
rect 23952 13317 23980 13348
rect 24578 13336 24584 13348
rect 24636 13376 24642 13388
rect 24762 13376 24768 13388
rect 24636 13348 24768 13376
rect 24636 13336 24642 13348
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 25133 13379 25191 13385
rect 25133 13345 25145 13379
rect 25179 13376 25191 13379
rect 26418 13376 26424 13388
rect 25179 13348 26424 13376
rect 25179 13345 25191 13348
rect 25133 13339 25191 13345
rect 26418 13336 26424 13348
rect 26476 13336 26482 13388
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 27062 13376 27068 13388
rect 26568 13348 27068 13376
rect 26568 13336 26574 13348
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 27338 13336 27344 13388
rect 27396 13336 27402 13388
rect 28534 13336 28540 13388
rect 28592 13376 28598 13388
rect 28902 13376 28908 13388
rect 28592 13348 28908 13376
rect 28592 13336 28598 13348
rect 28902 13336 28908 13348
rect 28960 13376 28966 13388
rect 30392 13376 30420 13416
rect 30466 13404 30472 13456
rect 30524 13444 30530 13456
rect 30561 13447 30619 13453
rect 30561 13444 30573 13447
rect 30524 13416 30573 13444
rect 30524 13404 30530 13416
rect 30561 13413 30573 13416
rect 30607 13413 30619 13447
rect 32232 13444 32260 13472
rect 33410 13444 33416 13456
rect 32232 13416 33416 13444
rect 30561 13407 30619 13413
rect 33410 13404 33416 13416
rect 33468 13444 33474 13456
rect 33870 13444 33876 13456
rect 33468 13416 33876 13444
rect 33468 13404 33474 13416
rect 33870 13404 33876 13416
rect 33928 13404 33934 13456
rect 33042 13376 33048 13388
rect 28960 13348 29592 13376
rect 30392 13348 33048 13376
rect 28960 13336 28966 13348
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13277 23995 13311
rect 23937 13271 23995 13277
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13308 24363 13311
rect 24486 13308 24492 13320
rect 24351 13280 24492 13308
rect 24351 13277 24363 13280
rect 24305 13271 24363 13277
rect 24486 13268 24492 13280
rect 24544 13268 24550 13320
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 26878 13308 26884 13320
rect 26266 13280 26884 13308
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 26970 13268 26976 13320
rect 27028 13268 27034 13320
rect 27608 13311 27666 13317
rect 27608 13277 27620 13311
rect 27654 13308 27666 13311
rect 28074 13308 28080 13320
rect 27654 13280 28080 13308
rect 27654 13277 27666 13280
rect 27608 13271 27666 13277
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 28626 13268 28632 13320
rect 28684 13308 28690 13320
rect 29181 13311 29239 13317
rect 29181 13308 29193 13311
rect 28684 13280 29193 13308
rect 28684 13268 28690 13280
rect 29181 13277 29193 13280
rect 29227 13277 29239 13311
rect 29181 13271 29239 13277
rect 29273 13311 29331 13317
rect 29273 13277 29285 13311
rect 29319 13277 29331 13311
rect 29273 13271 29331 13277
rect 21542 13240 21548 13252
rect 21390 13212 21548 13240
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 23198 13200 23204 13252
rect 23256 13240 23262 13252
rect 23256 13212 25544 13240
rect 23256 13200 23262 13212
rect 20346 13172 20352 13184
rect 19904 13144 20352 13172
rect 20346 13132 20352 13144
rect 20404 13172 20410 13184
rect 20806 13172 20812 13184
rect 20404 13144 20812 13172
rect 20404 13132 20410 13144
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 22462 13132 22468 13184
rect 22520 13132 22526 13184
rect 23109 13175 23167 13181
rect 23109 13141 23121 13175
rect 23155 13172 23167 13175
rect 23474 13172 23480 13184
rect 23155 13144 23480 13172
rect 23155 13141 23167 13144
rect 23109 13135 23167 13141
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24670 13172 24676 13184
rect 24084 13144 24676 13172
rect 24084 13132 24090 13144
rect 24670 13132 24676 13144
rect 24728 13132 24734 13184
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 25130 13172 25136 13184
rect 24912 13144 25136 13172
rect 24912 13132 24918 13144
rect 25130 13132 25136 13144
rect 25188 13172 25194 13184
rect 25406 13172 25412 13184
rect 25188 13144 25412 13172
rect 25188 13132 25194 13144
rect 25406 13132 25412 13144
rect 25464 13132 25470 13184
rect 25516 13172 25544 13212
rect 26418 13200 26424 13252
rect 26476 13240 26482 13252
rect 26697 13243 26755 13249
rect 26697 13240 26709 13243
rect 26476 13212 26709 13240
rect 26476 13200 26482 13212
rect 26697 13209 26709 13212
rect 26743 13240 26755 13243
rect 26988 13240 27016 13268
rect 26743 13212 27016 13240
rect 27632 13212 28856 13240
rect 26743 13209 26755 13212
rect 26697 13203 26755 13209
rect 27632 13184 27660 13212
rect 26786 13172 26792 13184
rect 25516 13144 26792 13172
rect 26786 13132 26792 13144
rect 26844 13172 26850 13184
rect 26897 13175 26955 13181
rect 26897 13172 26909 13175
rect 26844 13144 26909 13172
rect 26844 13132 26850 13144
rect 26897 13141 26909 13144
rect 26943 13141 26955 13175
rect 26897 13135 26955 13141
rect 27614 13132 27620 13184
rect 27672 13132 27678 13184
rect 27890 13132 27896 13184
rect 27948 13172 27954 13184
rect 28074 13172 28080 13184
rect 27948 13144 28080 13172
rect 27948 13132 27954 13144
rect 28074 13132 28080 13144
rect 28132 13172 28138 13184
rect 28626 13172 28632 13184
rect 28132 13144 28632 13172
rect 28132 13132 28138 13144
rect 28626 13132 28632 13144
rect 28684 13132 28690 13184
rect 28718 13132 28724 13184
rect 28776 13132 28782 13184
rect 28828 13172 28856 13212
rect 29086 13200 29092 13252
rect 29144 13240 29150 13252
rect 29288 13240 29316 13271
rect 29362 13268 29368 13320
rect 29420 13268 29426 13320
rect 29564 13317 29592 13348
rect 33042 13336 33048 13348
rect 33100 13376 33106 13388
rect 33137 13379 33195 13385
rect 33137 13376 33149 13379
rect 33100 13348 33149 13376
rect 33100 13336 33106 13348
rect 33137 13345 33149 13348
rect 33183 13345 33195 13379
rect 33137 13339 33195 13345
rect 33226 13336 33232 13388
rect 33284 13336 33290 13388
rect 33318 13336 33324 13388
rect 33376 13376 33382 13388
rect 34057 13379 34115 13385
rect 34057 13376 34069 13379
rect 33376 13348 34069 13376
rect 33376 13336 33382 13348
rect 34057 13345 34069 13348
rect 34103 13345 34115 13379
rect 34057 13339 34115 13345
rect 29549 13311 29607 13317
rect 29549 13277 29561 13311
rect 29595 13277 29607 13311
rect 29549 13271 29607 13277
rect 29730 13268 29736 13320
rect 29788 13308 29794 13320
rect 29825 13311 29883 13317
rect 29825 13308 29837 13311
rect 29788 13280 29837 13308
rect 29788 13268 29794 13280
rect 29825 13277 29837 13280
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 30466 13268 30472 13320
rect 30524 13268 30530 13320
rect 30558 13268 30564 13320
rect 30616 13308 30622 13320
rect 30745 13311 30803 13317
rect 30745 13308 30757 13311
rect 30616 13280 30757 13308
rect 30616 13268 30622 13280
rect 30745 13277 30757 13280
rect 30791 13277 30803 13311
rect 30745 13271 30803 13277
rect 30834 13268 30840 13320
rect 30892 13268 30898 13320
rect 33689 13311 33747 13317
rect 33689 13277 33701 13311
rect 33735 13308 33747 13311
rect 33962 13308 33968 13320
rect 33735 13280 33968 13308
rect 33735 13277 33747 13280
rect 33689 13271 33747 13277
rect 33962 13268 33968 13280
rect 34020 13268 34026 13320
rect 35544 13308 35572 13484
rect 35894 13472 35900 13524
rect 35952 13472 35958 13524
rect 35986 13472 35992 13524
rect 36044 13512 36050 13524
rect 36354 13512 36360 13524
rect 36044 13484 36360 13512
rect 36044 13472 36050 13484
rect 36354 13472 36360 13484
rect 36412 13512 36418 13524
rect 36412 13484 37228 13512
rect 36412 13472 36418 13484
rect 35912 13444 35940 13472
rect 37200 13444 37228 13484
rect 37366 13472 37372 13524
rect 37424 13512 37430 13524
rect 37737 13515 37795 13521
rect 37737 13512 37749 13515
rect 37424 13484 37749 13512
rect 37424 13472 37430 13484
rect 37737 13481 37749 13484
rect 37783 13481 37795 13515
rect 37737 13475 37795 13481
rect 38010 13472 38016 13524
rect 38068 13512 38074 13524
rect 38105 13515 38163 13521
rect 38105 13512 38117 13515
rect 38068 13484 38117 13512
rect 38068 13472 38074 13484
rect 38105 13481 38117 13484
rect 38151 13481 38163 13515
rect 38105 13475 38163 13481
rect 39298 13472 39304 13524
rect 39356 13472 39362 13524
rect 40218 13472 40224 13524
rect 40276 13512 40282 13524
rect 40276 13484 40908 13512
rect 40276 13472 40282 13484
rect 39022 13444 39028 13456
rect 35912 13416 36032 13444
rect 37200 13416 39028 13444
rect 35618 13336 35624 13388
rect 35676 13376 35682 13388
rect 35897 13379 35955 13385
rect 35897 13376 35909 13379
rect 35676 13348 35909 13376
rect 35676 13336 35682 13348
rect 35897 13345 35909 13348
rect 35943 13345 35955 13379
rect 36004 13376 36032 13416
rect 36173 13379 36231 13385
rect 36173 13376 36185 13379
rect 36004 13348 36185 13376
rect 35897 13339 35955 13345
rect 36173 13345 36185 13348
rect 36219 13345 36231 13379
rect 36173 13339 36231 13345
rect 36538 13336 36544 13388
rect 36596 13376 36602 13388
rect 37645 13379 37703 13385
rect 37645 13376 37657 13379
rect 36596 13348 37657 13376
rect 36596 13336 36602 13348
rect 37645 13345 37657 13348
rect 37691 13345 37703 13379
rect 38194 13376 38200 13388
rect 37645 13339 37703 13345
rect 37844 13348 38200 13376
rect 35544 13280 35664 13308
rect 29144 13212 29316 13240
rect 30484 13240 30512 13268
rect 31113 13243 31171 13249
rect 31113 13240 31125 13243
rect 30484 13212 31125 13240
rect 29144 13200 29150 13212
rect 31113 13209 31125 13212
rect 31159 13209 31171 13243
rect 31113 13203 31171 13209
rect 31386 13200 31392 13252
rect 31444 13240 31450 13252
rect 31444 13212 31602 13240
rect 32416 13212 32720 13240
rect 31444 13200 31450 13212
rect 28905 13175 28963 13181
rect 28905 13172 28917 13175
rect 28828 13144 28917 13172
rect 28905 13141 28917 13144
rect 28951 13172 28963 13175
rect 30926 13172 30932 13184
rect 28951 13144 30932 13172
rect 28951 13141 28963 13144
rect 28905 13135 28963 13141
rect 30926 13132 30932 13144
rect 30984 13132 30990 13184
rect 31478 13132 31484 13184
rect 31536 13172 31542 13184
rect 32416 13172 32444 13212
rect 32692 13181 32720 13212
rect 33870 13200 33876 13252
rect 33928 13200 33934 13252
rect 34330 13200 34336 13252
rect 34388 13200 34394 13252
rect 35636 13240 35664 13280
rect 37550 13268 37556 13320
rect 37608 13308 37614 13320
rect 37737 13311 37795 13317
rect 37737 13308 37749 13311
rect 37608 13280 37749 13308
rect 37608 13268 37614 13280
rect 37737 13277 37749 13280
rect 37783 13277 37795 13311
rect 37737 13271 37795 13277
rect 37642 13240 37648 13252
rect 34440 13212 34822 13240
rect 35636 13212 35940 13240
rect 37398 13212 37648 13240
rect 31536 13144 32444 13172
rect 32677 13175 32735 13181
rect 31536 13132 31542 13144
rect 32677 13141 32689 13175
rect 32723 13141 32735 13175
rect 32677 13135 32735 13141
rect 33042 13132 33048 13184
rect 33100 13132 33106 13184
rect 33502 13132 33508 13184
rect 33560 13132 33566 13184
rect 33888 13172 33916 13200
rect 34440 13172 34468 13212
rect 34716 13184 34744 13212
rect 33888 13144 34468 13172
rect 34698 13132 34704 13184
rect 34756 13132 34762 13184
rect 35066 13132 35072 13184
rect 35124 13172 35130 13184
rect 35805 13175 35863 13181
rect 35805 13172 35817 13175
rect 35124 13144 35817 13172
rect 35124 13132 35130 13144
rect 35805 13141 35817 13144
rect 35851 13141 35863 13175
rect 35912 13172 35940 13212
rect 37642 13200 37648 13212
rect 37700 13240 37706 13252
rect 37844 13240 37872 13348
rect 38194 13336 38200 13348
rect 38252 13336 38258 13388
rect 38764 13385 38792 13416
rect 39022 13404 39028 13416
rect 39080 13444 39086 13456
rect 39316 13444 39344 13472
rect 39080 13416 39344 13444
rect 39080 13404 39086 13416
rect 38749 13379 38807 13385
rect 38749 13345 38761 13379
rect 38795 13345 38807 13379
rect 40770 13376 40776 13388
rect 38749 13339 38807 13345
rect 38948 13348 40776 13376
rect 37921 13311 37979 13317
rect 37921 13277 37933 13311
rect 37967 13308 37979 13311
rect 38948 13308 38976 13348
rect 40770 13336 40776 13348
rect 40828 13336 40834 13388
rect 37967 13280 38976 13308
rect 37967 13277 37979 13280
rect 37921 13271 37979 13277
rect 39022 13268 39028 13320
rect 39080 13308 39086 13320
rect 39209 13311 39267 13317
rect 39209 13308 39221 13311
rect 39080 13280 39221 13308
rect 39080 13268 39086 13280
rect 39209 13277 39221 13280
rect 39255 13277 39267 13311
rect 39209 13271 39267 13277
rect 37700 13212 37872 13240
rect 38473 13243 38531 13249
rect 37700 13200 37706 13212
rect 38473 13209 38485 13243
rect 38519 13240 38531 13243
rect 38519 13212 38976 13240
rect 38519 13209 38531 13212
rect 38473 13203 38531 13209
rect 38565 13175 38623 13181
rect 38565 13172 38577 13175
rect 35912 13144 38577 13172
rect 35805 13135 35863 13141
rect 38565 13141 38577 13144
rect 38611 13172 38623 13175
rect 38838 13172 38844 13184
rect 38611 13144 38844 13172
rect 38611 13141 38623 13144
rect 38565 13135 38623 13141
rect 38838 13132 38844 13144
rect 38896 13132 38902 13184
rect 38948 13172 38976 13212
rect 39482 13200 39488 13252
rect 39540 13200 39546 13252
rect 39758 13200 39764 13252
rect 39816 13200 39822 13252
rect 40218 13200 40224 13252
rect 40276 13200 40282 13252
rect 40880 13240 40908 13484
rect 41322 13472 41328 13524
rect 41380 13472 41386 13524
rect 40954 13404 40960 13456
rect 41012 13444 41018 13456
rect 41601 13447 41659 13453
rect 41601 13444 41613 13447
rect 41012 13416 41613 13444
rect 41012 13404 41018 13416
rect 41601 13413 41613 13416
rect 41647 13444 41659 13447
rect 42337 13447 42395 13453
rect 42337 13444 42349 13447
rect 41647 13416 42349 13444
rect 41647 13413 41659 13416
rect 41601 13407 41659 13413
rect 42337 13413 42349 13416
rect 42383 13444 42395 13447
rect 43070 13444 43076 13456
rect 42383 13416 43076 13444
rect 42383 13413 42395 13416
rect 42337 13407 42395 13413
rect 43070 13404 43076 13416
rect 43128 13444 43134 13456
rect 43441 13447 43499 13453
rect 43441 13444 43453 13447
rect 43128 13416 43453 13444
rect 43128 13404 43134 13416
rect 43441 13413 43453 13416
rect 43487 13413 43499 13447
rect 43441 13407 43499 13413
rect 45005 13243 45063 13249
rect 45005 13240 45017 13243
rect 40880 13212 42012 13240
rect 39206 13172 39212 13184
rect 38948 13144 39212 13172
rect 39206 13132 39212 13144
rect 39264 13132 39270 13184
rect 39776 13172 39804 13200
rect 41984 13184 42012 13212
rect 43824 13212 45017 13240
rect 40957 13175 41015 13181
rect 40957 13172 40969 13175
rect 39776 13144 40969 13172
rect 40957 13141 40969 13144
rect 41003 13141 41015 13175
rect 40957 13135 41015 13141
rect 41966 13132 41972 13184
rect 42024 13172 42030 13184
rect 42705 13175 42763 13181
rect 42705 13172 42717 13175
rect 42024 13144 42717 13172
rect 42024 13132 42030 13144
rect 42705 13141 42717 13144
rect 42751 13172 42763 13175
rect 43346 13172 43352 13184
rect 42751 13144 43352 13172
rect 42751 13141 42763 13144
rect 42705 13135 42763 13141
rect 43346 13132 43352 13144
rect 43404 13172 43410 13184
rect 43824 13181 43852 13212
rect 45005 13209 45017 13212
rect 45051 13209 45063 13243
rect 45005 13203 45063 13209
rect 43809 13175 43867 13181
rect 43809 13172 43821 13175
rect 43404 13144 43821 13172
rect 43404 13132 43410 13144
rect 43809 13141 43821 13144
rect 43855 13141 43867 13175
rect 43809 13135 43867 13141
rect 44542 13132 44548 13184
rect 44600 13132 44606 13184
rect 460 13082 45540 13104
rect 460 13030 6070 13082
rect 6122 13030 6134 13082
rect 6186 13030 6198 13082
rect 6250 13030 6262 13082
rect 6314 13030 6326 13082
rect 6378 13030 11070 13082
rect 11122 13030 11134 13082
rect 11186 13030 11198 13082
rect 11250 13030 11262 13082
rect 11314 13030 11326 13082
rect 11378 13030 16070 13082
rect 16122 13030 16134 13082
rect 16186 13030 16198 13082
rect 16250 13030 16262 13082
rect 16314 13030 16326 13082
rect 16378 13030 21070 13082
rect 21122 13030 21134 13082
rect 21186 13030 21198 13082
rect 21250 13030 21262 13082
rect 21314 13030 21326 13082
rect 21378 13030 26070 13082
rect 26122 13030 26134 13082
rect 26186 13030 26198 13082
rect 26250 13030 26262 13082
rect 26314 13030 26326 13082
rect 26378 13030 31070 13082
rect 31122 13030 31134 13082
rect 31186 13030 31198 13082
rect 31250 13030 31262 13082
rect 31314 13030 31326 13082
rect 31378 13030 36070 13082
rect 36122 13030 36134 13082
rect 36186 13030 36198 13082
rect 36250 13030 36262 13082
rect 36314 13030 36326 13082
rect 36378 13030 41070 13082
rect 41122 13030 41134 13082
rect 41186 13030 41198 13082
rect 41250 13030 41262 13082
rect 41314 13030 41326 13082
rect 41378 13030 45540 13082
rect 460 13008 45540 13030
rect 5902 12968 5908 12980
rect 4724 12940 5908 12968
rect 4724 12841 4752 12940
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7282 12968 7288 12980
rect 6972 12940 7288 12968
rect 6972 12928 6978 12940
rect 7282 12928 7288 12940
rect 7340 12968 7346 12980
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 7340 12940 7481 12968
rect 7340 12928 7346 12940
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 7469 12931 7527 12937
rect 8478 12928 8484 12980
rect 8536 12928 8542 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10008 12940 11376 12968
rect 10008 12928 10014 12940
rect 4801 12903 4859 12909
rect 4801 12869 4813 12903
rect 4847 12900 4859 12903
rect 5997 12903 6055 12909
rect 5997 12900 6009 12903
rect 4847 12872 6009 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 5997 12869 6009 12872
rect 6043 12869 6055 12903
rect 5997 12863 6055 12869
rect 6638 12860 6644 12912
rect 6696 12860 6702 12912
rect 8496 12900 8524 12928
rect 9033 12903 9091 12909
rect 9033 12900 9045 12903
rect 8496 12872 9045 12900
rect 9033 12869 9045 12872
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 10965 12903 11023 12909
rect 10965 12869 10977 12903
rect 11011 12869 11023 12903
rect 11348 12900 11376 12940
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11480 12940 12173 12968
rect 11480 12928 11486 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12894 12968 12900 12980
rect 12299 12940 12900 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12894 12928 12900 12940
rect 12952 12968 12958 12980
rect 13541 12971 13599 12977
rect 13541 12968 13553 12971
rect 12952 12940 13553 12968
rect 12952 12928 12958 12940
rect 13541 12937 13553 12940
rect 13587 12937 13599 12971
rect 13541 12931 13599 12937
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13906 12968 13912 12980
rect 13679 12940 13912 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17862 12977 17868 12980
rect 17819 12971 17868 12977
rect 17819 12968 17831 12971
rect 17000 12940 17831 12968
rect 17000 12928 17006 12940
rect 17819 12937 17831 12940
rect 17865 12937 17868 12971
rect 17819 12931 17868 12937
rect 17862 12928 17868 12931
rect 17920 12928 17926 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 19150 12968 19156 12980
rect 18012 12940 19156 12968
rect 18012 12928 18018 12940
rect 11701 12903 11759 12909
rect 11348 12872 11652 12900
rect 10965 12863 11023 12869
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 5169 12838 5227 12841
rect 5169 12835 5396 12838
rect 5169 12801 5181 12835
rect 5215 12832 5396 12835
rect 5626 12832 5632 12844
rect 5215 12810 5632 12832
rect 5215 12801 5227 12810
rect 5368 12804 5632 12810
rect 5169 12795 5227 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8757 12835 8815 12841
rect 8757 12832 8769 12835
rect 8260 12804 8769 12832
rect 8260 12792 8266 12804
rect 8757 12801 8769 12804
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 10134 12792 10140 12844
rect 10192 12792 10198 12844
rect 10980 12832 11008 12863
rect 11330 12832 11336 12844
rect 10980 12804 11336 12832
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 4908 12764 4936 12792
rect 5074 12764 5080 12776
rect 4908 12736 5080 12764
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5258 12724 5264 12776
rect 5316 12724 5322 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5736 12696 5764 12727
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6638 12764 6644 12776
rect 6052 12736 6644 12764
rect 6052 12724 6058 12736
rect 6638 12724 6644 12736
rect 6696 12764 6702 12776
rect 8018 12764 8024 12776
rect 6696 12736 8024 12764
rect 6696 12724 6702 12736
rect 8018 12724 8024 12736
rect 8076 12764 8082 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8076 12736 8585 12764
rect 8076 12724 8082 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9766 12764 9772 12776
rect 9180 12736 9772 12764
rect 9180 12724 9186 12736
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 9824 12736 10517 12764
rect 9824 12724 9830 12736
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10551 12736 11529 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 5684 12668 5764 12696
rect 8297 12699 8355 12705
rect 5684 12656 5690 12668
rect 8297 12665 8309 12699
rect 8343 12696 8355 12699
rect 10965 12699 11023 12705
rect 8343 12668 8892 12696
rect 8343 12665 8355 12668
rect 8297 12659 8355 12665
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5445 12631 5503 12637
rect 5445 12628 5457 12631
rect 5224 12600 5457 12628
rect 5224 12588 5230 12600
rect 5445 12597 5457 12600
rect 5491 12597 5503 12631
rect 5445 12591 5503 12597
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8202 12628 8208 12640
rect 7892 12600 8208 12628
rect 7892 12588 7898 12600
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8864 12628 8892 12668
rect 10965 12665 10977 12699
rect 11011 12665 11023 12699
rect 11624 12696 11652 12872
rect 11701 12869 11713 12903
rect 11747 12900 11759 12903
rect 13170 12900 13176 12912
rect 11747 12872 13176 12900
rect 11747 12869 11759 12872
rect 11701 12863 11759 12869
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13354 12860 13360 12912
rect 13412 12860 13418 12912
rect 13725 12903 13783 12909
rect 13725 12869 13737 12903
rect 13771 12900 13783 12903
rect 14016 12900 14044 12928
rect 13771 12872 14044 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 18156 12900 18184 12940
rect 19150 12928 19156 12940
rect 19208 12968 19214 12980
rect 19208 12940 19473 12968
rect 19208 12928 19214 12940
rect 14424 12872 14766 12900
rect 17434 12872 18184 12900
rect 14424 12860 14430 12872
rect 18230 12860 18236 12912
rect 18288 12860 18294 12912
rect 19445 12872 19473 12940
rect 19610 12928 19616 12980
rect 19668 12968 19674 12980
rect 20257 12971 20315 12977
rect 20257 12968 20269 12971
rect 19668 12940 20269 12968
rect 19668 12928 19674 12940
rect 20257 12937 20269 12940
rect 20303 12937 20315 12971
rect 20257 12931 20315 12937
rect 20717 12971 20775 12977
rect 20717 12937 20729 12971
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 20809 12971 20867 12977
rect 20809 12937 20821 12971
rect 20855 12968 20867 12971
rect 20898 12968 20904 12980
rect 20855 12940 20904 12968
rect 20855 12937 20867 12940
rect 20809 12931 20867 12937
rect 20349 12903 20407 12909
rect 20349 12869 20361 12903
rect 20395 12900 20407 12903
rect 20438 12900 20444 12912
rect 20395 12872 20444 12900
rect 20395 12869 20407 12872
rect 20349 12863 20407 12869
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 20565 12903 20623 12909
rect 20565 12869 20577 12903
rect 20611 12900 20623 12903
rect 20611 12872 20694 12900
rect 20611 12869 20623 12872
rect 20565 12863 20623 12869
rect 12618 12792 12624 12844
rect 12676 12792 12682 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12768 12804 12817 12832
rect 12768 12792 12774 12804
rect 12805 12801 12817 12804
rect 12851 12832 12863 12835
rect 13262 12832 13268 12844
rect 12851 12804 13268 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 16482 12832 16488 12844
rect 16040 12804 16488 12832
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 12636 12764 12664 12792
rect 12986 12764 12992 12776
rect 12636 12736 12992 12764
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 13998 12724 14004 12776
rect 14056 12724 14062 12776
rect 14274 12764 14280 12776
rect 14108 12736 14280 12764
rect 14108 12696 14136 12736
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 16040 12773 16068 12804
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 17586 12792 17592 12844
rect 17644 12832 17650 12844
rect 17957 12835 18015 12841
rect 17957 12832 17969 12835
rect 17644 12804 17969 12832
rect 17644 12792 17650 12804
rect 17957 12801 17969 12804
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 19978 12832 19984 12844
rect 19852 12804 19984 12832
rect 19852 12792 19858 12804
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20162 12832 20168 12844
rect 20119 12804 20168 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 16025 12767 16083 12773
rect 16025 12764 16037 12767
rect 15528 12736 16037 12764
rect 15528 12724 15534 12736
rect 16025 12733 16037 12736
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 16393 12767 16451 12773
rect 16393 12733 16405 12767
rect 16439 12764 16451 12767
rect 17770 12764 17776 12776
rect 16439 12736 17776 12764
rect 16439 12733 16451 12736
rect 16393 12727 16451 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18874 12764 18880 12776
rect 18288 12736 18880 12764
rect 18288 12724 18294 12736
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19242 12764 19248 12776
rect 19024 12736 19248 12764
rect 19024 12724 19030 12736
rect 19242 12724 19248 12736
rect 19300 12724 19306 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 11624 12668 14136 12696
rect 10965 12659 11023 12665
rect 9398 12628 9404 12640
rect 8864 12600 9404 12628
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10980 12628 11008 12659
rect 19610 12656 19616 12708
rect 19668 12696 19674 12708
rect 19904 12696 19932 12727
rect 19668 12668 19932 12696
rect 19668 12656 19674 12668
rect 20666 12640 20694 12872
rect 20732 12832 20760 12931
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 22925 12971 22983 12977
rect 22925 12968 22937 12971
rect 22796 12940 22937 12968
rect 22796 12928 22802 12940
rect 22925 12937 22937 12940
rect 22971 12937 22983 12971
rect 22925 12931 22983 12937
rect 23109 12971 23167 12977
rect 23109 12937 23121 12971
rect 23155 12968 23167 12971
rect 24489 12971 24547 12977
rect 24489 12968 24501 12971
rect 23155 12940 24501 12968
rect 23155 12937 23167 12940
rect 23109 12931 23167 12937
rect 24489 12937 24501 12940
rect 24535 12937 24547 12971
rect 24489 12931 24547 12937
rect 24578 12928 24584 12980
rect 24636 12928 24642 12980
rect 25685 12971 25743 12977
rect 25685 12937 25697 12971
rect 25731 12968 25743 12971
rect 25731 12940 27200 12968
rect 25731 12937 25743 12940
rect 25685 12931 25743 12937
rect 24596 12900 24624 12928
rect 24946 12900 24952 12912
rect 23584 12872 24624 12900
rect 24688 12872 24952 12900
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20732 12804 21005 12832
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22520 12804 22586 12832
rect 22520 12792 22526 12804
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23584 12841 23612 12872
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 23348 12804 23489 12832
rect 23348 12792 23354 12804
rect 23477 12801 23489 12804
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12801 23627 12835
rect 23569 12795 23627 12801
rect 23750 12792 23756 12844
rect 23808 12792 23814 12844
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12832 23903 12835
rect 24305 12835 24363 12841
rect 23891 12804 24261 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 21177 12767 21235 12773
rect 21177 12764 21189 12767
rect 20864 12736 21189 12764
rect 20864 12724 20870 12736
rect 21177 12733 21189 12736
rect 21223 12733 21235 12767
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 21177 12727 21235 12733
rect 21284 12736 21465 12764
rect 20898 12656 20904 12708
rect 20956 12696 20962 12708
rect 21284 12696 21312 12736
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 21542 12724 21548 12776
rect 21600 12764 21606 12776
rect 22480 12764 22508 12792
rect 21600 12736 22508 12764
rect 21600 12724 21606 12736
rect 20956 12668 21312 12696
rect 20956 12656 20962 12668
rect 23198 12656 23204 12708
rect 23256 12656 23262 12708
rect 23290 12656 23296 12708
rect 23348 12696 23354 12708
rect 23860 12696 23888 12795
rect 24026 12724 24032 12776
rect 24084 12764 24090 12776
rect 24121 12767 24179 12773
rect 24121 12764 24133 12767
rect 24084 12736 24133 12764
rect 24084 12724 24090 12736
rect 24121 12733 24133 12736
rect 24167 12733 24179 12767
rect 24233 12764 24261 12804
rect 24305 12801 24317 12835
rect 24351 12832 24363 12835
rect 24394 12832 24400 12844
rect 24351 12804 24400 12832
rect 24351 12801 24363 12804
rect 24305 12795 24363 12801
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 24688 12832 24716 12872
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 25314 12900 25320 12912
rect 25056 12872 25320 12900
rect 25056 12832 25084 12872
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 25406 12860 25412 12912
rect 25464 12900 25470 12912
rect 25777 12903 25835 12909
rect 25777 12900 25789 12903
rect 25464 12872 25789 12900
rect 25464 12860 25470 12872
rect 25777 12869 25789 12872
rect 25823 12869 25835 12903
rect 26329 12903 26387 12909
rect 26329 12900 26341 12903
rect 25777 12863 25835 12869
rect 25976 12872 26341 12900
rect 25976 12832 26004 12872
rect 26329 12869 26341 12872
rect 26375 12900 26387 12903
rect 26418 12900 26424 12912
rect 26375 12872 26424 12900
rect 26375 12869 26387 12872
rect 26329 12863 26387 12869
rect 26418 12860 26424 12872
rect 26476 12860 26482 12912
rect 26545 12903 26603 12909
rect 26545 12869 26557 12903
rect 26591 12900 26603 12903
rect 26786 12900 26792 12912
rect 26591 12872 26792 12900
rect 26591 12869 26603 12872
rect 26545 12863 26603 12869
rect 26786 12860 26792 12872
rect 26844 12860 26850 12912
rect 27172 12844 27200 12940
rect 27614 12928 27620 12980
rect 27672 12968 27678 12980
rect 27801 12971 27859 12977
rect 27801 12968 27813 12971
rect 27672 12940 27813 12968
rect 27672 12928 27678 12940
rect 27801 12937 27813 12940
rect 27847 12937 27859 12971
rect 27801 12931 27859 12937
rect 28261 12971 28319 12977
rect 28261 12937 28273 12971
rect 28307 12968 28319 12971
rect 28350 12968 28356 12980
rect 28307 12940 28356 12968
rect 28307 12937 28319 12940
rect 28261 12931 28319 12937
rect 28350 12928 28356 12940
rect 28408 12928 28414 12980
rect 28997 12971 29055 12977
rect 28997 12937 29009 12971
rect 29043 12968 29055 12971
rect 29362 12968 29368 12980
rect 29043 12940 29368 12968
rect 29043 12937 29055 12940
rect 28997 12931 29055 12937
rect 29362 12928 29368 12940
rect 29420 12928 29426 12980
rect 29546 12928 29552 12980
rect 29604 12928 29610 12980
rect 29822 12928 29828 12980
rect 29880 12968 29886 12980
rect 29880 12940 30236 12968
rect 29880 12928 29886 12940
rect 28074 12900 28080 12912
rect 27264 12872 28080 12900
rect 24504 12804 24716 12832
rect 24857 12815 24915 12821
rect 24504 12764 24532 12804
rect 24857 12781 24869 12815
rect 24903 12812 24915 12815
rect 24964 12812 25084 12832
rect 24903 12804 25084 12812
rect 25332 12804 26004 12832
rect 24903 12784 24992 12804
rect 24903 12781 24915 12784
rect 24857 12775 24915 12781
rect 24766 12767 24824 12773
rect 24766 12764 24778 12767
rect 24233 12736 24532 12764
rect 24688 12736 24778 12764
rect 24121 12727 24179 12733
rect 23348 12668 23888 12696
rect 23348 12656 23354 12668
rect 9732 12600 11008 12628
rect 9732 12588 9738 12600
rect 11790 12588 11796 12640
rect 11848 12588 11854 12640
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12628 13967 12631
rect 14090 12628 14096 12640
rect 13955 12600 14096 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15344 12600 15761 12628
rect 15344 12588 15350 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 19702 12588 19708 12640
rect 19760 12588 19766 12640
rect 19886 12588 19892 12640
rect 19944 12628 19950 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19944 12600 20085 12628
rect 19944 12588 19950 12600
rect 20073 12597 20085 12600
rect 20119 12628 20131 12631
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20119 12600 20545 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 20533 12597 20545 12600
rect 20579 12597 20591 12631
rect 20533 12591 20591 12597
rect 20622 12588 20628 12640
rect 20680 12628 20694 12640
rect 23216 12628 23244 12656
rect 20680 12600 23244 12628
rect 20680 12588 20686 12600
rect 24118 12588 24124 12640
rect 24176 12588 24182 12640
rect 24578 12588 24584 12640
rect 24636 12588 24642 12640
rect 24688 12628 24716 12736
rect 24766 12733 24778 12736
rect 24812 12733 24824 12767
rect 24766 12727 24824 12733
rect 25133 12767 25191 12773
rect 25133 12733 25145 12767
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 24854 12656 24860 12708
rect 24912 12696 24918 12708
rect 25148 12696 25176 12727
rect 25222 12724 25228 12776
rect 25280 12764 25286 12776
rect 25332 12764 25360 12804
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 27264 12841 27292 12872
rect 28074 12860 28080 12872
rect 28132 12860 28138 12912
rect 28169 12903 28227 12909
rect 28169 12869 28181 12903
rect 28215 12900 28227 12903
rect 28215 12872 28663 12900
rect 28215 12869 28227 12872
rect 28169 12863 28227 12869
rect 28635 12844 28663 12872
rect 28902 12860 28908 12912
rect 28960 12900 28966 12912
rect 29181 12903 29239 12909
rect 28960 12872 29132 12900
rect 28960 12860 28966 12872
rect 27249 12835 27307 12841
rect 27249 12801 27261 12835
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27341 12835 27399 12841
rect 27341 12801 27353 12835
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27522 12832 27528 12844
rect 27479 12804 27528 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 25280 12736 25360 12764
rect 25280 12724 25286 12736
rect 25682 12724 25688 12776
rect 25740 12764 25746 12776
rect 25961 12767 26019 12773
rect 25961 12764 25973 12767
rect 25740 12736 25973 12764
rect 25740 12724 25746 12736
rect 25961 12733 25973 12736
rect 26007 12764 26019 12767
rect 26510 12764 26516 12776
rect 26007 12736 26516 12764
rect 26007 12733 26019 12736
rect 25961 12727 26019 12733
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 26602 12724 26608 12776
rect 26660 12764 26666 12776
rect 27356 12764 27384 12795
rect 27522 12792 27528 12804
rect 27580 12792 27586 12844
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12832 27675 12835
rect 28534 12832 28540 12844
rect 27663 12804 28540 12832
rect 27663 12801 27675 12804
rect 27617 12795 27675 12801
rect 27632 12764 27660 12795
rect 28534 12792 28540 12804
rect 28592 12792 28598 12844
rect 28626 12792 28632 12844
rect 28684 12832 28690 12844
rect 29104 12841 29132 12872
rect 29181 12869 29193 12903
rect 29227 12900 29239 12903
rect 29564 12900 29592 12928
rect 30006 12900 30012 12912
rect 29227 12872 29592 12900
rect 29656 12872 30012 12900
rect 29227 12869 29239 12872
rect 29181 12863 29239 12869
rect 28813 12835 28871 12841
rect 28684 12804 28729 12832
rect 28684 12792 28690 12804
rect 28813 12801 28825 12835
rect 28859 12801 28871 12835
rect 28813 12795 28871 12801
rect 29089 12835 29147 12841
rect 29089 12801 29101 12835
rect 29135 12832 29147 12835
rect 29656 12832 29684 12872
rect 30006 12860 30012 12872
rect 30064 12900 30070 12912
rect 30101 12903 30159 12909
rect 30101 12900 30113 12903
rect 30064 12872 30113 12900
rect 30064 12860 30070 12872
rect 30101 12869 30113 12872
rect 30147 12869 30159 12903
rect 30208 12900 30236 12940
rect 30466 12928 30472 12980
rect 30524 12968 30530 12980
rect 30742 12968 30748 12980
rect 30524 12940 30748 12968
rect 30524 12928 30530 12940
rect 30742 12928 30748 12940
rect 30800 12928 30806 12980
rect 31113 12971 31171 12977
rect 31113 12937 31125 12971
rect 31159 12968 31171 12971
rect 31159 12940 31800 12968
rect 31159 12937 31171 12940
rect 31113 12931 31171 12937
rect 30653 12903 30711 12909
rect 30653 12900 30665 12903
rect 30208 12872 30665 12900
rect 30101 12863 30159 12869
rect 30653 12869 30665 12872
rect 30699 12869 30711 12903
rect 31478 12900 31484 12912
rect 30653 12863 30711 12869
rect 31312 12872 31484 12900
rect 29135 12804 29684 12832
rect 29135 12801 29147 12804
rect 29089 12795 29147 12801
rect 26660 12736 27384 12764
rect 27448 12736 27660 12764
rect 26660 12724 26666 12736
rect 26418 12696 26424 12708
rect 24912 12668 25176 12696
rect 25240 12668 26424 12696
rect 24912 12656 24918 12668
rect 25240 12628 25268 12668
rect 26418 12656 26424 12668
rect 26476 12656 26482 12708
rect 26528 12668 26832 12696
rect 24688 12600 25268 12628
rect 25317 12631 25375 12637
rect 25317 12597 25329 12631
rect 25363 12628 25375 12631
rect 25774 12628 25780 12640
rect 25363 12600 25780 12628
rect 25363 12597 25375 12600
rect 25317 12591 25375 12597
rect 25774 12588 25780 12600
rect 25832 12588 25838 12640
rect 26528 12637 26556 12668
rect 26804 12640 26832 12668
rect 26970 12656 26976 12708
rect 27028 12656 27034 12708
rect 27448 12696 27476 12736
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28353 12767 28411 12773
rect 28353 12764 28365 12767
rect 27856 12736 28365 12764
rect 27856 12724 27862 12736
rect 28353 12733 28365 12736
rect 28399 12733 28411 12767
rect 28828 12764 28856 12795
rect 29730 12792 29736 12844
rect 29788 12792 29794 12844
rect 30282 12792 30288 12844
rect 30340 12792 30346 12844
rect 31312 12841 31340 12872
rect 31478 12860 31484 12872
rect 31536 12860 31542 12912
rect 31772 12909 31800 12940
rect 33244 12940 34928 12968
rect 33244 12912 33272 12940
rect 31757 12903 31815 12909
rect 31757 12869 31769 12903
rect 31803 12869 31815 12903
rect 31757 12863 31815 12869
rect 32214 12860 32220 12912
rect 32272 12860 32278 12912
rect 33226 12860 33232 12912
rect 33284 12860 33290 12912
rect 33502 12860 33508 12912
rect 33560 12900 33566 12912
rect 33597 12903 33655 12909
rect 33597 12900 33609 12903
rect 33560 12872 33609 12900
rect 33560 12860 33566 12872
rect 33597 12869 33609 12872
rect 33643 12869 33655 12903
rect 33597 12863 33655 12869
rect 33870 12860 33876 12912
rect 33928 12900 33934 12912
rect 34900 12900 34928 12940
rect 34974 12928 34980 12980
rect 35032 12968 35038 12980
rect 35069 12971 35127 12977
rect 35069 12968 35081 12971
rect 35032 12940 35081 12968
rect 35032 12928 35038 12940
rect 35069 12937 35081 12940
rect 35115 12937 35127 12971
rect 35069 12931 35127 12937
rect 35253 12971 35311 12977
rect 35253 12937 35265 12971
rect 35299 12968 35311 12971
rect 35802 12968 35808 12980
rect 35299 12940 35808 12968
rect 35299 12937 35311 12940
rect 35253 12931 35311 12937
rect 35802 12928 35808 12940
rect 35860 12928 35866 12980
rect 35897 12971 35955 12977
rect 35897 12937 35909 12971
rect 35943 12968 35955 12971
rect 36538 12968 36544 12980
rect 35943 12940 36544 12968
rect 35943 12937 35955 12940
rect 35897 12931 35955 12937
rect 36538 12928 36544 12940
rect 36596 12928 36602 12980
rect 37274 12928 37280 12980
rect 37332 12968 37338 12980
rect 37642 12968 37648 12980
rect 37332 12940 37648 12968
rect 37332 12928 37338 12940
rect 37642 12928 37648 12940
rect 37700 12968 37706 12980
rect 38381 12971 38439 12977
rect 38381 12968 38393 12971
rect 37700 12940 38393 12968
rect 37700 12928 37706 12940
rect 38381 12937 38393 12940
rect 38427 12937 38439 12971
rect 38381 12931 38439 12937
rect 38930 12928 38936 12980
rect 38988 12928 38994 12980
rect 39482 12928 39488 12980
rect 39540 12968 39546 12980
rect 40037 12971 40095 12977
rect 40037 12968 40049 12971
rect 39540 12940 40049 12968
rect 39540 12928 39546 12940
rect 40037 12937 40049 12940
rect 40083 12937 40095 12971
rect 40037 12931 40095 12937
rect 40126 12928 40132 12980
rect 40184 12928 40190 12980
rect 42426 12928 42432 12980
rect 42484 12928 42490 12980
rect 35342 12900 35348 12912
rect 33928 12872 34086 12900
rect 34900 12872 35348 12900
rect 33928 12860 33934 12872
rect 35342 12860 35348 12872
rect 35400 12900 35406 12912
rect 35989 12903 36047 12909
rect 35989 12900 36001 12903
rect 35400 12872 36001 12900
rect 35400 12860 35406 12872
rect 35989 12869 36001 12872
rect 36035 12869 36047 12903
rect 38194 12900 38200 12912
rect 38134 12872 38200 12900
rect 35989 12863 36047 12869
rect 38194 12860 38200 12872
rect 38252 12860 38258 12912
rect 30377 12835 30435 12841
rect 30377 12801 30389 12835
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 31297 12835 31355 12841
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 28353 12727 28411 12733
rect 28736 12736 28856 12764
rect 27080 12668 27476 12696
rect 26513 12631 26571 12637
rect 26513 12597 26525 12631
rect 26559 12597 26571 12631
rect 26513 12591 26571 12597
rect 26694 12588 26700 12640
rect 26752 12588 26758 12640
rect 26786 12588 26792 12640
rect 26844 12628 26850 12640
rect 27080 12628 27108 12668
rect 26844 12600 27108 12628
rect 26844 12588 26850 12600
rect 27430 12588 27436 12640
rect 27488 12628 27494 12640
rect 27890 12628 27896 12640
rect 27488 12600 27896 12628
rect 27488 12588 27494 12600
rect 27890 12588 27896 12600
rect 27948 12628 27954 12640
rect 28736 12628 28764 12736
rect 29270 12724 29276 12776
rect 29328 12764 29334 12776
rect 29549 12767 29607 12773
rect 29549 12764 29561 12767
rect 29328 12736 29561 12764
rect 29328 12724 29334 12736
rect 29549 12733 29561 12736
rect 29595 12733 29607 12767
rect 29549 12727 29607 12733
rect 30098 12724 30104 12776
rect 30156 12724 30162 12776
rect 30392 12764 30420 12795
rect 33318 12792 33324 12844
rect 33376 12792 33382 12844
rect 35437 12835 35495 12841
rect 35437 12801 35449 12835
rect 35483 12832 35495 12835
rect 35483 12804 35572 12832
rect 35483 12801 35495 12804
rect 35437 12795 35495 12801
rect 30392 12736 30788 12764
rect 28810 12656 28816 12708
rect 28868 12696 28874 12708
rect 30116 12696 30144 12724
rect 28868 12668 30144 12696
rect 28868 12656 28874 12668
rect 30760 12640 30788 12736
rect 30834 12724 30840 12776
rect 30892 12764 30898 12776
rect 31478 12764 31484 12776
rect 30892 12736 31484 12764
rect 30892 12724 30898 12736
rect 31478 12724 31484 12736
rect 31536 12764 31542 12776
rect 33336 12764 33364 12792
rect 31536 12736 33364 12764
rect 31536 12724 31542 12736
rect 35544 12705 35572 12804
rect 35618 12792 35624 12844
rect 35676 12832 35682 12844
rect 36633 12835 36691 12841
rect 36633 12832 36645 12835
rect 35676 12804 36645 12832
rect 35676 12792 35682 12804
rect 36633 12801 36645 12804
rect 36679 12801 36691 12835
rect 38948 12832 38976 12928
rect 39209 12903 39267 12909
rect 39209 12869 39221 12903
rect 39255 12869 39267 12903
rect 39209 12863 39267 12869
rect 39025 12835 39083 12841
rect 39025 12832 39037 12835
rect 38948 12804 39037 12832
rect 36633 12795 36691 12801
rect 39025 12801 39037 12804
rect 39071 12801 39083 12835
rect 39224 12832 39252 12863
rect 39666 12860 39672 12912
rect 39724 12860 39730 12912
rect 39758 12860 39764 12912
rect 39816 12860 39822 12912
rect 39850 12860 39856 12912
rect 39908 12900 39914 12912
rect 39945 12903 40003 12909
rect 39945 12900 39957 12903
rect 39908 12872 39957 12900
rect 39908 12860 39914 12872
rect 39945 12869 39957 12872
rect 39991 12869 40003 12903
rect 39945 12863 40003 12869
rect 40034 12832 40040 12844
rect 39224 12804 40040 12832
rect 39025 12795 39083 12801
rect 40034 12792 40040 12804
rect 40092 12792 40098 12844
rect 40144 12832 40172 12928
rect 40221 12835 40279 12841
rect 40221 12832 40233 12835
rect 40144 12804 40233 12832
rect 40221 12801 40233 12804
rect 40267 12801 40279 12835
rect 40221 12795 40279 12801
rect 35986 12724 35992 12776
rect 36044 12764 36050 12776
rect 36081 12767 36139 12773
rect 36081 12764 36093 12767
rect 36044 12736 36093 12764
rect 36044 12724 36050 12736
rect 36081 12733 36093 12736
rect 36127 12733 36139 12767
rect 36081 12727 36139 12733
rect 36906 12724 36912 12776
rect 36964 12724 36970 12776
rect 39574 12764 39580 12776
rect 38856 12736 39580 12764
rect 38856 12705 38884 12736
rect 39574 12724 39580 12736
rect 39632 12724 39638 12776
rect 40954 12764 40960 12776
rect 40512 12736 40960 12764
rect 35529 12699 35587 12705
rect 35529 12665 35541 12699
rect 35575 12665 35587 12699
rect 35529 12659 35587 12665
rect 38841 12699 38899 12705
rect 38841 12665 38853 12699
rect 38887 12665 38899 12699
rect 38841 12659 38899 12665
rect 39206 12656 39212 12708
rect 39264 12656 39270 12708
rect 40512 12640 40540 12736
rect 40954 12724 40960 12736
rect 41012 12764 41018 12776
rect 41969 12767 42027 12773
rect 41969 12764 41981 12767
rect 41012 12736 41981 12764
rect 41012 12724 41018 12736
rect 41969 12733 41981 12736
rect 42015 12764 42027 12767
rect 42705 12767 42763 12773
rect 42705 12764 42717 12767
rect 42015 12736 42717 12764
rect 42015 12733 42027 12736
rect 41969 12727 42027 12733
rect 42705 12733 42717 12736
rect 42751 12764 42763 12767
rect 42886 12764 42892 12776
rect 42751 12736 42892 12764
rect 42751 12733 42763 12736
rect 42705 12727 42763 12733
rect 42886 12724 42892 12736
rect 42944 12764 42950 12776
rect 43441 12767 43499 12773
rect 43441 12764 43453 12767
rect 42944 12736 43453 12764
rect 42944 12724 42950 12736
rect 43441 12733 43453 12736
rect 43487 12764 43499 12767
rect 43809 12767 43867 12773
rect 43809 12764 43821 12767
rect 43487 12736 43821 12764
rect 43487 12733 43499 12736
rect 43441 12727 43499 12733
rect 43809 12733 43821 12736
rect 43855 12764 43867 12767
rect 44177 12767 44235 12773
rect 44177 12764 44189 12767
rect 43855 12736 44189 12764
rect 43855 12733 43867 12736
rect 43809 12727 43867 12733
rect 44177 12733 44189 12736
rect 44223 12764 44235 12767
rect 44545 12767 44603 12773
rect 44545 12764 44557 12767
rect 44223 12736 44557 12764
rect 44223 12733 44235 12736
rect 44177 12727 44235 12733
rect 44545 12733 44557 12736
rect 44591 12733 44603 12767
rect 44545 12727 44603 12733
rect 40589 12699 40647 12705
rect 40589 12665 40601 12699
rect 40635 12696 40647 12699
rect 41233 12699 41291 12705
rect 41233 12696 41245 12699
rect 40635 12668 41245 12696
rect 40635 12665 40647 12668
rect 40589 12659 40647 12665
rect 41233 12665 41245 12668
rect 41279 12696 41291 12699
rect 41279 12668 41414 12696
rect 41279 12665 41291 12668
rect 41233 12659 41291 12665
rect 27948 12600 28764 12628
rect 27948 12588 27954 12600
rect 29086 12588 29092 12640
rect 29144 12628 29150 12640
rect 29822 12628 29828 12640
rect 29144 12600 29828 12628
rect 29144 12588 29150 12600
rect 29822 12588 29828 12600
rect 29880 12588 29886 12640
rect 29914 12588 29920 12640
rect 29972 12588 29978 12640
rect 30101 12631 30159 12637
rect 30101 12597 30113 12631
rect 30147 12628 30159 12631
rect 30374 12628 30380 12640
rect 30147 12600 30380 12628
rect 30147 12597 30159 12600
rect 30101 12591 30159 12597
rect 30374 12588 30380 12600
rect 30432 12588 30438 12640
rect 30742 12588 30748 12640
rect 30800 12588 30806 12640
rect 32306 12588 32312 12640
rect 32364 12628 32370 12640
rect 32766 12628 32772 12640
rect 32364 12600 32772 12628
rect 32364 12588 32370 12600
rect 32766 12588 32772 12600
rect 32824 12588 32830 12640
rect 32858 12588 32864 12640
rect 32916 12628 32922 12640
rect 33042 12628 33048 12640
rect 32916 12600 33048 12628
rect 32916 12588 32922 12600
rect 33042 12588 33048 12600
rect 33100 12628 33106 12640
rect 33229 12631 33287 12637
rect 33229 12628 33241 12631
rect 33100 12600 33241 12628
rect 33100 12588 33106 12600
rect 33229 12597 33241 12600
rect 33275 12597 33287 12631
rect 33229 12591 33287 12597
rect 33410 12588 33416 12640
rect 33468 12628 33474 12640
rect 34146 12628 34152 12640
rect 33468 12600 34152 12628
rect 33468 12588 33474 12600
rect 34146 12588 34152 12600
rect 34204 12588 34210 12640
rect 38749 12631 38807 12637
rect 38749 12597 38761 12631
rect 38795 12628 38807 12631
rect 39022 12628 39028 12640
rect 38795 12600 39028 12628
rect 38795 12597 38807 12600
rect 38749 12591 38807 12597
rect 39022 12588 39028 12600
rect 39080 12628 39086 12640
rect 40494 12628 40500 12640
rect 39080 12600 40500 12628
rect 39080 12588 39086 12600
rect 40494 12588 40500 12600
rect 40552 12628 40558 12640
rect 40865 12631 40923 12637
rect 40865 12628 40877 12631
rect 40552 12600 40877 12628
rect 40552 12588 40558 12600
rect 40865 12597 40877 12600
rect 40911 12597 40923 12631
rect 41386 12628 41414 12668
rect 41966 12628 41972 12640
rect 41386 12600 41972 12628
rect 40865 12591 40923 12597
rect 41966 12588 41972 12600
rect 42024 12628 42030 12640
rect 42610 12628 42616 12640
rect 42024 12600 42616 12628
rect 42024 12588 42030 12600
rect 42610 12588 42616 12600
rect 42668 12628 42674 12640
rect 43073 12631 43131 12637
rect 43073 12628 43085 12631
rect 42668 12600 43085 12628
rect 42668 12588 42674 12600
rect 43073 12597 43085 12600
rect 43119 12597 43131 12631
rect 43073 12591 43131 12597
rect 44358 12588 44364 12640
rect 44416 12628 44422 12640
rect 44913 12631 44971 12637
rect 44913 12628 44925 12631
rect 44416 12600 44925 12628
rect 44416 12588 44422 12600
rect 44913 12597 44925 12600
rect 44959 12597 44971 12631
rect 44913 12591 44971 12597
rect 460 12538 45540 12560
rect 460 12486 3570 12538
rect 3622 12486 3634 12538
rect 3686 12486 3698 12538
rect 3750 12486 3762 12538
rect 3814 12486 3826 12538
rect 3878 12486 8570 12538
rect 8622 12486 8634 12538
rect 8686 12486 8698 12538
rect 8750 12486 8762 12538
rect 8814 12486 8826 12538
rect 8878 12486 13570 12538
rect 13622 12486 13634 12538
rect 13686 12486 13698 12538
rect 13750 12486 13762 12538
rect 13814 12486 13826 12538
rect 13878 12486 18570 12538
rect 18622 12486 18634 12538
rect 18686 12486 18698 12538
rect 18750 12486 18762 12538
rect 18814 12486 18826 12538
rect 18878 12486 23570 12538
rect 23622 12486 23634 12538
rect 23686 12486 23698 12538
rect 23750 12486 23762 12538
rect 23814 12486 23826 12538
rect 23878 12486 28570 12538
rect 28622 12486 28634 12538
rect 28686 12486 28698 12538
rect 28750 12486 28762 12538
rect 28814 12486 28826 12538
rect 28878 12486 33570 12538
rect 33622 12486 33634 12538
rect 33686 12486 33698 12538
rect 33750 12486 33762 12538
rect 33814 12486 33826 12538
rect 33878 12486 38570 12538
rect 38622 12486 38634 12538
rect 38686 12486 38698 12538
rect 38750 12486 38762 12538
rect 38814 12486 38826 12538
rect 38878 12486 43570 12538
rect 43622 12486 43634 12538
rect 43686 12486 43698 12538
rect 43750 12486 43762 12538
rect 43814 12486 43826 12538
rect 43878 12486 45540 12538
rect 460 12464 45540 12486
rect 5169 12427 5227 12433
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5258 12424 5264 12436
rect 5215 12396 5264 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5368 12396 6592 12424
rect 5074 12316 5080 12368
rect 5132 12356 5138 12368
rect 5368 12356 5396 12396
rect 5132 12328 5396 12356
rect 6564 12356 6592 12396
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 7064 12396 7113 12424
rect 7064 12384 7070 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7101 12387 7159 12393
rect 8018 12384 8024 12436
rect 8076 12384 8082 12436
rect 8772 12396 10916 12424
rect 8772 12365 8800 12396
rect 7561 12359 7619 12365
rect 7561 12356 7573 12359
rect 6564 12328 7573 12356
rect 5132 12316 5138 12328
rect 7561 12325 7573 12328
rect 7607 12325 7619 12359
rect 7561 12319 7619 12325
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12325 8815 12359
rect 10888 12356 10916 12396
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 11698 12424 11704 12436
rect 11655 12396 11704 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12434 12384 12440 12436
rect 12492 12384 12498 12436
rect 15381 12427 15439 12433
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 17126 12424 17132 12436
rect 15427 12396 17132 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 17126 12384 17132 12396
rect 17184 12424 17190 12436
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 17184 12396 17693 12424
rect 17184 12384 17190 12396
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 17770 12384 17776 12436
rect 17828 12384 17834 12436
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 18874 12424 18880 12436
rect 17920 12396 18880 12424
rect 17920 12384 17926 12396
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19337 12427 19395 12433
rect 19337 12424 19349 12427
rect 19116 12396 19349 12424
rect 19116 12384 19122 12396
rect 19337 12393 19349 12396
rect 19383 12393 19395 12427
rect 19337 12387 19395 12393
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 19886 12424 19892 12436
rect 19843 12396 19892 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 19886 12384 19892 12396
rect 19944 12424 19950 12436
rect 20346 12424 20352 12436
rect 19944 12396 20352 12424
rect 19944 12384 19950 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 23382 12424 23388 12436
rect 22980 12396 23388 12424
rect 22980 12384 22986 12396
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23569 12427 23627 12433
rect 23569 12393 23581 12427
rect 23615 12424 23627 12427
rect 23934 12424 23940 12436
rect 23615 12396 23940 12424
rect 23615 12393 23627 12396
rect 23569 12387 23627 12393
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 24210 12384 24216 12436
rect 24268 12384 24274 12436
rect 24486 12384 24492 12436
rect 24544 12424 24550 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24544 12396 24593 12424
rect 24544 12384 24550 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 10888 12328 13032 12356
rect 8757 12319 8815 12325
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5534 12288 5540 12300
rect 5307 12260 5540 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 7098 12288 7104 12300
rect 6052 12260 7104 12288
rect 6052 12248 6058 12260
rect 6656 12206 6684 12260
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 13004 12232 13032 12328
rect 16850 12316 16856 12368
rect 16908 12356 16914 12368
rect 16908 12328 17372 12356
rect 16908 12316 16914 12328
rect 14734 12248 14740 12300
rect 14792 12248 14798 12300
rect 17344 12288 17372 12328
rect 17402 12316 17408 12368
rect 17460 12316 17466 12368
rect 17788 12356 17816 12384
rect 19245 12359 19303 12365
rect 19245 12356 19257 12359
rect 17788 12328 19257 12356
rect 19245 12325 19257 12328
rect 19291 12325 19303 12359
rect 19518 12356 19524 12368
rect 19245 12319 19303 12325
rect 19352 12328 19524 12356
rect 17678 12288 17684 12300
rect 17344 12260 17684 12288
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 18414 12288 18420 12300
rect 18156 12260 18420 12288
rect 7374 12180 7380 12232
rect 7432 12180 7438 12232
rect 9582 12220 9588 12232
rect 9416 12192 9588 12220
rect 4801 12155 4859 12161
rect 4801 12121 4813 12155
rect 4847 12121 4859 12155
rect 4801 12115 4859 12121
rect 4816 12084 4844 12115
rect 4982 12112 4988 12164
rect 5040 12112 5046 12164
rect 5074 12112 5080 12164
rect 5132 12112 5138 12164
rect 5537 12155 5595 12161
rect 5537 12121 5549 12155
rect 5583 12121 5595 12155
rect 5537 12115 5595 12121
rect 5092 12084 5120 12112
rect 4816 12056 5120 12084
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 5552 12084 5580 12115
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7101 12155 7159 12161
rect 7101 12152 7113 12155
rect 6880 12124 7113 12152
rect 6880 12112 6886 12124
rect 7101 12121 7113 12124
rect 7147 12121 7159 12155
rect 7101 12115 7159 12121
rect 5316 12056 5580 12084
rect 5316 12044 5322 12056
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9416 12093 9444 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 11790 12180 11796 12232
rect 11848 12180 11854 12232
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 13044 12192 13737 12220
rect 13044 12180 13050 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 14001 12223 14059 12229
rect 14001 12189 14013 12223
rect 14047 12220 14059 12223
rect 14274 12220 14280 12232
rect 14047 12192 14280 12220
rect 14047 12189 14059 12192
rect 14001 12183 14059 12189
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12220 14979 12223
rect 15286 12220 15292 12232
rect 14967 12192 15292 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 15729 12223 15787 12229
rect 15729 12220 15741 12223
rect 15620 12192 15741 12220
rect 15620 12180 15626 12192
rect 15729 12189 15741 12192
rect 15775 12189 15787 12223
rect 15729 12183 15787 12189
rect 17862 12180 17868 12232
rect 17920 12180 17926 12232
rect 18156 12229 18184 12260
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 18764 12260 19288 12288
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18322 12180 18328 12232
rect 18380 12220 18386 12232
rect 18764 12229 18792 12260
rect 19260 12232 19288 12260
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18380 12192 18613 12220
rect 18380 12180 18386 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18749 12223 18807 12229
rect 18749 12189 18761 12223
rect 18795 12189 18807 12223
rect 18749 12183 18807 12189
rect 18966 12180 18972 12232
rect 19024 12180 19030 12232
rect 19058 12180 19064 12232
rect 19116 12229 19122 12232
rect 19116 12183 19124 12229
rect 19116 12180 19122 12183
rect 19242 12180 19248 12232
rect 19300 12180 19306 12232
rect 19352 12229 19380 12328
rect 19518 12316 19524 12328
rect 19576 12316 19582 12368
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20027 12328 21220 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20346 12288 20352 12300
rect 20272 12260 20352 12288
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19567 12192 20050 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10192 12124 10350 12152
rect 10192 12112 10198 12124
rect 15010 12112 15016 12164
rect 15068 12152 15074 12164
rect 15488 12152 15516 12180
rect 15068 12124 15516 12152
rect 15068 12112 15074 12124
rect 18046 12112 18052 12164
rect 18104 12112 18110 12164
rect 18248 12152 18276 12180
rect 18877 12155 18935 12161
rect 18877 12152 18889 12155
rect 18248 12124 18736 12152
rect 18708 12096 18736 12124
rect 18800 12124 18889 12152
rect 9401 12087 9459 12093
rect 9401 12084 9413 12087
rect 9088 12056 9413 12084
rect 9088 12044 9094 12056
rect 9401 12053 9413 12056
rect 9447 12053 9459 12087
rect 9401 12047 9459 12053
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 12216 12056 12265 12084
rect 12216 12044 12222 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 12676 12056 13185 12084
rect 12676 12044 12682 12056
rect 13173 12053 13185 12056
rect 13219 12053 13231 12087
rect 13173 12047 13231 12053
rect 13814 12044 13820 12096
rect 13872 12044 13878 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17954 12084 17960 12096
rect 16632 12056 17960 12084
rect 16632 12044 16638 12056
rect 17954 12044 17960 12056
rect 18012 12084 18018 12096
rect 18230 12084 18236 12096
rect 18012 12056 18236 12084
rect 18012 12044 18018 12056
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 18414 12044 18420 12096
rect 18472 12044 18478 12096
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 18800 12084 18828 12124
rect 18877 12121 18889 12124
rect 18923 12121 18935 12155
rect 18877 12115 18935 12121
rect 19150 12112 19156 12164
rect 19208 12152 19214 12164
rect 19536 12152 19564 12183
rect 19208 12124 19564 12152
rect 19208 12112 19214 12124
rect 19610 12112 19616 12164
rect 19668 12112 19674 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 19813 12155 19871 12161
rect 19813 12152 19825 12155
rect 19760 12124 19825 12152
rect 19760 12112 19766 12124
rect 19813 12121 19825 12124
rect 19859 12121 19871 12155
rect 20022 12152 20050 12192
rect 20162 12180 20168 12232
rect 20220 12180 20226 12232
rect 20272 12229 20300 12260
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 21192 12288 21220 12328
rect 22830 12316 22836 12368
rect 22888 12316 22894 12368
rect 23753 12359 23811 12365
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 24228 12356 24256 12384
rect 23799 12328 24256 12356
rect 24596 12356 24624 12387
rect 24670 12384 24676 12436
rect 24728 12424 24734 12436
rect 25041 12427 25099 12433
rect 25041 12424 25053 12427
rect 24728 12396 25053 12424
rect 24728 12384 24734 12396
rect 25041 12393 25053 12396
rect 25087 12393 25099 12427
rect 25041 12387 25099 12393
rect 25590 12384 25596 12436
rect 25648 12424 25654 12436
rect 26881 12427 26939 12433
rect 25648 12396 26464 12424
rect 25648 12384 25654 12396
rect 26436 12356 26464 12396
rect 26881 12393 26893 12427
rect 26927 12424 26939 12427
rect 27154 12424 27160 12436
rect 26927 12396 27160 12424
rect 26927 12393 26939 12396
rect 26881 12387 26939 12393
rect 27154 12384 27160 12396
rect 27212 12424 27218 12436
rect 28902 12424 28908 12436
rect 27212 12396 28908 12424
rect 27212 12384 27218 12396
rect 28902 12384 28908 12396
rect 28960 12384 28966 12436
rect 29104 12396 30620 12424
rect 28353 12359 28411 12365
rect 28353 12356 28365 12359
rect 24596 12328 25084 12356
rect 26436 12328 28365 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 25056 12300 25084 12328
rect 28353 12325 28365 12328
rect 28399 12356 28411 12359
rect 29104 12356 29132 12396
rect 28399 12328 29132 12356
rect 30592 12356 30620 12396
rect 30650 12384 30656 12436
rect 30708 12424 30714 12436
rect 30834 12424 30840 12436
rect 30708 12396 30840 12424
rect 30708 12384 30714 12396
rect 30834 12384 30840 12396
rect 30892 12424 30898 12436
rect 30929 12427 30987 12433
rect 30929 12424 30941 12427
rect 30892 12396 30941 12424
rect 30892 12384 30898 12396
rect 30929 12393 30941 12396
rect 30975 12393 30987 12427
rect 30929 12387 30987 12393
rect 33229 12427 33287 12433
rect 33229 12393 33241 12427
rect 33275 12424 33287 12427
rect 33318 12424 33324 12436
rect 33275 12396 33324 12424
rect 33275 12393 33287 12396
rect 33229 12387 33287 12393
rect 33318 12384 33324 12396
rect 33376 12384 33382 12436
rect 33870 12384 33876 12436
rect 33928 12384 33934 12436
rect 34054 12384 34060 12436
rect 34112 12384 34118 12436
rect 34364 12396 34560 12424
rect 34364 12356 34392 12396
rect 30592 12328 34392 12356
rect 28399 12325 28411 12328
rect 28353 12319 28411 12325
rect 34422 12316 34428 12368
rect 34480 12316 34486 12368
rect 34532 12356 34560 12396
rect 34606 12384 34612 12436
rect 34664 12424 34670 12436
rect 34885 12427 34943 12433
rect 34885 12424 34897 12427
rect 34664 12396 34897 12424
rect 34664 12384 34670 12396
rect 34885 12393 34897 12396
rect 34931 12393 34943 12427
rect 35710 12424 35716 12436
rect 34885 12387 34943 12393
rect 35452 12396 35716 12424
rect 34790 12356 34796 12368
rect 34532 12328 34796 12356
rect 34790 12316 34796 12328
rect 34848 12316 34854 12368
rect 21192 12260 22692 12288
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20487 12192 20545 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 20533 12189 20545 12192
rect 20579 12220 20591 12223
rect 20622 12220 20628 12232
rect 20579 12192 20628 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 20732 12152 20760 12183
rect 20806 12180 20812 12232
rect 20864 12220 20870 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 20864 12192 21097 12220
rect 20864 12180 20870 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 20022 12124 20760 12152
rect 21361 12155 21419 12161
rect 19813 12115 19871 12121
rect 21361 12121 21373 12155
rect 21407 12152 21419 12155
rect 21450 12152 21456 12164
rect 21407 12124 21456 12152
rect 21407 12121 21419 12124
rect 21361 12115 21419 12121
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 19426 12084 19432 12096
rect 18800 12056 19432 12084
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20622 12044 20628 12096
rect 20680 12044 20686 12096
rect 22664 12084 22692 12260
rect 22756 12260 24256 12288
rect 22756 12232 22784 12260
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 22830 12180 22836 12232
rect 22888 12180 22894 12232
rect 23106 12180 23112 12232
rect 23164 12180 23170 12232
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 24026 12220 24032 12232
rect 23440 12192 24032 12220
rect 23440 12180 23446 12192
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 24228 12229 24256 12260
rect 24762 12248 24768 12300
rect 24820 12248 24826 12300
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 25409 12291 25467 12297
rect 25409 12257 25421 12291
rect 25455 12288 25467 12291
rect 25958 12288 25964 12300
rect 25455 12260 25964 12288
rect 25455 12257 25467 12260
rect 25409 12251 25467 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 26878 12288 26884 12300
rect 26528 12260 26884 12288
rect 26528 12232 26556 12260
rect 26878 12248 26884 12260
rect 26936 12288 26942 12300
rect 27706 12288 27712 12300
rect 26936 12260 27712 12288
rect 26936 12248 26942 12260
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 27890 12248 27896 12300
rect 27948 12248 27954 12300
rect 28442 12248 28448 12300
rect 28500 12248 28506 12300
rect 28997 12291 29055 12297
rect 28997 12257 29009 12291
rect 29043 12288 29055 12291
rect 29638 12288 29644 12300
rect 29043 12260 29644 12288
rect 29043 12257 29055 12260
rect 28997 12251 29055 12257
rect 29638 12248 29644 12260
rect 29696 12248 29702 12300
rect 29822 12248 29828 12300
rect 29880 12288 29886 12300
rect 32585 12291 32643 12297
rect 29880 12260 30512 12288
rect 29880 12248 29886 12260
rect 24121 12223 24179 12229
rect 24121 12189 24133 12223
rect 24167 12189 24179 12223
rect 24121 12183 24179 12189
rect 24213 12223 24271 12229
rect 24213 12189 24225 12223
rect 24259 12189 24271 12223
rect 24213 12183 24271 12189
rect 22848 12152 22876 12180
rect 24136 12152 24164 12183
rect 24302 12180 24308 12232
rect 24360 12180 24366 12232
rect 24394 12180 24400 12232
rect 24452 12180 24458 12232
rect 24489 12223 24547 12229
rect 24489 12189 24501 12223
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 22848 12124 24164 12152
rect 24320 12152 24348 12180
rect 24504 12152 24532 12183
rect 25130 12180 25136 12232
rect 25188 12180 25194 12232
rect 26510 12180 26516 12232
rect 26568 12180 26574 12232
rect 26694 12180 26700 12232
rect 26752 12220 26758 12232
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 26752 12192 27169 12220
rect 26752 12180 26758 12192
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 28460 12220 28488 12248
rect 27157 12183 27215 12189
rect 27586 12192 28488 12220
rect 24320 12124 24532 12152
rect 25148 12152 25176 12180
rect 25682 12152 25688 12164
rect 25148 12124 25688 12152
rect 25682 12112 25688 12124
rect 25740 12112 25746 12164
rect 27586 12152 27614 12192
rect 26912 12124 27614 12152
rect 27709 12155 27767 12161
rect 26912 12084 26940 12124
rect 27709 12121 27721 12155
rect 27755 12152 27767 12155
rect 27890 12152 27896 12164
rect 27755 12124 27896 12152
rect 27755 12121 27767 12124
rect 27709 12115 27767 12121
rect 27890 12112 27896 12124
rect 27948 12112 27954 12164
rect 29273 12155 29331 12161
rect 29273 12121 29285 12155
rect 29319 12121 29331 12155
rect 30484 12152 30512 12260
rect 31128 12260 31708 12288
rect 30650 12180 30656 12232
rect 30708 12220 30714 12232
rect 31128 12229 31156 12260
rect 31680 12232 31708 12260
rect 32585 12257 32597 12291
rect 32631 12288 32643 12291
rect 32858 12288 32864 12300
rect 32631 12260 32864 12288
rect 32631 12257 32643 12260
rect 32585 12251 32643 12257
rect 32858 12248 32864 12260
rect 32916 12248 32922 12300
rect 33318 12248 33324 12300
rect 33376 12248 33382 12300
rect 34440 12288 34468 12316
rect 34609 12291 34667 12297
rect 34609 12288 34621 12291
rect 34440 12260 34621 12288
rect 34609 12257 34621 12260
rect 34655 12257 34667 12291
rect 34609 12251 34667 12257
rect 31113 12223 31171 12229
rect 31113 12220 31125 12223
rect 30708 12192 31125 12220
rect 30708 12180 30714 12192
rect 31113 12189 31125 12192
rect 31159 12189 31171 12223
rect 31113 12183 31171 12189
rect 31570 12180 31576 12232
rect 31628 12180 31634 12232
rect 31662 12180 31668 12232
rect 31720 12180 31726 12232
rect 32490 12180 32496 12232
rect 32548 12180 32554 12232
rect 33689 12223 33747 12229
rect 33689 12189 33701 12223
rect 33735 12189 33747 12223
rect 33689 12183 33747 12189
rect 33704 12152 33732 12183
rect 33870 12180 33876 12232
rect 33928 12180 33934 12232
rect 34425 12223 34483 12229
rect 34425 12189 34437 12223
rect 34471 12220 34483 12223
rect 34900 12220 34928 12387
rect 34974 12248 34980 12300
rect 35032 12248 35038 12300
rect 35452 12297 35480 12396
rect 35710 12384 35716 12396
rect 35768 12384 35774 12436
rect 37090 12384 37096 12436
rect 37148 12384 37154 12436
rect 37182 12384 37188 12436
rect 37240 12384 37246 12436
rect 43438 12384 43444 12436
rect 43496 12424 43502 12436
rect 43533 12427 43591 12433
rect 43533 12424 43545 12427
rect 43496 12396 43545 12424
rect 43496 12384 43502 12396
rect 43533 12393 43545 12396
rect 43579 12393 43591 12427
rect 43533 12387 43591 12393
rect 37108 12356 37136 12384
rect 37108 12328 37872 12356
rect 35437 12291 35495 12297
rect 35437 12257 35449 12291
rect 35483 12257 35495 12291
rect 35437 12251 35495 12257
rect 35713 12291 35771 12297
rect 35713 12257 35725 12291
rect 35759 12288 35771 12291
rect 36446 12288 36452 12300
rect 35759 12260 36452 12288
rect 35759 12257 35771 12260
rect 35713 12251 35771 12257
rect 36446 12248 36452 12260
rect 36504 12248 36510 12300
rect 37734 12248 37740 12300
rect 37792 12248 37798 12300
rect 34471 12192 34928 12220
rect 34471 12189 34483 12192
rect 34425 12183 34483 12189
rect 35158 12180 35164 12232
rect 35216 12180 35222 12232
rect 37550 12220 37556 12232
rect 36846 12192 37556 12220
rect 37550 12180 37556 12192
rect 37608 12180 37614 12232
rect 37642 12180 37648 12232
rect 37700 12180 37706 12232
rect 37844 12220 37872 12328
rect 37936 12328 38700 12356
rect 37936 12297 37964 12328
rect 37921 12291 37979 12297
rect 37921 12257 37933 12291
rect 37967 12257 37979 12291
rect 37921 12251 37979 12257
rect 38562 12248 38568 12300
rect 38620 12248 38626 12300
rect 38672 12297 38700 12328
rect 38746 12316 38752 12368
rect 38804 12356 38810 12368
rect 41417 12359 41475 12365
rect 41417 12356 41429 12359
rect 38804 12328 41429 12356
rect 38804 12316 38810 12328
rect 41417 12325 41429 12328
rect 41463 12356 41475 12359
rect 42242 12356 42248 12368
rect 41463 12328 42248 12356
rect 41463 12325 41475 12328
rect 41417 12319 41475 12325
rect 42242 12316 42248 12328
rect 42300 12356 42306 12368
rect 44542 12356 44548 12368
rect 42300 12328 44548 12356
rect 42300 12316 42306 12328
rect 44542 12316 44548 12328
rect 44600 12316 44606 12368
rect 38657 12291 38715 12297
rect 38657 12257 38669 12291
rect 38703 12288 38715 12291
rect 39298 12288 39304 12300
rect 38703 12260 39304 12288
rect 38703 12257 38715 12260
rect 38657 12251 38715 12257
rect 39298 12248 39304 12260
rect 39356 12288 39362 12300
rect 39761 12291 39819 12297
rect 39761 12288 39773 12291
rect 39356 12260 39773 12288
rect 39356 12248 39362 12260
rect 39761 12257 39773 12260
rect 39807 12257 39819 12291
rect 39761 12251 39819 12257
rect 40313 12291 40371 12297
rect 40313 12257 40325 12291
rect 40359 12288 40371 12291
rect 40957 12291 41015 12297
rect 40957 12288 40969 12291
rect 40359 12260 40969 12288
rect 40359 12257 40371 12260
rect 40313 12251 40371 12257
rect 40957 12257 40969 12260
rect 41003 12288 41015 12291
rect 41598 12288 41604 12300
rect 41003 12260 41604 12288
rect 41003 12257 41015 12260
rect 40957 12251 41015 12257
rect 41598 12248 41604 12260
rect 41656 12248 41662 12300
rect 38286 12220 38292 12232
rect 37844 12192 38292 12220
rect 38286 12180 38292 12192
rect 38344 12220 38350 12232
rect 38473 12223 38531 12229
rect 38473 12220 38485 12223
rect 38344 12192 38485 12220
rect 38344 12180 38350 12192
rect 38473 12189 38485 12192
rect 38519 12189 38531 12223
rect 38473 12183 38531 12189
rect 39114 12180 39120 12232
rect 39172 12180 39178 12232
rect 41414 12220 41420 12232
rect 41386 12180 41420 12220
rect 41472 12180 41478 12232
rect 30484 12138 31984 12152
rect 30498 12124 31984 12138
rect 29273 12115 29331 12121
rect 22664 12056 26940 12084
rect 26970 12044 26976 12096
rect 27028 12044 27034 12096
rect 27341 12087 27399 12093
rect 27341 12053 27353 12087
rect 27387 12084 27399 12087
rect 27614 12084 27620 12096
rect 27387 12056 27620 12084
rect 27387 12053 27399 12056
rect 27341 12047 27399 12053
rect 27614 12044 27620 12056
rect 27672 12044 27678 12096
rect 27801 12087 27859 12093
rect 27801 12053 27813 12087
rect 27847 12084 27859 12087
rect 28074 12084 28080 12096
rect 27847 12056 28080 12084
rect 27847 12053 27859 12056
rect 27801 12047 27859 12053
rect 28074 12044 28080 12056
rect 28132 12044 28138 12096
rect 29288 12084 29316 12115
rect 30006 12084 30012 12096
rect 29288 12056 30012 12084
rect 30006 12044 30012 12056
rect 30064 12044 30070 12096
rect 30190 12044 30196 12096
rect 30248 12084 30254 12096
rect 31956 12093 31984 12124
rect 32876 12124 33732 12152
rect 33888 12152 33916 12180
rect 34885 12155 34943 12161
rect 33888 12124 34652 12152
rect 30745 12087 30803 12093
rect 30745 12084 30757 12087
rect 30248 12056 30757 12084
rect 30248 12044 30254 12056
rect 30745 12053 30757 12056
rect 30791 12053 30803 12087
rect 30745 12047 30803 12053
rect 31941 12087 31999 12093
rect 31941 12053 31953 12087
rect 31987 12084 31999 12087
rect 32306 12084 32312 12096
rect 31987 12056 32312 12084
rect 31987 12053 31999 12056
rect 31941 12047 31999 12053
rect 32306 12044 32312 12056
rect 32364 12044 32370 12096
rect 32876 12093 32904 12124
rect 32861 12087 32919 12093
rect 32861 12053 32873 12087
rect 32907 12053 32919 12087
rect 32861 12047 32919 12053
rect 33134 12044 33140 12096
rect 33192 12084 33198 12096
rect 33318 12084 33324 12096
rect 33192 12056 33324 12084
rect 33192 12044 33198 12056
rect 33318 12044 33324 12056
rect 33376 12044 33382 12096
rect 33502 12044 33508 12096
rect 33560 12044 33566 12096
rect 34238 12044 34244 12096
rect 34296 12084 34302 12096
rect 34517 12087 34575 12093
rect 34517 12084 34529 12087
rect 34296 12056 34529 12084
rect 34296 12044 34302 12056
rect 34517 12053 34529 12056
rect 34563 12053 34575 12087
rect 34624 12084 34652 12124
rect 34885 12121 34897 12155
rect 34931 12152 34943 12155
rect 34931 12124 36124 12152
rect 34931 12121 34943 12124
rect 34885 12115 34943 12121
rect 35345 12087 35403 12093
rect 35345 12084 35357 12087
rect 34624 12056 35357 12084
rect 34517 12047 34575 12053
rect 35345 12053 35357 12056
rect 35391 12053 35403 12087
rect 36096 12084 36124 12124
rect 37090 12112 37096 12164
rect 37148 12152 37154 12164
rect 37148 12124 38148 12152
rect 37148 12112 37154 12124
rect 36446 12084 36452 12096
rect 36096 12056 36452 12084
rect 35345 12047 35403 12053
rect 36446 12044 36452 12056
rect 36504 12044 36510 12096
rect 37274 12044 37280 12096
rect 37332 12044 37338 12096
rect 38120 12093 38148 12124
rect 38194 12112 38200 12164
rect 38252 12152 38258 12164
rect 39132 12152 39160 12180
rect 39577 12155 39635 12161
rect 38252 12124 39344 12152
rect 38252 12112 38258 12124
rect 38105 12087 38163 12093
rect 38105 12053 38117 12087
rect 38151 12053 38163 12087
rect 38105 12047 38163 12053
rect 39114 12044 39120 12096
rect 39172 12084 39178 12096
rect 39209 12087 39267 12093
rect 39209 12084 39221 12087
rect 39172 12056 39221 12084
rect 39172 12044 39178 12056
rect 39209 12053 39221 12056
rect 39255 12053 39267 12087
rect 39316 12084 39344 12124
rect 39577 12121 39589 12155
rect 39623 12152 39635 12155
rect 41386 12152 41414 12180
rect 39623 12124 41414 12152
rect 42521 12155 42579 12161
rect 39623 12121 39635 12124
rect 39577 12115 39635 12121
rect 42521 12121 42533 12155
rect 42567 12152 42579 12155
rect 43070 12152 43076 12164
rect 42567 12124 43076 12152
rect 42567 12121 42579 12124
rect 42521 12115 42579 12121
rect 43070 12112 43076 12124
rect 43128 12152 43134 12164
rect 43165 12155 43223 12161
rect 43165 12152 43177 12155
rect 43128 12124 43177 12152
rect 43128 12112 43134 12124
rect 43165 12121 43177 12124
rect 43211 12121 43223 12155
rect 43165 12115 43223 12121
rect 39669 12087 39727 12093
rect 39669 12084 39681 12087
rect 39316 12056 39681 12084
rect 39209 12047 39267 12053
rect 39669 12053 39681 12056
rect 39715 12084 39727 12087
rect 39942 12084 39948 12096
rect 39715 12056 39948 12084
rect 39715 12053 39727 12056
rect 39669 12047 39727 12053
rect 39942 12044 39948 12056
rect 40000 12044 40006 12096
rect 40494 12044 40500 12096
rect 40552 12084 40558 12096
rect 40681 12087 40739 12093
rect 40681 12084 40693 12087
rect 40552 12056 40693 12084
rect 40552 12044 40558 12056
rect 40681 12053 40693 12056
rect 40727 12084 40739 12087
rect 40954 12084 40960 12096
rect 40727 12056 40960 12084
rect 40727 12053 40739 12056
rect 40681 12047 40739 12053
rect 40954 12044 40960 12056
rect 41012 12044 41018 12096
rect 41782 12044 41788 12096
rect 41840 12084 41846 12096
rect 42061 12087 42119 12093
rect 42061 12084 42073 12087
rect 41840 12056 42073 12084
rect 41840 12044 41846 12056
rect 42061 12053 42073 12056
rect 42107 12084 42119 12087
rect 42610 12084 42616 12096
rect 42107 12056 42616 12084
rect 42107 12053 42119 12056
rect 42061 12047 42119 12053
rect 42610 12044 42616 12056
rect 42668 12084 42674 12096
rect 42797 12087 42855 12093
rect 42797 12084 42809 12087
rect 42668 12056 42809 12084
rect 42668 12044 42674 12056
rect 42797 12053 42809 12056
rect 42843 12084 42855 12087
rect 43901 12087 43959 12093
rect 43901 12084 43913 12087
rect 42843 12056 43913 12084
rect 42843 12053 42855 12056
rect 42797 12047 42855 12053
rect 43901 12053 43913 12056
rect 43947 12084 43959 12087
rect 44358 12084 44364 12096
rect 43947 12056 44364 12084
rect 43947 12053 43959 12056
rect 43901 12047 43959 12053
rect 44358 12044 44364 12056
rect 44416 12084 44422 12096
rect 44545 12087 44603 12093
rect 44545 12084 44557 12087
rect 44416 12056 44557 12084
rect 44416 12044 44422 12056
rect 44545 12053 44557 12056
rect 44591 12053 44603 12087
rect 44545 12047 44603 12053
rect 44634 12044 44640 12096
rect 44692 12084 44698 12096
rect 44913 12087 44971 12093
rect 44913 12084 44925 12087
rect 44692 12056 44925 12084
rect 44692 12044 44698 12056
rect 44913 12053 44925 12056
rect 44959 12053 44971 12087
rect 44913 12047 44971 12053
rect 460 11994 45540 12016
rect 460 11942 6070 11994
rect 6122 11942 6134 11994
rect 6186 11942 6198 11994
rect 6250 11942 6262 11994
rect 6314 11942 6326 11994
rect 6378 11942 11070 11994
rect 11122 11942 11134 11994
rect 11186 11942 11198 11994
rect 11250 11942 11262 11994
rect 11314 11942 11326 11994
rect 11378 11942 16070 11994
rect 16122 11942 16134 11994
rect 16186 11942 16198 11994
rect 16250 11942 16262 11994
rect 16314 11942 16326 11994
rect 16378 11942 21070 11994
rect 21122 11942 21134 11994
rect 21186 11942 21198 11994
rect 21250 11942 21262 11994
rect 21314 11942 21326 11994
rect 21378 11942 26070 11994
rect 26122 11942 26134 11994
rect 26186 11942 26198 11994
rect 26250 11942 26262 11994
rect 26314 11942 26326 11994
rect 26378 11942 31070 11994
rect 31122 11942 31134 11994
rect 31186 11942 31198 11994
rect 31250 11942 31262 11994
rect 31314 11942 31326 11994
rect 31378 11942 36070 11994
rect 36122 11942 36134 11994
rect 36186 11942 36198 11994
rect 36250 11942 36262 11994
rect 36314 11942 36326 11994
rect 36378 11942 41070 11994
rect 41122 11942 41134 11994
rect 41186 11942 41198 11994
rect 41250 11942 41262 11994
rect 41314 11942 41326 11994
rect 41378 11942 45540 11994
rect 460 11920 45540 11942
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4120 11852 4905 11880
rect 4120 11840 4126 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 4908 11540 4936 11843
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5902 11880 5908 11892
rect 5132 11852 5908 11880
rect 5132 11840 5138 11852
rect 5166 11772 5172 11824
rect 5224 11772 5230 11824
rect 5644 11812 5672 11852
rect 5902 11840 5908 11852
rect 5960 11880 5966 11892
rect 6822 11880 6828 11892
rect 5960 11852 6828 11880
rect 5960 11840 5966 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 8076 11852 8217 11880
rect 8076 11840 8082 11852
rect 8205 11849 8217 11852
rect 8251 11880 8263 11883
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8251 11852 8953 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 8941 11849 8953 11852
rect 8987 11849 8999 11883
rect 8941 11843 8999 11849
rect 9490 11840 9496 11892
rect 9548 11840 9554 11892
rect 9674 11840 9680 11892
rect 9732 11840 9738 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9824 11852 9965 11880
rect 9824 11840 9830 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10192 11852 11161 11880
rect 10192 11840 10198 11852
rect 11149 11849 11161 11852
rect 11195 11880 11207 11883
rect 12158 11880 12164 11892
rect 11195 11852 12164 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 13872 11852 14412 11880
rect 13872 11840 13878 11852
rect 5460 11784 5672 11812
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 5092 11676 5120 11707
rect 5266 11704 5272 11756
rect 5324 11704 5330 11756
rect 5359 11747 5417 11753
rect 5359 11713 5371 11747
rect 5405 11744 5417 11747
rect 5460 11744 5488 11784
rect 5718 11772 5724 11824
rect 5776 11812 5782 11824
rect 5997 11815 6055 11821
rect 5997 11812 6009 11815
rect 5776 11784 6009 11812
rect 5776 11772 5782 11784
rect 5997 11781 6009 11784
rect 6043 11781 6055 11815
rect 9692 11812 9720 11840
rect 9861 11815 9919 11821
rect 9861 11812 9873 11815
rect 9692 11784 9873 11812
rect 5997 11775 6055 11781
rect 9861 11781 9873 11784
rect 9907 11781 9919 11815
rect 12176 11812 12204 11840
rect 12986 11812 12992 11824
rect 12176 11784 12992 11812
rect 9861 11775 9919 11781
rect 12986 11772 12992 11784
rect 13044 11772 13050 11824
rect 14384 11821 14412 11852
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15804 11852 16037 11880
rect 15804 11840 15810 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16025 11843 16083 11849
rect 16393 11883 16451 11889
rect 16393 11849 16405 11883
rect 16439 11880 16451 11883
rect 16850 11880 16856 11892
rect 16439 11852 16856 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18414 11880 18420 11892
rect 17788 11852 18420 11880
rect 14369 11815 14427 11821
rect 14369 11781 14381 11815
rect 14415 11781 14427 11815
rect 14369 11775 14427 11781
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 17788 11821 17816 11852
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 19150 11840 19156 11892
rect 19208 11840 19214 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 20346 11880 20352 11892
rect 19475 11852 20352 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20898 11880 20904 11892
rect 20487 11852 20904 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21177 11883 21235 11889
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21450 11880 21456 11892
rect 21223 11852 21456 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 22186 11840 22192 11892
rect 22244 11840 22250 11892
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 22888 11852 23704 11880
rect 22888 11840 22894 11852
rect 16485 11815 16543 11821
rect 14516 11784 14858 11812
rect 14516 11772 14522 11784
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 17313 11815 17371 11821
rect 17313 11812 17325 11815
rect 16531 11784 17325 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 17313 11781 17325 11784
rect 17359 11781 17371 11815
rect 17313 11775 17371 11781
rect 17773 11815 17831 11821
rect 17773 11781 17785 11815
rect 17819 11781 17831 11815
rect 17773 11775 17831 11781
rect 18230 11772 18236 11824
rect 18288 11772 18294 11824
rect 19168 11812 19196 11840
rect 19613 11815 19671 11821
rect 19168 11784 19288 11812
rect 5405 11716 5488 11744
rect 5405 11713 5417 11716
rect 5359 11707 5417 11713
rect 5534 11702 5540 11754
rect 5592 11702 5598 11754
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 11882 11744 11888 11756
rect 11563 11716 11888 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 15804 11716 16711 11744
rect 15804 11704 15810 11716
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 5092 11648 5212 11676
rect 5184 11608 5212 11648
rect 5368 11648 5457 11676
rect 5368 11608 5396 11648
rect 5445 11645 5457 11648
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5718 11636 5724 11688
rect 5776 11636 5782 11688
rect 7374 11676 7380 11688
rect 5828 11648 7380 11676
rect 5184 11580 5396 11608
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5828 11608 5856 11648
rect 7374 11636 7380 11648
rect 7432 11676 7438 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7432 11648 7481 11676
rect 7432 11636 7438 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10226 11676 10232 11688
rect 10183 11648 10232 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 11606 11676 11612 11688
rect 11379 11648 11612 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 5592 11580 5856 11608
rect 9324 11580 10609 11608
rect 5592 11568 5598 11580
rect 7650 11540 7656 11552
rect 4908 11512 7656 11540
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 7892 11512 8585 11540
rect 7892 11500 7898 11512
rect 8573 11509 8585 11512
rect 8619 11540 8631 11543
rect 9030 11540 9036 11552
rect 8619 11512 9036 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9030 11500 9036 11512
rect 9088 11540 9094 11552
rect 9324 11549 9352 11580
rect 10597 11577 10609 11580
rect 10643 11608 10655 11611
rect 11514 11608 11520 11620
rect 10643 11580 11520 11608
rect 10643 11577 10655 11580
rect 10597 11571 10655 11577
rect 11514 11568 11520 11580
rect 11572 11608 11578 11620
rect 12069 11611 12127 11617
rect 12069 11608 12081 11611
rect 11572 11580 12081 11608
rect 11572 11568 11578 11580
rect 12069 11577 12081 11580
rect 12115 11608 12127 11611
rect 12268 11608 12296 11639
rect 12526 11636 12532 11688
rect 12584 11636 12590 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 14056 11648 14105 11676
rect 14056 11636 14062 11648
rect 14093 11645 14105 11648
rect 14139 11676 14151 11679
rect 15010 11676 15016 11688
rect 14139 11648 15016 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16574 11676 16580 11688
rect 15896 11648 16580 11676
rect 15896 11636 15902 11648
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16683 11676 16711 11716
rect 16942 11704 16948 11756
rect 17000 11704 17006 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11713 17279 11747
rect 19260 11750 19288 11784
rect 19613 11781 19625 11815
rect 19659 11812 19671 11815
rect 19702 11812 19708 11824
rect 19659 11784 19708 11812
rect 19659 11781 19671 11784
rect 19613 11775 19671 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 22204 11812 22232 11840
rect 19843 11781 19901 11787
rect 19843 11778 19855 11781
rect 19329 11753 19387 11759
rect 19828 11756 19855 11778
rect 19329 11750 19341 11753
rect 19260 11722 19341 11750
rect 19329 11719 19341 11722
rect 19375 11719 19387 11753
rect 19794 11744 19800 11756
rect 19329 11713 19387 11719
rect 19445 11716 19800 11744
rect 17221 11707 17279 11713
rect 17236 11676 17264 11707
rect 16683 11648 17264 11676
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 19245 11679 19303 11685
rect 19245 11645 19257 11679
rect 19291 11676 19303 11679
rect 19445 11676 19473 11716
rect 19794 11704 19800 11716
rect 19852 11747 19855 11756
rect 19889 11747 19901 11781
rect 20732 11784 22232 11812
rect 19852 11741 19901 11747
rect 19852 11704 19858 11741
rect 19978 11704 19984 11756
rect 20036 11744 20042 11756
rect 20073 11747 20131 11753
rect 20073 11744 20085 11747
rect 20036 11716 20085 11744
rect 20036 11704 20042 11716
rect 20073 11713 20085 11716
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 20257 11747 20315 11753
rect 20257 11744 20269 11747
rect 20220 11716 20269 11744
rect 20220 11704 20226 11716
rect 20257 11713 20269 11716
rect 20303 11744 20315 11747
rect 20530 11744 20536 11756
rect 20303 11716 20536 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20622 11704 20628 11756
rect 20680 11704 20686 11756
rect 20732 11753 20760 11784
rect 22462 11772 22468 11824
rect 22520 11772 22526 11824
rect 23676 11821 23704 11852
rect 28074 11840 28080 11892
rect 28132 11840 28138 11892
rect 28368 11852 29763 11880
rect 23661 11815 23719 11821
rect 23661 11781 23673 11815
rect 23707 11781 23719 11815
rect 23661 11775 23719 11781
rect 24397 11815 24455 11821
rect 24397 11781 24409 11815
rect 24443 11812 24455 11815
rect 24486 11812 24492 11824
rect 24443 11784 24492 11812
rect 24443 11781 24455 11784
rect 24397 11775 24455 11781
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 26510 11812 26516 11824
rect 25622 11784 26516 11812
rect 26510 11772 26516 11784
rect 26568 11772 26574 11824
rect 26602 11772 26608 11824
rect 26660 11772 26666 11824
rect 28368 11812 28396 11852
rect 28184 11784 28396 11812
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 19291 11648 19473 11676
rect 19291 11645 19303 11648
rect 19245 11639 19303 11645
rect 17512 11608 17540 11639
rect 19518 11636 19524 11688
rect 19576 11676 19582 11688
rect 21008 11676 21036 11707
rect 21358 11704 21364 11756
rect 21416 11704 21422 11756
rect 21634 11704 21640 11756
rect 21692 11704 21698 11756
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 25740 11716 26280 11744
rect 25740 11704 25746 11716
rect 21652 11676 21680 11704
rect 26252 11688 26280 11716
rect 27706 11704 27712 11756
rect 27764 11742 27770 11756
rect 28184 11744 28212 11784
rect 28442 11772 28448 11824
rect 28500 11772 28506 11824
rect 29735 11812 29763 11852
rect 30006 11840 30012 11892
rect 30064 11840 30070 11892
rect 30098 11840 30104 11892
rect 30156 11880 30162 11892
rect 30156 11852 30328 11880
rect 30156 11840 30162 11852
rect 29822 11812 29828 11824
rect 29670 11784 29828 11812
rect 29822 11772 29828 11784
rect 29880 11772 29886 11824
rect 30024 11812 30052 11840
rect 30300 11812 30328 11852
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 30558 11880 30564 11892
rect 30432 11852 30564 11880
rect 30432 11840 30438 11852
rect 30558 11840 30564 11852
rect 30616 11840 30622 11892
rect 30742 11840 30748 11892
rect 30800 11880 30806 11892
rect 31021 11883 31079 11889
rect 31021 11880 31033 11883
rect 30800 11852 31033 11880
rect 30800 11840 30806 11852
rect 31021 11849 31033 11852
rect 31067 11849 31079 11883
rect 31665 11883 31723 11889
rect 31665 11880 31677 11883
rect 31021 11843 31079 11849
rect 31312 11852 31677 11880
rect 30024 11784 30236 11812
rect 30300 11784 30788 11812
rect 30009 11747 30067 11753
rect 30009 11744 30021 11747
rect 27908 11742 28212 11744
rect 27764 11716 28212 11742
rect 29656 11716 30021 11744
rect 27764 11714 27936 11716
rect 27764 11704 27770 11714
rect 19576 11648 20208 11676
rect 21008 11648 21680 11676
rect 21729 11679 21787 11685
rect 19576 11636 19582 11648
rect 19886 11608 19892 11620
rect 12115 11580 12296 11608
rect 12115 11577 12127 11580
rect 12069 11571 12127 11577
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9088 11512 9321 11540
rect 9088 11500 9094 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 11698 11500 11704 11552
rect 11756 11500 11762 11552
rect 12268 11540 12296 11580
rect 17236 11580 17540 11608
rect 19812 11580 19892 11608
rect 17236 11552 17264 11580
rect 12618 11540 12624 11552
rect 12268 11512 12624 11540
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13964 11512 14013 11540
rect 13964 11500 13970 11512
rect 14001 11509 14013 11512
rect 14047 11509 14059 11543
rect 14001 11503 14059 11509
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15712 11512 15853 11540
rect 15712 11500 15718 11512
rect 15841 11509 15853 11512
rect 15887 11509 15899 11543
rect 15841 11503 15899 11509
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 15988 11512 17049 11540
rect 15988 11500 15994 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 17218 11500 17224 11552
rect 17276 11500 17282 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 19812 11549 19840 11580
rect 19886 11568 19892 11580
rect 19944 11568 19950 11620
rect 19978 11568 19984 11620
rect 20036 11568 20042 11620
rect 20180 11617 20208 11648
rect 21729 11645 21741 11679
rect 21775 11645 21787 11679
rect 21729 11639 21787 11645
rect 20165 11611 20223 11617
rect 20165 11577 20177 11611
rect 20211 11608 20223 11611
rect 20254 11608 20260 11620
rect 20211 11580 20260 11608
rect 20211 11577 20223 11580
rect 20165 11571 20223 11577
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 20714 11568 20720 11620
rect 20772 11608 20778 11620
rect 21744 11608 21772 11639
rect 22002 11636 22008 11688
rect 22060 11636 22066 11688
rect 24121 11679 24179 11685
rect 24121 11645 24133 11679
rect 24167 11676 24179 11679
rect 25130 11676 25136 11688
rect 24167 11648 25136 11676
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 25130 11636 25136 11648
rect 25188 11636 25194 11688
rect 25406 11636 25412 11688
rect 25464 11676 25470 11688
rect 25774 11676 25780 11688
rect 25464 11648 25780 11676
rect 25464 11636 25470 11648
rect 25774 11636 25780 11648
rect 25832 11676 25838 11688
rect 26145 11679 26203 11685
rect 26145 11676 26157 11679
rect 25832 11648 26157 11676
rect 25832 11636 25838 11648
rect 26145 11645 26157 11648
rect 26191 11645 26203 11679
rect 26145 11639 26203 11645
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 26329 11679 26387 11685
rect 26329 11676 26341 11679
rect 26292 11648 26341 11676
rect 26292 11636 26298 11648
rect 26329 11645 26341 11648
rect 26375 11676 26387 11679
rect 28074 11676 28080 11688
rect 26375 11648 28080 11676
rect 26375 11645 26387 11648
rect 26329 11639 26387 11645
rect 28074 11636 28080 11648
rect 28132 11676 28138 11688
rect 28169 11679 28227 11685
rect 28169 11676 28181 11679
rect 28132 11648 28181 11676
rect 28132 11636 28138 11648
rect 28169 11645 28181 11648
rect 28215 11676 28227 11679
rect 28215 11648 29592 11676
rect 28215 11645 28227 11648
rect 28169 11639 28227 11645
rect 29564 11620 29592 11648
rect 20772 11580 21772 11608
rect 23477 11611 23535 11617
rect 20772 11568 20778 11580
rect 23477 11577 23489 11611
rect 23523 11608 23535 11611
rect 23523 11580 24256 11608
rect 23523 11577 23535 11580
rect 23477 11571 23535 11577
rect 19797 11543 19855 11549
rect 19797 11540 19809 11543
rect 19024 11512 19809 11540
rect 19024 11500 19030 11512
rect 19797 11509 19809 11512
rect 19843 11509 19855 11543
rect 19797 11503 19855 11509
rect 20898 11500 20904 11552
rect 20956 11500 20962 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 23106 11540 23112 11552
rect 21600 11512 23112 11540
rect 21600 11500 21606 11512
rect 23106 11500 23112 11512
rect 23164 11540 23170 11552
rect 23753 11543 23811 11549
rect 23753 11540 23765 11543
rect 23164 11512 23765 11540
rect 23164 11500 23170 11512
rect 23753 11509 23765 11512
rect 23799 11540 23811 11543
rect 24118 11540 24124 11552
rect 23799 11512 24124 11540
rect 23799 11509 23811 11512
rect 23753 11503 23811 11509
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24228 11540 24256 11580
rect 29546 11568 29552 11620
rect 29604 11568 29610 11620
rect 29656 11608 29684 11716
rect 30009 11713 30021 11716
rect 30055 11713 30067 11747
rect 30208 11744 30236 11784
rect 30561 11747 30619 11753
rect 30208 11716 30420 11744
rect 30009 11707 30067 11713
rect 29730 11636 29736 11688
rect 29788 11676 29794 11688
rect 29917 11679 29975 11685
rect 29917 11676 29929 11679
rect 29788 11648 29929 11676
rect 29788 11636 29794 11648
rect 29917 11645 29929 11648
rect 29963 11676 29975 11679
rect 29963 11648 30328 11676
rect 29963 11645 29975 11648
rect 29917 11639 29975 11645
rect 30190 11608 30196 11620
rect 29656 11580 30196 11608
rect 30190 11568 30196 11580
rect 30248 11568 30254 11620
rect 24394 11540 24400 11552
rect 24228 11512 24400 11540
rect 24394 11500 24400 11512
rect 24452 11500 24458 11552
rect 25682 11500 25688 11552
rect 25740 11540 25746 11552
rect 29822 11540 29828 11552
rect 25740 11512 29828 11540
rect 25740 11500 25746 11512
rect 29822 11500 29828 11512
rect 29880 11500 29886 11552
rect 30006 11500 30012 11552
rect 30064 11540 30070 11552
rect 30101 11543 30159 11549
rect 30101 11540 30113 11543
rect 30064 11512 30113 11540
rect 30064 11500 30070 11512
rect 30101 11509 30113 11512
rect 30147 11509 30159 11543
rect 30300 11540 30328 11648
rect 30392 11608 30420 11716
rect 30561 11713 30573 11747
rect 30607 11744 30619 11747
rect 30650 11744 30656 11756
rect 30607 11716 30656 11744
rect 30607 11713 30619 11716
rect 30561 11707 30619 11713
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 30760 11744 30788 11784
rect 30834 11772 30840 11824
rect 30892 11812 30898 11824
rect 31312 11812 31340 11852
rect 31665 11849 31677 11852
rect 31711 11849 31723 11883
rect 31665 11843 31723 11849
rect 32122 11840 32128 11892
rect 32180 11840 32186 11892
rect 32306 11840 32312 11892
rect 32364 11840 32370 11892
rect 32493 11883 32551 11889
rect 32493 11849 32505 11883
rect 32539 11880 32551 11883
rect 33226 11880 33232 11892
rect 32539 11852 33232 11880
rect 32539 11849 32551 11852
rect 32493 11843 32551 11849
rect 33226 11840 33232 11852
rect 33284 11840 33290 11892
rect 33318 11840 33324 11892
rect 33376 11880 33382 11892
rect 33613 11883 33671 11889
rect 33613 11880 33625 11883
rect 33376 11852 33625 11880
rect 33376 11840 33382 11852
rect 33613 11849 33625 11852
rect 33659 11849 33671 11883
rect 33613 11843 33671 11849
rect 33781 11883 33839 11889
rect 33781 11849 33793 11883
rect 33827 11880 33839 11883
rect 34606 11880 34612 11892
rect 33827 11852 34612 11880
rect 33827 11849 33839 11852
rect 33781 11843 33839 11849
rect 34606 11840 34612 11852
rect 34664 11840 34670 11892
rect 35434 11840 35440 11892
rect 35492 11880 35498 11892
rect 35621 11883 35679 11889
rect 35621 11880 35633 11883
rect 35492 11852 35633 11880
rect 35492 11840 35498 11852
rect 35621 11849 35633 11852
rect 35667 11880 35679 11883
rect 35710 11880 35716 11892
rect 35667 11852 35716 11880
rect 35667 11849 35679 11852
rect 35621 11843 35679 11849
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 37090 11880 37096 11892
rect 36096 11852 37096 11880
rect 30892 11784 31340 11812
rect 30892 11772 30898 11784
rect 31481 11747 31539 11753
rect 31481 11744 31493 11747
rect 30760 11716 31493 11744
rect 31481 11713 31493 11716
rect 31527 11713 31539 11747
rect 31481 11707 31539 11713
rect 31757 11747 31815 11753
rect 31757 11713 31769 11747
rect 31803 11713 31815 11747
rect 31757 11707 31815 11713
rect 31941 11747 31999 11753
rect 31941 11713 31953 11747
rect 31987 11713 31999 11747
rect 31941 11707 31999 11713
rect 30469 11679 30527 11685
rect 30469 11645 30481 11679
rect 30515 11676 30527 11679
rect 31772 11676 31800 11707
rect 30515 11648 31800 11676
rect 30515 11645 30527 11648
rect 30469 11639 30527 11645
rect 31481 11611 31539 11617
rect 31481 11608 31493 11611
rect 30392 11580 31493 11608
rect 31481 11577 31493 11580
rect 31527 11577 31539 11611
rect 31481 11571 31539 11577
rect 30837 11543 30895 11549
rect 30837 11540 30849 11543
rect 30300 11512 30849 11540
rect 30101 11503 30159 11509
rect 30837 11509 30849 11512
rect 30883 11540 30895 11543
rect 31956 11540 31984 11707
rect 30883 11512 31984 11540
rect 32033 11543 32091 11549
rect 30883 11509 30895 11512
rect 30837 11503 30895 11509
rect 32033 11509 32045 11543
rect 32079 11540 32091 11543
rect 32140 11540 32168 11840
rect 32214 11772 32220 11824
rect 32272 11772 32278 11824
rect 32324 11812 32352 11840
rect 32582 11812 32588 11824
rect 32324 11784 32588 11812
rect 32582 11772 32588 11784
rect 32640 11812 32646 11824
rect 32769 11815 32827 11821
rect 32769 11812 32781 11815
rect 32640 11784 32781 11812
rect 32640 11772 32646 11784
rect 32769 11781 32781 11784
rect 32815 11781 32827 11815
rect 33413 11815 33471 11821
rect 33413 11812 33425 11815
rect 32769 11775 32827 11781
rect 33060 11784 33425 11812
rect 32232 11744 32260 11772
rect 33060 11744 33088 11784
rect 33413 11781 33425 11784
rect 33459 11781 33471 11815
rect 34333 11815 34391 11821
rect 34333 11812 34345 11815
rect 33413 11775 33471 11781
rect 33888 11784 34345 11812
rect 32232 11716 33088 11744
rect 33318 11704 33324 11756
rect 33376 11704 33382 11756
rect 32858 11636 32864 11688
rect 32916 11676 32922 11688
rect 32916 11648 33364 11676
rect 32916 11636 32922 11648
rect 32674 11568 32680 11620
rect 32732 11608 32738 11620
rect 33336 11608 33364 11648
rect 33888 11608 33916 11784
rect 34333 11781 34345 11784
rect 34379 11812 34391 11815
rect 34514 11812 34520 11824
rect 34379 11784 34520 11812
rect 34379 11781 34391 11784
rect 34333 11775 34391 11781
rect 34514 11772 34520 11784
rect 34572 11772 34578 11824
rect 35728 11812 35756 11840
rect 35728 11784 36032 11812
rect 34241 11747 34299 11753
rect 34241 11713 34253 11747
rect 34287 11744 34299 11747
rect 34287 11716 34560 11744
rect 34287 11713 34299 11716
rect 34241 11707 34299 11713
rect 34532 11688 34560 11716
rect 34698 11704 34704 11756
rect 34756 11704 34762 11756
rect 35253 11747 35311 11753
rect 35253 11713 35265 11747
rect 35299 11744 35311 11747
rect 35894 11744 35900 11756
rect 35299 11716 35900 11744
rect 35299 11713 35311 11716
rect 35253 11707 35311 11713
rect 35894 11704 35900 11716
rect 35952 11704 35958 11756
rect 33962 11636 33968 11688
rect 34020 11636 34026 11688
rect 34422 11636 34428 11688
rect 34480 11636 34486 11688
rect 34514 11636 34520 11688
rect 34572 11636 34578 11688
rect 36004 11676 36032 11784
rect 36096 11753 36124 11852
rect 37090 11840 37096 11852
rect 37148 11840 37154 11892
rect 37274 11840 37280 11892
rect 37332 11840 37338 11892
rect 37642 11840 37648 11892
rect 37700 11880 37706 11892
rect 37700 11852 38240 11880
rect 37700 11840 37706 11852
rect 37292 11812 37320 11840
rect 36372 11784 37320 11812
rect 36372 11753 36400 11784
rect 37458 11772 37464 11824
rect 37516 11772 37522 11824
rect 38212 11812 38240 11852
rect 38286 11840 38292 11892
rect 38344 11880 38350 11892
rect 38381 11883 38439 11889
rect 38381 11880 38393 11883
rect 38344 11852 38393 11880
rect 38344 11840 38350 11852
rect 38381 11849 38393 11852
rect 38427 11849 38439 11883
rect 38381 11843 38439 11849
rect 40770 11840 40776 11892
rect 40828 11840 40834 11892
rect 41509 11883 41567 11889
rect 41509 11849 41521 11883
rect 41555 11880 41567 11883
rect 41598 11880 41604 11892
rect 41555 11852 41604 11880
rect 41555 11849 41567 11852
rect 41509 11843 41567 11849
rect 41598 11840 41604 11852
rect 41656 11880 41662 11892
rect 42334 11880 42340 11892
rect 41656 11852 42340 11880
rect 41656 11840 41662 11852
rect 42334 11840 42340 11852
rect 42392 11880 42398 11892
rect 42705 11883 42763 11889
rect 42705 11880 42717 11883
rect 42392 11852 42717 11880
rect 42392 11840 42398 11852
rect 42705 11849 42717 11852
rect 42751 11849 42763 11883
rect 42705 11843 42763 11849
rect 39206 11812 39212 11824
rect 38212 11784 39212 11812
rect 39206 11772 39212 11784
rect 39264 11772 39270 11824
rect 44726 11812 44732 11824
rect 44482 11784 44732 11812
rect 44726 11772 44732 11784
rect 44784 11772 44790 11824
rect 36081 11747 36139 11753
rect 36081 11713 36093 11747
rect 36127 11713 36139 11747
rect 36081 11707 36139 11713
rect 36357 11747 36415 11753
rect 36357 11713 36369 11747
rect 36403 11713 36415 11747
rect 36357 11707 36415 11713
rect 40313 11747 40371 11753
rect 40313 11713 40325 11747
rect 40359 11713 40371 11747
rect 40313 11707 40371 11713
rect 40589 11747 40647 11753
rect 40589 11713 40601 11747
rect 40635 11744 40647 11747
rect 41414 11744 41420 11756
rect 40635 11716 41420 11744
rect 40635 11713 40647 11716
rect 40589 11707 40647 11713
rect 36538 11676 36544 11688
rect 36004 11648 36544 11676
rect 36538 11636 36544 11648
rect 36596 11676 36602 11688
rect 36633 11679 36691 11685
rect 36633 11676 36645 11679
rect 36596 11648 36645 11676
rect 36596 11636 36602 11648
rect 36633 11645 36645 11648
rect 36679 11645 36691 11679
rect 36909 11679 36967 11685
rect 36909 11676 36921 11679
rect 36633 11639 36691 11645
rect 36740 11648 36921 11676
rect 32732 11580 33272 11608
rect 33336 11580 33916 11608
rect 33980 11608 34008 11636
rect 34440 11608 34468 11636
rect 33980 11580 34468 11608
rect 34885 11611 34943 11617
rect 32732 11568 32738 11580
rect 33244 11552 33272 11580
rect 34885 11577 34897 11611
rect 34931 11608 34943 11611
rect 35710 11608 35716 11620
rect 34931 11580 35716 11608
rect 34931 11577 34943 11580
rect 34885 11571 34943 11577
rect 35710 11568 35716 11580
rect 35768 11568 35774 11620
rect 35897 11611 35955 11617
rect 35897 11577 35909 11611
rect 35943 11608 35955 11611
rect 36740 11608 36768 11648
rect 36909 11645 36921 11648
rect 36955 11645 36967 11679
rect 36909 11639 36967 11645
rect 36998 11636 37004 11688
rect 37056 11676 37062 11688
rect 38194 11676 38200 11688
rect 37056 11648 38200 11676
rect 37056 11636 37062 11648
rect 38194 11636 38200 11648
rect 38252 11636 38258 11688
rect 38470 11636 38476 11688
rect 38528 11636 38534 11688
rect 38749 11679 38807 11685
rect 38749 11676 38761 11679
rect 38580 11648 38761 11676
rect 35943 11580 36768 11608
rect 35943 11577 35955 11580
rect 35897 11571 35955 11577
rect 37918 11568 37924 11620
rect 37976 11608 37982 11620
rect 38580 11608 38608 11648
rect 38749 11645 38761 11648
rect 38795 11645 38807 11679
rect 38749 11639 38807 11645
rect 39758 11636 39764 11688
rect 39816 11676 39822 11688
rect 40328 11676 40356 11707
rect 41414 11704 41420 11716
rect 41472 11704 41478 11756
rect 43070 11704 43076 11756
rect 43128 11704 43134 11756
rect 43441 11747 43499 11753
rect 43441 11713 43453 11747
rect 43487 11713 43499 11747
rect 45002 11744 45008 11756
rect 43441 11707 43499 11713
rect 44744 11716 45008 11744
rect 39816 11648 40356 11676
rect 39816 11636 39822 11648
rect 40402 11636 40408 11688
rect 40460 11636 40466 11688
rect 41598 11636 41604 11688
rect 41656 11676 41662 11688
rect 42061 11679 42119 11685
rect 42061 11676 42073 11679
rect 41656 11648 42073 11676
rect 41656 11636 41662 11648
rect 42061 11645 42073 11648
rect 42107 11676 42119 11679
rect 42426 11676 42432 11688
rect 42107 11648 42432 11676
rect 42107 11645 42119 11648
rect 42061 11639 42119 11645
rect 42426 11636 42432 11648
rect 42484 11676 42490 11688
rect 42702 11676 42708 11688
rect 42484 11648 42708 11676
rect 42484 11636 42490 11648
rect 42702 11636 42708 11648
rect 42760 11636 42766 11688
rect 43456 11676 43484 11707
rect 44744 11676 44772 11716
rect 45002 11704 45008 11716
rect 45060 11704 45066 11756
rect 43456 11648 44772 11676
rect 44818 11636 44824 11688
rect 44876 11636 44882 11688
rect 37976 11580 38608 11608
rect 37976 11568 37982 11580
rect 33042 11540 33048 11552
rect 32079 11512 33048 11540
rect 32079 11509 32091 11512
rect 32033 11503 32091 11509
rect 33042 11500 33048 11512
rect 33100 11500 33106 11552
rect 33134 11500 33140 11552
rect 33192 11500 33198 11552
rect 33226 11500 33232 11552
rect 33284 11540 33290 11552
rect 33597 11543 33655 11549
rect 33597 11540 33609 11543
rect 33284 11512 33609 11540
rect 33284 11500 33290 11512
rect 33597 11509 33609 11512
rect 33643 11509 33655 11543
rect 33597 11503 33655 11509
rect 33873 11543 33931 11549
rect 33873 11509 33885 11543
rect 33919 11540 33931 11543
rect 34054 11540 34060 11552
rect 33919 11512 34060 11540
rect 33919 11509 33931 11512
rect 33873 11503 33931 11509
rect 34054 11500 34060 11512
rect 34112 11500 34118 11552
rect 35066 11500 35072 11552
rect 35124 11500 35130 11552
rect 36173 11543 36231 11549
rect 36173 11509 36185 11543
rect 36219 11540 36231 11543
rect 36906 11540 36912 11552
rect 36219 11512 36912 11540
rect 36219 11509 36231 11512
rect 36173 11503 36231 11509
rect 36906 11500 36912 11512
rect 36964 11500 36970 11552
rect 37090 11500 37096 11552
rect 37148 11540 37154 11552
rect 38746 11540 38752 11552
rect 37148 11512 38752 11540
rect 37148 11500 37154 11512
rect 38746 11500 38752 11512
rect 38804 11500 38810 11552
rect 38930 11500 38936 11552
rect 38988 11540 38994 11552
rect 40221 11543 40279 11549
rect 40221 11540 40233 11543
rect 38988 11512 40233 11540
rect 38988 11500 38994 11512
rect 40221 11509 40233 11512
rect 40267 11540 40279 11543
rect 40313 11543 40371 11549
rect 40313 11540 40325 11543
rect 40267 11512 40325 11540
rect 40267 11509 40279 11512
rect 40221 11503 40279 11509
rect 40313 11509 40325 11512
rect 40359 11509 40371 11543
rect 40313 11503 40371 11509
rect 40954 11500 40960 11552
rect 41012 11540 41018 11552
rect 41049 11543 41107 11549
rect 41049 11540 41061 11543
rect 41012 11512 41061 11540
rect 41012 11500 41018 11512
rect 41049 11509 41061 11512
rect 41095 11509 41107 11543
rect 41049 11503 41107 11509
rect 460 11450 45540 11472
rect 460 11398 3570 11450
rect 3622 11398 3634 11450
rect 3686 11398 3698 11450
rect 3750 11398 3762 11450
rect 3814 11398 3826 11450
rect 3878 11398 8570 11450
rect 8622 11398 8634 11450
rect 8686 11398 8698 11450
rect 8750 11398 8762 11450
rect 8814 11398 8826 11450
rect 8878 11398 13570 11450
rect 13622 11398 13634 11450
rect 13686 11398 13698 11450
rect 13750 11398 13762 11450
rect 13814 11398 13826 11450
rect 13878 11398 18570 11450
rect 18622 11398 18634 11450
rect 18686 11398 18698 11450
rect 18750 11398 18762 11450
rect 18814 11398 18826 11450
rect 18878 11398 23570 11450
rect 23622 11398 23634 11450
rect 23686 11398 23698 11450
rect 23750 11398 23762 11450
rect 23814 11398 23826 11450
rect 23878 11398 28570 11450
rect 28622 11398 28634 11450
rect 28686 11398 28698 11450
rect 28750 11398 28762 11450
rect 28814 11398 28826 11450
rect 28878 11398 33570 11450
rect 33622 11398 33634 11450
rect 33686 11398 33698 11450
rect 33750 11398 33762 11450
rect 33814 11398 33826 11450
rect 33878 11398 38570 11450
rect 38622 11398 38634 11450
rect 38686 11398 38698 11450
rect 38750 11398 38762 11450
rect 38814 11398 38826 11450
rect 38878 11398 43570 11450
rect 43622 11398 43634 11450
rect 43686 11398 43698 11450
rect 43750 11398 43762 11450
rect 43814 11398 43826 11450
rect 43878 11398 45540 11450
rect 460 11376 45540 11398
rect 5445 11339 5503 11345
rect 5445 11305 5457 11339
rect 5491 11336 5503 11339
rect 7009 11339 7067 11345
rect 7009 11336 7021 11339
rect 5491 11308 7021 11336
rect 5491 11305 5503 11308
rect 5445 11299 5503 11305
rect 7009 11305 7021 11308
rect 7055 11336 7067 11339
rect 7098 11336 7104 11348
rect 7055 11308 7104 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 7098 11296 7104 11308
rect 7156 11336 7162 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7156 11308 7757 11336
rect 7156 11296 7162 11308
rect 7745 11305 7757 11308
rect 7791 11336 7803 11339
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7791 11308 8125 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8113 11305 8125 11308
rect 8159 11336 8171 11339
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8159 11308 8861 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 8849 11305 8861 11308
rect 8895 11336 8907 11339
rect 10134 11336 10140 11348
rect 8895 11308 10140 11336
rect 8895 11305 8907 11308
rect 8849 11299 8907 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 12584 11308 13461 11336
rect 12584 11296 12590 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 11716 11268 11744 11296
rect 11471 11240 11744 11268
rect 11900 11240 12572 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 11900 11200 11928 11240
rect 5123 11172 5396 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5368 11144 5396 11172
rect 10428 11172 11928 11200
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 4982 11132 4988 11144
rect 4939 11104 4988 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4816 11064 4844 11095
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9324 11104 9413 11132
rect 4212 11036 5212 11064
rect 4212 11024 4218 11036
rect 5184 11008 5212 11036
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8444 11036 8953 11064
rect 8444 11024 8450 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 9088 11036 9137 11064
rect 9088 11024 9094 11036
rect 9125 11033 9137 11036
rect 9171 11033 9183 11067
rect 9125 11027 9183 11033
rect 9324 11008 9352 11104
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 9674 11132 9680 11144
rect 9631 11104 9680 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 10428 11141 10456 11172
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 11256 11141 11284 11172
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11422 11132 11428 11144
rect 11379 11104 11428 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 9490 11024 9496 11076
rect 9548 11024 9554 11076
rect 10704 11064 10732 11095
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11900 11141 11928 11172
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 12023 11172 12449 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12437 11169 12449 11172
rect 12483 11169 12495 11203
rect 12544 11200 12572 11240
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 12805 11271 12863 11277
rect 12805 11268 12817 11271
rect 12676 11240 12817 11268
rect 12676 11228 12682 11240
rect 12805 11237 12817 11240
rect 12851 11268 12863 11271
rect 12986 11268 12992 11280
rect 12851 11240 12992 11268
rect 12851 11237 12863 11240
rect 12805 11231 12863 11237
rect 12986 11228 12992 11240
rect 13044 11228 13050 11280
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 13136 11240 13185 11268
rect 13136 11228 13142 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 12544 11172 13676 11200
rect 12437 11163 12495 11169
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11532 11064 11560 11095
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12176 11064 12204 11095
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 13648 11141 13676 11172
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 14108 11200 14136 11299
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 17000 11308 18245 11336
rect 17000 11296 17006 11308
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18233 11299 18291 11305
rect 18785 11339 18843 11345
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 19058 11336 19064 11348
rect 18831 11308 19064 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 19521 11339 19579 11345
rect 19521 11305 19533 11339
rect 19567 11336 19579 11339
rect 20714 11336 20720 11348
rect 19567 11308 20720 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20956 11308 21005 11336
rect 20956 11296 20962 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21358 11336 21364 11348
rect 21223 11308 21364 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22002 11296 22008 11348
rect 22060 11296 22066 11348
rect 23290 11296 23296 11348
rect 23348 11296 23354 11348
rect 24118 11296 24124 11348
rect 24176 11296 24182 11348
rect 24949 11339 25007 11345
rect 24949 11305 24961 11339
rect 24995 11336 25007 11339
rect 25958 11336 25964 11348
rect 24995 11308 25964 11336
rect 24995 11305 25007 11308
rect 24949 11299 25007 11305
rect 25958 11296 25964 11308
rect 26016 11296 26022 11348
rect 26234 11296 26240 11348
rect 26292 11296 26298 11348
rect 27614 11296 27620 11348
rect 27672 11296 27678 11348
rect 27890 11296 27896 11348
rect 27948 11296 27954 11348
rect 27985 11339 28043 11345
rect 27985 11305 27997 11339
rect 28031 11336 28043 11339
rect 28442 11336 28448 11348
rect 28031 11308 28448 11336
rect 28031 11305 28043 11308
rect 27985 11299 28043 11305
rect 28442 11296 28448 11308
rect 28500 11296 28506 11348
rect 29638 11296 29644 11348
rect 29696 11336 29702 11348
rect 29696 11308 30144 11336
rect 29696 11296 29702 11308
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 14645 11271 14703 11277
rect 14645 11268 14657 11271
rect 14424 11240 14657 11268
rect 14424 11228 14430 11240
rect 14645 11237 14657 11240
rect 14691 11237 14703 11271
rect 14645 11231 14703 11237
rect 17589 11271 17647 11277
rect 17589 11237 17601 11271
rect 17635 11268 17647 11271
rect 17678 11268 17684 11280
rect 17635 11240 17684 11268
rect 17635 11237 17647 11240
rect 17589 11231 17647 11237
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 21634 11268 21640 11280
rect 17828 11240 21640 11268
rect 17828 11228 17834 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 23382 11268 23388 11280
rect 22664 11240 23388 11268
rect 22664 11212 22692 11240
rect 23382 11228 23388 11240
rect 23440 11268 23446 11280
rect 24136 11268 24164 11296
rect 25317 11271 25375 11277
rect 25317 11268 25329 11271
rect 23440 11240 23704 11268
rect 24136 11240 25329 11268
rect 23440 11228 23446 11240
rect 19334 11200 19340 11212
rect 13872 11172 14136 11200
rect 17788 11172 19340 11200
rect 13872 11160 13878 11172
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 13722 11132 13728 11144
rect 13679 11104 13728 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13832 11073 13860 11160
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 10704 11036 12204 11064
rect 4338 10956 4344 11008
rect 4396 10996 4402 11008
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 4396 10968 5089 10996
rect 4396 10956 4402 10968
rect 5077 10965 5089 10968
rect 5123 10965 5135 10999
rect 5077 10959 5135 10965
rect 5166 10956 5172 11008
rect 5224 10956 5230 11008
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5718 10996 5724 11008
rect 5592 10968 5724 10996
rect 5592 10956 5598 10968
rect 5718 10956 5724 10968
rect 5776 10996 5782 11008
rect 5994 10996 6000 11008
rect 5776 10968 6000 10996
rect 5776 10956 5782 10968
rect 5994 10956 6000 10968
rect 6052 10996 6058 11008
rect 6181 10999 6239 11005
rect 6181 10996 6193 10999
rect 6052 10968 6193 10996
rect 6052 10956 6058 10968
rect 6181 10965 6193 10968
rect 6227 10996 6239 10999
rect 6549 10999 6607 11005
rect 6549 10996 6561 10999
rect 6227 10968 6561 10996
rect 6227 10965 6239 10968
rect 6181 10959 6239 10965
rect 6549 10965 6561 10968
rect 6595 10996 6607 10999
rect 7285 10999 7343 11005
rect 7285 10996 7297 10999
rect 6595 10968 7297 10996
rect 6595 10965 6607 10968
rect 6549 10959 6607 10965
rect 7285 10965 7297 10968
rect 7331 10965 7343 10999
rect 7285 10959 7343 10965
rect 9306 10956 9312 11008
rect 9364 10956 9370 11008
rect 10226 10956 10232 11008
rect 10284 10956 10290 11008
rect 11057 10999 11115 11005
rect 11057 10965 11069 10999
rect 11103 10996 11115 10999
rect 11422 10996 11428 11008
rect 11103 10968 11428 10996
rect 11103 10965 11115 10968
rect 11057 10959 11115 10965
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 11698 10956 11704 11008
rect 11756 10956 11762 11008
rect 12176 10996 12204 11036
rect 13817 11067 13875 11073
rect 13817 11033 13829 11067
rect 13863 11033 13875 11067
rect 13817 11027 13875 11033
rect 13924 11008 13952 11095
rect 13998 11092 14004 11144
rect 14056 11092 14062 11144
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14108 11064 14136 11095
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 17788 11141 17816 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 19576 11172 20085 11200
rect 19576 11160 19582 11172
rect 20073 11169 20085 11172
rect 20119 11169 20131 11203
rect 20254 11200 20260 11212
rect 20073 11163 20131 11169
rect 20180 11172 20260 11200
rect 15105 11135 15163 11141
rect 15105 11132 15117 11135
rect 15068 11104 15117 11132
rect 15068 11092 15074 11104
rect 15105 11101 15117 11104
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 18693 11135 18751 11141
rect 17972 11104 18644 11132
rect 14016 11036 14136 11064
rect 15381 11067 15439 11073
rect 14016 11008 14044 11036
rect 15381 11033 15393 11067
rect 15427 11064 15439 11067
rect 15654 11064 15660 11076
rect 15427 11036 15660 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 15654 11024 15660 11036
rect 15712 11024 15718 11076
rect 15838 11024 15844 11076
rect 15896 11024 15902 11076
rect 17497 11067 17555 11073
rect 17497 11033 17509 11067
rect 17543 11064 17555 11067
rect 17972 11064 18000 11104
rect 17543 11036 18000 11064
rect 18049 11067 18107 11073
rect 17543 11033 17555 11036
rect 17497 11027 17555 11033
rect 18049 11033 18061 11067
rect 18095 11033 18107 11067
rect 18616 11064 18644 11104
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 19242 11132 19248 11144
rect 18739 11104 19248 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20180 11141 20208 11172
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 21729 11203 21787 11209
rect 21729 11169 21741 11203
rect 21775 11169 21787 11203
rect 21729 11163 21787 11169
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20404 11104 20668 11132
rect 20404 11092 20410 11104
rect 20640 11064 20668 11104
rect 20898 11092 20904 11144
rect 20956 11092 20962 11144
rect 21744 11064 21772 11163
rect 22462 11160 22468 11212
rect 22520 11160 22526 11212
rect 22646 11160 22652 11212
rect 22704 11160 22710 11212
rect 22830 11160 22836 11212
rect 22888 11160 22894 11212
rect 23676 11200 23704 11240
rect 25317 11237 25329 11240
rect 25363 11268 25375 11271
rect 25682 11268 25688 11280
rect 25363 11240 25688 11268
rect 25363 11237 25375 11240
rect 25317 11231 25375 11237
rect 25682 11228 25688 11240
rect 25740 11228 25746 11280
rect 24213 11203 24271 11209
rect 24213 11200 24225 11203
rect 23676 11172 24225 11200
rect 24213 11169 24225 11172
rect 24259 11200 24271 11203
rect 24578 11200 24584 11212
rect 24259 11172 24584 11200
rect 24259 11169 24271 11172
rect 24213 11163 24271 11169
rect 24578 11160 24584 11172
rect 24636 11160 24642 11212
rect 25958 11160 25964 11212
rect 26016 11200 26022 11212
rect 26145 11203 26203 11209
rect 26145 11200 26157 11203
rect 26016 11172 26157 11200
rect 26016 11160 26022 11172
rect 26145 11169 26157 11172
rect 26191 11200 26203 11203
rect 26252 11200 26280 11296
rect 26191 11172 26280 11200
rect 26421 11203 26479 11209
rect 26191 11169 26203 11172
rect 26145 11163 26203 11169
rect 26421 11169 26433 11203
rect 26467 11200 26479 11203
rect 26970 11200 26976 11212
rect 26467 11172 26976 11200
rect 26467 11169 26479 11172
rect 26421 11163 26479 11169
rect 26970 11160 26976 11172
rect 27028 11160 27034 11212
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22278 11092 22284 11144
rect 22336 11092 22342 11144
rect 22557 11135 22615 11141
rect 22557 11101 22569 11135
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 18616 11036 20592 11064
rect 20640 11036 21772 11064
rect 18049 11027 18107 11033
rect 13630 10996 13636 11008
rect 12176 10968 13636 10996
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 13906 10956 13912 11008
rect 13964 10956 13970 11008
rect 13998 10956 14004 11008
rect 14056 10956 14062 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 14332 10968 14381 10996
rect 14332 10956 14338 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 14369 10959 14427 10965
rect 16850 10956 16856 11008
rect 16908 10956 16914 11008
rect 18064 10996 18092 11027
rect 18966 10996 18972 11008
rect 18064 10968 18972 10996
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 19889 10999 19947 11005
rect 19889 10965 19901 10999
rect 19935 10996 19947 10999
rect 20254 10996 20260 11008
rect 19935 10968 20260 10996
rect 19935 10965 19947 10968
rect 19889 10959 19947 10965
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 20564 10996 20592 11036
rect 21542 10996 21548 11008
rect 20564 10968 21548 10996
rect 21542 10956 21548 10968
rect 21600 10956 21606 11008
rect 21634 10956 21640 11008
rect 21692 10996 21698 11008
rect 21910 10996 21916 11008
rect 21692 10968 21916 10996
rect 21692 10956 21698 10968
rect 21910 10956 21916 10968
rect 21968 10996 21974 11008
rect 22572 10996 22600 11095
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 22848 11132 22876 11160
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 22848 11104 22937 11132
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 24026 11092 24032 11144
rect 24084 11092 24090 11144
rect 24394 11092 24400 11144
rect 24452 11132 24458 11144
rect 24673 11135 24731 11141
rect 24673 11132 24685 11135
rect 24452 11104 24685 11132
rect 24452 11092 24458 11104
rect 24673 11101 24685 11104
rect 24719 11101 24731 11135
rect 27632 11132 27660 11296
rect 29454 11268 29460 11280
rect 28552 11240 29460 11268
rect 28552 11141 28580 11240
rect 29454 11228 29460 11240
rect 29512 11228 29518 11280
rect 29178 11160 29184 11212
rect 29236 11200 29242 11212
rect 29273 11203 29331 11209
rect 29273 11200 29285 11203
rect 29236 11172 29285 11200
rect 29236 11160 29242 11172
rect 29273 11169 29285 11172
rect 29319 11200 29331 11203
rect 29638 11200 29644 11212
rect 29319 11172 29644 11200
rect 29319 11169 29331 11172
rect 29273 11163 29331 11169
rect 29638 11160 29644 11172
rect 29696 11160 29702 11212
rect 30116 11209 30144 11308
rect 31754 11296 31760 11348
rect 31812 11336 31818 11348
rect 32401 11339 32459 11345
rect 32401 11336 32413 11339
rect 31812 11308 32413 11336
rect 31812 11296 31818 11308
rect 32401 11305 32413 11308
rect 32447 11336 32459 11339
rect 32674 11336 32680 11348
rect 32447 11308 32680 11336
rect 32447 11305 32459 11308
rect 32401 11299 32459 11305
rect 32674 11296 32680 11308
rect 32732 11336 32738 11348
rect 32861 11339 32919 11345
rect 32861 11336 32873 11339
rect 32732 11308 32873 11336
rect 32732 11296 32738 11308
rect 32861 11305 32873 11308
rect 32907 11305 32919 11339
rect 33318 11336 33324 11348
rect 32861 11299 32919 11305
rect 33244 11308 33324 11336
rect 31846 11228 31852 11280
rect 31904 11268 31910 11280
rect 32585 11271 32643 11277
rect 31904 11240 32444 11268
rect 31904 11228 31910 11240
rect 30101 11203 30159 11209
rect 30101 11169 30113 11203
rect 30147 11200 30159 11203
rect 30742 11200 30748 11212
rect 30147 11172 30748 11200
rect 30147 11169 30159 11172
rect 30101 11163 30159 11169
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 31662 11160 31668 11212
rect 31720 11200 31726 11212
rect 32125 11203 32183 11209
rect 32125 11200 32137 11203
rect 31720 11172 32137 11200
rect 31720 11160 31726 11172
rect 32125 11169 32137 11172
rect 32171 11169 32183 11203
rect 32125 11163 32183 11169
rect 28169 11135 28227 11141
rect 28169 11132 28181 11135
rect 27632 11104 28181 11132
rect 24673 11095 24731 11101
rect 28169 11101 28181 11104
rect 28215 11101 28227 11135
rect 28169 11095 28227 11101
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28997 11135 29055 11141
rect 28997 11101 29009 11135
rect 29043 11132 29055 11135
rect 29730 11132 29736 11144
rect 29043 11104 29736 11132
rect 29043 11101 29055 11104
rect 28997 11095 29055 11101
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 32030 11132 32036 11144
rect 31510 11104 32036 11132
rect 32030 11092 32036 11104
rect 32088 11132 32094 11144
rect 32306 11132 32312 11144
rect 32088 11104 32312 11132
rect 32088 11092 32094 11104
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 32416 11132 32444 11240
rect 32585 11237 32597 11271
rect 32631 11268 32643 11271
rect 33045 11271 33103 11277
rect 33045 11268 33057 11271
rect 32631 11240 32720 11268
rect 32631 11237 32643 11240
rect 32585 11231 32643 11237
rect 32692 11212 32720 11240
rect 32876 11240 33057 11268
rect 32876 11212 32904 11240
rect 33045 11237 33057 11240
rect 33091 11237 33103 11271
rect 33045 11231 33103 11237
rect 33137 11271 33195 11277
rect 33137 11237 33149 11271
rect 33183 11268 33195 11271
rect 33244 11268 33272 11308
rect 33318 11296 33324 11308
rect 33376 11296 33382 11348
rect 36998 11336 37004 11348
rect 33628 11308 37004 11336
rect 33183 11240 33272 11268
rect 33183 11237 33195 11240
rect 33137 11231 33195 11237
rect 32674 11160 32680 11212
rect 32732 11160 32738 11212
rect 32858 11160 32864 11212
rect 32916 11160 32922 11212
rect 32950 11160 32956 11212
rect 33008 11200 33014 11212
rect 33628 11209 33656 11308
rect 36998 11296 37004 11308
rect 37056 11296 37062 11348
rect 37185 11339 37243 11345
rect 37185 11305 37197 11339
rect 37231 11336 37243 11339
rect 37918 11336 37924 11348
rect 37231 11308 37924 11336
rect 37231 11305 37243 11308
rect 37185 11299 37243 11305
rect 37918 11296 37924 11308
rect 37976 11296 37982 11348
rect 38838 11336 38844 11348
rect 38028 11308 38844 11336
rect 33597 11203 33656 11209
rect 33597 11200 33609 11203
rect 33008 11172 33609 11200
rect 33008 11160 33014 11172
rect 33597 11169 33609 11172
rect 33643 11172 33656 11203
rect 33781 11203 33839 11209
rect 33643 11169 33655 11172
rect 33597 11163 33655 11169
rect 33781 11169 33793 11203
rect 33827 11200 33839 11203
rect 33962 11200 33968 11212
rect 33827 11172 33968 11200
rect 33827 11169 33839 11172
rect 33781 11163 33839 11169
rect 33962 11160 33968 11172
rect 34020 11160 34026 11212
rect 34054 11160 34060 11212
rect 34112 11160 34118 11212
rect 34422 11160 34428 11212
rect 34480 11200 34486 11212
rect 35434 11200 35440 11212
rect 34480 11172 35440 11200
rect 34480 11160 34486 11172
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 35710 11160 35716 11212
rect 35768 11200 35774 11212
rect 38028 11209 38056 11308
rect 38838 11296 38844 11308
rect 38896 11336 38902 11348
rect 39298 11336 39304 11348
rect 38896 11308 39304 11336
rect 38896 11296 38902 11308
rect 39298 11296 39304 11308
rect 39356 11296 39362 11348
rect 39942 11296 39948 11348
rect 40000 11336 40006 11348
rect 42613 11339 42671 11345
rect 40000 11308 42288 11336
rect 40000 11296 40006 11308
rect 38289 11271 38347 11277
rect 38289 11237 38301 11271
rect 38335 11237 38347 11271
rect 41141 11271 41199 11277
rect 38289 11231 38347 11237
rect 38764 11240 38976 11268
rect 38013 11203 38071 11209
rect 38013 11200 38025 11203
rect 35768 11172 38025 11200
rect 35768 11160 35774 11172
rect 38013 11169 38025 11172
rect 38059 11169 38071 11203
rect 38013 11163 38071 11169
rect 34072 11132 34100 11160
rect 34241 11135 34299 11141
rect 34241 11132 34253 11135
rect 32416 11104 32812 11132
rect 34072 11104 34253 11132
rect 22756 11064 22784 11092
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 22756 11036 23121 11064
rect 23109 11033 23121 11036
rect 23155 11033 23167 11067
rect 27706 11064 27712 11076
rect 27646 11036 27712 11064
rect 23109 11027 23167 11033
rect 27706 11024 27712 11036
rect 27764 11024 27770 11076
rect 29362 11024 29368 11076
rect 29420 11024 29426 11076
rect 29546 11024 29552 11076
rect 29604 11024 29610 11076
rect 30377 11067 30435 11073
rect 30377 11033 30389 11067
rect 30423 11064 30435 11067
rect 30650 11064 30656 11076
rect 30423 11036 30656 11064
rect 30423 11033 30435 11036
rect 30377 11027 30435 11033
rect 30650 11024 30656 11036
rect 30708 11024 30714 11076
rect 32217 11067 32275 11073
rect 32217 11033 32229 11067
rect 32263 11064 32275 11067
rect 32677 11067 32735 11073
rect 32263 11036 32536 11064
rect 32263 11033 32275 11036
rect 32217 11027 32275 11033
rect 22922 10996 22928 11008
rect 21968 10968 22928 10996
rect 21968 10956 21974 10968
rect 22922 10956 22928 10968
rect 22980 10956 22986 11008
rect 25590 10956 25596 11008
rect 25648 10996 25654 11008
rect 25685 10999 25743 11005
rect 25685 10996 25697 10999
rect 25648 10968 25697 10996
rect 25648 10956 25654 10968
rect 25685 10965 25697 10968
rect 25731 10965 25743 10999
rect 25685 10959 25743 10965
rect 28442 10956 28448 11008
rect 28500 10996 28506 11008
rect 28629 10999 28687 11005
rect 28629 10996 28641 10999
rect 28500 10968 28641 10996
rect 28500 10956 28506 10968
rect 28629 10965 28641 10968
rect 28675 10965 28687 10999
rect 29380 10996 29408 11024
rect 32324 11008 32352 11036
rect 29641 10999 29699 11005
rect 29641 10996 29653 10999
rect 29380 10968 29653 10996
rect 28629 10959 28687 10965
rect 29641 10965 29653 10968
rect 29687 10965 29699 10999
rect 29641 10959 29699 10965
rect 32306 10956 32312 11008
rect 32364 10956 32370 11008
rect 32398 10956 32404 11008
rect 32456 11005 32462 11008
rect 32456 10999 32480 11005
rect 32468 10965 32480 10999
rect 32508 10996 32536 11036
rect 32677 11033 32689 11067
rect 32723 11033 32735 11067
rect 32677 11027 32735 11033
rect 32692 10996 32720 11027
rect 32508 10968 32720 10996
rect 32784 10996 32812 11104
rect 34241 11101 34253 11104
rect 34287 11101 34299 11135
rect 36541 11135 36599 11141
rect 36541 11132 36553 11135
rect 35834 11118 36553 11132
rect 34241 11095 34299 11101
rect 35820 11104 36553 11118
rect 33505 11067 33563 11073
rect 33505 11033 33517 11067
rect 33551 11064 33563 11067
rect 34330 11064 34336 11076
rect 33551 11036 34336 11064
rect 33551 11033 33563 11036
rect 33505 11027 33563 11033
rect 34330 11024 34336 11036
rect 34388 11024 34394 11076
rect 34701 11067 34759 11073
rect 34701 11033 34713 11067
rect 34747 11064 34759 11067
rect 34974 11064 34980 11076
rect 34747 11036 34980 11064
rect 34747 11033 34759 11036
rect 34701 11027 34759 11033
rect 34974 11024 34980 11036
rect 35032 11024 35038 11076
rect 35084 11036 35190 11064
rect 32887 10999 32945 11005
rect 32887 10996 32899 10999
rect 32784 10968 32899 10996
rect 32456 10959 32480 10965
rect 32887 10965 32899 10968
rect 32933 10996 32945 10999
rect 33318 10996 33324 11008
rect 32933 10968 33324 10996
rect 32933 10965 32945 10968
rect 32887 10959 32945 10965
rect 32456 10956 32462 10959
rect 33318 10956 33324 10968
rect 33376 10956 33382 11008
rect 33870 10956 33876 11008
rect 33928 10996 33934 11008
rect 34057 10999 34115 11005
rect 34057 10996 34069 10999
rect 33928 10968 34069 10996
rect 33928 10956 33934 10968
rect 34057 10965 34069 10968
rect 34103 10965 34115 10999
rect 34057 10959 34115 10965
rect 34882 10956 34888 11008
rect 34940 10996 34946 11008
rect 35084 10996 35112 11036
rect 35820 10996 35848 11104
rect 36541 11101 36553 11104
rect 36587 11101 36599 11135
rect 36541 11095 36599 11101
rect 34940 10968 35848 10996
rect 34940 10956 34946 10968
rect 36078 10956 36084 11008
rect 36136 10996 36142 11008
rect 36173 10999 36231 11005
rect 36173 10996 36185 10999
rect 36136 10968 36185 10996
rect 36136 10956 36142 10968
rect 36173 10965 36185 10968
rect 36219 10965 36231 10999
rect 36556 10996 36584 11095
rect 36630 11092 36636 11144
rect 36688 11092 36694 11144
rect 37369 11135 37427 11141
rect 37369 11101 37381 11135
rect 37415 11132 37427 11135
rect 38304 11132 38332 11231
rect 38764 11209 38792 11240
rect 38749 11203 38807 11209
rect 38749 11169 38761 11203
rect 38795 11169 38807 11203
rect 38749 11163 38807 11169
rect 38838 11160 38844 11212
rect 38896 11160 38902 11212
rect 38948 11200 38976 11240
rect 41141 11237 41153 11271
rect 41187 11268 41199 11271
rect 41966 11268 41972 11280
rect 41187 11240 41972 11268
rect 41187 11237 41199 11240
rect 41141 11231 41199 11237
rect 41966 11228 41972 11240
rect 42024 11228 42030 11280
rect 39022 11200 39028 11212
rect 38948 11172 39028 11200
rect 39022 11160 39028 11172
rect 39080 11200 39086 11212
rect 41598 11200 41604 11212
rect 39080 11172 41604 11200
rect 39080 11160 39086 11172
rect 41598 11160 41604 11172
rect 41656 11160 41662 11212
rect 41785 11203 41843 11209
rect 41785 11169 41797 11203
rect 41831 11200 41843 11203
rect 42058 11200 42064 11212
rect 41831 11172 42064 11200
rect 41831 11169 41843 11172
rect 41785 11163 41843 11169
rect 42058 11160 42064 11172
rect 42116 11160 42122 11212
rect 37415 11104 38332 11132
rect 37415 11101 37427 11104
rect 37369 11095 37427 11101
rect 38654 11092 38660 11144
rect 38712 11092 38718 11144
rect 39209 11135 39267 11141
rect 39209 11132 39221 11135
rect 38948 11104 39221 11132
rect 36648 11064 36676 11092
rect 37090 11064 37096 11076
rect 36648 11036 37096 11064
rect 37090 11024 37096 11036
rect 37148 11064 37154 11076
rect 37829 11067 37887 11073
rect 37148 11036 37780 11064
rect 37148 11024 37154 11036
rect 36817 10999 36875 11005
rect 36817 10996 36829 10999
rect 36556 10968 36829 10996
rect 36173 10959 36231 10965
rect 36817 10965 36829 10968
rect 36863 10965 36875 10999
rect 36817 10959 36875 10965
rect 37458 10956 37464 11008
rect 37516 10956 37522 11008
rect 37752 10996 37780 11036
rect 37829 11033 37841 11067
rect 37875 11064 37887 11067
rect 38562 11064 38568 11076
rect 37875 11036 38568 11064
rect 37875 11033 37887 11036
rect 37829 11027 37887 11033
rect 38562 11024 38568 11036
rect 38620 11024 38626 11076
rect 37921 10999 37979 11005
rect 37921 10996 37933 10999
rect 37752 10968 37933 10996
rect 37921 10965 37933 10968
rect 37967 10965 37979 10999
rect 37921 10959 37979 10965
rect 38470 10956 38476 11008
rect 38528 10996 38534 11008
rect 38948 10996 38976 11104
rect 39209 11101 39221 11104
rect 39255 11101 39267 11135
rect 39209 11095 39267 11101
rect 41506 11092 41512 11144
rect 41564 11092 41570 11144
rect 42260 11141 42288 11308
rect 42613 11305 42625 11339
rect 42659 11336 42671 11339
rect 42794 11336 42800 11348
rect 42659 11308 42800 11336
rect 42659 11305 42671 11308
rect 42613 11299 42671 11305
rect 42794 11296 42800 11308
rect 42852 11296 42858 11348
rect 43349 11339 43407 11345
rect 43349 11305 43361 11339
rect 43395 11336 43407 11339
rect 44542 11336 44548 11348
rect 43395 11308 44548 11336
rect 43395 11305 43407 11308
rect 43349 11299 43407 11305
rect 44542 11296 44548 11308
rect 44600 11296 44606 11348
rect 42702 11228 42708 11280
rect 42760 11268 42766 11280
rect 43625 11271 43683 11277
rect 43625 11268 43637 11271
rect 42760 11240 43637 11268
rect 42760 11228 42766 11240
rect 43625 11237 43637 11240
rect 43671 11237 43683 11271
rect 43625 11231 43683 11237
rect 42245 11135 42303 11141
rect 42245 11101 42257 11135
rect 42291 11132 42303 11135
rect 43438 11132 43444 11144
rect 42291 11104 43444 11132
rect 42291 11101 42303 11104
rect 42245 11095 42303 11101
rect 43438 11092 43444 11104
rect 43496 11092 43502 11144
rect 39022 11024 39028 11076
rect 39080 11064 39086 11076
rect 39485 11067 39543 11073
rect 39485 11064 39497 11067
rect 39080 11036 39497 11064
rect 39080 11024 39086 11036
rect 39485 11033 39497 11036
rect 39531 11033 39543 11067
rect 39485 11027 39543 11033
rect 39942 11024 39948 11076
rect 40000 11024 40006 11076
rect 40770 11024 40776 11076
rect 40828 11064 40834 11076
rect 42794 11064 42800 11076
rect 40828 11036 42800 11064
rect 40828 11024 40834 11036
rect 42794 11024 42800 11036
rect 42852 11024 42858 11076
rect 44085 11067 44143 11073
rect 44085 11033 44097 11067
rect 44131 11064 44143 11067
rect 44131 11036 44772 11064
rect 44131 11033 44143 11036
rect 44085 11027 44143 11033
rect 44744 11008 44772 11036
rect 39666 10996 39672 11008
rect 38528 10968 39672 10996
rect 38528 10956 38534 10968
rect 39666 10956 39672 10968
rect 39724 10956 39730 11008
rect 40310 10956 40316 11008
rect 40368 10996 40374 11008
rect 40957 10999 41015 11005
rect 40957 10996 40969 10999
rect 40368 10968 40969 10996
rect 40368 10956 40374 10968
rect 40957 10965 40969 10968
rect 41003 10965 41015 10999
rect 40957 10959 41015 10965
rect 41601 10999 41659 11005
rect 41601 10965 41613 10999
rect 41647 10996 41659 10999
rect 41874 10996 41880 11008
rect 41647 10968 41880 10996
rect 41647 10965 41659 10968
rect 41601 10959 41659 10965
rect 41874 10956 41880 10968
rect 41932 10956 41938 11008
rect 42978 10956 42984 11008
rect 43036 10956 43042 11008
rect 44542 10956 44548 11008
rect 44600 10956 44606 11008
rect 44726 10956 44732 11008
rect 44784 10996 44790 11008
rect 44913 10999 44971 11005
rect 44913 10996 44925 10999
rect 44784 10968 44925 10996
rect 44784 10956 44790 10968
rect 44913 10965 44925 10968
rect 44959 10965 44971 10999
rect 44913 10959 44971 10965
rect 460 10906 45540 10928
rect 460 10854 6070 10906
rect 6122 10854 6134 10906
rect 6186 10854 6198 10906
rect 6250 10854 6262 10906
rect 6314 10854 6326 10906
rect 6378 10854 11070 10906
rect 11122 10854 11134 10906
rect 11186 10854 11198 10906
rect 11250 10854 11262 10906
rect 11314 10854 11326 10906
rect 11378 10854 16070 10906
rect 16122 10854 16134 10906
rect 16186 10854 16198 10906
rect 16250 10854 16262 10906
rect 16314 10854 16326 10906
rect 16378 10854 21070 10906
rect 21122 10854 21134 10906
rect 21186 10854 21198 10906
rect 21250 10854 21262 10906
rect 21314 10854 21326 10906
rect 21378 10854 26070 10906
rect 26122 10854 26134 10906
rect 26186 10854 26198 10906
rect 26250 10854 26262 10906
rect 26314 10854 26326 10906
rect 26378 10854 31070 10906
rect 31122 10854 31134 10906
rect 31186 10854 31198 10906
rect 31250 10854 31262 10906
rect 31314 10854 31326 10906
rect 31378 10854 36070 10906
rect 36122 10854 36134 10906
rect 36186 10854 36198 10906
rect 36250 10854 36262 10906
rect 36314 10854 36326 10906
rect 36378 10854 41070 10906
rect 41122 10854 41134 10906
rect 41186 10854 41198 10906
rect 41250 10854 41262 10906
rect 41314 10854 41326 10906
rect 41378 10854 45540 10906
rect 460 10832 45540 10854
rect 7098 10792 7104 10804
rect 5644 10764 7104 10792
rect 5644 10724 5672 10764
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 9306 10792 9312 10804
rect 8527 10764 9312 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 11514 10792 11520 10804
rect 10643 10764 11520 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 11848 10764 12633 10792
rect 11848 10752 11854 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 13078 10752 13084 10804
rect 13136 10752 13142 10804
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 14332 10764 14872 10792
rect 14332 10752 14338 10764
rect 6089 10727 6147 10733
rect 6089 10724 6101 10727
rect 4554 10696 5672 10724
rect 5736 10696 6101 10724
rect 5736 10665 5764 10696
rect 6089 10693 6101 10696
rect 6135 10693 6147 10727
rect 9030 10724 9036 10736
rect 6089 10687 6147 10693
rect 8220 10696 9036 10724
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5721 10659 5779 10665
rect 5123 10628 5396 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5368 10600 5396 10628
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5902 10616 5908 10668
rect 5960 10616 5966 10668
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3068 10452 3096 10551
rect 3326 10548 3332 10600
rect 3384 10548 3390 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10588 4859 10591
rect 5166 10588 5172 10600
rect 4847 10560 5172 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 6012 10588 6040 10619
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 8220 10665 8248 10696
rect 9030 10684 9036 10696
rect 9088 10684 9094 10736
rect 10226 10684 10232 10736
rect 10284 10684 10290 10736
rect 11149 10727 11207 10733
rect 11149 10693 11161 10727
rect 11195 10724 11207 10727
rect 11422 10724 11428 10736
rect 11195 10696 11428 10724
rect 11195 10693 11207 10696
rect 11149 10687 11207 10693
rect 11422 10684 11428 10696
rect 11480 10684 11486 10736
rect 12158 10684 12164 10736
rect 12216 10684 12222 10736
rect 13096 10724 13124 10752
rect 14844 10733 14872 10764
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17770 10792 17776 10804
rect 17184 10764 17776 10792
rect 17184 10752 17190 10764
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 18966 10752 18972 10804
rect 19024 10752 19030 10804
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 21821 10795 21879 10801
rect 19300 10764 21772 10792
rect 19300 10752 19306 10764
rect 14829 10727 14887 10733
rect 13096 10696 13754 10724
rect 14829 10693 14841 10727
rect 14875 10693 14887 10727
rect 14829 10687 14887 10693
rect 15013 10727 15071 10733
rect 15013 10693 15025 10727
rect 15059 10724 15071 10727
rect 15102 10724 15108 10736
rect 15059 10696 15108 10724
rect 15059 10693 15071 10696
rect 15013 10687 15071 10693
rect 15102 10684 15108 10696
rect 15160 10724 15166 10736
rect 15930 10724 15936 10736
rect 15160 10696 15936 10724
rect 15160 10684 15166 10696
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 16025 10727 16083 10733
rect 16025 10693 16037 10727
rect 16071 10724 16083 10727
rect 16850 10724 16856 10736
rect 16071 10696 16856 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 18230 10684 18236 10736
rect 18288 10684 18294 10736
rect 20254 10684 20260 10736
rect 20312 10684 20318 10736
rect 21634 10684 21640 10736
rect 21692 10684 21698 10736
rect 21744 10724 21772 10764
rect 21821 10761 21833 10795
rect 21867 10792 21879 10795
rect 22186 10792 22192 10804
rect 21867 10764 22192 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 22186 10752 22192 10764
rect 22244 10752 22250 10804
rect 22373 10795 22431 10801
rect 22373 10761 22385 10795
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 22388 10724 22416 10755
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22557 10795 22615 10801
rect 22557 10792 22569 10795
rect 22520 10764 22569 10792
rect 22520 10752 22526 10764
rect 22557 10761 22569 10764
rect 22603 10761 22615 10795
rect 22557 10755 22615 10761
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25314 10792 25320 10804
rect 24912 10764 25320 10792
rect 24912 10752 24918 10764
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 25682 10752 25688 10804
rect 25740 10752 25746 10804
rect 27614 10752 27620 10804
rect 27672 10792 27678 10804
rect 28074 10792 28080 10804
rect 27672 10764 28080 10792
rect 27672 10752 27678 10764
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 28261 10795 28319 10801
rect 28261 10792 28273 10795
rect 28224 10764 28273 10792
rect 28224 10752 28230 10764
rect 28261 10761 28273 10764
rect 28307 10792 28319 10795
rect 28350 10792 28356 10804
rect 28307 10764 28356 10792
rect 28307 10761 28319 10764
rect 28261 10755 28319 10761
rect 28350 10752 28356 10764
rect 28408 10752 28414 10804
rect 29362 10752 29368 10804
rect 29420 10801 29426 10804
rect 29420 10795 29439 10801
rect 29427 10761 29439 10795
rect 29420 10755 29439 10761
rect 29420 10752 29426 10755
rect 29546 10752 29552 10804
rect 29604 10792 29610 10804
rect 30009 10795 30067 10801
rect 30009 10792 30021 10795
rect 29604 10764 30021 10792
rect 29604 10752 29610 10764
rect 30009 10761 30021 10764
rect 30055 10761 30067 10795
rect 30009 10755 30067 10761
rect 30190 10752 30196 10804
rect 30248 10752 30254 10804
rect 30745 10795 30803 10801
rect 30745 10761 30757 10795
rect 30791 10792 30803 10795
rect 30791 10764 31800 10792
rect 30791 10761 30803 10764
rect 30745 10755 30803 10761
rect 25590 10724 25596 10736
rect 21744 10696 22416 10724
rect 24426 10696 25596 10724
rect 25590 10684 25596 10696
rect 25648 10684 25654 10736
rect 29178 10684 29184 10736
rect 29236 10684 29242 10736
rect 29638 10684 29644 10736
rect 29696 10724 29702 10736
rect 29914 10724 29920 10736
rect 29696 10696 29920 10724
rect 29696 10684 29702 10696
rect 29914 10684 29920 10696
rect 29972 10724 29978 10736
rect 30101 10727 30159 10733
rect 30101 10724 30113 10727
rect 29972 10696 30113 10724
rect 29972 10684 29978 10696
rect 30101 10693 30113 10696
rect 30147 10693 30159 10727
rect 30101 10687 30159 10693
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8478 10656 8484 10668
rect 8343 10628 8484 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 5460 10560 6040 10588
rect 5460 10529 5488 10560
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 4724 10492 5457 10520
rect 3418 10452 3424 10464
rect 3068 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4724 10452 4752 10492
rect 5445 10489 5457 10492
rect 5491 10489 5503 10523
rect 5445 10483 5503 10489
rect 5994 10480 6000 10532
rect 6052 10520 6058 10532
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 6052 10492 6745 10520
rect 6052 10480 6058 10492
rect 6733 10489 6745 10492
rect 6779 10520 6791 10523
rect 7469 10523 7527 10529
rect 7469 10520 7481 10523
rect 6779 10492 7481 10520
rect 6779 10489 6791 10492
rect 6733 10483 6791 10489
rect 7469 10489 7481 10492
rect 7515 10520 7527 10523
rect 7834 10520 7840 10532
rect 7515 10492 7840 10520
rect 7515 10489 7527 10492
rect 7469 10483 7527 10489
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 8036 10520 8064 10619
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8588 10588 8616 10619
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 8159 10560 8616 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8662 10548 8668 10600
rect 8720 10548 8726 10600
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 10244 10588 10272 10684
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 8987 10560 10272 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 8036 10492 8432 10520
rect 8404 10464 8432 10492
rect 4028 10424 4752 10452
rect 4028 10412 4034 10424
rect 5074 10412 5080 10464
rect 5132 10412 5138 10464
rect 5810 10412 5816 10464
rect 5868 10412 5874 10464
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 8938 10452 8944 10464
rect 8536 10424 8944 10452
rect 8536 10412 8542 10424
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 10410 10412 10416 10464
rect 10468 10412 10474 10464
rect 10520 10452 10548 10619
rect 10704 10520 10732 10619
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10836 10560 10885 10588
rect 10836 10548 10842 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 11606 10588 11612 10600
rect 10873 10551 10931 10557
rect 10980 10560 11612 10588
rect 10980 10520 11008 10560
rect 11606 10548 11612 10560
rect 11664 10588 11670 10600
rect 11790 10588 11796 10600
rect 11664 10560 11796 10588
rect 11664 10548 11670 10560
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 10704 10492 11008 10520
rect 12728 10464 12756 10619
rect 11882 10452 11888 10464
rect 10520 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 12710 10412 12716 10464
rect 12768 10412 12774 10464
rect 12802 10412 12808 10464
rect 12860 10412 12866 10464
rect 12912 10452 12940 10619
rect 12986 10616 12992 10668
rect 13044 10616 13050 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 15746 10656 15752 10668
rect 15243 10628 15752 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13354 10588 13360 10600
rect 13311 10560 13360 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13630 10548 13636 10600
rect 13688 10588 13694 10600
rect 15212 10588 15240 10619
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 16761 10659 16819 10665
rect 16761 10625 16773 10659
rect 16807 10625 16819 10659
rect 16761 10619 16819 10625
rect 13688 10560 15240 10588
rect 16485 10591 16543 10597
rect 13688 10548 13694 10560
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16776 10588 16804 10619
rect 19518 10616 19524 10668
rect 19576 10616 19582 10668
rect 21910 10616 21916 10668
rect 21968 10616 21974 10668
rect 22462 10616 22468 10668
rect 22520 10616 22526 10668
rect 25038 10616 25044 10668
rect 25096 10616 25102 10668
rect 25958 10616 25964 10668
rect 26016 10656 26022 10668
rect 26142 10656 26148 10668
rect 26016 10628 26148 10656
rect 26016 10616 26022 10628
rect 26142 10616 26148 10628
rect 26200 10656 26206 10668
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 26200 10628 26341 10656
rect 26200 10616 26206 10628
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 27706 10616 27712 10668
rect 27764 10616 27770 10668
rect 28258 10616 28264 10668
rect 28316 10616 28322 10668
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10656 28687 10659
rect 29270 10656 29276 10668
rect 28675 10628 29276 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 16531 10560 16804 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 17184 10560 17233 10588
rect 17184 10548 17190 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 15712 10492 16313 10520
rect 15712 10480 15718 10492
rect 16301 10489 16313 10492
rect 16347 10489 16359 10523
rect 16301 10483 16359 10489
rect 13998 10452 14004 10464
rect 12912 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10452 14062 10464
rect 14550 10452 14556 10464
rect 14056 10424 14556 10452
rect 14056 10412 14062 10424
rect 14550 10412 14556 10424
rect 14608 10452 14614 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14608 10424 14749 10452
rect 14608 10412 14614 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 15838 10412 15844 10464
rect 15896 10412 15902 10464
rect 16574 10412 16580 10464
rect 16632 10412 16638 10464
rect 17236 10452 17264 10551
rect 17494 10548 17500 10600
rect 17552 10548 17558 10600
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10557 19211 10591
rect 22925 10591 22983 10597
rect 19153 10551 19211 10557
rect 21192 10560 21864 10588
rect 19168 10452 19196 10551
rect 21192 10464 21220 10560
rect 21269 10523 21327 10529
rect 21269 10489 21281 10523
rect 21315 10489 21327 10523
rect 21836 10520 21864 10560
rect 22925 10557 22937 10591
rect 22971 10557 22983 10591
rect 22925 10551 22983 10557
rect 22189 10523 22247 10529
rect 22189 10520 22201 10523
rect 21836 10492 22201 10520
rect 21269 10483 21327 10489
rect 22189 10489 22201 10492
rect 22235 10489 22247 10523
rect 22189 10483 22247 10489
rect 17236 10424 19196 10452
rect 19978 10412 19984 10464
rect 20036 10452 20042 10464
rect 20806 10452 20812 10464
rect 20036 10424 20812 10452
rect 20036 10412 20042 10424
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 20901 10455 20959 10461
rect 20901 10421 20913 10455
rect 20947 10452 20959 10455
rect 21174 10452 21180 10464
rect 20947 10424 21180 10452
rect 20947 10421 20959 10424
rect 20901 10415 20959 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21284 10452 21312 10483
rect 21542 10452 21548 10464
rect 21284 10424 21548 10452
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 21637 10455 21695 10461
rect 21637 10421 21649 10455
rect 21683 10452 21695 10455
rect 22002 10452 22008 10464
rect 21683 10424 22008 10452
rect 21683 10421 21695 10424
rect 21637 10415 21695 10421
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 22940 10452 22968 10551
rect 23198 10548 23204 10600
rect 23256 10548 23262 10600
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 23992 10560 24685 10588
rect 23992 10548 23998 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 25590 10548 25596 10600
rect 25648 10588 25654 10600
rect 25976 10588 26004 10616
rect 25648 10560 26004 10588
rect 26605 10591 26663 10597
rect 25648 10548 25654 10560
rect 26605 10557 26617 10591
rect 26651 10588 26663 10591
rect 28644 10588 28672 10619
rect 29270 10616 29276 10628
rect 29328 10616 29334 10668
rect 29730 10616 29736 10668
rect 29788 10616 29794 10668
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10656 29883 10659
rect 30208 10656 30236 10752
rect 29871 10628 30236 10656
rect 30331 10693 30389 10699
rect 30331 10659 30343 10693
rect 30377 10659 30389 10693
rect 30926 10684 30932 10736
rect 30984 10724 30990 10736
rect 31662 10724 31668 10736
rect 30984 10696 31156 10724
rect 30984 10684 30990 10696
rect 30331 10656 30389 10659
rect 30466 10656 30472 10668
rect 30331 10653 30472 10656
rect 30332 10628 30472 10653
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 30466 10616 30472 10628
rect 30524 10656 30530 10668
rect 30834 10656 30840 10668
rect 30524 10628 30840 10656
rect 30524 10616 30530 10628
rect 30834 10616 30840 10628
rect 30892 10616 30898 10668
rect 31128 10665 31156 10696
rect 31220 10696 31668 10724
rect 31113 10659 31171 10665
rect 31113 10625 31125 10659
rect 31159 10625 31171 10659
rect 31113 10619 31171 10625
rect 26651 10560 28672 10588
rect 26651 10557 26663 10560
rect 26605 10551 26663 10557
rect 30282 10548 30288 10600
rect 30340 10588 30346 10600
rect 31220 10597 31248 10696
rect 31662 10684 31668 10696
rect 31720 10684 31726 10736
rect 31772 10733 31800 10764
rect 32582 10752 32588 10804
rect 32640 10792 32646 10804
rect 34422 10792 34428 10804
rect 32640 10764 33088 10792
rect 32640 10752 32646 10764
rect 31757 10727 31815 10733
rect 31757 10693 31769 10727
rect 31803 10693 31815 10727
rect 33060 10724 33088 10764
rect 32982 10696 33088 10724
rect 31757 10687 31815 10693
rect 31478 10616 31484 10668
rect 31536 10616 31542 10668
rect 30929 10591 30987 10597
rect 30340 10560 30788 10588
rect 30340 10548 30346 10560
rect 28258 10480 28264 10532
rect 28316 10520 28322 10532
rect 29270 10520 29276 10532
rect 28316 10492 29276 10520
rect 28316 10480 28322 10492
rect 29270 10480 29276 10492
rect 29328 10480 29334 10532
rect 29822 10520 29828 10532
rect 29380 10492 29828 10520
rect 23934 10452 23940 10464
rect 22940 10424 23940 10452
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24854 10412 24860 10464
rect 24912 10412 24918 10464
rect 25774 10412 25780 10464
rect 25832 10452 25838 10464
rect 26053 10455 26111 10461
rect 26053 10452 26065 10455
rect 25832 10424 26065 10452
rect 25832 10412 25838 10424
rect 26053 10421 26065 10424
rect 26099 10421 26111 10455
rect 26053 10415 26111 10421
rect 28074 10412 28080 10464
rect 28132 10412 28138 10464
rect 29380 10461 29408 10492
rect 29822 10480 29828 10492
rect 29880 10520 29886 10532
rect 30760 10520 30788 10560
rect 30929 10557 30941 10591
rect 30975 10557 30987 10591
rect 30929 10551 30987 10557
rect 31021 10591 31079 10597
rect 31021 10557 31033 10591
rect 31067 10557 31079 10591
rect 31021 10551 31079 10557
rect 31205 10591 31263 10597
rect 31205 10557 31217 10591
rect 31251 10557 31263 10591
rect 32490 10588 32496 10600
rect 31205 10551 31263 10557
rect 31588 10560 32496 10588
rect 30944 10520 30972 10551
rect 29880 10492 30328 10520
rect 30760 10492 30972 10520
rect 31036 10520 31064 10551
rect 31588 10520 31616 10560
rect 32490 10548 32496 10560
rect 32548 10588 32554 10600
rect 33060 10588 33088 10696
rect 33336 10764 34428 10792
rect 33336 10665 33364 10764
rect 34422 10752 34428 10764
rect 34480 10752 34486 10804
rect 34514 10752 34520 10804
rect 34572 10792 34578 10804
rect 35069 10795 35127 10801
rect 35069 10792 35081 10795
rect 34572 10764 35081 10792
rect 34572 10752 34578 10764
rect 33597 10727 33655 10733
rect 33597 10693 33609 10727
rect 33643 10724 33655 10727
rect 33870 10724 33876 10736
rect 33643 10696 33876 10724
rect 33643 10693 33655 10696
rect 33597 10687 33655 10693
rect 33870 10684 33876 10696
rect 33928 10684 33934 10736
rect 33321 10659 33379 10665
rect 33321 10625 33333 10659
rect 33367 10625 33379 10659
rect 34900 10656 34928 10764
rect 35069 10761 35081 10764
rect 35115 10761 35127 10795
rect 35069 10755 35127 10761
rect 35529 10795 35587 10801
rect 35529 10761 35541 10795
rect 35575 10792 35587 10795
rect 35986 10792 35992 10804
rect 35575 10764 35992 10792
rect 35575 10761 35587 10764
rect 35529 10755 35587 10761
rect 35986 10752 35992 10764
rect 36044 10752 36050 10804
rect 36446 10752 36452 10804
rect 36504 10752 36510 10804
rect 36633 10795 36691 10801
rect 36633 10761 36645 10795
rect 36679 10761 36691 10795
rect 36633 10755 36691 10761
rect 34974 10684 34980 10736
rect 35032 10724 35038 10736
rect 36648 10724 36676 10755
rect 37458 10752 37464 10804
rect 37516 10752 37522 10804
rect 37553 10795 37611 10801
rect 37553 10761 37565 10795
rect 37599 10792 37611 10795
rect 37599 10764 38148 10792
rect 37599 10761 37611 10764
rect 37553 10755 37611 10761
rect 37093 10727 37151 10733
rect 37093 10724 37105 10727
rect 35032 10696 36676 10724
rect 36740 10696 37105 10724
rect 35032 10684 35038 10696
rect 35989 10659 36047 10665
rect 35989 10656 36001 10659
rect 33321 10619 33379 10625
rect 34716 10588 34744 10642
rect 34900 10628 36001 10656
rect 35989 10625 36001 10628
rect 36035 10625 36047 10659
rect 35989 10619 36047 10625
rect 36262 10616 36268 10668
rect 36320 10616 36326 10668
rect 36538 10616 36544 10668
rect 36596 10656 36602 10668
rect 36740 10656 36768 10696
rect 37093 10693 37105 10696
rect 37139 10693 37151 10727
rect 37093 10687 37151 10693
rect 36596 10628 36768 10656
rect 36817 10659 36875 10665
rect 36596 10616 36602 10628
rect 36817 10625 36829 10659
rect 36863 10625 36875 10659
rect 36817 10619 36875 10625
rect 34882 10588 34888 10600
rect 32548 10560 32812 10588
rect 33060 10560 34888 10588
rect 32548 10548 32554 10560
rect 31036 10492 31616 10520
rect 32784 10520 32812 10560
rect 34882 10548 34888 10560
rect 34940 10548 34946 10600
rect 35618 10548 35624 10600
rect 35676 10548 35682 10600
rect 35710 10548 35716 10600
rect 35768 10548 35774 10600
rect 35802 10548 35808 10600
rect 35860 10588 35866 10600
rect 36081 10591 36139 10597
rect 36081 10588 36093 10591
rect 35860 10560 36093 10588
rect 35860 10548 35866 10560
rect 36081 10557 36093 10560
rect 36127 10557 36139 10591
rect 36081 10551 36139 10557
rect 33229 10523 33287 10529
rect 33229 10520 33241 10523
rect 32784 10492 33241 10520
rect 29880 10480 29886 10492
rect 29365 10455 29423 10461
rect 29365 10421 29377 10455
rect 29411 10421 29423 10455
rect 29365 10415 29423 10421
rect 29549 10455 29607 10461
rect 29549 10421 29561 10455
rect 29595 10452 29607 10455
rect 29638 10452 29644 10464
rect 29595 10424 29644 10452
rect 29595 10421 29607 10424
rect 29549 10415 29607 10421
rect 29638 10412 29644 10424
rect 29696 10412 29702 10464
rect 30300 10461 30328 10492
rect 33229 10489 33241 10492
rect 33275 10489 33287 10523
rect 33229 10483 33287 10489
rect 35161 10523 35219 10529
rect 35161 10489 35173 10523
rect 35207 10520 35219 10523
rect 36832 10520 36860 10619
rect 37108 10600 37136 10687
rect 37476 10656 37504 10752
rect 38120 10733 38148 10764
rect 38746 10752 38752 10804
rect 38804 10792 38810 10804
rect 39577 10795 39635 10801
rect 39577 10792 39589 10795
rect 38804 10764 39589 10792
rect 38804 10752 38810 10764
rect 39577 10761 39589 10764
rect 39623 10792 39635 10795
rect 39758 10792 39764 10804
rect 39623 10764 39764 10792
rect 39623 10761 39635 10764
rect 39577 10755 39635 10761
rect 39758 10752 39764 10764
rect 39816 10752 39822 10804
rect 40328 10764 41092 10792
rect 38105 10727 38163 10733
rect 38105 10693 38117 10727
rect 38151 10693 38163 10727
rect 39942 10724 39948 10736
rect 38105 10687 38163 10693
rect 39684 10696 39948 10724
rect 37737 10659 37795 10665
rect 37737 10656 37749 10659
rect 37476 10628 37749 10656
rect 37737 10625 37749 10628
rect 37783 10625 37795 10659
rect 37737 10619 37795 10625
rect 39206 10616 39212 10668
rect 39264 10656 39270 10668
rect 39684 10656 39712 10696
rect 39942 10684 39948 10696
rect 40000 10724 40006 10736
rect 40328 10724 40356 10764
rect 40000 10696 40434 10724
rect 40000 10684 40006 10696
rect 39264 10628 39712 10656
rect 39264 10616 39270 10628
rect 37090 10548 37096 10600
rect 37148 10588 37154 10600
rect 37829 10591 37887 10597
rect 37829 10588 37841 10591
rect 37148 10560 37841 10588
rect 37148 10548 37154 10560
rect 37829 10557 37841 10560
rect 37875 10557 37887 10591
rect 37829 10551 37887 10557
rect 39666 10548 39672 10600
rect 39724 10548 39730 10600
rect 39942 10548 39948 10600
rect 40000 10548 40006 10600
rect 41064 10588 41092 10764
rect 41414 10752 41420 10804
rect 41472 10752 41478 10804
rect 42334 10752 42340 10804
rect 42392 10792 42398 10804
rect 43073 10795 43131 10801
rect 43073 10792 43085 10795
rect 42392 10764 43085 10792
rect 42392 10752 42398 10764
rect 43073 10761 43085 10764
rect 43119 10792 43131 10795
rect 43254 10792 43260 10804
rect 43119 10764 43260 10792
rect 43119 10761 43131 10764
rect 43073 10755 43131 10761
rect 43254 10752 43260 10764
rect 43312 10752 43318 10804
rect 43809 10795 43867 10801
rect 43809 10761 43821 10795
rect 43855 10792 43867 10795
rect 44266 10792 44272 10804
rect 43855 10764 44272 10792
rect 43855 10761 43867 10764
rect 43809 10755 43867 10761
rect 44266 10752 44272 10764
rect 44324 10752 44330 10804
rect 44542 10752 44548 10804
rect 44600 10752 44606 10804
rect 42705 10727 42763 10733
rect 42705 10693 42717 10727
rect 42751 10724 42763 10727
rect 42978 10724 42984 10736
rect 42751 10696 42984 10724
rect 42751 10693 42763 10696
rect 42705 10687 42763 10693
rect 42978 10684 42984 10696
rect 43036 10724 43042 10736
rect 43441 10727 43499 10733
rect 43441 10724 43453 10727
rect 43036 10696 43453 10724
rect 43036 10684 43042 10696
rect 43441 10693 43453 10696
rect 43487 10724 43499 10727
rect 44177 10727 44235 10733
rect 44177 10724 44189 10727
rect 43487 10696 44189 10724
rect 43487 10693 43499 10696
rect 43441 10687 43499 10693
rect 44177 10693 44189 10696
rect 44223 10724 44235 10727
rect 44560 10724 44588 10752
rect 44223 10696 44588 10724
rect 44223 10693 44235 10696
rect 44177 10687 44235 10693
rect 41966 10616 41972 10668
rect 42024 10616 42030 10668
rect 41782 10588 41788 10600
rect 41064 10560 41788 10588
rect 41782 10548 41788 10560
rect 41840 10588 41846 10600
rect 42518 10588 42524 10600
rect 41840 10560 42524 10588
rect 41840 10548 41846 10560
rect 42518 10548 42524 10560
rect 42576 10548 42582 10600
rect 35207 10492 36860 10520
rect 35207 10489 35219 10492
rect 35161 10483 35219 10489
rect 30285 10455 30343 10461
rect 30285 10421 30297 10455
rect 30331 10421 30343 10455
rect 30285 10415 30343 10421
rect 30469 10455 30527 10461
rect 30469 10421 30481 10455
rect 30515 10452 30527 10455
rect 30558 10452 30564 10464
rect 30515 10424 30564 10452
rect 30515 10421 30527 10424
rect 30469 10415 30527 10421
rect 30558 10412 30564 10424
rect 30616 10412 30622 10464
rect 30742 10412 30748 10464
rect 30800 10452 30806 10464
rect 31478 10452 31484 10464
rect 30800 10424 31484 10452
rect 30800 10412 30806 10424
rect 31478 10412 31484 10424
rect 31536 10412 31542 10464
rect 32122 10412 32128 10464
rect 32180 10452 32186 10464
rect 35986 10452 35992 10464
rect 32180 10424 35992 10452
rect 32180 10412 32186 10424
rect 35986 10412 35992 10424
rect 36044 10412 36050 10464
rect 36078 10412 36084 10464
rect 36136 10412 36142 10464
rect 41782 10412 41788 10464
rect 41840 10412 41846 10464
rect 44545 10455 44603 10461
rect 44545 10421 44557 10455
rect 44591 10452 44603 10455
rect 44726 10452 44732 10464
rect 44591 10424 44732 10452
rect 44591 10421 44603 10424
rect 44545 10415 44603 10421
rect 44726 10412 44732 10424
rect 44784 10412 44790 10464
rect 44818 10412 44824 10464
rect 44876 10412 44882 10464
rect 460 10362 45540 10384
rect 460 10310 3570 10362
rect 3622 10310 3634 10362
rect 3686 10310 3698 10362
rect 3750 10310 3762 10362
rect 3814 10310 3826 10362
rect 3878 10310 8570 10362
rect 8622 10310 8634 10362
rect 8686 10310 8698 10362
rect 8750 10310 8762 10362
rect 8814 10310 8826 10362
rect 8878 10310 13570 10362
rect 13622 10310 13634 10362
rect 13686 10310 13698 10362
rect 13750 10310 13762 10362
rect 13814 10310 13826 10362
rect 13878 10310 18570 10362
rect 18622 10310 18634 10362
rect 18686 10310 18698 10362
rect 18750 10310 18762 10362
rect 18814 10310 18826 10362
rect 18878 10310 23570 10362
rect 23622 10310 23634 10362
rect 23686 10310 23698 10362
rect 23750 10310 23762 10362
rect 23814 10310 23826 10362
rect 23878 10310 28570 10362
rect 28622 10310 28634 10362
rect 28686 10310 28698 10362
rect 28750 10310 28762 10362
rect 28814 10310 28826 10362
rect 28878 10310 33570 10362
rect 33622 10310 33634 10362
rect 33686 10310 33698 10362
rect 33750 10310 33762 10362
rect 33814 10310 33826 10362
rect 33878 10310 38570 10362
rect 38622 10310 38634 10362
rect 38686 10310 38698 10362
rect 38750 10310 38762 10362
rect 38814 10310 38826 10362
rect 38878 10310 43570 10362
rect 43622 10310 43634 10362
rect 43686 10310 43698 10362
rect 43750 10310 43762 10362
rect 43814 10310 43826 10362
rect 43878 10310 45540 10362
rect 460 10288 45540 10310
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3384 10220 3433 10248
rect 3384 10208 3390 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3421 10211 3479 10217
rect 4338 10208 4344 10260
rect 4396 10208 4402 10260
rect 5534 10248 5540 10260
rect 4540 10220 5540 10248
rect 4356 10180 4384 10208
rect 3620 10152 4384 10180
rect 3620 10053 3648 10152
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10081 4215 10115
rect 4157 10075 4215 10081
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 3878 10044 3884 10056
rect 3835 10016 3884 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 3344 9976 3372 10007
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4080 9976 4108 10004
rect 3344 9948 4108 9976
rect 4172 9976 4200 10075
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4540 10053 4568 10220
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5810 10208 5816 10260
rect 5868 10208 5874 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 9732 10220 10057 10248
rect 9732 10208 9738 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10502 10248 10508 10260
rect 10275 10220 10508 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 11698 10208 11704 10260
rect 11756 10208 11762 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 11848 10220 12265 10248
rect 11848 10208 11854 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12253 10211 12311 10217
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12621 10251 12679 10257
rect 12621 10248 12633 10251
rect 12400 10220 12633 10248
rect 12400 10208 12406 10220
rect 12621 10217 12633 10220
rect 12667 10217 12679 10251
rect 12621 10211 12679 10217
rect 12802 10208 12808 10260
rect 12860 10208 12866 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 13412 10220 13461 10248
rect 13412 10208 13418 10220
rect 13449 10217 13461 10220
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 5828 10112 5856 10208
rect 4847 10084 5856 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6052 10084 6377 10112
rect 6052 10072 6058 10084
rect 6365 10081 6377 10084
rect 6411 10112 6423 10115
rect 7006 10112 7012 10124
rect 6411 10084 7012 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 9030 10112 9036 10124
rect 8312 10084 9036 10112
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4396 10016 4537 10044
rect 4396 10004 4402 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8312 10053 8340 10084
rect 9030 10072 9036 10084
rect 9088 10112 9094 10124
rect 10689 10115 10747 10121
rect 9088 10084 10456 10112
rect 9088 10072 9094 10084
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8076 10016 8309 10044
rect 8076 10004 8082 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 10042 10044 10048 10056
rect 9706 10016 10048 10044
rect 8297 10007 8355 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 10428 10053 10456 10084
rect 10689 10081 10701 10115
rect 10735 10112 10747 10115
rect 11716 10112 11744 10208
rect 12158 10140 12164 10192
rect 12216 10140 12222 10192
rect 12176 10112 12204 10140
rect 10735 10084 11744 10112
rect 11808 10084 12204 10112
rect 12820 10112 12848 10208
rect 12989 10183 13047 10189
rect 12989 10149 13001 10183
rect 13035 10180 13047 10183
rect 13078 10180 13084 10192
rect 13035 10152 13084 10180
rect 13035 10149 13047 10152
rect 12989 10143 13047 10149
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 14016 10180 14044 10211
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14148 10220 14289 10248
rect 14148 10208 14154 10220
rect 14277 10217 14289 10220
rect 14323 10248 14335 10251
rect 14458 10248 14464 10260
rect 14323 10220 14464 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15102 10208 15108 10260
rect 15160 10208 15166 10260
rect 16574 10208 16580 10260
rect 16632 10208 16638 10260
rect 17402 10208 17408 10260
rect 17460 10208 17466 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17552 10220 17693 10248
rect 17552 10208 17558 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 19242 10248 19248 10260
rect 18104 10220 19248 10248
rect 18104 10208 18110 10220
rect 15120 10180 15148 10208
rect 13228 10152 13860 10180
rect 14016 10152 15148 10180
rect 13228 10140 13234 10152
rect 13832 10112 13860 10152
rect 14366 10112 14372 10124
rect 12820 10084 13768 10112
rect 13832 10084 14372 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10013 10471 10047
rect 11808 10030 11836 10084
rect 10413 10007 10471 10013
rect 5074 9976 5080 9988
rect 4172 9948 5080 9976
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 6641 9979 6699 9985
rect 6026 9948 6592 9976
rect 6564 9920 6592 9948
rect 6641 9945 6653 9979
rect 6687 9976 6699 9979
rect 6914 9976 6920 9988
rect 6687 9948 6920 9976
rect 6687 9945 6699 9948
rect 6641 9939 6699 9945
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 8573 9979 8631 9985
rect 8573 9976 8585 9979
rect 8536 9948 8585 9976
rect 8536 9936 8542 9948
rect 8573 9945 8585 9948
rect 8619 9945 8631 9979
rect 10428 9976 10456 10007
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12032 10016 12265 10044
rect 12032 10004 12038 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 10778 9976 10784 9988
rect 10428 9948 10784 9976
rect 8573 9939 8631 9945
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 12360 9976 12388 10007
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 13170 10044 13176 10056
rect 13044 10016 13176 10044
rect 13044 10004 13050 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13740 10053 13768 10084
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 15381 10115 15439 10121
rect 15381 10081 15393 10115
rect 15427 10112 15439 10115
rect 16592 10112 16620 10208
rect 17420 10180 17448 10208
rect 15427 10084 16620 10112
rect 17236 10152 17448 10180
rect 15427 10081 15439 10084
rect 15381 10075 15439 10081
rect 17236 10056 17264 10152
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10044 13875 10047
rect 14274 10044 14280 10056
rect 13863 10016 14280 10044
rect 13863 10013 13875 10016
rect 13817 10007 13875 10013
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16724 10016 17141 10044
rect 16724 10004 16730 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17218 10004 17224 10056
rect 17276 10004 17282 10056
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17770 10044 17776 10056
rect 17543 10016 17776 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 12176 9948 12388 9976
rect 13449 9979 13507 9985
rect 3789 9911 3847 9917
rect 3789 9877 3801 9911
rect 3835 9908 3847 9911
rect 4154 9908 4160 9920
rect 3835 9880 4160 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6178 9908 6184 9920
rect 5776 9880 6184 9908
rect 5776 9868 5782 9880
rect 6178 9868 6184 9880
rect 6236 9908 6242 9920
rect 6273 9911 6331 9917
rect 6273 9908 6285 9911
rect 6236 9880 6285 9908
rect 6236 9868 6242 9880
rect 6273 9877 6285 9880
rect 6319 9877 6331 9911
rect 6273 9871 6331 9877
rect 6546 9868 6552 9920
rect 6604 9868 6610 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8386 9908 8392 9920
rect 8159 9880 8392 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8386 9868 8392 9880
rect 8444 9908 8450 9920
rect 9582 9908 9588 9920
rect 8444 9880 9588 9908
rect 8444 9868 8450 9880
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 12176 9917 12204 9948
rect 13449 9945 13461 9979
rect 13495 9976 13507 9979
rect 14090 9976 14096 9988
rect 13495 9948 14096 9976
rect 13495 9945 13507 9948
rect 13449 9939 13507 9945
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 14369 9979 14427 9985
rect 14369 9976 14381 9979
rect 14240 9948 14381 9976
rect 14240 9936 14246 9948
rect 14369 9945 14381 9948
rect 14415 9945 14427 9979
rect 15838 9976 15844 9988
rect 14369 9939 14427 9945
rect 15028 9948 15844 9976
rect 15028 9920 15056 9948
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 11572 9880 12173 9908
rect 11572 9868 11578 9880
rect 12161 9877 12173 9880
rect 12207 9877 12219 9911
rect 12161 9871 12219 9877
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12768 9880 13185 9908
rect 12768 9868 12774 9880
rect 13173 9877 13185 9880
rect 13219 9908 13231 9911
rect 13538 9908 13544 9920
rect 13219 9880 13544 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13906 9908 13912 9920
rect 13679 9880 13912 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13906 9868 13912 9880
rect 13964 9908 13970 9920
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 13964 9880 14749 9908
rect 13964 9868 13970 9880
rect 14737 9877 14749 9880
rect 14783 9877 14795 9911
rect 14737 9871 14795 9877
rect 15010 9868 15016 9920
rect 15068 9868 15074 9920
rect 15764 9908 15792 9948
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 17512 9976 17540 10007
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18156 10053 18184 10220
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 20165 10251 20223 10257
rect 20165 10217 20177 10251
rect 20211 10217 20223 10251
rect 20165 10211 20223 10217
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 20622 10248 20628 10260
rect 20395 10220 20628 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 19610 10180 19616 10192
rect 18340 10152 19616 10180
rect 18340 10053 18368 10152
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 20180 10180 20208 10211
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 20898 10248 20904 10260
rect 20732 10220 20904 10248
rect 20441 10183 20499 10189
rect 20180 10152 20408 10180
rect 18966 10072 18972 10124
rect 19024 10112 19030 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 19024 10084 19257 10112
rect 19024 10072 19030 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 20162 10112 20168 10124
rect 19245 10075 19303 10081
rect 19536 10084 20168 10112
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 16776 9948 17540 9976
rect 17880 9976 17908 10007
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18874 10004 18880 10056
rect 18932 10044 18938 10056
rect 19536 10053 19564 10084
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 20380 10112 20408 10152
rect 20441 10149 20453 10183
rect 20487 10180 20499 10183
rect 20732 10180 20760 10220
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 22462 10248 22468 10260
rect 21315 10220 22468 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 23017 10251 23075 10257
rect 23017 10217 23029 10251
rect 23063 10248 23075 10251
rect 23198 10248 23204 10260
rect 23063 10220 23204 10248
rect 23063 10217 23075 10220
rect 23017 10211 23075 10217
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 24286 10251 24344 10257
rect 24286 10248 24298 10251
rect 23348 10220 24298 10248
rect 23348 10208 23354 10220
rect 24286 10217 24298 10220
rect 24332 10217 24344 10251
rect 24286 10211 24344 10217
rect 24854 10208 24860 10260
rect 24912 10248 24918 10260
rect 24912 10220 25728 10248
rect 24912 10208 24918 10220
rect 22002 10180 22008 10192
rect 20487 10152 20760 10180
rect 20916 10152 22008 10180
rect 20487 10149 20499 10152
rect 20441 10143 20499 10149
rect 20916 10112 20944 10152
rect 22002 10140 22008 10152
rect 22060 10140 22066 10192
rect 22664 10152 23980 10180
rect 20380 10084 20944 10112
rect 19061 10047 19119 10053
rect 19061 10044 19073 10047
rect 18932 10016 19073 10044
rect 18932 10004 18938 10016
rect 19061 10013 19073 10016
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10044 19855 10047
rect 20167 10044 20195 10072
rect 20622 10044 20628 10056
rect 19843 10016 20116 10044
rect 20167 10016 20628 10044
rect 19843 10013 19855 10016
rect 19797 10007 19855 10013
rect 17880 9948 18736 9976
rect 16776 9908 16804 9948
rect 15764 9880 16804 9908
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 18708 9917 18736 9948
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9877 18751 9911
rect 18693 9871 18751 9877
rect 19153 9911 19211 9917
rect 19153 9877 19165 9911
rect 19199 9908 19211 9911
rect 19426 9908 19432 9920
rect 19199 9880 19432 9908
rect 19199 9877 19211 9880
rect 19153 9871 19211 9877
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 20088 9908 20116 10016
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 20916 10053 20944 10084
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 20162 9936 20168 9988
rect 20220 9976 20226 9988
rect 21008 9976 21036 10075
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21634 10112 21640 10124
rect 21140 10084 21640 10112
rect 21140 10072 21146 10084
rect 21634 10072 21640 10084
rect 21692 10112 21698 10124
rect 21821 10115 21879 10121
rect 21821 10112 21833 10115
rect 21692 10084 21833 10112
rect 21692 10072 21698 10084
rect 21821 10081 21833 10084
rect 21867 10081 21879 10115
rect 21821 10075 21879 10081
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 21450 10044 21456 10056
rect 21232 10016 21456 10044
rect 21232 10004 21238 10016
rect 21450 10004 21456 10016
rect 21508 10044 21514 10056
rect 22097 10047 22155 10053
rect 22097 10044 22109 10047
rect 21508 10016 22109 10044
rect 21508 10004 21514 10016
rect 21542 9976 21548 9988
rect 20220 9948 21036 9976
rect 21100 9948 21548 9976
rect 20220 9936 20226 9948
rect 20809 9911 20867 9917
rect 20809 9908 20821 9911
rect 20088 9880 20821 9908
rect 20809 9877 20821 9880
rect 20855 9908 20867 9911
rect 21100 9908 21128 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 21652 9985 21680 10016
rect 22097 10013 22109 10016
rect 22143 10013 22155 10047
rect 22097 10007 22155 10013
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10044 22339 10047
rect 22327 10016 22508 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 21637 9979 21695 9985
rect 21637 9945 21649 9979
rect 21683 9945 21695 9979
rect 22112 9976 22140 10007
rect 22480 9976 22508 10016
rect 22554 10004 22560 10056
rect 22612 10004 22618 10056
rect 22664 10053 22692 10152
rect 22830 10072 22836 10124
rect 22888 10072 22894 10124
rect 23382 10112 23388 10124
rect 23308 10084 23388 10112
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22922 10044 22928 10056
rect 22649 10007 22707 10013
rect 22756 10016 22928 10044
rect 22756 9976 22784 10016
rect 22922 10004 22928 10016
rect 22980 10044 22986 10056
rect 22980 10016 23060 10044
rect 22980 10004 22986 10016
rect 22112 9948 22324 9976
rect 22480 9948 22784 9976
rect 23032 9976 23060 10016
rect 23198 10004 23204 10056
rect 23256 10004 23262 10056
rect 23308 10053 23336 10084
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 23477 10115 23535 10121
rect 23477 10081 23489 10115
rect 23523 10112 23535 10115
rect 23845 10115 23903 10121
rect 23845 10112 23857 10115
rect 23523 10084 23857 10112
rect 23523 10081 23535 10084
rect 23477 10075 23535 10081
rect 23845 10081 23857 10084
rect 23891 10081 23903 10115
rect 23952 10112 23980 10152
rect 25406 10140 25412 10192
rect 25464 10140 25470 10192
rect 24302 10112 24308 10124
rect 23952 10084 24308 10112
rect 23845 10075 23903 10081
rect 24302 10072 24308 10084
rect 24360 10112 24366 10124
rect 25424 10112 25452 10140
rect 25700 10112 25728 10220
rect 28442 10208 28448 10260
rect 28500 10248 28506 10260
rect 28537 10251 28595 10257
rect 28537 10248 28549 10251
rect 28500 10220 28549 10248
rect 28500 10208 28506 10220
rect 28537 10217 28549 10220
rect 28583 10217 28595 10251
rect 28537 10211 28595 10217
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 29086 10248 29092 10260
rect 29043 10220 29092 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29086 10208 29092 10220
rect 29144 10248 29150 10260
rect 29144 10220 30052 10248
rect 29144 10208 29150 10220
rect 29733 10183 29791 10189
rect 29733 10180 29745 10183
rect 28276 10152 29745 10180
rect 28276 10124 28304 10152
rect 29733 10149 29745 10152
rect 29779 10149 29791 10183
rect 29733 10143 29791 10149
rect 26421 10115 26479 10121
rect 26421 10112 26433 10115
rect 24360 10084 25544 10112
rect 25700 10084 26433 10112
rect 24360 10072 24366 10084
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10013 23351 10047
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 23293 10007 23351 10013
rect 23408 10016 23581 10044
rect 23408 9976 23436 10016
rect 23569 10013 23581 10016
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23750 10004 23756 10056
rect 23808 10004 23814 10056
rect 24026 10004 24032 10056
rect 24084 10004 24090 10056
rect 25516 10044 25544 10084
rect 26421 10081 26433 10084
rect 26467 10081 26479 10115
rect 26421 10075 26479 10081
rect 28258 10072 28264 10124
rect 28316 10072 28322 10124
rect 28534 10072 28540 10124
rect 28592 10112 28598 10124
rect 28721 10115 28779 10121
rect 28721 10112 28733 10115
rect 28592 10084 28733 10112
rect 28592 10072 28598 10084
rect 28721 10081 28733 10084
rect 28767 10081 28779 10115
rect 29914 10112 29920 10124
rect 28721 10075 28779 10081
rect 29104 10084 29920 10112
rect 26053 10047 26111 10053
rect 26053 10044 26065 10047
rect 25516 10016 26065 10044
rect 26053 10013 26065 10016
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 26142 10004 26148 10056
rect 26200 10004 26206 10056
rect 27706 10044 27712 10056
rect 27554 10016 27712 10044
rect 27706 10004 27712 10016
rect 27764 10044 27770 10056
rect 28350 10044 28356 10056
rect 27764 10016 28356 10044
rect 27764 10004 27770 10016
rect 28350 10004 28356 10016
rect 28408 10004 28414 10056
rect 28445 10047 28503 10053
rect 28445 10013 28457 10047
rect 28491 10044 28503 10047
rect 29104 10044 29132 10084
rect 28491 10016 29132 10044
rect 29181 10047 29239 10053
rect 28491 10013 28503 10016
rect 28445 10007 28503 10013
rect 29181 10013 29193 10047
rect 29227 10044 29239 10047
rect 29362 10044 29368 10056
rect 29227 10016 29368 10044
rect 29227 10013 29239 10016
rect 29181 10007 29239 10013
rect 29362 10004 29368 10016
rect 29420 10004 29426 10056
rect 29472 10053 29500 10084
rect 29914 10072 29920 10084
rect 29972 10072 29978 10124
rect 30024 10112 30052 10220
rect 30650 10208 30656 10260
rect 30708 10248 30714 10260
rect 33042 10248 33048 10260
rect 30708 10220 33048 10248
rect 30708 10208 30714 10220
rect 33042 10208 33048 10220
rect 33100 10208 33106 10260
rect 33134 10208 33140 10260
rect 33192 10208 33198 10260
rect 33226 10208 33232 10260
rect 33284 10248 33290 10260
rect 33597 10251 33655 10257
rect 33597 10248 33609 10251
rect 33284 10220 33609 10248
rect 33284 10208 33290 10220
rect 33597 10217 33609 10220
rect 33643 10248 33655 10251
rect 34054 10248 34060 10260
rect 33643 10220 34060 10248
rect 33643 10217 33655 10220
rect 33597 10211 33655 10217
rect 34054 10208 34060 10220
rect 34112 10208 34118 10260
rect 34330 10208 34336 10260
rect 34388 10248 34394 10260
rect 35802 10248 35808 10260
rect 34388 10220 35808 10248
rect 34388 10208 34394 10220
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 35894 10208 35900 10260
rect 35952 10208 35958 10260
rect 35986 10208 35992 10260
rect 36044 10248 36050 10260
rect 36538 10248 36544 10260
rect 36044 10220 36544 10248
rect 36044 10208 36050 10220
rect 36538 10208 36544 10220
rect 36596 10208 36602 10260
rect 38378 10208 38384 10260
rect 38436 10208 38442 10260
rect 38841 10251 38899 10257
rect 38841 10217 38853 10251
rect 38887 10248 38899 10251
rect 39942 10248 39948 10260
rect 38887 10220 39948 10248
rect 38887 10217 38899 10220
rect 38841 10211 38899 10217
rect 39942 10208 39948 10220
rect 40000 10208 40006 10260
rect 41782 10208 41788 10260
rect 41840 10208 41846 10260
rect 41874 10208 41880 10260
rect 41932 10248 41938 10260
rect 42245 10251 42303 10257
rect 42245 10248 42257 10251
rect 41932 10220 42257 10248
rect 41932 10208 41938 10220
rect 42245 10217 42257 10220
rect 42291 10217 42303 10251
rect 42245 10211 42303 10217
rect 42613 10251 42671 10257
rect 42613 10217 42625 10251
rect 42659 10248 42671 10251
rect 42978 10248 42984 10260
rect 42659 10220 42984 10248
rect 42659 10217 42671 10220
rect 42613 10211 42671 10217
rect 30101 10183 30159 10189
rect 30101 10149 30113 10183
rect 30147 10180 30159 10183
rect 32858 10180 32864 10192
rect 30147 10152 30696 10180
rect 30147 10149 30159 10152
rect 30101 10143 30159 10149
rect 30024 10084 30138 10112
rect 29457 10047 29515 10053
rect 29457 10013 29469 10047
rect 29503 10013 29515 10047
rect 29457 10007 29515 10013
rect 29546 10004 29552 10056
rect 29604 10044 29610 10056
rect 30009 10047 30067 10053
rect 30009 10044 30021 10047
rect 29604 10016 30021 10044
rect 29604 10004 29610 10016
rect 30009 10013 30021 10016
rect 30055 10013 30067 10047
rect 30009 10007 30067 10013
rect 25682 9976 25688 9988
rect 23032 9948 23436 9976
rect 25530 9948 25688 9976
rect 21637 9939 21695 9945
rect 22296 9920 22324 9948
rect 20855 9880 21128 9908
rect 20855 9877 20867 9880
rect 20809 9871 20867 9877
rect 21726 9868 21732 9920
rect 21784 9868 21790 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 22189 9911 22247 9917
rect 22189 9908 22201 9911
rect 21876 9880 22201 9908
rect 21876 9868 21882 9880
rect 22189 9877 22201 9880
rect 22235 9877 22247 9911
rect 22189 9871 22247 9877
rect 22278 9868 22284 9920
rect 22336 9868 22342 9920
rect 22373 9911 22431 9917
rect 22373 9877 22385 9911
rect 22419 9908 22431 9911
rect 23290 9908 23296 9920
rect 22419 9880 23296 9908
rect 22419 9877 22431 9880
rect 22373 9871 22431 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 23408 9908 23436 9948
rect 25682 9936 25688 9948
rect 25740 9936 25746 9988
rect 28169 9979 28227 9985
rect 28169 9976 28181 9979
rect 27724 9948 28181 9976
rect 23842 9908 23848 9920
rect 23408 9880 23848 9908
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 24394 9868 24400 9920
rect 24452 9908 24458 9920
rect 25130 9908 25136 9920
rect 24452 9880 25136 9908
rect 24452 9868 24458 9880
rect 25130 9868 25136 9880
rect 25188 9908 25194 9920
rect 27724 9908 27752 9948
rect 28169 9945 28181 9948
rect 28215 9976 28227 9979
rect 28994 9976 29000 9988
rect 28215 9948 29000 9976
rect 28215 9945 28227 9948
rect 28169 9939 28227 9945
rect 28994 9936 29000 9948
rect 29052 9936 29058 9988
rect 29270 9936 29276 9988
rect 29328 9976 29334 9988
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 29328 9948 29745 9976
rect 29328 9936 29334 9948
rect 29733 9945 29745 9948
rect 29779 9945 29791 9979
rect 29733 9939 29791 9945
rect 29917 9979 29975 9985
rect 29917 9945 29929 9979
rect 29963 9976 29975 9979
rect 30110 9976 30138 10084
rect 30282 10072 30288 10124
rect 30340 10072 30346 10124
rect 30668 10112 30696 10152
rect 32048 10152 32864 10180
rect 31021 10115 31079 10121
rect 31021 10112 31033 10115
rect 30668 10084 31033 10112
rect 31021 10081 31033 10084
rect 31067 10081 31079 10115
rect 31021 10075 31079 10081
rect 31754 10072 31760 10124
rect 31812 10112 31818 10124
rect 32048 10112 32076 10152
rect 32858 10140 32864 10152
rect 32916 10140 32922 10192
rect 33152 10180 33180 10208
rect 37553 10183 37611 10189
rect 33152 10152 33805 10180
rect 31812 10084 32076 10112
rect 32493 10115 32551 10121
rect 31812 10072 31818 10084
rect 32493 10081 32505 10115
rect 32539 10112 32551 10115
rect 33045 10115 33103 10121
rect 33045 10112 33057 10115
rect 32539 10084 33057 10112
rect 32539 10081 32551 10084
rect 32493 10075 32551 10081
rect 33045 10081 33057 10084
rect 33091 10081 33103 10115
rect 33045 10075 33103 10081
rect 33137 10115 33195 10121
rect 33137 10081 33149 10115
rect 33183 10081 33195 10115
rect 33594 10112 33600 10124
rect 33137 10075 33195 10081
rect 33428 10084 33600 10112
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30469 10047 30527 10053
rect 30469 10013 30481 10047
rect 30515 10013 30527 10047
rect 30469 10007 30527 10013
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10044 30619 10047
rect 30650 10044 30656 10056
rect 30607 10016 30656 10044
rect 30607 10013 30619 10016
rect 30561 10007 30619 10013
rect 30282 9976 30288 9988
rect 29963 9948 30288 9976
rect 29963 9945 29975 9948
rect 29917 9939 29975 9945
rect 30282 9936 30288 9948
rect 30340 9936 30346 9988
rect 25188 9880 27752 9908
rect 25188 9868 25194 9880
rect 27982 9868 27988 9920
rect 28040 9908 28046 9920
rect 28721 9911 28779 9917
rect 28721 9908 28733 9911
rect 28040 9880 28733 9908
rect 28040 9868 28046 9880
rect 28721 9877 28733 9880
rect 28767 9877 28779 9911
rect 30392 9908 30420 10007
rect 30484 9976 30512 10007
rect 30650 10004 30656 10016
rect 30708 10004 30714 10056
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 32030 10004 32036 10056
rect 32088 10044 32094 10056
rect 32088 10016 32154 10044
rect 32088 10004 32094 10016
rect 30926 9976 30932 9988
rect 30484 9948 30932 9976
rect 30926 9936 30932 9948
rect 30984 9936 30990 9988
rect 32508 9908 32536 10075
rect 32766 10004 32772 10056
rect 32824 10044 32830 10056
rect 33152 10044 33180 10075
rect 32824 10016 33180 10044
rect 32824 10004 32830 10016
rect 32858 9936 32864 9988
rect 32916 9976 32922 9988
rect 33428 9985 33456 10084
rect 33594 10072 33600 10084
rect 33652 10072 33658 10124
rect 33777 10112 33805 10152
rect 37553 10149 37565 10183
rect 37599 10149 37611 10183
rect 37553 10143 37611 10149
rect 34333 10115 34391 10121
rect 34333 10112 34345 10115
rect 33777 10084 34345 10112
rect 34333 10081 34345 10084
rect 34379 10081 34391 10115
rect 34333 10075 34391 10081
rect 35710 10072 35716 10124
rect 35768 10112 35774 10124
rect 36449 10115 36507 10121
rect 36449 10112 36461 10115
rect 35768 10084 36461 10112
rect 35768 10072 35774 10084
rect 36449 10081 36461 10084
rect 36495 10081 36507 10115
rect 37568 10112 37596 10143
rect 36449 10075 36507 10081
rect 37200 10084 37596 10112
rect 38197 10115 38255 10121
rect 34057 10047 34115 10053
rect 34057 10013 34069 10047
rect 34103 10013 34115 10047
rect 34057 10007 34115 10013
rect 33413 9979 33471 9985
rect 32916 9948 33088 9976
rect 32916 9936 32922 9948
rect 30392 9880 32536 9908
rect 28721 9871 28779 9877
rect 32582 9868 32588 9920
rect 32640 9868 32646 9920
rect 32950 9868 32956 9920
rect 33008 9868 33014 9920
rect 33060 9908 33088 9948
rect 33413 9945 33425 9979
rect 33459 9945 33471 9979
rect 33413 9939 33471 9945
rect 33502 9936 33508 9988
rect 33560 9976 33566 9988
rect 33613 9979 33671 9985
rect 33613 9976 33625 9979
rect 33560 9948 33625 9976
rect 33560 9936 33566 9948
rect 33613 9945 33625 9948
rect 33659 9945 33671 9979
rect 34072 9976 34100 10007
rect 36262 10004 36268 10056
rect 36320 10004 36326 10056
rect 36906 10004 36912 10056
rect 36964 10004 36970 10056
rect 37200 10053 37228 10084
rect 38197 10081 38209 10115
rect 38243 10112 38255 10115
rect 38396 10112 38424 10208
rect 38565 10183 38623 10189
rect 38565 10149 38577 10183
rect 38611 10180 38623 10183
rect 39022 10180 39028 10192
rect 38611 10152 39028 10180
rect 38611 10149 38623 10152
rect 38565 10143 38623 10149
rect 39022 10140 39028 10152
rect 39080 10140 39086 10192
rect 39209 10183 39267 10189
rect 39209 10149 39221 10183
rect 39255 10149 39267 10183
rect 39209 10143 39267 10149
rect 39316 10152 39804 10180
rect 39224 10112 39252 10143
rect 39316 10124 39344 10152
rect 38243 10084 38424 10112
rect 38764 10084 39252 10112
rect 38243 10081 38255 10084
rect 38197 10075 38255 10081
rect 37185 10047 37243 10053
rect 37185 10013 37197 10047
rect 37231 10013 37243 10047
rect 37185 10007 37243 10013
rect 37461 10047 37519 10053
rect 37461 10013 37473 10047
rect 37507 10044 37519 10047
rect 38654 10044 38660 10056
rect 37507 10016 38660 10044
rect 37507 10013 37519 10016
rect 37461 10007 37519 10013
rect 38654 10004 38660 10016
rect 38712 10004 38718 10056
rect 38764 10053 38792 10084
rect 39298 10072 39304 10124
rect 39356 10072 39362 10124
rect 39390 10072 39396 10124
rect 39448 10112 39454 10124
rect 39776 10121 39804 10152
rect 39669 10115 39727 10121
rect 39669 10112 39681 10115
rect 39448 10084 39681 10112
rect 39448 10072 39454 10084
rect 39669 10081 39681 10084
rect 39715 10081 39727 10115
rect 39669 10075 39727 10081
rect 39761 10115 39819 10121
rect 39761 10081 39773 10115
rect 39807 10081 39819 10115
rect 39761 10075 39819 10081
rect 40773 10115 40831 10121
rect 40773 10081 40785 10115
rect 40819 10112 40831 10115
rect 41800 10112 41828 10208
rect 40819 10084 41828 10112
rect 40819 10081 40831 10084
rect 40773 10075 40831 10081
rect 38749 10047 38807 10053
rect 38749 10013 38761 10047
rect 38795 10013 38807 10047
rect 38749 10007 38807 10013
rect 39025 10047 39083 10053
rect 39025 10013 39037 10047
rect 39071 10044 39083 10047
rect 39114 10044 39120 10056
rect 39071 10016 39120 10044
rect 39071 10013 39083 10016
rect 39025 10007 39083 10013
rect 39114 10004 39120 10016
rect 39172 10004 39178 10056
rect 39577 10047 39635 10053
rect 39577 10013 39589 10047
rect 39623 10044 39635 10047
rect 40310 10044 40316 10056
rect 39623 10016 40316 10044
rect 39623 10013 39635 10016
rect 39577 10007 39635 10013
rect 40310 10004 40316 10016
rect 40368 10004 40374 10056
rect 40402 10004 40408 10056
rect 40460 10044 40466 10056
rect 40497 10047 40555 10053
rect 40497 10044 40509 10047
rect 40460 10016 40509 10044
rect 40460 10004 40466 10016
rect 40497 10013 40509 10016
rect 40543 10013 40555 10047
rect 40497 10007 40555 10013
rect 34422 9976 34428 9988
rect 34072 9948 34428 9976
rect 33613 9939 33671 9945
rect 34422 9936 34428 9948
rect 34480 9936 34486 9988
rect 34882 9936 34888 9988
rect 34940 9936 34946 9988
rect 35618 9936 35624 9988
rect 35676 9976 35682 9988
rect 40770 9976 40776 9988
rect 35676 9948 40776 9976
rect 35676 9936 35682 9948
rect 40770 9936 40776 9948
rect 40828 9936 40834 9988
rect 42518 9976 42524 9988
rect 41998 9948 42524 9976
rect 42518 9936 42524 9948
rect 42576 9936 42582 9988
rect 33781 9911 33839 9917
rect 33781 9908 33793 9911
rect 33060 9880 33793 9908
rect 33781 9877 33793 9880
rect 33827 9877 33839 9911
rect 33781 9871 33839 9877
rect 35342 9868 35348 9920
rect 35400 9908 35406 9920
rect 36357 9911 36415 9917
rect 36357 9908 36369 9911
rect 35400 9880 36369 9908
rect 35400 9868 35406 9880
rect 36357 9877 36369 9880
rect 36403 9877 36415 9911
rect 36357 9871 36415 9877
rect 36722 9868 36728 9920
rect 36780 9868 36786 9920
rect 36998 9868 37004 9920
rect 37056 9868 37062 9920
rect 37274 9868 37280 9920
rect 37332 9868 37338 9920
rect 37918 9868 37924 9920
rect 37976 9868 37982 9920
rect 38010 9868 38016 9920
rect 38068 9868 38074 9920
rect 39666 9868 39672 9920
rect 39724 9908 39730 9920
rect 40221 9911 40279 9917
rect 40221 9908 40233 9911
rect 39724 9880 40233 9908
rect 39724 9868 39730 9880
rect 40221 9877 40233 9880
rect 40267 9908 40279 9911
rect 40402 9908 40408 9920
rect 40267 9880 40408 9908
rect 40267 9877 40279 9880
rect 40221 9871 40279 9877
rect 40402 9868 40408 9880
rect 40460 9908 40466 9920
rect 40954 9908 40960 9920
rect 40460 9880 40960 9908
rect 40460 9868 40466 9880
rect 40954 9868 40960 9880
rect 41012 9908 41018 9920
rect 42628 9908 42656 10211
rect 42978 10208 42984 10220
rect 43036 10248 43042 10260
rect 43717 10251 43775 10257
rect 43717 10248 43729 10251
rect 43036 10220 43729 10248
rect 43036 10208 43042 10220
rect 43717 10217 43729 10220
rect 43763 10248 43775 10251
rect 44542 10248 44548 10260
rect 43763 10220 44548 10248
rect 43763 10217 43775 10220
rect 43717 10211 43775 10217
rect 44542 10208 44548 10220
rect 44600 10208 44606 10260
rect 43254 10140 43260 10192
rect 43312 10180 43318 10192
rect 43993 10183 44051 10189
rect 43993 10180 44005 10183
rect 43312 10152 44005 10180
rect 43312 10140 43318 10152
rect 43993 10149 44005 10152
rect 44039 10180 44051 10183
rect 44818 10180 44824 10192
rect 44039 10152 44824 10180
rect 44039 10149 44051 10152
rect 43993 10143 44051 10149
rect 44818 10140 44824 10152
rect 44876 10180 44882 10192
rect 44913 10183 44971 10189
rect 44913 10180 44925 10183
rect 44876 10152 44925 10180
rect 44876 10140 44882 10152
rect 44913 10149 44925 10152
rect 44959 10149 44971 10183
rect 44913 10143 44971 10149
rect 41012 9880 42656 9908
rect 41012 9868 41018 9880
rect 460 9818 45540 9840
rect 460 9766 6070 9818
rect 6122 9766 6134 9818
rect 6186 9766 6198 9818
rect 6250 9766 6262 9818
rect 6314 9766 6326 9818
rect 6378 9766 11070 9818
rect 11122 9766 11134 9818
rect 11186 9766 11198 9818
rect 11250 9766 11262 9818
rect 11314 9766 11326 9818
rect 11378 9766 16070 9818
rect 16122 9766 16134 9818
rect 16186 9766 16198 9818
rect 16250 9766 16262 9818
rect 16314 9766 16326 9818
rect 16378 9766 21070 9818
rect 21122 9766 21134 9818
rect 21186 9766 21198 9818
rect 21250 9766 21262 9818
rect 21314 9766 21326 9818
rect 21378 9766 26070 9818
rect 26122 9766 26134 9818
rect 26186 9766 26198 9818
rect 26250 9766 26262 9818
rect 26314 9766 26326 9818
rect 26378 9766 31070 9818
rect 31122 9766 31134 9818
rect 31186 9766 31198 9818
rect 31250 9766 31262 9818
rect 31314 9766 31326 9818
rect 31378 9766 36070 9818
rect 36122 9766 36134 9818
rect 36186 9766 36198 9818
rect 36250 9766 36262 9818
rect 36314 9766 36326 9818
rect 36378 9766 41070 9818
rect 41122 9766 41134 9818
rect 41186 9766 41198 9818
rect 41250 9766 41262 9818
rect 41314 9766 41326 9818
rect 41378 9766 45540 9818
rect 460 9744 45540 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 4338 9704 4344 9716
rect 3476 9676 4344 9704
rect 3476 9664 3482 9676
rect 3804 9577 3832 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4430 9664 4436 9716
rect 4488 9664 4494 9716
rect 5644 9676 5856 9704
rect 4065 9639 4123 9645
rect 4065 9605 4077 9639
rect 4111 9636 4123 9639
rect 4448 9636 4476 9664
rect 5644 9636 5672 9676
rect 4111 9608 4476 9636
rect 5290 9608 5672 9636
rect 4111 9605 4123 9608
rect 4065 9599 4123 9605
rect 5718 9596 5724 9648
rect 5776 9596 5782 9648
rect 5828 9636 5856 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 5960 9676 6193 9704
rect 5960 9664 5966 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 8018 9704 8024 9716
rect 6181 9667 6239 9673
rect 7852 9676 8024 9704
rect 6638 9636 6644 9648
rect 5828 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 6696 9608 7389 9636
rect 6696 9596 6702 9608
rect 7377 9605 7389 9608
rect 7423 9636 7435 9639
rect 7742 9636 7748 9648
rect 7423 9608 7748 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 3789 9531 3847 9537
rect 5276 9540 6009 9568
rect 5276 9512 5304 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 5258 9460 5264 9512
rect 5316 9460 5322 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 7852 9509 7880 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 9180 9676 9597 9704
rect 9180 9664 9186 9676
rect 9585 9673 9597 9676
rect 9631 9673 9643 9707
rect 9585 9667 9643 9673
rect 8113 9639 8171 9645
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 8312 9636 8340 9664
rect 8159 9608 8340 9636
rect 9600 9636 9628 9667
rect 10134 9664 10140 9716
rect 10192 9664 10198 9716
rect 12989 9707 13047 9713
rect 12989 9673 13001 9707
rect 13035 9704 13047 9707
rect 13262 9704 13268 9716
rect 13035 9676 13268 9704
rect 13035 9673 13047 9676
rect 12989 9667 13047 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 13446 9664 13452 9716
rect 13504 9664 13510 9716
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 14182 9704 14188 9716
rect 13596 9676 14188 9704
rect 13596 9664 13602 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 15102 9664 15108 9716
rect 15160 9704 15166 9716
rect 15160 9676 15240 9704
rect 15160 9664 15166 9676
rect 9600 9608 9904 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 5408 9472 5917 9500
rect 5408 9460 5414 9472
rect 5905 9469 5917 9472
rect 5951 9500 5963 9503
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 5951 9472 6132 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 6104 9376 6132 9472
rect 7760 9472 7849 9500
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5132 9336 5549 9364
rect 5132 9324 5138 9336
rect 5537 9333 5549 9336
rect 5583 9364 5595 9367
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5583 9336 5733 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5721 9333 5733 9336
rect 5767 9333 5779 9367
rect 5721 9327 5779 9333
rect 6086 9324 6092 9376
rect 6144 9324 6150 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7760 9373 7788 9472
rect 7837 9469 7849 9472
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 9232 9500 9260 9554
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 9876 9577 9904 9608
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 10652 9608 10701 9636
rect 10652 9596 10658 9608
rect 10689 9605 10701 9608
rect 10735 9605 10747 9639
rect 10689 9599 10747 9605
rect 11333 9639 11391 9645
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 12066 9636 12072 9648
rect 11379 9608 12072 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12176 9608 12449 9636
rect 9677 9571 9735 9577
rect 9677 9568 9689 9571
rect 9640 9540 9689 9568
rect 9640 9528 9646 9540
rect 9677 9537 9689 9540
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10410 9568 10416 9580
rect 9999 9540 10416 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11790 9528 11796 9580
rect 11848 9528 11854 9580
rect 12176 9577 12204 9608
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 12437 9599 12495 9605
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12452 9568 12480 9599
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12584 9608 13124 9636
rect 12584 9596 12590 9608
rect 12710 9568 12716 9580
rect 12452 9540 12716 9568
rect 12253 9531 12311 9537
rect 10042 9500 10048 9512
rect 8260 9472 10048 9500
rect 8260 9460 8266 9472
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 11992 9500 12020 9531
rect 12268 9500 12296 9531
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 12894 9528 12900 9580
rect 12952 9566 12958 9580
rect 13096 9577 13124 9608
rect 13354 9596 13360 9648
rect 13412 9596 13418 9648
rect 13464 9636 13492 9664
rect 15212 9636 15240 9676
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17126 9704 17132 9716
rect 16632 9676 17132 9704
rect 16632 9664 16638 9676
rect 17126 9664 17132 9676
rect 17184 9704 17190 9716
rect 17184 9676 17540 9704
rect 17184 9664 17190 9676
rect 16292 9639 16350 9645
rect 13464 9608 13846 9636
rect 15212 9608 16068 9636
rect 12989 9571 13047 9577
rect 12989 9566 13001 9571
rect 12952 9538 13001 9566
rect 12952 9528 12958 9538
rect 12989 9537 13001 9538
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13088 9571 13146 9577
rect 13088 9537 13100 9571
rect 13134 9537 13146 9571
rect 13088 9531 13146 9537
rect 15396 9512 15424 9608
rect 16040 9577 16068 9608
rect 16292 9605 16304 9639
rect 16338 9636 16350 9639
rect 16942 9636 16948 9648
rect 16338 9608 16948 9636
rect 16338 9605 16350 9608
rect 16292 9599 16350 9605
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 16025 9571 16083 9577
rect 15519 9540 15976 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 12342 9500 12348 9512
rect 11992 9472 12348 9500
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 13412 9472 14964 9500
rect 13412 9460 13418 9472
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 7064 9336 7757 9364
rect 7064 9324 7070 9336
rect 7745 9333 7757 9336
rect 7791 9333 7803 9367
rect 7745 9327 7803 9333
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 11238 9324 11244 9376
rect 11296 9324 11302 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11572 9336 11713 9364
rect 11572 9324 11578 9336
rect 11701 9333 11713 9336
rect 11747 9364 11759 9367
rect 11974 9364 11980 9376
rect 11747 9336 11980 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 12618 9324 12624 9376
rect 12676 9324 12682 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13998 9364 14004 9376
rect 12952 9336 14004 9364
rect 12952 9324 12958 9336
rect 13998 9324 14004 9336
rect 14056 9364 14062 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 14056 9336 14841 9364
rect 14056 9324 14062 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14936 9364 14964 9472
rect 15378 9460 15384 9512
rect 15436 9460 15442 9512
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15948 9500 15976 9540
rect 16025 9537 16037 9571
rect 16071 9537 16083 9571
rect 16850 9568 16856 9580
rect 16025 9531 16083 9537
rect 16132 9540 16856 9568
rect 16132 9500 16160 9540
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17512 9577 17540 9676
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 18472 9676 19196 9704
rect 18472 9664 18478 9676
rect 19168 9648 19196 9676
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21818 9704 21824 9716
rect 20864 9676 21824 9704
rect 20864 9664 20870 9676
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 17773 9639 17831 9645
rect 17773 9636 17785 9639
rect 17736 9608 17785 9636
rect 17736 9596 17742 9608
rect 17773 9605 17785 9608
rect 17819 9605 17831 9639
rect 17773 9599 17831 9605
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18104 9608 18262 9636
rect 18104 9596 18110 9608
rect 19150 9596 19156 9648
rect 19208 9636 19214 9648
rect 19797 9639 19855 9645
rect 19797 9636 19809 9639
rect 19208 9608 19809 9636
rect 19208 9596 19214 9608
rect 19797 9605 19809 9608
rect 19843 9605 19855 9639
rect 19797 9599 19855 9605
rect 20346 9596 20352 9648
rect 20404 9596 20410 9648
rect 21266 9636 21272 9648
rect 20640 9608 21272 9636
rect 20640 9577 20668 9608
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 20625 9571 20683 9577
rect 19751 9540 20392 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 15948 9472 16160 9500
rect 15565 9463 15623 9469
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15105 9435 15163 9441
rect 15105 9432 15117 9435
rect 15068 9404 15117 9432
rect 15068 9392 15074 9404
rect 15105 9401 15117 9404
rect 15151 9401 15163 9435
rect 15580 9432 15608 9463
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19720 9500 19748 9531
rect 19300 9472 19748 9500
rect 19300 9460 19306 9472
rect 19886 9460 19892 9512
rect 19944 9460 19950 9512
rect 20364 9500 20392 9540
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 20714 9528 20720 9580
rect 20772 9528 20778 9580
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9537 21051 9571
rect 21284 9568 21312 9596
rect 21542 9577 21600 9583
rect 21652 9580 21680 9676
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 21928 9676 22094 9704
rect 21453 9571 21511 9577
rect 21376 9568 21465 9571
rect 21284 9543 21465 9568
rect 21284 9540 21404 9543
rect 20993 9531 21051 9537
rect 21453 9537 21465 9543
rect 21499 9537 21511 9571
rect 21542 9543 21554 9577
rect 21588 9543 21600 9577
rect 21542 9537 21600 9543
rect 21637 9574 21695 9580
rect 21637 9540 21649 9574
rect 21683 9540 21695 9574
rect 21453 9531 21511 9537
rect 20916 9500 20944 9528
rect 20364 9472 20944 9500
rect 15580 9404 16068 9432
rect 15105 9395 15163 9401
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 14936 9336 15853 9364
rect 14829 9327 14887 9333
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 16040 9364 16068 9404
rect 19334 9392 19340 9444
rect 19392 9392 19398 9444
rect 17402 9364 17408 9376
rect 16040 9336 17408 9364
rect 15841 9327 15899 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 19904 9364 19932 9460
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 21008 9432 21036 9531
rect 21557 9444 21585 9537
rect 21637 9534 21695 9540
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 21836 9500 21864 9531
rect 21784 9472 21864 9500
rect 21784 9460 21790 9472
rect 20036 9404 21036 9432
rect 20036 9392 20042 9404
rect 21174 9392 21180 9444
rect 21232 9392 21238 9444
rect 21542 9392 21548 9444
rect 21600 9392 21606 9444
rect 19024 9336 19932 9364
rect 19024 9324 19030 9336
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 21818 9364 21824 9376
rect 20496 9336 21824 9364
rect 20496 9324 20502 9336
rect 21818 9324 21824 9336
rect 21876 9364 21882 9376
rect 21928 9364 21956 9676
rect 22066 9636 22094 9676
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 22373 9707 22431 9713
rect 22373 9704 22385 9707
rect 22336 9676 22385 9704
rect 22336 9664 22342 9676
rect 22373 9673 22385 9676
rect 22419 9704 22431 9707
rect 22833 9707 22891 9713
rect 22419 9676 22692 9704
rect 22419 9673 22431 9676
rect 22373 9667 22431 9673
rect 22465 9639 22523 9645
rect 22465 9636 22477 9639
rect 22066 9608 22477 9636
rect 22465 9605 22477 9608
rect 22511 9605 22523 9639
rect 22664 9636 22692 9676
rect 22833 9673 22845 9707
rect 22879 9704 22891 9707
rect 23750 9704 23756 9716
rect 22879 9676 23756 9704
rect 22879 9673 22891 9676
rect 22833 9667 22891 9673
rect 23750 9664 23756 9676
rect 23808 9664 23814 9716
rect 24394 9664 24400 9716
rect 24452 9664 24458 9716
rect 24578 9664 24584 9716
rect 24636 9704 24642 9716
rect 24946 9704 24952 9716
rect 24636 9676 24952 9704
rect 24636 9664 24642 9676
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 25406 9664 25412 9716
rect 25464 9704 25470 9716
rect 27706 9704 27712 9716
rect 25464 9676 26556 9704
rect 25464 9664 25470 9676
rect 23106 9636 23112 9648
rect 22664 9608 23112 9636
rect 22465 9599 22523 9605
rect 23106 9596 23112 9608
rect 23164 9636 23170 9648
rect 23164 9608 23796 9636
rect 23164 9596 23170 9608
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 23768 9577 23796 9608
rect 23842 9596 23848 9648
rect 23900 9636 23906 9648
rect 24489 9639 24547 9645
rect 24489 9636 24501 9639
rect 23900 9608 24501 9636
rect 23900 9596 23906 9608
rect 24489 9605 24501 9608
rect 24535 9636 24547 9639
rect 24535 9608 25268 9636
rect 24535 9605 24547 9608
rect 24489 9599 24547 9605
rect 23201 9571 23259 9577
rect 22060 9540 23060 9568
rect 22060 9528 22066 9540
rect 23032 9512 23060 9540
rect 23201 9537 23213 9571
rect 23247 9568 23259 9571
rect 23753 9571 23811 9577
rect 23247 9540 23520 9568
rect 23247 9537 23259 9540
rect 23201 9531 23259 9537
rect 22370 9460 22376 9512
rect 22428 9500 22434 9512
rect 22557 9503 22615 9509
rect 22557 9500 22569 9503
rect 22428 9472 22569 9500
rect 22428 9460 22434 9472
rect 22557 9469 22569 9472
rect 22603 9469 22615 9503
rect 22557 9463 22615 9469
rect 23014 9460 23020 9512
rect 23072 9500 23078 9512
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 23072 9472 23305 9500
rect 23072 9460 23078 9472
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 23385 9503 23443 9509
rect 23385 9469 23397 9503
rect 23431 9469 23443 9503
rect 23492 9500 23520 9540
rect 23753 9537 23765 9571
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 24949 9571 25007 9577
rect 24949 9537 24961 9571
rect 24995 9537 25007 9571
rect 24949 9531 25007 9537
rect 23934 9500 23940 9512
rect 23492 9472 23940 9500
rect 23385 9463 23443 9469
rect 23198 9432 23204 9444
rect 22020 9404 23204 9432
rect 22020 9373 22048 9404
rect 23198 9392 23204 9404
rect 23256 9392 23262 9444
rect 21876 9336 21956 9364
rect 22005 9367 22063 9373
rect 21876 9324 21882 9336
rect 22005 9333 22017 9367
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 22830 9364 22836 9376
rect 22244 9336 22836 9364
rect 22244 9324 22250 9336
rect 22830 9324 22836 9336
rect 22888 9364 22894 9376
rect 23400 9364 23428 9463
rect 23934 9460 23940 9472
rect 23992 9460 23998 9512
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 23474 9392 23480 9444
rect 23532 9432 23538 9444
rect 24596 9432 24624 9463
rect 24762 9460 24768 9512
rect 24820 9500 24826 9512
rect 24964 9500 24992 9531
rect 25240 9512 25268 9608
rect 25590 9596 25596 9648
rect 25648 9596 25654 9648
rect 25682 9596 25688 9648
rect 25740 9636 25746 9648
rect 26528 9645 26556 9676
rect 26611 9676 27712 9704
rect 25961 9639 26019 9645
rect 25961 9636 25973 9639
rect 25740 9608 25973 9636
rect 25740 9596 25746 9608
rect 25961 9605 25973 9608
rect 26007 9605 26019 9639
rect 25961 9599 26019 9605
rect 26513 9639 26571 9645
rect 26513 9605 26525 9639
rect 26559 9605 26571 9639
rect 26513 9599 26571 9605
rect 25976 9568 26004 9599
rect 26611 9568 26639 9676
rect 27706 9664 27712 9676
rect 27764 9664 27770 9716
rect 29730 9664 29736 9716
rect 29788 9704 29794 9716
rect 31691 9707 31749 9713
rect 29788 9676 30236 9704
rect 29788 9664 29794 9676
rect 30208 9648 30236 9676
rect 30944 9676 31524 9704
rect 29026 9608 29500 9636
rect 25976 9540 26639 9568
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9568 27031 9571
rect 27019 9540 27936 9568
rect 27019 9537 27031 9540
rect 26973 9531 27031 9537
rect 24820 9472 24992 9500
rect 24820 9460 24826 9472
rect 25038 9460 25044 9512
rect 25096 9460 25102 9512
rect 25222 9460 25228 9512
rect 25280 9460 25286 9512
rect 26694 9460 26700 9512
rect 26752 9460 26758 9512
rect 27614 9460 27620 9512
rect 27672 9460 27678 9512
rect 27908 9500 27936 9540
rect 27982 9528 27988 9580
rect 28040 9528 28046 9580
rect 28166 9500 28172 9512
rect 27908 9472 28172 9500
rect 28166 9460 28172 9472
rect 28224 9460 28230 9512
rect 29362 9460 29368 9512
rect 29420 9460 29426 9512
rect 29472 9500 29500 9608
rect 29932 9580 30144 9602
rect 30190 9596 30196 9648
rect 30248 9596 30254 9648
rect 30374 9596 30380 9648
rect 30432 9596 30438 9648
rect 30466 9596 30472 9648
rect 30524 9636 30530 9648
rect 30577 9639 30635 9645
rect 30577 9636 30589 9639
rect 30524 9608 30589 9636
rect 30524 9596 30530 9608
rect 30577 9605 30589 9608
rect 30623 9605 30635 9639
rect 30837 9639 30895 9645
rect 30837 9636 30849 9639
rect 30577 9599 30635 9605
rect 30668 9608 30849 9636
rect 29822 9528 29828 9580
rect 29880 9528 29886 9580
rect 29914 9528 29920 9580
rect 29972 9577 30144 9580
rect 29972 9574 30159 9577
rect 29972 9528 29978 9574
rect 30101 9571 30159 9574
rect 30101 9537 30113 9571
rect 30147 9537 30159 9571
rect 30101 9531 30159 9537
rect 30006 9500 30012 9512
rect 29472 9472 30012 9500
rect 30006 9460 30012 9472
rect 30064 9460 30070 9512
rect 25056 9432 25084 9460
rect 23532 9404 24624 9432
rect 24688 9404 25084 9432
rect 23532 9392 23538 9404
rect 22888 9336 23428 9364
rect 23845 9367 23903 9373
rect 22888 9324 22894 9336
rect 23845 9333 23857 9367
rect 23891 9364 23903 9367
rect 23934 9364 23940 9376
rect 23891 9336 23940 9364
rect 23891 9333 23903 9336
rect 23845 9327 23903 9333
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24029 9367 24087 9373
rect 24029 9333 24041 9367
rect 24075 9364 24087 9367
rect 24688 9364 24716 9404
rect 24075 9336 24716 9364
rect 24075 9333 24087 9336
rect 24029 9327 24087 9333
rect 25038 9324 25044 9376
rect 25096 9324 25102 9376
rect 29380 9373 29408 9460
rect 29914 9392 29920 9444
rect 29972 9432 29978 9444
rect 30374 9432 30380 9444
rect 29972 9404 30380 9432
rect 29972 9392 29978 9404
rect 30374 9392 30380 9404
rect 30432 9432 30438 9444
rect 30668 9432 30696 9608
rect 30837 9605 30849 9608
rect 30883 9636 30895 9639
rect 30944 9636 30972 9676
rect 31496 9645 31524 9676
rect 31691 9673 31703 9707
rect 31737 9704 31749 9707
rect 31938 9704 31944 9716
rect 31737 9676 31944 9704
rect 31737 9673 31749 9676
rect 31691 9667 31749 9673
rect 31938 9664 31944 9676
rect 31996 9664 32002 9716
rect 32490 9664 32496 9716
rect 32548 9664 32554 9716
rect 32950 9664 32956 9716
rect 33008 9664 33014 9716
rect 33042 9664 33048 9716
rect 33100 9704 33106 9716
rect 34149 9707 34207 9713
rect 34149 9704 34161 9707
rect 33100 9676 34161 9704
rect 33100 9664 33106 9676
rect 34149 9673 34161 9676
rect 34195 9673 34207 9707
rect 34149 9667 34207 9673
rect 34514 9664 34520 9716
rect 34572 9704 34578 9716
rect 34882 9704 34888 9716
rect 34572 9676 34888 9704
rect 34572 9664 34578 9676
rect 34882 9664 34888 9676
rect 34940 9704 34946 9716
rect 36265 9707 36323 9713
rect 34940 9676 35204 9704
rect 34940 9664 34946 9676
rect 30883 9608 30972 9636
rect 31481 9639 31539 9645
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 31067 9605 31125 9611
rect 31067 9571 31079 9605
rect 31113 9571 31125 9605
rect 31481 9605 31493 9639
rect 31527 9636 31539 9639
rect 31570 9636 31576 9648
rect 31527 9608 31576 9636
rect 31527 9605 31539 9608
rect 31481 9599 31539 9605
rect 31570 9596 31576 9608
rect 31628 9636 31634 9648
rect 33781 9639 33839 9645
rect 33781 9636 33793 9639
rect 31628 9608 33793 9636
rect 31628 9596 31634 9608
rect 33781 9605 33793 9608
rect 33827 9605 33839 9639
rect 33781 9599 33839 9605
rect 33962 9596 33968 9648
rect 34020 9645 34026 9648
rect 34020 9639 34039 9645
rect 34027 9605 34039 9639
rect 34020 9599 34039 9605
rect 34793 9639 34851 9645
rect 34793 9605 34805 9639
rect 34839 9636 34851 9639
rect 35066 9636 35072 9648
rect 34839 9608 35072 9636
rect 34839 9605 34851 9608
rect 34793 9599 34851 9605
rect 34020 9596 34026 9599
rect 35066 9596 35072 9608
rect 35124 9596 35130 9648
rect 35176 9636 35204 9676
rect 36265 9673 36277 9707
rect 36311 9704 36323 9707
rect 36446 9704 36452 9716
rect 36311 9676 36452 9704
rect 36311 9673 36323 9676
rect 36265 9667 36323 9673
rect 36446 9664 36452 9676
rect 36504 9664 36510 9716
rect 38654 9664 38660 9716
rect 38712 9704 38718 9716
rect 38933 9707 38991 9713
rect 38933 9704 38945 9707
rect 38712 9676 38945 9704
rect 38712 9664 38718 9676
rect 38933 9673 38945 9676
rect 38979 9673 38991 9707
rect 38933 9667 38991 9673
rect 40402 9664 40408 9716
rect 40460 9704 40466 9716
rect 40773 9707 40831 9713
rect 40773 9704 40785 9707
rect 40460 9676 40785 9704
rect 40460 9664 40466 9676
rect 40773 9673 40785 9676
rect 40819 9673 40831 9707
rect 41782 9704 41788 9716
rect 40773 9667 40831 9673
rect 41386 9676 41788 9704
rect 36633 9639 36691 9645
rect 36633 9636 36645 9639
rect 35176 9608 35282 9636
rect 36096 9608 36645 9636
rect 31067 9568 31125 9571
rect 32030 9568 32036 9580
rect 31067 9565 32036 9568
rect 31082 9540 32036 9565
rect 32030 9528 32036 9540
rect 32088 9528 32094 9580
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9568 32459 9571
rect 33226 9568 33232 9580
rect 32447 9540 33232 9568
rect 32447 9537 32459 9540
rect 32401 9531 32459 9537
rect 33226 9528 33232 9540
rect 33284 9528 33290 9580
rect 33318 9528 33324 9580
rect 33376 9528 33382 9580
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9568 33471 9571
rect 33459 9540 34468 9568
rect 33459 9537 33471 9540
rect 33413 9531 33471 9537
rect 32677 9503 32735 9509
rect 32677 9469 32689 9503
rect 32723 9500 32735 9503
rect 32766 9500 32772 9512
rect 32723 9472 32772 9500
rect 32723 9469 32735 9472
rect 32677 9463 32735 9469
rect 32766 9460 32772 9472
rect 32824 9460 32830 9512
rect 33597 9503 33655 9509
rect 33597 9469 33609 9503
rect 33643 9500 33655 9503
rect 34330 9500 34336 9512
rect 33643 9472 34336 9500
rect 33643 9469 33655 9472
rect 33597 9463 33655 9469
rect 34330 9460 34336 9472
rect 34388 9460 34394 9512
rect 30432 9404 30696 9432
rect 30432 9392 30438 9404
rect 30742 9392 30748 9444
rect 30800 9392 30806 9444
rect 31202 9392 31208 9444
rect 31260 9392 31266 9444
rect 31680 9404 34008 9432
rect 29365 9367 29423 9373
rect 29365 9333 29377 9367
rect 29411 9333 29423 9367
rect 29365 9327 29423 9333
rect 29641 9367 29699 9373
rect 29641 9333 29653 9367
rect 29687 9364 29699 9367
rect 29730 9364 29736 9376
rect 29687 9336 29736 9364
rect 29687 9333 29699 9336
rect 29641 9327 29699 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 29822 9324 29828 9376
rect 29880 9364 29886 9376
rect 31680 9373 31708 9404
rect 33980 9376 34008 9404
rect 30561 9367 30619 9373
rect 30561 9364 30573 9367
rect 29880 9336 30573 9364
rect 29880 9324 29886 9336
rect 30561 9333 30573 9336
rect 30607 9364 30619 9367
rect 31021 9367 31079 9373
rect 31021 9364 31033 9367
rect 30607 9336 31033 9364
rect 30607 9333 30619 9336
rect 30561 9327 30619 9333
rect 31021 9333 31033 9336
rect 31067 9364 31079 9367
rect 31665 9367 31723 9373
rect 31665 9364 31677 9367
rect 31067 9336 31677 9364
rect 31067 9333 31079 9336
rect 31021 9327 31079 9333
rect 31665 9333 31677 9336
rect 31711 9333 31723 9367
rect 31665 9327 31723 9333
rect 31846 9324 31852 9376
rect 31904 9324 31910 9376
rect 32030 9324 32036 9376
rect 32088 9324 32094 9376
rect 32122 9324 32128 9376
rect 32180 9364 32186 9376
rect 32858 9364 32864 9376
rect 32180 9336 32864 9364
rect 32180 9324 32186 9336
rect 32858 9324 32864 9336
rect 32916 9324 32922 9376
rect 33962 9324 33968 9376
rect 34020 9324 34026 9376
rect 34440 9364 34468 9540
rect 34517 9503 34575 9509
rect 34517 9469 34529 9503
rect 34563 9500 34575 9503
rect 34790 9500 34796 9512
rect 34563 9472 34796 9500
rect 34563 9469 34575 9472
rect 34517 9463 34575 9469
rect 34790 9460 34796 9472
rect 34848 9460 34854 9512
rect 34882 9460 34888 9512
rect 34940 9500 34946 9512
rect 35802 9500 35808 9512
rect 34940 9472 35808 9500
rect 34940 9460 34946 9472
rect 35802 9460 35808 9472
rect 35860 9500 35866 9512
rect 36096 9500 36124 9608
rect 36633 9605 36645 9608
rect 36679 9605 36691 9639
rect 36633 9599 36691 9605
rect 36814 9596 36820 9648
rect 36872 9645 36878 9648
rect 36872 9639 36891 9645
rect 36879 9605 36891 9639
rect 36872 9599 36891 9605
rect 36872 9596 36878 9599
rect 37274 9596 37280 9648
rect 37332 9636 37338 9648
rect 37369 9639 37427 9645
rect 37369 9636 37381 9639
rect 37332 9608 37381 9636
rect 37332 9596 37338 9608
rect 37369 9605 37381 9608
rect 37415 9605 37427 9639
rect 37369 9599 37427 9605
rect 37458 9596 37464 9648
rect 37516 9636 37522 9648
rect 39301 9639 39359 9645
rect 37516 9608 37858 9636
rect 37516 9596 37522 9608
rect 39301 9605 39313 9639
rect 39347 9636 39359 9639
rect 40129 9639 40187 9645
rect 40129 9636 40141 9639
rect 39347 9608 40141 9636
rect 39347 9605 39359 9608
rect 39301 9599 39359 9605
rect 40129 9605 40141 9608
rect 40175 9636 40187 9639
rect 41386 9636 41414 9676
rect 41782 9664 41788 9676
rect 41840 9664 41846 9716
rect 42978 9664 42984 9716
rect 43036 9664 43042 9716
rect 43254 9664 43260 9716
rect 43312 9664 43318 9716
rect 40175 9608 41414 9636
rect 40175 9605 40187 9608
rect 40129 9599 40187 9605
rect 41506 9596 41512 9648
rect 41564 9636 41570 9648
rect 42613 9639 42671 9645
rect 42613 9636 42625 9639
rect 41564 9608 42625 9636
rect 41564 9596 41570 9608
rect 42613 9605 42625 9608
rect 42659 9636 42671 9639
rect 43272 9636 43300 9664
rect 42659 9608 43300 9636
rect 42659 9605 42671 9608
rect 42613 9599 42671 9605
rect 37090 9528 37096 9580
rect 37148 9528 37154 9580
rect 39592 9540 40448 9568
rect 35860 9472 36124 9500
rect 35860 9460 35866 9472
rect 36630 9460 36636 9512
rect 36688 9500 36694 9512
rect 37108 9500 37136 9528
rect 39592 9509 39620 9540
rect 38841 9503 38899 9509
rect 38841 9500 38853 9503
rect 36688 9472 37136 9500
rect 37200 9472 38853 9500
rect 36688 9460 36694 9472
rect 37200 9432 37228 9472
rect 38841 9469 38853 9472
rect 38887 9500 38899 9503
rect 39393 9503 39451 9509
rect 39393 9500 39405 9503
rect 38887 9472 39405 9500
rect 38887 9469 38899 9472
rect 38841 9463 38899 9469
rect 39393 9469 39405 9472
rect 39439 9469 39451 9503
rect 39393 9463 39451 9469
rect 39577 9503 39635 9509
rect 39577 9469 39589 9503
rect 39623 9469 39635 9503
rect 39577 9463 39635 9469
rect 40126 9460 40132 9512
rect 40184 9500 40190 9512
rect 40221 9503 40279 9509
rect 40221 9500 40233 9503
rect 40184 9472 40233 9500
rect 40184 9460 40190 9472
rect 40221 9469 40233 9472
rect 40267 9469 40279 9503
rect 40221 9463 40279 9469
rect 40313 9503 40371 9509
rect 40313 9469 40325 9503
rect 40359 9469 40371 9503
rect 40420 9500 40448 9540
rect 40862 9528 40868 9580
rect 40920 9568 40926 9580
rect 41141 9571 41199 9577
rect 41141 9568 41153 9571
rect 40920 9540 41153 9568
rect 40920 9528 40926 9540
rect 41141 9537 41153 9540
rect 41187 9537 41199 9571
rect 41141 9531 41199 9537
rect 41785 9571 41843 9577
rect 41785 9537 41797 9571
rect 41831 9568 41843 9571
rect 42702 9568 42708 9580
rect 41831 9540 42708 9568
rect 41831 9537 41843 9540
rect 41785 9531 41843 9537
rect 42702 9528 42708 9540
rect 42760 9528 42766 9580
rect 43441 9571 43499 9577
rect 43441 9537 43453 9571
rect 43487 9568 43499 9571
rect 44634 9568 44640 9580
rect 43487 9540 44640 9568
rect 43487 9537 43499 9540
rect 43441 9531 43499 9537
rect 44634 9528 44640 9540
rect 44692 9528 44698 9580
rect 41417 9503 41475 9509
rect 41417 9500 41429 9503
rect 40420 9472 41429 9500
rect 40313 9463 40371 9469
rect 41417 9469 41429 9472
rect 41463 9500 41475 9503
rect 41690 9500 41696 9512
rect 41463 9472 41696 9500
rect 41463 9469 41475 9472
rect 41417 9463 41475 9469
rect 35820 9404 37228 9432
rect 35820 9364 35848 9404
rect 38470 9392 38476 9444
rect 38528 9432 38534 9444
rect 40328 9432 40356 9463
rect 41690 9460 41696 9472
rect 41748 9460 41754 9512
rect 41966 9460 41972 9512
rect 42024 9500 42030 9512
rect 42610 9500 42616 9512
rect 42024 9472 42616 9500
rect 42024 9460 42030 9472
rect 42610 9460 42616 9472
rect 42668 9500 42674 9512
rect 42668 9472 42932 9500
rect 42668 9460 42674 9472
rect 42058 9432 42064 9444
rect 38528 9404 42064 9432
rect 38528 9392 38534 9404
rect 42058 9392 42064 9404
rect 42116 9392 42122 9444
rect 34440 9336 35848 9364
rect 35894 9324 35900 9376
rect 35952 9364 35958 9376
rect 36817 9367 36875 9373
rect 36817 9364 36829 9367
rect 35952 9336 36829 9364
rect 35952 9324 35958 9336
rect 36817 9333 36829 9336
rect 36863 9333 36875 9367
rect 36817 9327 36875 9333
rect 37001 9367 37059 9373
rect 37001 9333 37013 9367
rect 37047 9364 37059 9367
rect 37182 9364 37188 9376
rect 37047 9336 37188 9364
rect 37047 9333 37059 9336
rect 37001 9327 37059 9333
rect 37182 9324 37188 9336
rect 37240 9324 37246 9376
rect 39758 9324 39764 9376
rect 39816 9324 39822 9376
rect 42904 9364 42932 9472
rect 44726 9392 44732 9444
rect 44784 9392 44790 9444
rect 43349 9367 43407 9373
rect 43349 9364 43361 9367
rect 42904 9336 43361 9364
rect 43349 9333 43361 9336
rect 43395 9364 43407 9367
rect 44542 9364 44548 9376
rect 43395 9336 44548 9364
rect 43395 9333 43407 9336
rect 43349 9327 43407 9333
rect 44542 9324 44548 9336
rect 44600 9324 44606 9376
rect 460 9274 45540 9296
rect 460 9222 3570 9274
rect 3622 9222 3634 9274
rect 3686 9222 3698 9274
rect 3750 9222 3762 9274
rect 3814 9222 3826 9274
rect 3878 9222 8570 9274
rect 8622 9222 8634 9274
rect 8686 9222 8698 9274
rect 8750 9222 8762 9274
rect 8814 9222 8826 9274
rect 8878 9222 13570 9274
rect 13622 9222 13634 9274
rect 13686 9222 13698 9274
rect 13750 9222 13762 9274
rect 13814 9222 13826 9274
rect 13878 9222 18570 9274
rect 18622 9222 18634 9274
rect 18686 9222 18698 9274
rect 18750 9222 18762 9274
rect 18814 9222 18826 9274
rect 18878 9222 23570 9274
rect 23622 9222 23634 9274
rect 23686 9222 23698 9274
rect 23750 9222 23762 9274
rect 23814 9222 23826 9274
rect 23878 9222 28570 9274
rect 28622 9222 28634 9274
rect 28686 9222 28698 9274
rect 28750 9222 28762 9274
rect 28814 9222 28826 9274
rect 28878 9222 33570 9274
rect 33622 9222 33634 9274
rect 33686 9222 33698 9274
rect 33750 9222 33762 9274
rect 33814 9222 33826 9274
rect 33878 9222 38570 9274
rect 38622 9222 38634 9274
rect 38686 9222 38698 9274
rect 38750 9222 38762 9274
rect 38814 9222 38826 9274
rect 38878 9222 43570 9274
rect 43622 9222 43634 9274
rect 43686 9222 43698 9274
rect 43750 9222 43762 9274
rect 43814 9222 43826 9274
rect 43878 9222 45540 9274
rect 460 9200 45540 9222
rect 6086 9120 6092 9172
rect 6144 9120 6150 9172
rect 6638 9120 6644 9172
rect 6696 9120 6702 9172
rect 6914 9120 6920 9172
rect 6972 9120 6978 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8202 9160 8208 9172
rect 7800 9132 8208 9160
rect 7800 9120 7806 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8849 9163 8907 9169
rect 8849 9160 8861 9163
rect 8536 9132 8861 9160
rect 8536 9120 8542 9132
rect 8849 9129 8861 9132
rect 8895 9129 8907 9163
rect 8849 9123 8907 9129
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9585 9163 9643 9169
rect 9585 9160 9597 9163
rect 9088 9132 9597 9160
rect 9088 9120 9094 9132
rect 9585 9129 9597 9132
rect 9631 9160 9643 9163
rect 10502 9160 10508 9172
rect 9631 9132 10508 9160
rect 9631 9129 9643 9132
rect 9585 9123 9643 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11974 9160 11980 9172
rect 11112 9132 11980 9160
rect 11112 9120 11118 9132
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12768 9132 12909 9160
rect 12768 9120 12774 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 13354 9120 13360 9172
rect 13412 9120 13418 9172
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 6932 9092 6960 9120
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 6932 9064 8585 9092
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8573 9055 8631 9061
rect 8956 9064 9674 9092
rect 8956 9024 8984 9064
rect 768 8996 8984 9024
rect 9646 9024 9674 9064
rect 9950 9052 9956 9104
rect 10008 9052 10014 9104
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10318 9092 10324 9104
rect 10100 9064 10324 9092
rect 10100 9052 10106 9064
rect 10318 9052 10324 9064
rect 10376 9092 10382 9104
rect 10597 9095 10655 9101
rect 10597 9092 10609 9095
rect 10376 9064 10609 9092
rect 10376 9052 10382 9064
rect 10597 9061 10609 9064
rect 10643 9061 10655 9095
rect 10597 9055 10655 9061
rect 12986 9052 12992 9104
rect 13044 9052 13050 9104
rect 13372 9092 13400 9120
rect 13096 9064 13400 9092
rect 13096 9024 13124 9064
rect 13464 9036 13492 9123
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 15068 9132 15301 9160
rect 15068 9120 15074 9132
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 19242 9120 19248 9172
rect 19300 9120 19306 9172
rect 21542 9160 21548 9172
rect 19536 9132 21548 9160
rect 14182 9052 14188 9104
rect 14240 9052 14246 9104
rect 19260 9092 19288 9120
rect 19168 9064 19288 9092
rect 9646 8996 13124 9024
rect 768 8965 796 8996
rect 13446 8984 13452 9036
rect 13504 8984 13510 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15194 9024 15200 9036
rect 13872 8996 15200 9024
rect 13872 8984 13878 8996
rect 15194 8984 15200 8996
rect 15252 9024 15258 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 15252 8996 16405 9024
rect 15252 8984 15258 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 16945 9027 17003 9033
rect 16945 8993 16957 9027
rect 16991 9024 17003 9027
rect 18230 9024 18236 9036
rect 16991 8996 18236 9024
rect 16991 8993 17003 8996
rect 16945 8987 17003 8993
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 18966 8984 18972 9036
rect 19024 8984 19030 9036
rect 19168 9033 19196 9064
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19245 9027 19303 9033
rect 19245 8993 19257 9027
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 753 8959 811 8965
rect 753 8925 765 8959
rect 799 8925 811 8959
rect 753 8919 811 8925
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4338 8916 4344 8968
rect 4396 8916 4402 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 4172 8888 4200 8916
rect 4617 8891 4675 8897
rect 4617 8888 4629 8891
rect 4172 8860 4629 8888
rect 4617 8857 4629 8860
rect 4663 8857 4675 8891
rect 5994 8888 6000 8900
rect 5842 8860 6000 8888
rect 4617 8851 4675 8857
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8588 8888 8616 8919
rect 8754 8916 8760 8968
rect 8812 8916 8818 8968
rect 8849 8925 8907 8931
rect 8444 8860 8616 8888
rect 8849 8891 8861 8925
rect 8895 8922 8907 8925
rect 8938 8922 8944 8968
rect 8895 8916 8944 8922
rect 8996 8916 9002 8968
rect 9030 8916 9036 8968
rect 9088 8916 9094 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 9490 8956 9496 8968
rect 9171 8928 9496 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9674 8916 9680 8968
rect 9732 8916 9738 8968
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 8895 8894 8984 8916
rect 8895 8891 8907 8894
rect 8849 8885 8907 8891
rect 8444 8848 8450 8860
rect 934 8780 940 8832
rect 992 8780 998 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7006 8820 7012 8832
rect 6963 8792 7012 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7006 8780 7012 8792
rect 7064 8820 7070 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 7064 8792 7297 8820
rect 7064 8780 7070 8792
rect 7285 8789 7297 8792
rect 7331 8820 7343 8823
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 7331 8792 8125 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 8113 8789 8125 8792
rect 8159 8820 8171 8823
rect 8478 8820 8484 8832
rect 8159 8792 8484 8820
rect 8159 8789 8171 8792
rect 8113 8783 8171 8789
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8588 8820 8616 8860
rect 8956 8820 8984 8894
rect 9217 8891 9275 8897
rect 9217 8857 9229 8891
rect 9263 8888 9275 8891
rect 9306 8888 9312 8900
rect 9263 8860 9312 8888
rect 9263 8857 9275 8860
rect 9217 8851 9275 8857
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 9401 8891 9459 8897
rect 9401 8857 9413 8891
rect 9447 8888 9459 8891
rect 9692 8888 9720 8916
rect 9447 8860 9720 8888
rect 9953 8891 10011 8897
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 9953 8857 9965 8891
rect 9999 8857 10011 8891
rect 9953 8851 10011 8857
rect 9582 8820 9588 8832
rect 8588 8792 9588 8820
rect 9582 8780 9588 8792
rect 9640 8820 9646 8832
rect 9968 8820 9996 8851
rect 9640 8792 9996 8820
rect 9640 8780 9646 8792
rect 10134 8780 10140 8832
rect 10192 8780 10198 8832
rect 11164 8820 11192 8919
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 12952 8928 13277 8956
rect 12952 8916 12958 8928
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13412 8928 13737 8956
rect 13412 8916 13418 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 13998 8916 14004 8968
rect 14056 8916 14062 8968
rect 16574 8956 16580 8968
rect 15672 8928 16580 8956
rect 11425 8891 11483 8897
rect 11425 8857 11437 8891
rect 11471 8888 11483 8891
rect 11698 8888 11704 8900
rect 11471 8860 11704 8888
rect 11471 8857 11483 8860
rect 11425 8851 11483 8857
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 11882 8848 11888 8900
rect 11940 8848 11946 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12989 8891 13047 8897
rect 12989 8888 13001 8891
rect 12768 8860 13001 8888
rect 12768 8848 12774 8860
rect 12989 8857 13001 8860
rect 13035 8888 13047 8891
rect 13078 8888 13084 8900
rect 13035 8860 13084 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13170 8848 13176 8900
rect 13228 8848 13234 8900
rect 13449 8891 13507 8897
rect 13449 8857 13461 8891
rect 13495 8888 13507 8891
rect 13538 8888 13544 8900
rect 13495 8860 13544 8888
rect 13495 8857 13507 8860
rect 13449 8851 13507 8857
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 13633 8891 13691 8897
rect 13633 8857 13645 8891
rect 13679 8888 13691 8891
rect 13817 8891 13875 8897
rect 13817 8888 13829 8891
rect 13679 8860 13829 8888
rect 13679 8857 13691 8860
rect 13633 8851 13691 8857
rect 13817 8857 13829 8860
rect 13863 8888 13875 8891
rect 13863 8860 15148 8888
rect 13863 8857 13875 8860
rect 13817 8851 13875 8857
rect 12434 8820 12440 8832
rect 11164 8792 12440 8820
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13648 8820 13676 8851
rect 15120 8832 15148 8860
rect 12860 8792 13676 8820
rect 12860 8780 12866 8792
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 14553 8823 14611 8829
rect 14553 8820 14565 8823
rect 14516 8792 14565 8820
rect 14516 8780 14522 8792
rect 14553 8789 14565 8792
rect 14599 8820 14611 8823
rect 14921 8823 14979 8829
rect 14921 8820 14933 8823
rect 14599 8792 14933 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 14921 8789 14933 8792
rect 14967 8820 14979 8823
rect 15010 8820 15016 8832
rect 14967 8792 15016 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 15672 8829 15700 8928
rect 16574 8916 16580 8928
rect 16632 8956 16638 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16632 8928 16681 8956
rect 16632 8916 16638 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 18984 8956 19012 8984
rect 19260 8956 19288 8987
rect 18984 8928 19288 8956
rect 16669 8919 16727 8925
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 19536 8965 19564 9132
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 22649 9163 22707 9169
rect 22649 9129 22661 9163
rect 22695 9160 22707 9163
rect 22922 9160 22928 9172
rect 22695 9132 22928 9160
rect 22695 9129 22707 9132
rect 22649 9123 22707 9129
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 23014 9120 23020 9172
rect 23072 9160 23078 9172
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 23072 9132 23121 9160
rect 23072 9120 23078 9132
rect 23109 9129 23121 9132
rect 23155 9160 23167 9163
rect 23477 9163 23535 9169
rect 23155 9132 23428 9160
rect 23155 9129 23167 9132
rect 23109 9123 23167 9129
rect 19610 9052 19616 9104
rect 19668 9052 19674 9104
rect 23290 9052 23296 9104
rect 23348 9052 23354 9104
rect 23400 9092 23428 9132
rect 23477 9129 23489 9163
rect 23523 9160 23535 9163
rect 23658 9160 23664 9172
rect 23523 9132 23664 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24762 9160 24768 9172
rect 24167 9132 24768 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24136 9092 24164 9123
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 25958 9160 25964 9172
rect 25372 9132 25964 9160
rect 25372 9120 25378 9132
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26145 9163 26203 9169
rect 26145 9129 26157 9163
rect 26191 9160 26203 9163
rect 26694 9160 26700 9172
rect 26191 9132 26700 9160
rect 26191 9129 26203 9132
rect 26145 9123 26203 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 27522 9120 27528 9172
rect 27580 9160 27586 9172
rect 27890 9160 27896 9172
rect 27580 9132 27896 9160
rect 27580 9120 27586 9132
rect 27890 9120 27896 9132
rect 27948 9120 27954 9172
rect 29178 9120 29184 9172
rect 29236 9120 29242 9172
rect 29365 9163 29423 9169
rect 29365 9129 29377 9163
rect 29411 9160 29423 9163
rect 29546 9160 29552 9172
rect 29411 9132 29552 9160
rect 29411 9129 29423 9132
rect 29365 9123 29423 9129
rect 29546 9120 29552 9132
rect 29604 9120 29610 9172
rect 29720 9163 29778 9169
rect 29720 9129 29732 9163
rect 29766 9160 29778 9163
rect 29914 9160 29920 9172
rect 29766 9132 29920 9160
rect 29766 9129 29778 9132
rect 29720 9123 29778 9129
rect 29914 9120 29920 9132
rect 29972 9120 29978 9172
rect 30466 9120 30472 9172
rect 30524 9160 30530 9172
rect 31570 9160 31576 9172
rect 30524 9132 31576 9160
rect 30524 9120 30530 9132
rect 31570 9120 31576 9132
rect 31628 9120 31634 9172
rect 32766 9160 32772 9172
rect 32140 9132 32772 9160
rect 23400 9064 24164 9092
rect 25130 9052 25136 9104
rect 25188 9092 25194 9104
rect 25188 9064 25820 9092
rect 25188 9052 25194 9064
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19484 8928 19533 8956
rect 19484 8916 19490 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19628 8956 19656 9052
rect 25792 9036 25820 9064
rect 31662 9052 31668 9104
rect 31720 9092 31726 9104
rect 32030 9092 32036 9104
rect 31720 9064 32036 9092
rect 31720 9052 31726 9064
rect 32030 9052 32036 9064
rect 32088 9052 32094 9104
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 20119 8996 22293 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 22281 8987 22339 8993
rect 22756 8996 23765 9024
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19628 8928 19717 8956
rect 19521 8919 19579 8925
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19794 8916 19800 8968
rect 19852 8916 19858 8968
rect 21542 8956 21548 8968
rect 21206 8928 21548 8956
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8956 22155 8959
rect 22370 8956 22376 8968
rect 22143 8928 22376 8956
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 22646 8916 22652 8968
rect 22704 8956 22710 8968
rect 22756 8965 22784 8996
rect 23753 8993 23765 8996
rect 23799 9024 23811 9027
rect 23934 9024 23940 9036
rect 23799 8996 23940 9024
rect 23799 8993 23811 8996
rect 23753 8987 23811 8993
rect 23934 8984 23940 8996
rect 23992 9024 23998 9036
rect 24397 9027 24455 9033
rect 24397 9024 24409 9027
rect 23992 8996 24409 9024
rect 23992 8984 23998 8996
rect 24397 8993 24409 8996
rect 24443 8993 24455 9027
rect 24397 8987 24455 8993
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 25501 9027 25559 9033
rect 25501 9024 25513 9027
rect 24912 8996 25513 9024
rect 24912 8984 24918 8996
rect 25501 8993 25513 8996
rect 25547 8993 25559 9027
rect 25501 8987 25559 8993
rect 25774 8984 25780 9036
rect 25832 9024 25838 9036
rect 26789 9027 26847 9033
rect 26789 9024 26801 9027
rect 25832 8996 26801 9024
rect 25832 8984 25838 8996
rect 26789 8993 26801 8996
rect 26835 9024 26847 9027
rect 27430 9024 27436 9036
rect 26835 8996 27436 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 27430 8984 27436 8996
rect 27488 8984 27494 9036
rect 28074 8984 28080 9036
rect 28132 8984 28138 9036
rect 29822 9024 29828 9036
rect 28920 8996 29828 9024
rect 22741 8959 22799 8965
rect 22741 8956 22753 8959
rect 22704 8928 22753 8956
rect 22704 8916 22710 8928
rect 22741 8925 22753 8928
rect 22787 8925 22799 8959
rect 22741 8919 22799 8925
rect 22830 8916 22836 8968
rect 22888 8956 22894 8968
rect 22888 8928 23152 8956
rect 22888 8916 22894 8928
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 16850 8888 16856 8900
rect 16347 8860 16856 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 17494 8848 17500 8900
rect 17552 8848 17558 8900
rect 19061 8891 19119 8897
rect 19061 8888 19073 8891
rect 18432 8860 19073 8888
rect 15657 8823 15715 8829
rect 15657 8820 15669 8823
rect 15436 8792 15669 8820
rect 15436 8780 15442 8792
rect 15657 8789 15669 8792
rect 15703 8789 15715 8823
rect 15657 8783 15715 8789
rect 15838 8780 15844 8832
rect 15896 8780 15902 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 18432 8829 18460 8860
rect 19061 8857 19073 8860
rect 19107 8888 19119 8891
rect 20162 8888 20168 8900
rect 19107 8860 20168 8888
rect 19107 8857 19119 8860
rect 19061 8851 19119 8857
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 21637 8891 21695 8897
rect 21637 8888 21649 8891
rect 21376 8860 21649 8888
rect 16209 8823 16267 8829
rect 16209 8820 16221 8823
rect 15988 8792 16221 8820
rect 15988 8780 15994 8792
rect 16209 8789 16221 8792
rect 16255 8789 16267 8823
rect 16209 8783 16267 8789
rect 18417 8823 18475 8829
rect 18417 8789 18429 8823
rect 18463 8789 18475 8823
rect 18417 8783 18475 8789
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 18564 8792 18705 8820
rect 18564 8780 18570 8792
rect 18693 8789 18705 8792
rect 18739 8789 18751 8823
rect 18693 8783 18751 8789
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 21376 8820 21404 8860
rect 21637 8857 21649 8860
rect 21683 8888 21695 8891
rect 21726 8888 21732 8900
rect 21683 8860 21732 8888
rect 21683 8857 21695 8860
rect 21637 8851 21695 8857
rect 21726 8848 21732 8860
rect 21784 8848 21790 8900
rect 19751 8792 21404 8820
rect 22572 8820 22600 8916
rect 23124 8897 23152 8928
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 23385 8959 23443 8965
rect 23385 8956 23397 8959
rect 23256 8928 23397 8956
rect 23256 8916 23262 8928
rect 23385 8925 23397 8928
rect 23431 8925 23443 8959
rect 23385 8919 23443 8925
rect 25222 8916 25228 8968
rect 25280 8916 25286 8968
rect 25317 8959 25375 8965
rect 25317 8925 25329 8959
rect 25363 8956 25375 8959
rect 25593 8959 25651 8965
rect 25363 8928 25544 8956
rect 25363 8925 25375 8928
rect 25317 8919 25375 8925
rect 25516 8900 25544 8928
rect 25593 8925 25605 8959
rect 25639 8956 25651 8959
rect 26605 8959 26663 8965
rect 25639 8928 26096 8956
rect 25639 8925 25651 8928
rect 25593 8919 25651 8925
rect 23109 8891 23167 8897
rect 23109 8857 23121 8891
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 23308 8860 24348 8888
rect 23308 8820 23336 8860
rect 22572 8792 23336 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 23382 8780 23388 8832
rect 23440 8820 23446 8832
rect 24320 8829 24348 8860
rect 24486 8848 24492 8900
rect 24544 8888 24550 8900
rect 25041 8891 25099 8897
rect 25041 8888 25053 8891
rect 24544 8860 25053 8888
rect 24544 8848 24550 8860
rect 25041 8857 25053 8860
rect 25087 8857 25099 8891
rect 25041 8851 25099 8857
rect 25498 8848 25504 8900
rect 25556 8848 25562 8900
rect 24121 8823 24179 8829
rect 24121 8820 24133 8823
rect 23440 8792 24133 8820
rect 23440 8780 23446 8792
rect 24121 8789 24133 8792
rect 24167 8789 24179 8823
rect 24121 8783 24179 8789
rect 24305 8823 24363 8829
rect 24305 8789 24317 8823
rect 24351 8789 24363 8823
rect 24305 8783 24363 8789
rect 24394 8780 24400 8832
rect 24452 8820 24458 8832
rect 24765 8823 24823 8829
rect 24765 8820 24777 8823
rect 24452 8792 24777 8820
rect 24452 8780 24458 8792
rect 24765 8789 24777 8792
rect 24811 8789 24823 8823
rect 24765 8783 24823 8789
rect 24946 8780 24952 8832
rect 25004 8780 25010 8832
rect 25314 8780 25320 8832
rect 25372 8820 25378 8832
rect 25608 8820 25636 8919
rect 25372 8792 25636 8820
rect 25372 8780 25378 8792
rect 25958 8780 25964 8832
rect 26016 8780 26022 8832
rect 26068 8820 26096 8928
rect 26605 8925 26617 8959
rect 26651 8956 26663 8959
rect 28092 8956 28120 8984
rect 28920 8965 28948 8996
rect 29822 8984 29828 8996
rect 29880 8984 29886 9036
rect 30282 8984 30288 9036
rect 30340 9024 30346 9036
rect 31294 9024 31300 9036
rect 30340 8996 31300 9024
rect 30340 8984 30346 8996
rect 31294 8984 31300 8996
rect 31352 8984 31358 9036
rect 31478 8984 31484 9036
rect 31536 9024 31542 9036
rect 31846 9024 31852 9036
rect 31536 8996 31852 9024
rect 31536 8984 31542 8996
rect 31846 8984 31852 8996
rect 31904 8984 31910 9036
rect 31941 9027 31999 9033
rect 31941 8993 31953 9027
rect 31987 9024 31999 9027
rect 32140 9024 32168 9132
rect 32766 9120 32772 9132
rect 32824 9120 32830 9172
rect 33134 9120 33140 9172
rect 33192 9160 33198 9172
rect 33410 9160 33416 9172
rect 33192 9132 33416 9160
rect 33192 9120 33198 9132
rect 33410 9120 33416 9132
rect 33468 9160 33474 9172
rect 33597 9163 33655 9169
rect 33597 9160 33609 9163
rect 33468 9132 33609 9160
rect 33468 9120 33474 9132
rect 33597 9129 33609 9132
rect 33643 9129 33655 9163
rect 33597 9123 33655 9129
rect 33962 9120 33968 9172
rect 34020 9160 34026 9172
rect 35894 9160 35900 9172
rect 34020 9132 35900 9160
rect 34020 9120 34026 9132
rect 35894 9120 35900 9132
rect 35952 9120 35958 9172
rect 35986 9120 35992 9172
rect 36044 9160 36050 9172
rect 36081 9163 36139 9169
rect 36081 9160 36093 9163
rect 36044 9132 36093 9160
rect 36044 9120 36050 9132
rect 36081 9129 36093 9132
rect 36127 9129 36139 9163
rect 36081 9123 36139 9129
rect 36170 9120 36176 9172
rect 36228 9160 36234 9172
rect 36357 9163 36415 9169
rect 36357 9160 36369 9163
rect 36228 9132 36369 9160
rect 36228 9120 36234 9132
rect 36357 9129 36369 9132
rect 36403 9129 36415 9163
rect 38010 9160 38016 9172
rect 36357 9123 36415 9129
rect 36832 9132 38016 9160
rect 32214 9052 32220 9104
rect 32272 9092 32278 9104
rect 34330 9092 34336 9104
rect 32272 9064 32904 9092
rect 32272 9052 32278 9064
rect 31987 8996 32168 9024
rect 31987 8993 31999 8996
rect 31941 8987 31999 8993
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 32876 9033 32904 9064
rect 32968 9064 34336 9092
rect 32968 9033 32996 9064
rect 34330 9052 34336 9064
rect 34388 9052 34394 9104
rect 34882 9052 34888 9104
rect 34940 9052 34946 9104
rect 34974 9052 34980 9104
rect 35032 9092 35038 9104
rect 36541 9095 36599 9101
rect 36541 9092 36553 9095
rect 35032 9064 36553 9092
rect 35032 9052 35038 9064
rect 36541 9061 36553 9064
rect 36587 9061 36599 9095
rect 36541 9055 36599 9061
rect 32677 9027 32735 9033
rect 32677 9024 32689 9027
rect 32456 8996 32689 9024
rect 32456 8984 32462 8996
rect 32677 8993 32689 8996
rect 32723 8993 32735 9027
rect 32677 8987 32735 8993
rect 32861 9027 32919 9033
rect 32861 8993 32873 9027
rect 32907 8993 32919 9027
rect 32861 8987 32919 8993
rect 32953 9027 33011 9033
rect 32953 8993 32965 9027
rect 32999 8993 33011 9027
rect 32953 8987 33011 8993
rect 26651 8928 28120 8956
rect 28905 8959 28963 8965
rect 26651 8925 26663 8928
rect 26605 8919 26663 8925
rect 28905 8925 28917 8959
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 29457 8959 29515 8965
rect 29457 8925 29469 8959
rect 29503 8925 29515 8959
rect 29457 8919 29515 8925
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8956 31723 8959
rect 32217 8959 32275 8965
rect 31711 8928 32168 8956
rect 31711 8925 31723 8928
rect 31665 8919 31723 8925
rect 26510 8848 26516 8900
rect 26568 8848 26574 8900
rect 26878 8848 26884 8900
rect 26936 8848 26942 8900
rect 26970 8848 26976 8900
rect 27028 8888 27034 8900
rect 27982 8888 27988 8900
rect 27028 8860 27988 8888
rect 27028 8848 27034 8860
rect 27982 8848 27988 8860
rect 28040 8848 28046 8900
rect 29472 8888 29500 8919
rect 28368 8860 29500 8888
rect 26896 8820 26924 8848
rect 26068 8792 26924 8820
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 28368 8820 28396 8860
rect 30006 8848 30012 8900
rect 30064 8888 30070 8900
rect 31757 8891 31815 8897
rect 31757 8888 31769 8891
rect 30064 8860 30222 8888
rect 31220 8860 31769 8888
rect 30064 8848 30070 8860
rect 27672 8792 28396 8820
rect 27672 8780 27678 8792
rect 28442 8780 28448 8832
rect 28500 8820 28506 8832
rect 28718 8820 28724 8832
rect 28500 8792 28724 8820
rect 28500 8780 28506 8792
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 29178 8780 29184 8832
rect 29236 8820 29242 8832
rect 30098 8820 30104 8832
rect 29236 8792 30104 8820
rect 29236 8780 29242 8792
rect 30098 8780 30104 8792
rect 30156 8780 30162 8832
rect 30374 8780 30380 8832
rect 30432 8820 30438 8832
rect 31220 8829 31248 8860
rect 31757 8857 31769 8860
rect 31803 8857 31815 8891
rect 32140 8888 32168 8928
rect 32217 8925 32229 8959
rect 32263 8956 32275 8959
rect 32582 8956 32588 8968
rect 32263 8928 32588 8956
rect 32263 8925 32275 8928
rect 32217 8919 32275 8925
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 32769 8959 32827 8965
rect 32769 8925 32781 8959
rect 32815 8925 32827 8959
rect 32876 8956 32904 8987
rect 33226 8984 33232 9036
rect 33284 9024 33290 9036
rect 33594 9024 33600 9036
rect 33284 8996 33600 9024
rect 33284 8984 33290 8996
rect 33594 8984 33600 8996
rect 33652 8984 33658 9036
rect 34422 8984 34428 9036
rect 34480 9024 34486 9036
rect 34701 9027 34759 9033
rect 34701 9024 34713 9027
rect 34480 8996 34713 9024
rect 34480 8984 34486 8996
rect 34701 8993 34713 8996
rect 34747 9024 34759 9027
rect 35526 9024 35532 9036
rect 34747 8996 35532 9024
rect 34747 8993 34759 8996
rect 34701 8987 34759 8993
rect 35526 8984 35532 8996
rect 35584 8984 35590 9036
rect 36832 9024 36860 9132
rect 38010 9120 38016 9132
rect 38068 9160 38074 9172
rect 38473 9163 38531 9169
rect 38473 9160 38485 9163
rect 38068 9132 38485 9160
rect 38068 9120 38074 9132
rect 38473 9129 38485 9132
rect 38519 9129 38531 9163
rect 38473 9123 38531 9129
rect 39758 9120 39764 9172
rect 39816 9120 39822 9172
rect 43165 9163 43223 9169
rect 43165 9129 43177 9163
rect 43211 9160 43223 9163
rect 43254 9160 43260 9172
rect 43211 9132 43260 9160
rect 43211 9129 43223 9132
rect 43165 9123 43223 9129
rect 43254 9120 43260 9132
rect 43312 9160 43318 9172
rect 43717 9163 43775 9169
rect 43717 9160 43729 9163
rect 43312 9132 43729 9160
rect 43312 9120 43318 9132
rect 43717 9129 43729 9132
rect 43763 9129 43775 9163
rect 43717 9123 43775 9129
rect 38565 9095 38623 9101
rect 38565 9061 38577 9095
rect 38611 9061 38623 9095
rect 38565 9055 38623 9061
rect 35636 8996 36860 9024
rect 33505 8959 33563 8965
rect 33505 8956 33517 8959
rect 32876 8928 33517 8956
rect 32769 8919 32827 8925
rect 33505 8925 33517 8928
rect 33551 8925 33563 8959
rect 33505 8919 33563 8925
rect 35345 8959 35403 8965
rect 35345 8925 35357 8959
rect 35391 8956 35403 8959
rect 35434 8956 35440 8968
rect 35391 8928 35440 8956
rect 35391 8925 35403 8928
rect 35345 8919 35403 8925
rect 32784 8888 32812 8919
rect 35434 8916 35440 8928
rect 35492 8916 35498 8968
rect 33042 8888 33048 8900
rect 32140 8860 32720 8888
rect 32784 8860 33048 8888
rect 31757 8851 31815 8857
rect 31205 8823 31263 8829
rect 31205 8820 31217 8823
rect 30432 8792 31217 8820
rect 30432 8780 30438 8792
rect 31205 8789 31217 8792
rect 31251 8789 31263 8823
rect 31205 8783 31263 8789
rect 31297 8823 31355 8829
rect 31297 8789 31309 8823
rect 31343 8820 31355 8823
rect 31478 8820 31484 8832
rect 31343 8792 31484 8820
rect 31343 8789 31355 8792
rect 31297 8783 31355 8789
rect 31478 8780 31484 8792
rect 31536 8780 31542 8832
rect 32122 8780 32128 8832
rect 32180 8820 32186 8832
rect 32309 8823 32367 8829
rect 32309 8820 32321 8823
rect 32180 8792 32321 8820
rect 32180 8780 32186 8792
rect 32309 8789 32321 8792
rect 32355 8789 32367 8823
rect 32309 8783 32367 8789
rect 32490 8780 32496 8832
rect 32548 8780 32554 8832
rect 32692 8820 32720 8860
rect 33042 8848 33048 8860
rect 33100 8848 33106 8900
rect 33594 8848 33600 8900
rect 33652 8848 33658 8900
rect 34330 8848 34336 8900
rect 34388 8888 34394 8900
rect 34974 8888 34980 8900
rect 34388 8860 34980 8888
rect 34388 8848 34394 8860
rect 34974 8848 34980 8860
rect 35032 8848 35038 8900
rect 35636 8888 35664 8996
rect 36998 8984 37004 9036
rect 37056 8984 37062 9036
rect 37090 8984 37096 9036
rect 37148 9024 37154 9036
rect 38580 9024 38608 9055
rect 39776 9024 39804 9120
rect 37148 8996 38608 9024
rect 39040 8996 39804 9024
rect 37148 8984 37154 8996
rect 36538 8956 36544 8968
rect 36096 8928 36544 8956
rect 35176 8860 35664 8888
rect 35713 8891 35771 8897
rect 33226 8820 33232 8832
rect 32692 8792 33232 8820
rect 33226 8780 33232 8792
rect 33284 8780 33290 8832
rect 33612 8820 33640 8848
rect 34057 8823 34115 8829
rect 34057 8820 34069 8823
rect 33612 8792 34069 8820
rect 34057 8789 34069 8792
rect 34103 8789 34115 8823
rect 34057 8783 34115 8789
rect 34422 8780 34428 8832
rect 34480 8780 34486 8832
rect 34517 8823 34575 8829
rect 34517 8789 34529 8823
rect 34563 8820 34575 8823
rect 35176 8820 35204 8860
rect 35713 8857 35725 8891
rect 35759 8888 35771 8891
rect 35802 8888 35808 8900
rect 35759 8860 35808 8888
rect 35759 8857 35771 8860
rect 35713 8851 35771 8857
rect 35802 8848 35808 8860
rect 35860 8848 35866 8900
rect 35929 8891 35987 8897
rect 35929 8857 35941 8891
rect 35975 8888 35987 8891
rect 36096 8888 36124 8928
rect 36538 8916 36544 8928
rect 36596 8916 36602 8968
rect 36630 8916 36636 8968
rect 36688 8956 36694 8968
rect 36725 8959 36783 8965
rect 36725 8956 36737 8959
rect 36688 8928 36737 8956
rect 36688 8916 36694 8928
rect 36725 8925 36737 8928
rect 36771 8925 36783 8959
rect 36725 8919 36783 8925
rect 38286 8916 38292 8968
rect 38344 8956 38350 8968
rect 39040 8965 39068 8996
rect 40586 8984 40592 9036
rect 40644 9024 40650 9036
rect 40644 8996 41276 9024
rect 40644 8984 40650 8996
rect 38749 8959 38807 8965
rect 38749 8956 38761 8959
rect 38344 8928 38761 8956
rect 38344 8916 38350 8928
rect 38749 8925 38761 8928
rect 38795 8925 38807 8959
rect 38749 8919 38807 8925
rect 39025 8959 39083 8965
rect 39025 8925 39037 8959
rect 39071 8925 39083 8959
rect 39025 8919 39083 8925
rect 39666 8916 39672 8968
rect 39724 8916 39730 8968
rect 39758 8916 39764 8968
rect 39816 8916 39822 8968
rect 39853 8959 39911 8965
rect 39853 8925 39865 8959
rect 39899 8925 39911 8959
rect 41248 8956 41276 8996
rect 41506 8956 41512 8968
rect 41248 8942 41512 8956
rect 41262 8928 41512 8942
rect 39853 8919 39911 8925
rect 35975 8860 36124 8888
rect 35975 8857 35987 8860
rect 35929 8851 35987 8857
rect 36170 8848 36176 8900
rect 36228 8848 36234 8900
rect 36389 8891 36447 8897
rect 36389 8857 36401 8891
rect 36435 8888 36447 8891
rect 36556 8888 36584 8916
rect 36435 8860 36584 8888
rect 36435 8857 36447 8860
rect 36389 8851 36447 8857
rect 37458 8848 37464 8900
rect 37516 8848 37522 8900
rect 39684 8888 39712 8916
rect 39868 8888 39896 8919
rect 41506 8916 41512 8928
rect 41564 8916 41570 8968
rect 38304 8860 39436 8888
rect 39684 8860 39896 8888
rect 40129 8891 40187 8897
rect 34563 8792 35204 8820
rect 35253 8823 35311 8829
rect 34563 8789 34575 8792
rect 34517 8783 34575 8789
rect 35253 8789 35265 8823
rect 35299 8820 35311 8823
rect 35618 8820 35624 8832
rect 35299 8792 35624 8820
rect 35299 8789 35311 8792
rect 35253 8783 35311 8789
rect 35618 8780 35624 8792
rect 35676 8780 35682 8832
rect 36538 8780 36544 8832
rect 36596 8820 36602 8832
rect 38304 8820 38332 8860
rect 36596 8792 38332 8820
rect 36596 8780 36602 8792
rect 38838 8780 38844 8832
rect 38896 8780 38902 8832
rect 39408 8829 39436 8860
rect 40129 8857 40141 8891
rect 40175 8857 40187 8891
rect 40129 8851 40187 8857
rect 41693 8891 41751 8897
rect 41693 8857 41705 8891
rect 41739 8888 41751 8891
rect 42518 8888 42524 8900
rect 41739 8860 42524 8888
rect 41739 8857 41751 8860
rect 41693 8851 41751 8857
rect 39393 8823 39451 8829
rect 39393 8789 39405 8823
rect 39439 8789 39451 8823
rect 39393 8783 39451 8789
rect 39577 8823 39635 8829
rect 39577 8789 39589 8823
rect 39623 8820 39635 8823
rect 40144 8820 40172 8851
rect 42518 8848 42524 8860
rect 42576 8848 42582 8900
rect 39623 8792 40172 8820
rect 39623 8789 39635 8792
rect 39577 8783 39635 8789
rect 40954 8780 40960 8832
rect 41012 8820 41018 8832
rect 41601 8823 41659 8829
rect 41601 8820 41613 8823
rect 41012 8792 41613 8820
rect 41012 8780 41018 8792
rect 41601 8789 41613 8792
rect 41647 8820 41659 8823
rect 41874 8820 41880 8832
rect 41647 8792 41880 8820
rect 41647 8789 41659 8792
rect 41601 8783 41659 8789
rect 41874 8780 41880 8792
rect 41932 8780 41938 8832
rect 44177 8823 44235 8829
rect 44177 8789 44189 8823
rect 44223 8820 44235 8823
rect 44542 8820 44548 8832
rect 44223 8792 44548 8820
rect 44223 8789 44235 8792
rect 44177 8783 44235 8789
rect 44542 8780 44548 8792
rect 44600 8780 44606 8832
rect 44910 8780 44916 8832
rect 44968 8780 44974 8832
rect 460 8730 45540 8752
rect 460 8678 6070 8730
rect 6122 8678 6134 8730
rect 6186 8678 6198 8730
rect 6250 8678 6262 8730
rect 6314 8678 6326 8730
rect 6378 8678 11070 8730
rect 11122 8678 11134 8730
rect 11186 8678 11198 8730
rect 11250 8678 11262 8730
rect 11314 8678 11326 8730
rect 11378 8678 16070 8730
rect 16122 8678 16134 8730
rect 16186 8678 16198 8730
rect 16250 8678 16262 8730
rect 16314 8678 16326 8730
rect 16378 8678 21070 8730
rect 21122 8678 21134 8730
rect 21186 8678 21198 8730
rect 21250 8678 21262 8730
rect 21314 8678 21326 8730
rect 21378 8678 26070 8730
rect 26122 8678 26134 8730
rect 26186 8678 26198 8730
rect 26250 8678 26262 8730
rect 26314 8678 26326 8730
rect 26378 8678 31070 8730
rect 31122 8678 31134 8730
rect 31186 8678 31198 8730
rect 31250 8678 31262 8730
rect 31314 8678 31326 8730
rect 31378 8678 36070 8730
rect 36122 8678 36134 8730
rect 36186 8678 36198 8730
rect 36250 8678 36262 8730
rect 36314 8678 36326 8730
rect 36378 8678 41070 8730
rect 41122 8678 41134 8730
rect 41186 8678 41198 8730
rect 41250 8678 41262 8730
rect 41314 8678 41326 8730
rect 41378 8678 45540 8730
rect 460 8656 45540 8678
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6052 8588 6469 8616
rect 6052 8576 6058 8588
rect 6457 8585 6469 8588
rect 6503 8616 6515 8619
rect 6638 8616 6644 8628
rect 6503 8588 6644 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7650 8576 7656 8628
rect 7708 8576 7714 8628
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8202 8616 8208 8628
rect 8159 8588 8208 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8202 8576 8208 8588
rect 8260 8616 8266 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 8260 8588 8769 8616
rect 8260 8576 8266 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 11057 8619 11115 8625
rect 10192 8588 11008 8616
rect 10192 8576 10198 8588
rect 8938 8508 8944 8560
rect 8996 8548 9002 8560
rect 9217 8551 9275 8557
rect 9217 8548 9229 8551
rect 8996 8520 9229 8548
rect 8996 8508 9002 8520
rect 9217 8517 9229 8520
rect 9263 8517 9275 8551
rect 9217 8511 9275 8517
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10980 8480 11008 8588
rect 11057 8585 11069 8619
rect 11103 8616 11115 8619
rect 11238 8616 11244 8628
rect 11103 8588 11244 8616
rect 11103 8585 11115 8588
rect 11057 8579 11115 8585
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 12066 8576 12072 8628
rect 12124 8576 12130 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13320 8588 15056 8616
rect 13320 8576 13326 8588
rect 11333 8551 11391 8557
rect 11333 8548 11345 8551
rect 11164 8520 11345 8548
rect 11164 8489 11192 8520
rect 11333 8517 11345 8520
rect 11379 8517 11391 8551
rect 11790 8548 11796 8560
rect 11333 8511 11391 8517
rect 11440 8520 11796 8548
rect 11440 8489 11468 8520
rect 11790 8508 11796 8520
rect 11848 8508 11854 8560
rect 12084 8548 12112 8576
rect 13078 8548 13084 8560
rect 12084 8520 12296 8548
rect 12268 8489 12296 8520
rect 12912 8520 13084 8548
rect 11149 8483 11207 8489
rect 10980 8452 11100 8480
rect 10873 8443 10931 8449
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 5583 8384 6837 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6871 8384 7389 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7377 8381 7389 8384
rect 7423 8412 7435 8415
rect 8478 8412 8484 8424
rect 7423 8384 8484 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 8478 8372 8484 8384
rect 8536 8412 8542 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8536 8384 8953 8412
rect 8536 8372 8542 8384
rect 8941 8381 8953 8384
rect 8987 8412 8999 8415
rect 9306 8412 9312 8424
rect 8987 8384 9312 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 10888 8412 10916 8443
rect 9640 8384 10916 8412
rect 11072 8412 11100 8452
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8449 11483 8483
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11425 8443 11483 8449
rect 11624 8452 11989 8480
rect 11256 8412 11284 8443
rect 11072 8384 11284 8412
rect 9640 8372 9646 8384
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10689 8347 10747 8353
rect 10689 8344 10701 8347
rect 10468 8316 10701 8344
rect 10468 8304 10474 8316
rect 10689 8313 10701 8316
rect 10735 8313 10747 8347
rect 10888 8344 10916 8384
rect 11624 8344 11652 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12434 8480 12440 8492
rect 12253 8443 12311 8449
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 11992 8412 12020 8443
rect 12176 8412 12204 8443
rect 12406 8440 12440 8480
rect 12492 8440 12498 8492
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8480 12679 8483
rect 12710 8480 12716 8492
rect 12667 8452 12716 8480
rect 12667 8449 12679 8452
rect 12621 8443 12679 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 12912 8480 12940 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 13180 8551 13238 8557
rect 13180 8517 13192 8551
rect 13226 8548 13238 8551
rect 13446 8548 13452 8560
rect 13226 8520 13452 8548
rect 13226 8517 13238 8520
rect 13180 8511 13238 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 13630 8508 13636 8560
rect 13688 8508 13694 8560
rect 15028 8548 15056 8588
rect 15102 8576 15108 8628
rect 15160 8576 15166 8628
rect 17218 8616 17224 8628
rect 15764 8588 17224 8616
rect 15764 8557 15792 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 18046 8616 18052 8628
rect 17359 8588 18052 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 18046 8576 18052 8588
rect 18104 8616 18110 8628
rect 18104 8588 19012 8616
rect 18104 8576 18110 8588
rect 15749 8551 15807 8557
rect 15749 8548 15761 8551
rect 15028 8520 15761 8548
rect 15749 8517 15761 8520
rect 15795 8517 15807 8551
rect 15749 8511 15807 8517
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 17681 8551 17739 8557
rect 16632 8520 17448 8548
rect 16632 8508 16638 8520
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 12851 8452 12940 8480
rect 14384 8452 14749 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12406 8412 12434 8440
rect 11992 8384 12112 8412
rect 12176 8384 12434 8412
rect 10888 8316 11652 8344
rect 11716 8344 11744 8372
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11716 8316 11989 8344
rect 10689 8307 10747 8313
rect 11977 8313 11989 8316
rect 12023 8313 12035 8347
rect 12084 8344 12112 8384
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12584 8384 12909 8412
rect 12584 8372 12590 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 14182 8412 14188 8424
rect 13688 8384 14188 8412
rect 13688 8372 13694 8384
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 12802 8344 12808 8356
rect 12084 8316 12808 8344
rect 11977 8307 12035 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 14384 8344 14412 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15344 8452 16313 8480
rect 15344 8440 15350 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16666 8480 16672 8492
rect 16531 8452 16672 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17218 8480 17224 8492
rect 16991 8452 17224 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17420 8489 17448 8520
rect 17681 8517 17693 8551
rect 17727 8548 17739 8551
rect 17954 8548 17960 8560
rect 17727 8520 17960 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 18984 8548 19012 8588
rect 19150 8576 19156 8628
rect 19208 8576 19214 8628
rect 20254 8616 20260 8628
rect 19260 8588 20260 8616
rect 19260 8548 19288 8588
rect 20254 8576 20260 8588
rect 20312 8616 20318 8628
rect 21542 8616 21548 8628
rect 20312 8588 21548 8616
rect 20312 8576 20318 8588
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 25222 8616 25228 8628
rect 21867 8588 25228 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 25222 8576 25228 8588
rect 25280 8576 25286 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27249 8619 27307 8625
rect 26568 8588 27200 8616
rect 26568 8576 26574 8588
rect 18906 8520 19288 8548
rect 19518 8508 19524 8560
rect 19576 8548 19582 8560
rect 19978 8548 19984 8560
rect 19576 8520 19984 8548
rect 19576 8508 19582 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 20364 8520 20729 8548
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 17368 8452 17417 8480
rect 17368 8440 17374 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19610 8480 19616 8492
rect 19475 8452 19616 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 14829 8415 14887 8421
rect 14829 8412 14841 8415
rect 14660 8384 14841 8412
rect 14660 8353 14688 8384
rect 14829 8381 14841 8384
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15930 8412 15936 8424
rect 15068 8384 15936 8412
rect 15068 8372 15074 8384
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 19260 8412 19288 8443
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 20364 8480 20392 8520
rect 20717 8517 20729 8520
rect 20763 8548 20775 8551
rect 20806 8548 20812 8560
rect 20763 8520 20812 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 21637 8551 21695 8557
rect 21637 8517 21649 8551
rect 21683 8548 21695 8551
rect 22094 8548 22100 8560
rect 21683 8520 22100 8548
rect 21683 8517 21695 8520
rect 21637 8511 21695 8517
rect 22094 8508 22100 8520
rect 22152 8548 22158 8560
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 22152 8520 22385 8548
rect 22152 8508 22158 8520
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 22462 8508 22468 8560
rect 22520 8548 22526 8560
rect 22520 8520 22968 8548
rect 22520 8508 22526 8520
rect 19720 8452 20392 8480
rect 19720 8412 19748 8452
rect 20622 8440 20628 8492
rect 20680 8440 20686 8492
rect 22940 8489 22968 8520
rect 23106 8508 23112 8560
rect 23164 8508 23170 8560
rect 24394 8548 24400 8560
rect 23676 8520 24400 8548
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22925 8483 22983 8489
rect 22327 8452 22416 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22388 8424 22416 8452
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 23124 8480 23152 8508
rect 23385 8483 23443 8489
rect 23385 8480 23397 8483
rect 23124 8452 23397 8480
rect 22925 8443 22983 8449
rect 23385 8449 23397 8452
rect 23431 8449 23443 8483
rect 23385 8443 23443 8449
rect 17512 8384 19196 8412
rect 19260 8384 19748 8412
rect 14200 8316 14412 8344
rect 14645 8347 14703 8353
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 10778 8276 10784 8288
rect 9272 8248 10784 8276
rect 9272 8236 9278 8248
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 10870 8236 10876 8288
rect 10928 8236 10934 8288
rect 11882 8236 11888 8288
rect 11940 8236 11946 8288
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 14200 8276 14228 8316
rect 14645 8313 14657 8347
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 13228 8248 14228 8276
rect 13228 8236 13234 8248
rect 14274 8236 14280 8288
rect 14332 8276 14338 8288
rect 14660 8276 14688 8307
rect 14734 8304 14740 8356
rect 14792 8344 14798 8356
rect 17512 8344 17540 8384
rect 14792 8316 17540 8344
rect 19168 8344 19196 8384
rect 19886 8372 19892 8424
rect 19944 8372 19950 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20162 8412 20168 8424
rect 20027 8384 20168 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20272 8384 20913 8412
rect 19610 8344 19616 8356
rect 19168 8316 19616 8344
rect 14792 8304 14798 8316
rect 19610 8304 19616 8316
rect 19668 8304 19674 8356
rect 19904 8344 19932 8372
rect 20272 8344 20300 8384
rect 20901 8381 20913 8384
rect 20947 8412 20959 8415
rect 22002 8412 22008 8424
rect 20947 8384 22008 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22370 8372 22376 8424
rect 22428 8372 22434 8424
rect 22465 8415 22523 8421
rect 22465 8381 22477 8415
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 20714 8344 20720 8356
rect 19904 8316 20300 8344
rect 20364 8316 20720 8344
rect 14332 8248 14688 8276
rect 14332 8236 14338 8248
rect 14918 8236 14924 8288
rect 14976 8236 14982 8288
rect 15378 8236 15384 8288
rect 15436 8236 15442 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 16080 8248 16405 8276
rect 16080 8236 16086 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16393 8239 16451 8245
rect 16758 8236 16764 8288
rect 16816 8236 16822 8288
rect 19337 8279 19395 8285
rect 19337 8245 19349 8279
rect 19383 8276 19395 8279
rect 19518 8276 19524 8288
rect 19383 8248 19524 8276
rect 19383 8245 19395 8248
rect 19337 8239 19395 8245
rect 19518 8236 19524 8248
rect 19576 8236 19582 8288
rect 20162 8236 20168 8288
rect 20220 8236 20226 8288
rect 20257 8279 20315 8285
rect 20257 8245 20269 8279
rect 20303 8276 20315 8279
rect 20364 8276 20392 8316
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 20990 8304 20996 8356
rect 21048 8344 21054 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 21048 8316 21281 8344
rect 21048 8304 21054 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21910 8304 21916 8356
rect 21968 8304 21974 8356
rect 22020 8344 22048 8372
rect 22480 8344 22508 8375
rect 23474 8372 23480 8424
rect 23532 8372 23538 8424
rect 23676 8421 23704 8520
rect 24394 8508 24400 8520
rect 24452 8508 24458 8560
rect 26421 8551 26479 8557
rect 26421 8517 26433 8551
rect 26467 8548 26479 8551
rect 26786 8548 26792 8560
rect 26467 8520 26792 8548
rect 26467 8517 26479 8520
rect 26421 8511 26479 8517
rect 26786 8508 26792 8520
rect 26844 8508 26850 8560
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8449 23903 8483
rect 25682 8480 25688 8492
rect 25530 8452 25688 8480
rect 23845 8443 23903 8449
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8381 23719 8415
rect 23661 8375 23719 8381
rect 22020 8316 22508 8344
rect 20303 8248 20392 8276
rect 21637 8279 21695 8285
rect 20303 8245 20315 8248
rect 20257 8239 20315 8245
rect 21637 8245 21649 8279
rect 21683 8276 21695 8279
rect 22020 8276 22048 8316
rect 22738 8304 22744 8356
rect 22796 8304 22802 8356
rect 23860 8344 23888 8443
rect 25682 8440 25688 8452
rect 25740 8480 25746 8492
rect 25740 8452 27016 8480
rect 25740 8440 25746 8452
rect 26988 8424 27016 8452
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 23032 8316 23888 8344
rect 23032 8285 23060 8316
rect 24136 8288 24164 8375
rect 24394 8372 24400 8424
rect 24452 8372 24458 8424
rect 24762 8372 24768 8424
rect 24820 8412 24826 8424
rect 25958 8412 25964 8424
rect 24820 8384 25964 8412
rect 24820 8372 24826 8384
rect 25958 8372 25964 8384
rect 26016 8412 26022 8424
rect 26145 8415 26203 8421
rect 26145 8412 26157 8415
rect 26016 8384 26157 8412
rect 26016 8372 26022 8384
rect 26145 8381 26157 8384
rect 26191 8381 26203 8415
rect 26145 8375 26203 8381
rect 26160 8344 26188 8375
rect 26970 8372 26976 8424
rect 27028 8372 27034 8424
rect 27172 8344 27200 8588
rect 27249 8585 27261 8619
rect 27295 8616 27307 8619
rect 27295 8588 29592 8616
rect 27295 8585 27307 8588
rect 27249 8579 27307 8585
rect 27985 8551 28043 8557
rect 27985 8517 27997 8551
rect 28031 8548 28043 8551
rect 28258 8548 28264 8560
rect 28031 8520 28264 8548
rect 28031 8517 28043 8520
rect 27985 8511 28043 8517
rect 28258 8508 28264 8520
rect 28316 8508 28322 8560
rect 29564 8548 29592 8588
rect 29914 8576 29920 8628
rect 29972 8616 29978 8628
rect 30101 8619 30159 8625
rect 30101 8616 30113 8619
rect 29972 8588 30113 8616
rect 29972 8576 29978 8588
rect 30101 8585 30113 8588
rect 30147 8585 30159 8619
rect 30101 8579 30159 8585
rect 30945 8619 31003 8625
rect 30945 8585 30957 8619
rect 30991 8585 31003 8619
rect 30945 8579 31003 8585
rect 30466 8548 30472 8560
rect 29564 8520 30472 8548
rect 30466 8508 30472 8520
rect 30524 8508 30530 8560
rect 30742 8508 30748 8560
rect 30800 8508 30806 8560
rect 30834 8508 30840 8560
rect 30892 8548 30898 8560
rect 30960 8548 30988 8579
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32548 8588 32812 8616
rect 32548 8576 32554 8588
rect 30892 8520 30988 8548
rect 31573 8551 31631 8557
rect 30892 8508 30898 8520
rect 31573 8517 31585 8551
rect 31619 8548 31631 8551
rect 31662 8548 31668 8560
rect 31619 8520 31668 8548
rect 31619 8517 31631 8520
rect 31573 8511 31631 8517
rect 31662 8508 31668 8520
rect 31720 8508 31726 8560
rect 31846 8508 31852 8560
rect 31904 8548 31910 8560
rect 32784 8557 32812 8588
rect 33042 8576 33048 8628
rect 33100 8616 33106 8628
rect 34146 8616 34152 8628
rect 33100 8588 34152 8616
rect 33100 8576 33106 8588
rect 34146 8576 34152 8588
rect 34204 8616 34210 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 34204 8588 34253 8616
rect 34204 8576 34210 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 34330 8576 34336 8628
rect 34388 8576 34394 8628
rect 34514 8576 34520 8628
rect 34572 8616 34578 8628
rect 34572 8588 35112 8616
rect 34572 8576 34578 8588
rect 32769 8551 32827 8557
rect 31904 8520 32536 8548
rect 31904 8508 31910 8520
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 27614 8480 27620 8492
rect 27387 8452 27620 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 29733 8483 29791 8489
rect 27430 8372 27436 8424
rect 27488 8372 27494 8424
rect 28350 8412 28356 8424
rect 27816 8384 28356 8412
rect 27816 8344 27844 8384
rect 28350 8372 28356 8384
rect 28408 8372 28414 8424
rect 28534 8372 28540 8424
rect 28592 8412 28598 8424
rect 29104 8412 29132 8466
rect 29733 8449 29745 8483
rect 29779 8480 29791 8483
rect 29822 8480 29828 8492
rect 29779 8452 29828 8480
rect 29779 8449 29791 8452
rect 29733 8443 29791 8449
rect 29822 8440 29828 8452
rect 29880 8440 29886 8492
rect 30006 8440 30012 8492
rect 30064 8440 30070 8492
rect 30374 8440 30380 8492
rect 30432 8440 30438 8492
rect 30561 8483 30619 8489
rect 30561 8449 30573 8483
rect 30607 8480 30619 8483
rect 30650 8480 30656 8492
rect 30607 8452 30656 8480
rect 30607 8449 30619 8452
rect 30561 8443 30619 8449
rect 30650 8440 30656 8452
rect 30708 8440 30714 8492
rect 31386 8440 31392 8492
rect 31444 8480 31450 8492
rect 32033 8483 32091 8489
rect 32033 8480 32045 8483
rect 31444 8452 32045 8480
rect 31444 8440 31450 8452
rect 32033 8449 32045 8452
rect 32079 8480 32091 8483
rect 32398 8480 32404 8492
rect 32079 8452 32404 8480
rect 32079 8449 32091 8452
rect 32033 8443 32091 8449
rect 32398 8440 32404 8452
rect 32456 8440 32462 8492
rect 32508 8489 32536 8520
rect 32769 8517 32781 8551
rect 32815 8517 32827 8551
rect 34054 8548 34060 8560
rect 33994 8520 34060 8548
rect 32769 8511 32827 8517
rect 34054 8508 34060 8520
rect 34112 8548 34118 8560
rect 34532 8548 34560 8576
rect 34790 8548 34796 8560
rect 34112 8520 34560 8548
rect 34624 8520 34796 8548
rect 34112 8508 34118 8520
rect 32493 8483 32551 8489
rect 32493 8449 32505 8483
rect 32539 8449 32551 8483
rect 32493 8443 32551 8449
rect 34514 8440 34520 8492
rect 34572 8440 34578 8492
rect 34624 8489 34652 8520
rect 34790 8508 34796 8520
rect 34848 8508 34854 8560
rect 34882 8508 34888 8560
rect 34940 8508 34946 8560
rect 35084 8548 35112 8588
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36357 8619 36415 8625
rect 36357 8616 36369 8619
rect 35860 8588 36369 8616
rect 35860 8576 35866 8588
rect 36357 8585 36369 8588
rect 36403 8585 36415 8619
rect 38746 8616 38752 8628
rect 36357 8579 36415 8585
rect 37292 8588 38752 8616
rect 35342 8548 35348 8560
rect 35084 8520 35348 8548
rect 35342 8508 35348 8520
rect 35400 8508 35406 8560
rect 36170 8508 36176 8560
rect 36228 8548 36234 8560
rect 37292 8548 37320 8588
rect 38746 8576 38752 8588
rect 38804 8576 38810 8628
rect 40865 8619 40923 8625
rect 40865 8585 40877 8619
rect 40911 8616 40923 8619
rect 40954 8616 40960 8628
rect 40911 8588 40960 8616
rect 40911 8585 40923 8588
rect 40865 8579 40923 8585
rect 40954 8576 40960 8588
rect 41012 8576 41018 8628
rect 41233 8619 41291 8625
rect 41233 8585 41245 8619
rect 41279 8616 41291 8619
rect 41279 8588 42104 8616
rect 41279 8585 41291 8588
rect 41233 8579 41291 8585
rect 37366 8548 37372 8560
rect 36228 8520 37372 8548
rect 36228 8508 36234 8520
rect 37366 8508 37372 8520
rect 37424 8508 37430 8560
rect 40034 8548 40040 8560
rect 39974 8520 40040 8548
rect 40034 8508 40040 8520
rect 40092 8548 40098 8560
rect 40092 8520 40172 8548
rect 40092 8508 40098 8520
rect 34609 8483 34667 8489
rect 34609 8449 34621 8483
rect 34655 8449 34667 8483
rect 34609 8443 34667 8449
rect 36630 8440 36636 8492
rect 36688 8440 36694 8492
rect 38473 8483 38531 8489
rect 38473 8480 38485 8483
rect 38212 8452 38485 8480
rect 30024 8412 30052 8440
rect 28592 8384 30052 8412
rect 28592 8372 28598 8384
rect 30282 8372 30288 8424
rect 30340 8372 30346 8424
rect 30469 8415 30527 8421
rect 30469 8381 30481 8415
rect 30515 8412 30527 8415
rect 30834 8412 30840 8424
rect 30515 8384 30840 8412
rect 30515 8381 30527 8384
rect 30469 8375 30527 8381
rect 30834 8372 30840 8384
rect 30892 8372 30898 8424
rect 31757 8415 31815 8421
rect 31757 8412 31769 8415
rect 31680 8384 31769 8412
rect 31680 8356 31708 8384
rect 31757 8381 31769 8384
rect 31803 8381 31815 8415
rect 31757 8375 31815 8381
rect 32125 8415 32183 8421
rect 32125 8381 32137 8415
rect 32171 8381 32183 8415
rect 32125 8375 32183 8381
rect 31113 8347 31171 8353
rect 31113 8344 31125 8347
rect 26160 8316 27016 8344
rect 27172 8316 27844 8344
rect 29012 8316 31125 8344
rect 21683 8248 22048 8276
rect 23017 8279 23075 8285
rect 21683 8245 21695 8248
rect 21637 8239 21695 8245
rect 23017 8245 23029 8279
rect 23063 8245 23075 8279
rect 23017 8239 23075 8245
rect 23937 8279 23995 8285
rect 23937 8245 23949 8279
rect 23983 8276 23995 8279
rect 24026 8276 24032 8288
rect 23983 8248 24032 8276
rect 23983 8245 23995 8248
rect 23937 8239 23995 8245
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 24118 8236 24124 8288
rect 24176 8276 24182 8288
rect 25038 8276 25044 8288
rect 24176 8248 25044 8276
rect 24176 8236 24182 8248
rect 25038 8236 25044 8248
rect 25096 8236 25102 8288
rect 26878 8236 26884 8288
rect 26936 8236 26942 8288
rect 26988 8276 27016 8316
rect 27246 8276 27252 8288
rect 26988 8248 27252 8276
rect 27246 8236 27252 8248
rect 27304 8236 27310 8288
rect 28442 8236 28448 8288
rect 28500 8276 28506 8288
rect 29012 8276 29040 8316
rect 31113 8313 31125 8316
rect 31159 8313 31171 8347
rect 31113 8307 31171 8313
rect 31662 8304 31668 8356
rect 31720 8304 31726 8356
rect 32140 8344 32168 8375
rect 32214 8372 32220 8424
rect 32272 8372 32278 8424
rect 32306 8372 32312 8424
rect 32364 8372 32370 8424
rect 32858 8412 32864 8424
rect 32600 8384 32864 8412
rect 32600 8344 32628 8384
rect 32858 8372 32864 8384
rect 32916 8372 32922 8424
rect 36078 8372 36084 8424
rect 36136 8372 36142 8424
rect 36648 8412 36676 8440
rect 38212 8424 38240 8452
rect 38473 8449 38485 8452
rect 38519 8449 38531 8483
rect 40144 8480 40172 8520
rect 40218 8508 40224 8560
rect 40276 8548 40282 8560
rect 42076 8557 42104 8588
rect 42061 8551 42119 8557
rect 40276 8520 40724 8548
rect 40276 8508 40282 8520
rect 40586 8480 40592 8492
rect 40144 8452 40592 8480
rect 38473 8443 38531 8449
rect 40586 8440 40592 8452
rect 40644 8440 40650 8492
rect 40696 8424 40724 8520
rect 42061 8517 42073 8551
rect 42107 8517 42119 8551
rect 42061 8511 42119 8517
rect 42518 8508 42524 8560
rect 42576 8508 42582 8560
rect 40770 8440 40776 8492
rect 40828 8440 40834 8492
rect 41414 8440 41420 8492
rect 41472 8440 41478 8492
rect 41785 8483 41843 8489
rect 41785 8449 41797 8483
rect 41831 8449 41843 8483
rect 41785 8443 41843 8449
rect 38194 8412 38200 8424
rect 36648 8384 38200 8412
rect 38194 8372 38200 8384
rect 38252 8372 38258 8424
rect 40126 8412 40132 8424
rect 38304 8384 40132 8412
rect 32140 8316 32628 8344
rect 28500 8248 29040 8276
rect 28500 8236 28506 8248
rect 29362 8236 29368 8288
rect 29420 8276 29426 8288
rect 30929 8279 30987 8285
rect 30929 8276 30941 8279
rect 29420 8248 30941 8276
rect 29420 8236 29426 8248
rect 30929 8245 30941 8248
rect 30975 8245 30987 8279
rect 30929 8239 30987 8245
rect 31202 8236 31208 8288
rect 31260 8276 31266 8288
rect 31754 8276 31760 8288
rect 31260 8248 31760 8276
rect 31260 8236 31266 8248
rect 31754 8236 31760 8248
rect 31812 8236 31818 8288
rect 31846 8236 31852 8288
rect 31904 8236 31910 8288
rect 31938 8236 31944 8288
rect 31996 8276 32002 8288
rect 36096 8276 36124 8372
rect 31996 8248 36124 8276
rect 36896 8279 36954 8285
rect 31996 8236 32002 8248
rect 36896 8245 36908 8279
rect 36942 8276 36954 8279
rect 37090 8276 37096 8288
rect 36942 8248 37096 8276
rect 36942 8245 36954 8248
rect 36896 8239 36954 8245
rect 37090 8236 37096 8248
rect 37148 8236 37154 8288
rect 37550 8236 37556 8288
rect 37608 8276 37614 8288
rect 37918 8276 37924 8288
rect 37608 8248 37924 8276
rect 37608 8236 37614 8248
rect 37918 8236 37924 8248
rect 37976 8276 37982 8288
rect 38304 8276 38332 8384
rect 40126 8372 40132 8384
rect 40184 8412 40190 8424
rect 40221 8415 40279 8421
rect 40221 8412 40233 8415
rect 40184 8384 40233 8412
rect 40184 8372 40190 8384
rect 40221 8381 40233 8384
rect 40267 8381 40279 8415
rect 40221 8375 40279 8381
rect 40678 8372 40684 8424
rect 40736 8412 40742 8424
rect 40957 8415 41015 8421
rect 40957 8412 40969 8415
rect 40736 8384 40969 8412
rect 40736 8372 40742 8384
rect 40957 8381 40969 8384
rect 41003 8381 41015 8415
rect 41800 8412 41828 8443
rect 43438 8412 43444 8424
rect 41800 8384 43444 8412
rect 40957 8375 41015 8381
rect 43438 8372 43444 8384
rect 43496 8412 43502 8424
rect 43809 8415 43867 8421
rect 43809 8412 43821 8415
rect 43496 8384 43821 8412
rect 43496 8372 43502 8384
rect 43809 8381 43821 8384
rect 43855 8412 43867 8415
rect 44177 8415 44235 8421
rect 44177 8412 44189 8415
rect 43855 8384 44189 8412
rect 43855 8381 43867 8384
rect 43809 8375 43867 8381
rect 44177 8381 44189 8384
rect 44223 8412 44235 8415
rect 44910 8412 44916 8424
rect 44223 8384 44916 8412
rect 44223 8381 44235 8384
rect 44177 8375 44235 8381
rect 44910 8372 44916 8384
rect 44968 8372 44974 8424
rect 39758 8304 39764 8356
rect 39816 8344 39822 8356
rect 40405 8347 40463 8353
rect 40405 8344 40417 8347
rect 39816 8316 40417 8344
rect 39816 8304 39822 8316
rect 40405 8313 40417 8316
rect 40451 8313 40463 8347
rect 40405 8307 40463 8313
rect 37976 8248 38332 8276
rect 37976 8236 37982 8248
rect 38378 8236 38384 8288
rect 38436 8236 38442 8288
rect 38736 8279 38794 8285
rect 38736 8245 38748 8279
rect 38782 8276 38794 8279
rect 38838 8276 38844 8288
rect 38782 8248 38844 8276
rect 38782 8245 38794 8248
rect 38736 8239 38794 8245
rect 38838 8236 38844 8248
rect 38896 8236 38902 8288
rect 42794 8236 42800 8288
rect 42852 8276 42858 8288
rect 43533 8279 43591 8285
rect 43533 8276 43545 8279
rect 42852 8248 43545 8276
rect 42852 8236 42858 8248
rect 43533 8245 43545 8248
rect 43579 8245 43591 8279
rect 43533 8239 43591 8245
rect 44542 8236 44548 8288
rect 44600 8276 44606 8288
rect 44637 8279 44695 8285
rect 44637 8276 44649 8279
rect 44600 8248 44649 8276
rect 44600 8236 44606 8248
rect 44637 8245 44649 8248
rect 44683 8245 44695 8279
rect 44637 8239 44695 8245
rect 460 8186 45540 8208
rect 460 8134 3570 8186
rect 3622 8134 3634 8186
rect 3686 8134 3698 8186
rect 3750 8134 3762 8186
rect 3814 8134 3826 8186
rect 3878 8134 8570 8186
rect 8622 8134 8634 8186
rect 8686 8134 8698 8186
rect 8750 8134 8762 8186
rect 8814 8134 8826 8186
rect 8878 8134 13570 8186
rect 13622 8134 13634 8186
rect 13686 8134 13698 8186
rect 13750 8134 13762 8186
rect 13814 8134 13826 8186
rect 13878 8134 18570 8186
rect 18622 8134 18634 8186
rect 18686 8134 18698 8186
rect 18750 8134 18762 8186
rect 18814 8134 18826 8186
rect 18878 8134 23570 8186
rect 23622 8134 23634 8186
rect 23686 8134 23698 8186
rect 23750 8134 23762 8186
rect 23814 8134 23826 8186
rect 23878 8134 28570 8186
rect 28622 8134 28634 8186
rect 28686 8134 28698 8186
rect 28750 8134 28762 8186
rect 28814 8134 28826 8186
rect 28878 8134 33570 8186
rect 33622 8134 33634 8186
rect 33686 8134 33698 8186
rect 33750 8134 33762 8186
rect 33814 8134 33826 8186
rect 33878 8134 38570 8186
rect 38622 8134 38634 8186
rect 38686 8134 38698 8186
rect 38750 8134 38762 8186
rect 38814 8134 38826 8186
rect 38878 8134 43570 8186
rect 43622 8134 43634 8186
rect 43686 8134 43698 8186
rect 43750 8134 43762 8186
rect 43814 8134 43826 8186
rect 43878 8134 45540 8186
rect 460 8112 45540 8134
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8478 8072 8484 8084
rect 8159 8044 8484 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 8938 8072 8944 8084
rect 8803 8044 8944 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9953 8075 10011 8081
rect 9048 8044 9904 8072
rect 9048 8004 9076 8044
rect 8496 7976 9168 8004
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8496 7877 8524 7976
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8619 7908 9076 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 9048 7877 9076 7908
rect 9140 7877 9168 7976
rect 9306 7964 9312 8016
rect 9364 8004 9370 8016
rect 9876 8004 9904 8044
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10134 8072 10140 8084
rect 9999 8044 10140 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 11882 8072 11888 8084
rect 10560 8044 11888 8072
rect 10560 8032 10566 8044
rect 10042 8004 10048 8016
rect 9364 7976 9628 8004
rect 9876 7976 10048 8004
rect 9364 7964 9370 7976
rect 9600 7948 9628 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 10321 7939 10379 7945
rect 9640 7908 10088 7936
rect 9640 7896 9646 7908
rect 10060 7877 10088 7908
rect 10321 7905 10333 7939
rect 10367 7936 10379 7939
rect 10870 7936 10876 7948
rect 10367 7908 10876 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 9033 7871 9091 7877
rect 8711 7840 8984 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8404 7800 8432 7828
rect 8757 7803 8815 7809
rect 8757 7800 8769 7803
rect 8404 7772 8769 7800
rect 8757 7769 8769 7772
rect 8803 7769 8815 7803
rect 8956 7800 8984 7840
rect 9033 7837 9045 7871
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 10045 7871 10103 7877
rect 9355 7840 9720 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9324 7800 9352 7831
rect 9585 7803 9643 7809
rect 9585 7800 9597 7803
rect 8956 7772 9352 7800
rect 9508 7772 9597 7800
rect 8757 7763 8815 7769
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 9508 7741 9536 7772
rect 9585 7769 9597 7772
rect 9631 7769 9643 7803
rect 9585 7763 9643 7769
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8987 7704 9505 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9692 7732 9720 7840
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 11440 7854 11468 8044
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 12894 8072 12900 8084
rect 12851 8044 12900 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13354 8072 13360 8084
rect 13219 8044 13360 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 14918 8072 14924 8084
rect 13464 8044 14924 8072
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 13464 8004 13492 8044
rect 14918 8032 14924 8044
rect 14976 8072 14982 8084
rect 15197 8075 15255 8081
rect 15197 8072 15209 8075
rect 14976 8044 15209 8072
rect 14976 8032 14982 8044
rect 15197 8041 15209 8044
rect 15243 8041 15255 8075
rect 15197 8035 15255 8041
rect 18230 8032 18236 8084
rect 18288 8032 18294 8084
rect 20622 8032 20628 8084
rect 20680 8072 20686 8084
rect 22186 8072 22192 8084
rect 20680 8044 22192 8072
rect 20680 8032 20686 8044
rect 22186 8032 22192 8044
rect 22244 8072 22250 8084
rect 23290 8072 23296 8084
rect 22244 8044 23296 8072
rect 22244 8032 22250 8044
rect 22480 8013 22508 8044
rect 23290 8032 23296 8044
rect 23348 8032 23354 8084
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 24854 8072 24860 8084
rect 23891 8044 24860 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 25498 8032 25504 8084
rect 25556 8032 25562 8084
rect 27614 8032 27620 8084
rect 27672 8072 27678 8084
rect 27985 8075 28043 8081
rect 27985 8072 27997 8075
rect 27672 8044 27997 8072
rect 27672 8032 27678 8044
rect 27985 8041 27997 8044
rect 28031 8041 28043 8075
rect 27985 8035 28043 8041
rect 12768 7976 13492 8004
rect 22465 8007 22523 8013
rect 12768 7964 12774 7976
rect 10045 7831 10103 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12618 7868 12624 7880
rect 12492 7840 12624 7868
rect 12492 7828 12498 7840
rect 12618 7828 12624 7840
rect 12676 7868 12682 7880
rect 13004 7877 13032 7976
rect 22465 7973 22477 8007
rect 22511 7973 22523 8007
rect 22465 7967 22523 7973
rect 22554 7964 22560 8016
rect 22612 7964 22618 8016
rect 22833 8007 22891 8013
rect 22833 7973 22845 8007
rect 22879 8004 22891 8007
rect 22879 7976 23796 8004
rect 22879 7973 22891 7976
rect 22833 7967 22891 7973
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13170 7936 13176 7948
rect 13127 7908 13176 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12676 7840 12725 7868
rect 12676 7828 12682 7840
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12943 7840 13001 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 9769 7803 9827 7809
rect 9769 7769 9781 7803
rect 9815 7800 9827 7803
rect 10594 7800 10600 7812
rect 9815 7772 10600 7800
rect 9815 7769 9827 7772
rect 9769 7763 9827 7769
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 12728 7800 12756 7831
rect 13096 7800 13124 7899
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 14274 7936 14280 7948
rect 13311 7908 14280 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 15396 7908 16129 7936
rect 15396 7880 15424 7908
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 16393 7939 16451 7945
rect 16393 7905 16405 7939
rect 16439 7936 16451 7939
rect 16758 7936 16764 7948
rect 16439 7908 16764 7936
rect 16439 7905 16451 7908
rect 16393 7899 16451 7905
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 18598 7936 18604 7948
rect 17420 7908 18604 7936
rect 17420 7880 17448 7908
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20680 7908 21005 7936
rect 20680 7896 20686 7908
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 21508 7908 22416 7936
rect 21508 7896 21514 7908
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 13188 7840 13461 7868
rect 13188 7812 13216 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 15378 7828 15384 7880
rect 15436 7828 15442 7880
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 17402 7828 17408 7880
rect 17460 7828 17466 7880
rect 17494 7828 17500 7880
rect 17552 7828 17558 7880
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 20717 7871 20775 7877
rect 20717 7868 20729 7871
rect 20588 7840 20729 7868
rect 20588 7828 20594 7840
rect 20717 7837 20729 7840
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 12728 7772 13124 7800
rect 13170 7760 13176 7812
rect 13228 7760 13234 7812
rect 13725 7803 13783 7809
rect 13725 7769 13737 7803
rect 13771 7769 13783 7803
rect 13725 7763 13783 7769
rect 10410 7732 10416 7744
rect 9692 7704 10416 7732
rect 9493 7695 9551 7701
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 11790 7692 11796 7744
rect 11848 7692 11854 7744
rect 12253 7735 12311 7741
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 12526 7732 12532 7744
rect 12299 7704 12532 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13740 7732 13768 7763
rect 14458 7760 14464 7812
rect 14516 7760 14522 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 15252 7772 15761 7800
rect 15252 7760 15258 7772
rect 15749 7769 15761 7772
rect 15795 7800 15807 7803
rect 16482 7800 16488 7812
rect 15795 7772 16488 7800
rect 15795 7769 15807 7772
rect 15749 7763 15807 7769
rect 16482 7760 16488 7772
rect 16540 7760 16546 7812
rect 13044 7704 13768 7732
rect 13044 7692 13050 7704
rect 15654 7692 15660 7744
rect 15712 7692 15718 7744
rect 15838 7732 15844 7744
rect 15896 7741 15902 7744
rect 15805 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7695 15905 7741
rect 15933 7735 15991 7741
rect 15933 7701 15945 7735
rect 15979 7732 15991 7735
rect 16758 7732 16764 7744
rect 15979 7704 16764 7732
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 15896 7692 15902 7695
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 17512 7732 17540 7828
rect 18874 7760 18880 7812
rect 18932 7760 18938 7812
rect 19886 7760 19892 7812
rect 19944 7760 19950 7812
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 20625 7803 20683 7809
rect 20625 7800 20637 7803
rect 20496 7772 20637 7800
rect 20496 7760 20502 7772
rect 20625 7769 20637 7772
rect 20671 7800 20683 7803
rect 20898 7800 20904 7812
rect 20671 7772 20904 7800
rect 20671 7769 20683 7772
rect 20625 7763 20683 7769
rect 20898 7760 20904 7772
rect 20956 7760 20962 7812
rect 22278 7800 22284 7812
rect 22218 7772 22284 7800
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 22388 7800 22416 7908
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7868 22799 7871
rect 22830 7868 22836 7880
rect 22787 7840 22836 7868
rect 22787 7837 22799 7840
rect 22741 7831 22799 7837
rect 22830 7828 22836 7840
rect 22888 7828 22894 7880
rect 23768 7877 23796 7976
rect 24118 7896 24124 7948
rect 24176 7896 24182 7948
rect 24397 7939 24455 7945
rect 24397 7905 24409 7939
rect 24443 7936 24455 7939
rect 24486 7936 24492 7948
rect 24443 7908 24492 7936
rect 24443 7905 24455 7908
rect 24397 7899 24455 7905
rect 24486 7896 24492 7908
rect 24544 7896 24550 7948
rect 25516 7936 25544 8032
rect 28000 8004 28028 8035
rect 28442 8032 28448 8084
rect 28500 8032 28506 8084
rect 31202 8072 31208 8084
rect 29380 8044 31208 8072
rect 28000 7976 28212 8004
rect 26145 7939 26203 7945
rect 26145 7936 26157 7939
rect 25516 7908 26157 7936
rect 26145 7905 26157 7908
rect 26191 7905 26203 7939
rect 26145 7899 26203 7905
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 26559 7908 28089 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28184 7936 28212 7976
rect 28353 7939 28411 7945
rect 28353 7936 28365 7939
rect 28184 7908 28365 7936
rect 28077 7899 28135 7905
rect 28353 7905 28365 7908
rect 28399 7905 28411 7939
rect 28460 7936 28488 8032
rect 29178 8004 29184 8016
rect 28644 7976 29184 8004
rect 28537 7939 28595 7945
rect 28537 7936 28549 7939
rect 28460 7908 28549 7936
rect 28353 7899 28411 7905
rect 28537 7905 28549 7908
rect 28583 7905 28595 7939
rect 28537 7899 28595 7905
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7837 23811 7871
rect 25682 7868 25688 7880
rect 25530 7854 25688 7868
rect 23753 7831 23811 7837
rect 25516 7840 25688 7854
rect 22646 7800 22652 7812
rect 22388 7772 22652 7800
rect 22646 7760 22652 7772
rect 22704 7800 22710 7812
rect 23201 7803 23259 7809
rect 23201 7800 23213 7803
rect 22704 7772 23213 7800
rect 22704 7760 22710 7772
rect 23201 7769 23213 7772
rect 23247 7769 23259 7803
rect 23201 7763 23259 7769
rect 17460 7704 17540 7732
rect 17865 7735 17923 7741
rect 17460 7692 17466 7704
rect 17865 7701 17877 7735
rect 17911 7732 17923 7735
rect 18046 7732 18052 7744
rect 17911 7704 18052 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 23014 7732 23020 7744
rect 21876 7704 23020 7732
rect 21876 7692 21882 7704
rect 23014 7692 23020 7704
rect 23072 7732 23078 7744
rect 23293 7735 23351 7741
rect 23293 7732 23305 7735
rect 23072 7704 23305 7732
rect 23072 7692 23078 7704
rect 23293 7701 23305 7704
rect 23339 7732 23351 7735
rect 23474 7732 23480 7744
rect 23339 7704 23480 7732
rect 23339 7701 23351 7704
rect 23293 7695 23351 7701
rect 23474 7692 23480 7704
rect 23532 7692 23538 7744
rect 24210 7692 24216 7744
rect 24268 7732 24274 7744
rect 25516 7732 25544 7840
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 24268 7704 25544 7732
rect 26160 7732 26188 7899
rect 26237 7871 26295 7877
rect 26237 7837 26249 7871
rect 26283 7837 26295 7871
rect 27982 7868 27988 7880
rect 27646 7840 27988 7868
rect 26237 7831 26295 7837
rect 26252 7800 26280 7831
rect 27982 7828 27988 7840
rect 28040 7828 28046 7880
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7837 28319 7871
rect 28261 7831 28319 7837
rect 28276 7800 28304 7831
rect 28442 7828 28448 7880
rect 28500 7868 28506 7880
rect 28644 7868 28672 7976
rect 29178 7964 29184 7976
rect 29236 7964 29242 8016
rect 28810 7896 28816 7948
rect 28868 7936 28874 7948
rect 28868 7908 28994 7936
rect 28868 7896 28874 7908
rect 28500 7840 28672 7868
rect 28966 7868 28994 7908
rect 29086 7896 29092 7948
rect 29144 7896 29150 7948
rect 29380 7945 29408 8044
rect 31202 8032 31208 8044
rect 31260 8032 31266 8084
rect 31481 8075 31539 8081
rect 31481 8041 31493 8075
rect 31527 8072 31539 8075
rect 31662 8072 31668 8084
rect 31527 8044 31668 8072
rect 31527 8041 31539 8044
rect 31481 8035 31539 8041
rect 31662 8032 31668 8044
rect 31720 8032 31726 8084
rect 31846 8032 31852 8084
rect 31904 8032 31910 8084
rect 32858 8032 32864 8084
rect 32916 8072 32922 8084
rect 33873 8075 33931 8081
rect 33873 8072 33885 8075
rect 32916 8044 33885 8072
rect 32916 8032 32922 8044
rect 33873 8041 33885 8044
rect 33919 8072 33931 8075
rect 34238 8072 34244 8084
rect 33919 8044 34244 8072
rect 33919 8041 33931 8044
rect 33873 8035 33931 8041
rect 34238 8032 34244 8044
rect 34296 8032 34302 8084
rect 36722 8032 36728 8084
rect 36780 8032 36786 8084
rect 36906 8032 36912 8084
rect 36964 8072 36970 8084
rect 37001 8075 37059 8081
rect 37001 8072 37013 8075
rect 36964 8044 37013 8072
rect 36964 8032 36970 8044
rect 37001 8041 37013 8044
rect 37047 8041 37059 8075
rect 37001 8035 37059 8041
rect 37458 8032 37464 8084
rect 37516 8072 37522 8084
rect 38013 8075 38071 8081
rect 38013 8072 38025 8075
rect 37516 8044 38025 8072
rect 37516 8032 37522 8044
rect 38013 8041 38025 8044
rect 38059 8072 38071 8075
rect 38381 8075 38439 8081
rect 38381 8072 38393 8075
rect 38059 8044 38393 8072
rect 38059 8041 38071 8044
rect 38013 8035 38071 8041
rect 38381 8041 38393 8044
rect 38427 8041 38439 8075
rect 38381 8035 38439 8041
rect 38470 8032 38476 8084
rect 38528 8032 38534 8084
rect 41414 8032 41420 8084
rect 41472 8072 41478 8084
rect 41509 8075 41567 8081
rect 41509 8072 41521 8075
rect 41472 8044 41521 8072
rect 41472 8032 41478 8044
rect 41509 8041 41521 8044
rect 41555 8041 41567 8075
rect 41509 8035 41567 8041
rect 43254 8032 43260 8084
rect 43312 8072 43318 8084
rect 43349 8075 43407 8081
rect 43349 8072 43361 8075
rect 43312 8044 43361 8072
rect 43312 8032 43318 8044
rect 43349 8041 43361 8044
rect 43395 8041 43407 8075
rect 43349 8035 43407 8041
rect 30374 8004 30380 8016
rect 30208 7976 30380 8004
rect 29365 7939 29423 7945
rect 29365 7905 29377 7939
rect 29411 7905 29423 7939
rect 29365 7899 29423 7905
rect 29638 7896 29644 7948
rect 29696 7936 29702 7948
rect 30009 7939 30067 7945
rect 30009 7936 30021 7939
rect 29696 7908 30021 7936
rect 29696 7896 29702 7908
rect 30009 7905 30021 7908
rect 30055 7905 30067 7939
rect 30208 7936 30236 7976
rect 30374 7964 30380 7976
rect 30432 8004 30438 8016
rect 30834 8004 30840 8016
rect 30432 7976 30840 8004
rect 30432 7964 30438 7976
rect 30834 7964 30840 7976
rect 30892 8004 30898 8016
rect 31754 8004 31760 8016
rect 30892 7976 30972 8004
rect 30892 7964 30898 7976
rect 30009 7899 30067 7905
rect 30116 7908 30236 7936
rect 29181 7871 29239 7877
rect 29181 7868 29193 7871
rect 28966 7840 29193 7868
rect 28500 7828 28506 7840
rect 29181 7837 29193 7840
rect 29227 7837 29239 7871
rect 29181 7831 29239 7837
rect 29270 7828 29276 7880
rect 29328 7828 29334 7880
rect 29730 7828 29736 7880
rect 29788 7828 29794 7880
rect 29822 7828 29828 7880
rect 29880 7828 29886 7880
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7868 29975 7871
rect 30116 7868 30144 7908
rect 30282 7896 30288 7948
rect 30340 7936 30346 7948
rect 30944 7945 30972 7976
rect 31036 7976 31760 8004
rect 31036 7945 31064 7976
rect 31754 7964 31760 7976
rect 31812 7964 31818 8016
rect 31864 8004 31892 8032
rect 31864 7976 32260 8004
rect 30929 7939 30987 7945
rect 30340 7908 30788 7936
rect 30340 7896 30346 7908
rect 30760 7880 30788 7908
rect 30929 7905 30941 7939
rect 30975 7905 30987 7939
rect 30929 7899 30987 7905
rect 31021 7939 31079 7945
rect 31021 7905 31033 7939
rect 31067 7905 31079 7939
rect 31021 7899 31079 7905
rect 31294 7896 31300 7948
rect 31352 7896 31358 7948
rect 31386 7896 31392 7948
rect 31444 7936 31450 7948
rect 32030 7936 32036 7948
rect 31444 7908 32036 7936
rect 31444 7896 31450 7908
rect 32030 7896 32036 7908
rect 32088 7936 32094 7948
rect 32125 7939 32183 7945
rect 32125 7936 32137 7939
rect 32088 7908 32137 7936
rect 32088 7896 32094 7908
rect 32125 7905 32137 7908
rect 32171 7905 32183 7939
rect 32232 7936 32260 7976
rect 34054 7964 34060 8016
rect 34112 7964 34118 8016
rect 32401 7939 32459 7945
rect 32401 7936 32413 7939
rect 32232 7908 32413 7936
rect 32125 7899 32183 7905
rect 32401 7905 32413 7908
rect 32447 7905 32459 7939
rect 32401 7899 32459 7905
rect 32950 7896 32956 7948
rect 33008 7936 33014 7948
rect 34072 7936 34100 7964
rect 33008 7908 34100 7936
rect 35437 7939 35495 7945
rect 33008 7896 33014 7908
rect 29963 7840 30144 7868
rect 29963 7837 29975 7840
rect 29917 7831 29975 7837
rect 30742 7828 30748 7880
rect 30800 7828 30806 7880
rect 30834 7828 30840 7880
rect 30892 7828 30898 7880
rect 31312 7868 31340 7896
rect 31665 7871 31723 7877
rect 31665 7868 31677 7871
rect 31312 7840 31677 7868
rect 31665 7837 31677 7840
rect 31711 7837 31723 7871
rect 31665 7831 31723 7837
rect 31754 7828 31760 7880
rect 31812 7828 31818 7880
rect 31849 7871 31907 7877
rect 31849 7837 31861 7871
rect 31895 7837 31907 7871
rect 31849 7831 31907 7837
rect 31942 7871 32000 7877
rect 31942 7837 31954 7871
rect 31988 7868 32000 7871
rect 31988 7840 32168 7868
rect 33520 7854 33548 7908
rect 35437 7905 35449 7939
rect 35483 7936 35495 7939
rect 36740 7936 36768 8032
rect 38488 8004 38516 8032
rect 42337 8007 42395 8013
rect 42337 8004 42349 8007
rect 37660 7976 38516 8004
rect 40972 7976 42349 8004
rect 37660 7948 37688 7976
rect 35483 7908 36768 7936
rect 35483 7905 35495 7908
rect 35437 7899 35495 7905
rect 36998 7896 37004 7948
rect 37056 7936 37062 7948
rect 37550 7936 37556 7948
rect 37056 7908 37556 7936
rect 37056 7896 37062 7908
rect 37550 7896 37556 7908
rect 37608 7896 37614 7948
rect 37642 7896 37648 7948
rect 37700 7896 37706 7948
rect 40972 7936 41000 7976
rect 42337 7973 42349 7976
rect 42383 7973 42395 8007
rect 42337 7967 42395 7973
rect 42720 7976 42932 8004
rect 42720 7948 42748 7976
rect 41417 7939 41475 7945
rect 41417 7936 41429 7939
rect 38488 7908 41000 7936
rect 41248 7908 41429 7936
rect 31988 7837 32000 7840
rect 31942 7831 32000 7837
rect 29086 7800 29092 7812
rect 26252 7772 26648 7800
rect 28276 7772 29092 7800
rect 26620 7744 26648 7772
rect 29086 7760 29092 7772
rect 29144 7760 29150 7812
rect 30285 7803 30343 7809
rect 30285 7769 30297 7803
rect 30331 7800 30343 7803
rect 31478 7800 31484 7812
rect 30331 7772 31484 7800
rect 30331 7769 30343 7772
rect 30285 7763 30343 7769
rect 31478 7760 31484 7772
rect 31536 7760 31542 7812
rect 31864 7800 31892 7831
rect 32030 7800 32036 7812
rect 31864 7772 32036 7800
rect 32030 7760 32036 7772
rect 32088 7760 32094 7812
rect 26418 7732 26424 7744
rect 26160 7704 26424 7732
rect 24268 7692 24274 7704
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 26602 7692 26608 7744
rect 26660 7692 26666 7744
rect 28166 7692 28172 7744
rect 28224 7732 28230 7744
rect 28905 7735 28963 7741
rect 28905 7732 28917 7735
rect 28224 7704 28917 7732
rect 28224 7692 28230 7704
rect 28905 7701 28917 7704
rect 28951 7701 28963 7735
rect 28905 7695 28963 7701
rect 29546 7692 29552 7744
rect 29604 7692 29610 7744
rect 30374 7692 30380 7744
rect 30432 7692 30438 7744
rect 30558 7692 30564 7744
rect 30616 7692 30622 7744
rect 32140 7732 32168 7840
rect 34054 7828 34060 7880
rect 34112 7828 34118 7880
rect 34333 7871 34391 7877
rect 34333 7837 34345 7871
rect 34379 7868 34391 7871
rect 34422 7868 34428 7880
rect 34379 7840 34428 7868
rect 34379 7837 34391 7840
rect 34333 7831 34391 7837
rect 34348 7800 34376 7831
rect 34422 7828 34428 7840
rect 34480 7828 34486 7880
rect 35066 7828 35072 7880
rect 35124 7868 35130 7880
rect 35161 7871 35219 7877
rect 35161 7868 35173 7871
rect 35124 7840 35173 7868
rect 35124 7828 35130 7840
rect 35161 7837 35173 7840
rect 35207 7837 35219 7871
rect 35161 7831 35219 7837
rect 37369 7871 37427 7877
rect 37369 7837 37381 7871
rect 37415 7868 37427 7871
rect 37458 7868 37464 7880
rect 37415 7840 37464 7868
rect 37415 7837 37427 7840
rect 37369 7831 37427 7837
rect 37458 7828 37464 7840
rect 37516 7868 37522 7880
rect 38378 7868 38384 7880
rect 37516 7840 38384 7868
rect 37516 7828 37522 7840
rect 38378 7828 38384 7840
rect 38436 7828 38442 7880
rect 34348 7772 35756 7800
rect 35728 7744 35756 7772
rect 35820 7772 35926 7800
rect 35820 7744 35848 7772
rect 37090 7760 37096 7812
rect 37148 7800 37154 7812
rect 38488 7800 38516 7908
rect 39574 7828 39580 7880
rect 39632 7828 39638 7880
rect 39666 7828 39672 7880
rect 39724 7828 39730 7880
rect 38841 7803 38899 7809
rect 38841 7800 38853 7803
rect 37148 7772 38516 7800
rect 38626 7772 38853 7800
rect 37148 7760 37154 7772
rect 34422 7732 34428 7744
rect 32140 7704 34428 7732
rect 34422 7692 34428 7704
rect 34480 7692 34486 7744
rect 35710 7692 35716 7744
rect 35768 7692 35774 7744
rect 35802 7692 35808 7744
rect 35860 7732 35866 7744
rect 36170 7732 36176 7744
rect 35860 7704 36176 7732
rect 35860 7692 35866 7704
rect 36170 7692 36176 7704
rect 36228 7692 36234 7744
rect 36722 7692 36728 7744
rect 36780 7732 36786 7744
rect 36909 7735 36967 7741
rect 36909 7732 36921 7735
rect 36780 7704 36921 7732
rect 36780 7692 36786 7704
rect 36909 7701 36921 7704
rect 36955 7732 36967 7735
rect 37461 7735 37519 7741
rect 37461 7732 37473 7735
rect 36955 7704 37473 7732
rect 36955 7701 36967 7704
rect 36909 7695 36967 7701
rect 37461 7701 37473 7704
rect 37507 7701 37519 7735
rect 37461 7695 37519 7701
rect 38194 7692 38200 7744
rect 38252 7732 38258 7744
rect 38626 7732 38654 7772
rect 38841 7769 38853 7772
rect 38887 7800 38899 7803
rect 39206 7800 39212 7812
rect 38887 7772 39212 7800
rect 38887 7769 38899 7772
rect 38841 7763 38899 7769
rect 39206 7760 39212 7772
rect 39264 7800 39270 7812
rect 39684 7800 39712 7828
rect 39264 7772 39712 7800
rect 39945 7803 40003 7809
rect 39264 7760 39270 7772
rect 39945 7769 39957 7803
rect 39991 7769 40003 7803
rect 39945 7763 40003 7769
rect 38252 7704 38654 7732
rect 39393 7735 39451 7741
rect 38252 7692 38258 7704
rect 39393 7701 39405 7735
rect 39439 7732 39451 7735
rect 39960 7732 39988 7763
rect 40586 7760 40592 7812
rect 40644 7760 40650 7812
rect 39439 7704 39988 7732
rect 39439 7701 39451 7704
rect 39393 7695 39451 7701
rect 40770 7692 40776 7744
rect 40828 7732 40834 7744
rect 41248 7732 41276 7908
rect 41417 7905 41429 7908
rect 41463 7905 41475 7939
rect 42058 7936 42064 7948
rect 41417 7899 41475 7905
rect 41800 7908 42064 7936
rect 41800 7868 41828 7908
rect 42058 7896 42064 7908
rect 42116 7896 42122 7948
rect 42702 7896 42708 7948
rect 42760 7896 42766 7948
rect 42794 7896 42800 7948
rect 42852 7896 42858 7948
rect 42904 7945 42932 7976
rect 42889 7939 42947 7945
rect 42889 7905 42901 7939
rect 42935 7905 42947 7939
rect 42889 7899 42947 7905
rect 41386 7840 41828 7868
rect 41386 7744 41414 7840
rect 41874 7828 41880 7880
rect 41932 7828 41938 7880
rect 41969 7871 42027 7877
rect 41969 7837 41981 7871
rect 42015 7868 42027 7871
rect 42812 7868 42840 7896
rect 42015 7840 42840 7868
rect 42015 7837 42027 7840
rect 41969 7831 42027 7837
rect 45002 7800 45008 7812
rect 40828 7704 41276 7732
rect 40828 7692 40834 7704
rect 41322 7692 41328 7744
rect 41380 7704 41414 7744
rect 42720 7772 45008 7800
rect 42720 7741 42748 7772
rect 45002 7760 45008 7772
rect 45060 7760 45066 7812
rect 42705 7735 42763 7741
rect 41380 7692 41386 7704
rect 42705 7701 42717 7735
rect 42751 7701 42763 7735
rect 42705 7695 42763 7701
rect 43438 7692 43444 7744
rect 43496 7732 43502 7744
rect 43717 7735 43775 7741
rect 43717 7732 43729 7735
rect 43496 7704 43729 7732
rect 43496 7692 43502 7704
rect 43717 7701 43729 7704
rect 43763 7701 43775 7735
rect 43717 7695 43775 7701
rect 44174 7692 44180 7744
rect 44232 7692 44238 7744
rect 44542 7692 44548 7744
rect 44600 7732 44606 7744
rect 44910 7732 44916 7744
rect 44600 7704 44916 7732
rect 44600 7692 44606 7704
rect 44910 7692 44916 7704
rect 44968 7692 44974 7744
rect 460 7642 45540 7664
rect 460 7590 6070 7642
rect 6122 7590 6134 7642
rect 6186 7590 6198 7642
rect 6250 7590 6262 7642
rect 6314 7590 6326 7642
rect 6378 7590 11070 7642
rect 11122 7590 11134 7642
rect 11186 7590 11198 7642
rect 11250 7590 11262 7642
rect 11314 7590 11326 7642
rect 11378 7590 16070 7642
rect 16122 7590 16134 7642
rect 16186 7590 16198 7642
rect 16250 7590 16262 7642
rect 16314 7590 16326 7642
rect 16378 7590 21070 7642
rect 21122 7590 21134 7642
rect 21186 7590 21198 7642
rect 21250 7590 21262 7642
rect 21314 7590 21326 7642
rect 21378 7590 26070 7642
rect 26122 7590 26134 7642
rect 26186 7590 26198 7642
rect 26250 7590 26262 7642
rect 26314 7590 26326 7642
rect 26378 7590 31070 7642
rect 31122 7590 31134 7642
rect 31186 7590 31198 7642
rect 31250 7590 31262 7642
rect 31314 7590 31326 7642
rect 31378 7590 36070 7642
rect 36122 7590 36134 7642
rect 36186 7590 36198 7642
rect 36250 7590 36262 7642
rect 36314 7590 36326 7642
rect 36378 7590 41070 7642
rect 41122 7590 41134 7642
rect 41186 7590 41198 7642
rect 41250 7590 41262 7642
rect 41314 7590 41326 7642
rect 41378 7590 45540 7642
rect 460 7568 45540 7590
rect 7650 7488 7656 7540
rect 7708 7488 7714 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9214 7528 9220 7540
rect 8536 7500 9220 7528
rect 8536 7488 8542 7500
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10100 7500 10548 7528
rect 10100 7488 10106 7500
rect 7668 7392 7696 7488
rect 7760 7460 7788 7488
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 7760 7432 8769 7460
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 10520 7460 10548 7500
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10652 7500 10701 7528
rect 10652 7488 10658 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11422 7528 11428 7540
rect 11379 7500 11428 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 11882 7528 11888 7540
rect 11839 7500 11888 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 11882 7488 11888 7500
rect 11940 7528 11946 7540
rect 12069 7531 12127 7537
rect 12069 7528 12081 7531
rect 11940 7500 12081 7528
rect 11940 7488 11946 7500
rect 12069 7497 12081 7500
rect 12115 7497 12127 7531
rect 12069 7491 12127 7497
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 13679 7500 14381 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 14369 7497 14381 7500
rect 14415 7528 14427 7531
rect 14458 7528 14464 7540
rect 14415 7500 14464 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 15672 7500 16620 7528
rect 15672 7469 15700 7500
rect 16592 7472 16620 7500
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 17586 7528 17592 7540
rect 16724 7500 17592 7528
rect 16724 7488 16730 7500
rect 17586 7488 17592 7500
rect 17644 7528 17650 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 17644 7500 17785 7528
rect 17644 7488 17650 7500
rect 17773 7497 17785 7500
rect 17819 7497 17831 7531
rect 17773 7491 17831 7497
rect 18417 7531 18475 7537
rect 18417 7497 18429 7531
rect 18463 7528 18475 7531
rect 18874 7528 18880 7540
rect 18463 7500 18880 7528
rect 18463 7497 18475 7500
rect 18417 7491 18475 7497
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 20162 7528 20168 7540
rect 19352 7500 20168 7528
rect 10873 7463 10931 7469
rect 10873 7460 10885 7463
rect 10520 7432 10885 7460
rect 8757 7423 8815 7429
rect 10873 7429 10885 7432
rect 10919 7429 10931 7463
rect 15657 7463 15715 7469
rect 15657 7460 15669 7463
rect 10873 7423 10931 7429
rect 15028 7432 15669 7460
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7668 7364 8033 7392
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 10502 7392 10508 7404
rect 10350 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11790 7392 11796 7404
rect 11195 7364 11796 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 15028 7401 15056 7432
rect 15657 7429 15669 7432
rect 15703 7429 15715 7463
rect 15657 7423 15715 7429
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 15896 7432 16313 7460
rect 15896 7420 15902 7432
rect 16301 7429 16313 7432
rect 16347 7429 16359 7463
rect 16301 7423 16359 7429
rect 16574 7420 16580 7472
rect 16632 7420 16638 7472
rect 17972 7432 18552 7460
rect 17972 7404 18000 7432
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15194 7392 15200 7404
rect 15151 7364 15200 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9950 7324 9956 7336
rect 9263 7296 9956 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10468 7296 10977 7324
rect 10468 7284 10474 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 13078 7216 13084 7268
rect 13136 7256 13142 7268
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 13136 7228 13277 7256
rect 13136 7216 13142 7228
rect 13265 7225 13277 7228
rect 13311 7256 13323 7259
rect 13909 7259 13967 7265
rect 13909 7256 13921 7259
rect 13311 7228 13921 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13909 7225 13921 7228
rect 13955 7225 13967 7259
rect 13909 7219 13967 7225
rect 14642 7216 14648 7268
rect 14700 7256 14706 7268
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14700 7228 14749 7256
rect 14700 7216 14706 7228
rect 14737 7225 14749 7228
rect 14783 7225 14795 7259
rect 14844 7256 14872 7355
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15473 7355 15531 7361
rect 15580 7364 16037 7392
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15396 7324 15424 7355
rect 14967 7296 15424 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15488 7256 15516 7355
rect 15580 7336 15608 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 17865 7395 17923 7401
rect 17865 7392 17877 7395
rect 17736 7364 17877 7392
rect 17736 7352 17742 7364
rect 17865 7361 17877 7364
rect 17911 7361 17923 7395
rect 17865 7355 17923 7361
rect 17954 7352 17960 7404
rect 18012 7352 18018 7404
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 18524 7401 18552 7432
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 19352 7469 19380 7500
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 20806 7488 20812 7540
rect 20864 7488 20870 7540
rect 21729 7531 21787 7537
rect 21729 7497 21741 7531
rect 21775 7528 21787 7531
rect 22462 7528 22468 7540
rect 21775 7500 22468 7528
rect 21775 7497 21787 7500
rect 21729 7491 21787 7497
rect 22462 7488 22468 7500
rect 22520 7488 22526 7540
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 24302 7488 24308 7540
rect 24360 7488 24366 7540
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 24946 7528 24952 7540
rect 24596 7500 24952 7528
rect 18969 7463 19027 7469
rect 18969 7460 18981 7463
rect 18656 7432 18981 7460
rect 18656 7420 18662 7432
rect 18969 7429 18981 7432
rect 19015 7429 19027 7463
rect 18969 7423 19027 7429
rect 19337 7463 19395 7469
rect 19337 7429 19349 7463
rect 19383 7429 19395 7463
rect 19337 7423 19395 7429
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7361 18383 7395
rect 18325 7355 18383 7361
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18984 7392 19012 7423
rect 20898 7420 20904 7472
rect 20956 7460 20962 7472
rect 21453 7463 21511 7469
rect 21453 7460 21465 7463
rect 20956 7432 21465 7460
rect 20956 7420 20962 7432
rect 21453 7429 21465 7432
rect 21499 7429 21511 7463
rect 21453 7423 21511 7429
rect 21637 7463 21695 7469
rect 21637 7429 21649 7463
rect 21683 7460 21695 7463
rect 21818 7460 21824 7472
rect 21683 7432 21824 7460
rect 21683 7429 21695 7432
rect 21637 7423 21695 7429
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 22002 7420 22008 7472
rect 22060 7460 22066 7472
rect 22572 7460 22600 7488
rect 22833 7463 22891 7469
rect 22833 7460 22845 7463
rect 22060 7432 22416 7460
rect 22572 7432 22845 7460
rect 22060 7420 22066 7432
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18984 7364 19073 7392
rect 18509 7355 18567 7361
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 15562 7284 15568 7336
rect 15620 7284 15626 7336
rect 15654 7284 15660 7336
rect 15712 7324 15718 7336
rect 17420 7324 17448 7352
rect 18064 7324 18092 7352
rect 15712 7296 17448 7324
rect 17696 7296 18092 7324
rect 15712 7284 15718 7296
rect 15930 7256 15936 7268
rect 14844 7228 15936 7256
rect 14737 7219 14795 7225
rect 15930 7216 15936 7228
rect 15988 7216 15994 7268
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 10873 7191 10931 7197
rect 10873 7188 10885 7191
rect 10652 7160 10885 7188
rect 10652 7148 10658 7160
rect 10873 7157 10885 7160
rect 10919 7157 10931 7191
rect 10873 7151 10931 7157
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12584 7160 12817 7188
rect 12584 7148 12590 7160
rect 12805 7157 12817 7160
rect 12851 7188 12863 7191
rect 13170 7188 13176 7200
rect 12851 7160 13176 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 15102 7148 15108 7200
rect 15160 7148 15166 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15838 7188 15844 7200
rect 15344 7160 15844 7188
rect 15344 7148 15350 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17696 7188 17724 7296
rect 18340 7200 18368 7355
rect 19076 7324 19104 7355
rect 19794 7324 19800 7336
rect 19076 7296 19800 7324
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 20456 7324 20484 7378
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22388 7392 22416 7432
rect 22833 7429 22845 7432
rect 22879 7429 22891 7463
rect 24210 7460 24216 7472
rect 24058 7432 24216 7460
rect 22833 7423 22891 7429
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 22462 7392 22468 7404
rect 22235 7364 22324 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 19944 7296 22140 7324
rect 19944 7284 19950 7296
rect 22112 7200 22140 7296
rect 22296 7256 22324 7364
rect 22388 7364 22468 7392
rect 22388 7333 22416 7364
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 24596 7401 24624 7500
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 25317 7531 25375 7537
rect 25317 7497 25329 7531
rect 25363 7528 25375 7531
rect 25406 7528 25412 7540
rect 25363 7500 25412 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 26510 7488 26516 7540
rect 26568 7488 26574 7540
rect 26878 7488 26884 7540
rect 26936 7488 26942 7540
rect 28166 7488 28172 7540
rect 28224 7488 28230 7540
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 28626 7528 28632 7540
rect 28408 7500 28632 7528
rect 28408 7488 28414 7500
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 29546 7528 29552 7540
rect 28736 7500 29552 7528
rect 25222 7460 25228 7472
rect 24946 7432 25228 7460
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7392 24731 7395
rect 24762 7392 24768 7404
rect 24719 7364 24768 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 24946 7401 24974 7432
rect 25222 7420 25228 7432
rect 25280 7420 25286 7472
rect 26896 7460 26924 7488
rect 26344 7432 26924 7460
rect 26344 7401 26372 7432
rect 24931 7395 24989 7401
rect 24931 7361 24943 7395
rect 24977 7361 24989 7395
rect 24931 7355 24989 7361
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 27982 7352 27988 7404
rect 28040 7352 28046 7404
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 23198 7324 23204 7336
rect 22664 7296 23204 7324
rect 22664 7256 22692 7296
rect 23198 7284 23204 7296
rect 23256 7284 23262 7336
rect 24026 7284 24032 7336
rect 24084 7284 24090 7336
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25222 7324 25228 7336
rect 25096 7296 25228 7324
rect 25096 7284 25102 7296
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25685 7327 25743 7333
rect 25685 7324 25697 7327
rect 25280 7296 25697 7324
rect 25280 7284 25286 7296
rect 25685 7293 25697 7296
rect 25731 7324 25743 7327
rect 26145 7327 26203 7333
rect 26145 7324 26157 7327
rect 25731 7296 26157 7324
rect 25731 7293 25743 7296
rect 25685 7287 25743 7293
rect 26145 7293 26157 7296
rect 26191 7324 26203 7327
rect 26602 7324 26608 7336
rect 26191 7296 26608 7324
rect 26191 7293 26203 7296
rect 26145 7287 26203 7293
rect 26602 7284 26608 7296
rect 26660 7284 26666 7336
rect 26881 7327 26939 7333
rect 26881 7293 26893 7327
rect 26927 7324 26939 7327
rect 28184 7324 28212 7488
rect 28736 7469 28764 7500
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 30374 7488 30380 7540
rect 30432 7488 30438 7540
rect 31662 7488 31668 7540
rect 31720 7528 31726 7540
rect 31720 7488 31754 7528
rect 31938 7488 31944 7540
rect 31996 7528 32002 7540
rect 32858 7528 32864 7540
rect 31996 7500 32864 7528
rect 31996 7488 32002 7500
rect 32858 7488 32864 7500
rect 32916 7528 32922 7540
rect 33321 7531 33379 7537
rect 33321 7528 33333 7531
rect 32916 7500 33333 7528
rect 32916 7488 32922 7500
rect 33321 7497 33333 7500
rect 33367 7497 33379 7531
rect 33321 7491 33379 7497
rect 33689 7531 33747 7537
rect 33689 7497 33701 7531
rect 33735 7528 33747 7531
rect 34054 7528 34060 7540
rect 33735 7500 34060 7528
rect 33735 7497 33747 7500
rect 33689 7491 33747 7497
rect 34054 7488 34060 7500
rect 34112 7488 34118 7540
rect 34146 7488 34152 7540
rect 34204 7488 34210 7540
rect 34238 7488 34244 7540
rect 34296 7488 34302 7540
rect 34514 7488 34520 7540
rect 34572 7528 34578 7540
rect 35529 7531 35587 7537
rect 35529 7528 35541 7531
rect 34572 7500 35541 7528
rect 34572 7488 34578 7500
rect 35529 7497 35541 7500
rect 35575 7497 35587 7531
rect 35529 7491 35587 7497
rect 35986 7488 35992 7540
rect 36044 7488 36050 7540
rect 36817 7531 36875 7537
rect 36817 7497 36829 7531
rect 36863 7528 36875 7531
rect 38286 7528 38292 7540
rect 36863 7500 38292 7528
rect 36863 7497 36875 7500
rect 36817 7491 36875 7497
rect 38286 7488 38292 7500
rect 38344 7488 38350 7540
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7497 38715 7531
rect 38657 7491 38715 7497
rect 28721 7463 28779 7469
rect 28721 7429 28733 7463
rect 28767 7429 28779 7463
rect 30098 7460 30104 7472
rect 29946 7432 30104 7460
rect 28721 7423 28779 7429
rect 30098 7420 30104 7432
rect 30156 7420 30162 7472
rect 30392 7392 30420 7488
rect 31726 7460 31754 7488
rect 31849 7463 31907 7469
rect 31849 7460 31861 7463
rect 31726 7432 31861 7460
rect 31849 7429 31861 7432
rect 31895 7429 31907 7463
rect 34256 7460 34284 7488
rect 34977 7463 35035 7469
rect 34977 7460 34989 7463
rect 34256 7432 34989 7460
rect 31849 7423 31907 7429
rect 34977 7429 34989 7432
rect 35023 7429 35035 7463
rect 34977 7423 35035 7429
rect 35897 7463 35955 7469
rect 35897 7429 35909 7463
rect 35943 7460 35955 7463
rect 35943 7432 37320 7460
rect 35943 7429 35955 7432
rect 35897 7423 35955 7429
rect 29932 7364 30420 7392
rect 26927 7296 28212 7324
rect 28445 7327 28503 7333
rect 26927 7293 26939 7296
rect 26881 7287 26939 7293
rect 28445 7293 28457 7327
rect 28491 7293 28503 7327
rect 29932 7324 29960 7364
rect 31478 7352 31484 7404
rect 31536 7392 31542 7404
rect 31573 7395 31631 7401
rect 31573 7392 31585 7395
rect 31536 7364 31585 7392
rect 31536 7352 31542 7364
rect 31573 7361 31585 7364
rect 31619 7361 31631 7395
rect 31573 7355 31631 7361
rect 32950 7352 32956 7404
rect 33008 7352 33014 7404
rect 34057 7395 34115 7401
rect 34057 7361 34069 7395
rect 34103 7392 34115 7395
rect 34103 7364 34836 7392
rect 34103 7361 34115 7364
rect 34057 7355 34115 7361
rect 28445 7287 28503 7293
rect 28552 7296 29960 7324
rect 30285 7327 30343 7333
rect 22296 7228 22692 7256
rect 17092 7160 17724 7188
rect 18233 7191 18291 7197
rect 17092 7148 17098 7160
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 18322 7188 18328 7200
rect 18279 7160 18328 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 22094 7148 22100 7200
rect 22152 7148 22158 7200
rect 22186 7148 22192 7200
rect 22244 7188 22250 7200
rect 23382 7188 23388 7200
rect 22244 7160 23388 7188
rect 22244 7148 22250 7160
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 24044 7188 24072 7284
rect 27982 7216 27988 7268
rect 28040 7256 28046 7268
rect 28460 7256 28488 7287
rect 28040 7228 28488 7256
rect 28040 7216 28046 7228
rect 24857 7191 24915 7197
rect 24857 7188 24869 7191
rect 24044 7160 24869 7188
rect 24857 7157 24869 7160
rect 24903 7157 24915 7191
rect 24857 7151 24915 7157
rect 25682 7148 25688 7200
rect 25740 7188 25746 7200
rect 28552 7188 28580 7296
rect 30285 7293 30297 7327
rect 30331 7293 30343 7327
rect 30285 7287 30343 7293
rect 30561 7327 30619 7333
rect 30561 7293 30573 7327
rect 30607 7324 30619 7327
rect 34146 7324 34152 7336
rect 30607 7296 30880 7324
rect 30607 7293 30619 7296
rect 30561 7287 30619 7293
rect 25740 7160 28580 7188
rect 25740 7148 25746 7160
rect 28902 7148 28908 7200
rect 28960 7188 28966 7200
rect 29822 7188 29828 7200
rect 28960 7160 29828 7188
rect 28960 7148 28966 7160
rect 29822 7148 29828 7160
rect 29880 7188 29886 7200
rect 30193 7191 30251 7197
rect 30193 7188 30205 7191
rect 29880 7160 30205 7188
rect 29880 7148 29886 7160
rect 30193 7157 30205 7160
rect 30239 7157 30251 7191
rect 30300 7188 30328 7287
rect 30852 7268 30880 7296
rect 31680 7296 34152 7324
rect 30834 7216 30840 7268
rect 30892 7216 30898 7268
rect 31110 7216 31116 7268
rect 31168 7256 31174 7268
rect 31680 7256 31708 7296
rect 34146 7284 34152 7296
rect 34204 7324 34210 7336
rect 34333 7327 34391 7333
rect 34333 7324 34345 7327
rect 34204 7296 34345 7324
rect 34204 7284 34210 7296
rect 34333 7293 34345 7296
rect 34379 7324 34391 7327
rect 34808 7324 34836 7364
rect 34882 7352 34888 7404
rect 34940 7352 34946 7404
rect 37090 7392 37096 7404
rect 34992 7364 37096 7392
rect 34992 7324 35020 7364
rect 37090 7352 37096 7364
rect 37148 7352 37154 7404
rect 37185 7395 37243 7401
rect 37185 7361 37197 7395
rect 37231 7361 37243 7395
rect 37185 7355 37243 7361
rect 34379 7296 34744 7324
rect 34808 7296 35020 7324
rect 34379 7293 34391 7296
rect 34333 7287 34391 7293
rect 34716 7256 34744 7296
rect 35158 7284 35164 7336
rect 35216 7284 35222 7336
rect 36081 7327 36139 7333
rect 36081 7293 36093 7327
rect 36127 7293 36139 7327
rect 36081 7287 36139 7293
rect 35176 7256 35204 7284
rect 31168 7228 31708 7256
rect 33152 7228 34560 7256
rect 34716 7228 35204 7256
rect 36096 7256 36124 7287
rect 36998 7284 37004 7336
rect 37056 7324 37062 7336
rect 37200 7324 37228 7355
rect 37292 7333 37320 7432
rect 37366 7420 37372 7472
rect 37424 7460 37430 7472
rect 38672 7460 38700 7491
rect 39574 7488 39580 7540
rect 39632 7528 39638 7540
rect 40129 7531 40187 7537
rect 40129 7528 40141 7531
rect 39632 7500 40141 7528
rect 39632 7488 39638 7500
rect 40129 7497 40141 7500
rect 40175 7497 40187 7531
rect 40129 7491 40187 7497
rect 40589 7531 40647 7537
rect 40589 7497 40601 7531
rect 40635 7528 40647 7531
rect 40770 7528 40776 7540
rect 40635 7500 40776 7528
rect 40635 7497 40647 7500
rect 40589 7491 40647 7497
rect 40770 7488 40776 7500
rect 40828 7528 40834 7540
rect 42153 7531 42211 7537
rect 42153 7528 42165 7531
rect 40828 7500 42165 7528
rect 40828 7488 40834 7500
rect 42153 7497 42165 7500
rect 42199 7497 42211 7531
rect 42153 7491 42211 7497
rect 43165 7531 43223 7537
rect 43165 7497 43177 7531
rect 43211 7528 43223 7531
rect 43254 7528 43260 7540
rect 43211 7500 43260 7528
rect 43211 7497 43223 7500
rect 43165 7491 43223 7497
rect 43254 7488 43260 7500
rect 43312 7528 43318 7540
rect 43993 7531 44051 7537
rect 43993 7528 44005 7531
rect 43312 7500 44005 7528
rect 43312 7488 43318 7500
rect 43993 7497 44005 7500
rect 44039 7528 44051 7531
rect 44542 7528 44548 7540
rect 44039 7500 44548 7528
rect 44039 7497 44051 7500
rect 43993 7491 44051 7497
rect 44542 7488 44548 7500
rect 44600 7528 44606 7540
rect 44637 7531 44695 7537
rect 44637 7528 44649 7531
rect 44600 7500 44649 7528
rect 44600 7488 44606 7500
rect 44637 7497 44649 7500
rect 44683 7497 44695 7531
rect 44637 7491 44695 7497
rect 39485 7463 39543 7469
rect 37424 7432 39068 7460
rect 37424 7420 37430 7432
rect 38013 7395 38071 7401
rect 38013 7361 38025 7395
rect 38059 7361 38071 7395
rect 38013 7355 38071 7361
rect 38565 7395 38623 7401
rect 38565 7361 38577 7395
rect 38611 7392 38623 7395
rect 38611 7364 38976 7392
rect 38611 7361 38623 7364
rect 38565 7355 38623 7361
rect 37056 7296 37228 7324
rect 37277 7327 37335 7333
rect 37056 7284 37062 7296
rect 37277 7293 37289 7327
rect 37323 7324 37335 7327
rect 37366 7324 37372 7336
rect 37323 7296 37372 7324
rect 37323 7293 37335 7296
rect 37277 7287 37335 7293
rect 37366 7284 37372 7296
rect 37424 7284 37430 7336
rect 37461 7327 37519 7333
rect 37461 7293 37473 7327
rect 37507 7324 37519 7327
rect 37642 7324 37648 7336
rect 37507 7296 37648 7324
rect 37507 7293 37519 7296
rect 37461 7287 37519 7293
rect 37642 7284 37648 7296
rect 37700 7284 37706 7336
rect 37734 7284 37740 7336
rect 37792 7324 37798 7336
rect 38028 7324 38056 7355
rect 37792 7296 38056 7324
rect 37792 7284 37798 7296
rect 36170 7256 36176 7268
rect 36096 7228 36176 7256
rect 31168 7216 31174 7228
rect 33152 7188 33180 7228
rect 30300 7160 33180 7188
rect 30193 7151 30251 7157
rect 33410 7148 33416 7200
rect 33468 7188 33474 7200
rect 34054 7188 34060 7200
rect 33468 7160 34060 7188
rect 33468 7148 33474 7160
rect 34054 7148 34060 7160
rect 34112 7148 34118 7200
rect 34532 7197 34560 7228
rect 36170 7216 36176 7228
rect 36228 7256 36234 7268
rect 36228 7228 38148 7256
rect 36228 7216 36234 7228
rect 34517 7191 34575 7197
rect 34517 7157 34529 7191
rect 34563 7157 34575 7191
rect 34517 7151 34575 7157
rect 34974 7148 34980 7200
rect 35032 7188 35038 7200
rect 37182 7188 37188 7200
rect 35032 7160 37188 7188
rect 35032 7148 35038 7160
rect 37182 7148 37188 7160
rect 37240 7148 37246 7200
rect 38120 7197 38148 7228
rect 38105 7191 38163 7197
rect 38105 7157 38117 7191
rect 38151 7188 38163 7191
rect 38194 7188 38200 7200
rect 38151 7160 38200 7188
rect 38151 7157 38163 7160
rect 38105 7151 38163 7157
rect 38194 7148 38200 7160
rect 38252 7148 38258 7200
rect 38948 7188 38976 7364
rect 39040 7324 39068 7432
rect 39485 7429 39497 7463
rect 39531 7460 39543 7463
rect 40494 7460 40500 7472
rect 39531 7432 40500 7460
rect 39531 7429 39543 7432
rect 39485 7423 39543 7429
rect 40494 7420 40500 7432
rect 40552 7420 40558 7472
rect 44174 7420 44180 7472
rect 44232 7460 44238 7472
rect 44726 7460 44732 7472
rect 44232 7432 44732 7460
rect 44232 7420 44238 7432
rect 44726 7420 44732 7432
rect 44784 7460 44790 7472
rect 45005 7463 45063 7469
rect 45005 7460 45017 7463
rect 44784 7432 45017 7460
rect 44784 7420 44790 7432
rect 45005 7429 45017 7432
rect 45051 7429 45063 7463
rect 45005 7423 45063 7429
rect 39114 7352 39120 7404
rect 39172 7392 39178 7404
rect 39393 7395 39451 7401
rect 39393 7392 39405 7395
rect 39172 7364 39405 7392
rect 39172 7352 39178 7364
rect 39393 7361 39405 7364
rect 39439 7361 39451 7395
rect 40037 7395 40095 7401
rect 40037 7392 40049 7395
rect 39393 7355 39451 7361
rect 39684 7364 40049 7392
rect 39574 7324 39580 7336
rect 39040 7296 39580 7324
rect 39574 7284 39580 7296
rect 39632 7284 39638 7336
rect 39025 7259 39083 7265
rect 39025 7225 39037 7259
rect 39071 7256 39083 7259
rect 39684 7256 39712 7364
rect 40037 7361 40049 7364
rect 40083 7361 40095 7395
rect 40037 7355 40095 7361
rect 41233 7395 41291 7401
rect 41233 7361 41245 7395
rect 41279 7392 41291 7395
rect 41414 7392 41420 7404
rect 41279 7364 41420 7392
rect 41279 7361 41291 7364
rect 41233 7355 41291 7361
rect 41414 7352 41420 7364
rect 41472 7352 41478 7404
rect 41506 7352 41512 7404
rect 41564 7352 41570 7404
rect 42245 7395 42303 7401
rect 42245 7361 42257 7395
rect 42291 7392 42303 7395
rect 43070 7392 43076 7404
rect 42291 7364 43076 7392
rect 42291 7361 42303 7364
rect 42245 7355 42303 7361
rect 43070 7352 43076 7364
rect 43128 7352 43134 7404
rect 40678 7284 40684 7336
rect 40736 7284 40742 7336
rect 42058 7284 42064 7336
rect 42116 7324 42122 7336
rect 42337 7327 42395 7333
rect 42337 7324 42349 7327
rect 42116 7296 42349 7324
rect 42116 7284 42122 7296
rect 42337 7293 42349 7296
rect 42383 7293 42395 7327
rect 42337 7287 42395 7293
rect 40696 7256 40724 7284
rect 44542 7256 44548 7268
rect 39071 7228 39712 7256
rect 39776 7228 44548 7256
rect 39071 7225 39083 7228
rect 39025 7219 39083 7225
rect 39776 7188 39804 7228
rect 44542 7216 44548 7228
rect 44600 7216 44606 7268
rect 38948 7160 39804 7188
rect 39850 7148 39856 7200
rect 39908 7148 39914 7200
rect 40954 7148 40960 7200
rect 41012 7188 41018 7200
rect 41049 7191 41107 7197
rect 41049 7188 41061 7191
rect 41012 7160 41061 7188
rect 41012 7148 41018 7160
rect 41049 7157 41061 7160
rect 41095 7157 41107 7191
rect 41049 7151 41107 7157
rect 41322 7148 41328 7200
rect 41380 7148 41386 7200
rect 41414 7148 41420 7200
rect 41472 7188 41478 7200
rect 41785 7191 41843 7197
rect 41785 7188 41797 7191
rect 41472 7160 41797 7188
rect 41472 7148 41478 7160
rect 41785 7157 41797 7160
rect 41831 7157 41843 7191
rect 41785 7151 41843 7157
rect 41874 7148 41880 7200
rect 41932 7188 41938 7200
rect 42797 7191 42855 7197
rect 42797 7188 42809 7191
rect 41932 7160 42809 7188
rect 41932 7148 41938 7160
rect 42797 7157 42809 7160
rect 42843 7188 42855 7191
rect 43438 7188 43444 7200
rect 42843 7160 43444 7188
rect 42843 7157 42855 7160
rect 42797 7151 42855 7157
rect 43438 7148 43444 7160
rect 43496 7188 43502 7200
rect 43533 7191 43591 7197
rect 43533 7188 43545 7191
rect 43496 7160 43545 7188
rect 43496 7148 43502 7160
rect 43533 7157 43545 7160
rect 43579 7188 43591 7191
rect 44269 7191 44327 7197
rect 44269 7188 44281 7191
rect 43579 7160 44281 7188
rect 43579 7157 43591 7160
rect 43533 7151 43591 7157
rect 44269 7157 44281 7160
rect 44315 7157 44327 7191
rect 44269 7151 44327 7157
rect 460 7098 45540 7120
rect 460 7046 3570 7098
rect 3622 7046 3634 7098
rect 3686 7046 3698 7098
rect 3750 7046 3762 7098
rect 3814 7046 3826 7098
rect 3878 7046 8570 7098
rect 8622 7046 8634 7098
rect 8686 7046 8698 7098
rect 8750 7046 8762 7098
rect 8814 7046 8826 7098
rect 8878 7046 13570 7098
rect 13622 7046 13634 7098
rect 13686 7046 13698 7098
rect 13750 7046 13762 7098
rect 13814 7046 13826 7098
rect 13878 7046 18570 7098
rect 18622 7046 18634 7098
rect 18686 7046 18698 7098
rect 18750 7046 18762 7098
rect 18814 7046 18826 7098
rect 18878 7046 23570 7098
rect 23622 7046 23634 7098
rect 23686 7046 23698 7098
rect 23750 7046 23762 7098
rect 23814 7046 23826 7098
rect 23878 7046 28570 7098
rect 28622 7046 28634 7098
rect 28686 7046 28698 7098
rect 28750 7046 28762 7098
rect 28814 7046 28826 7098
rect 28878 7046 33570 7098
rect 33622 7046 33634 7098
rect 33686 7046 33698 7098
rect 33750 7046 33762 7098
rect 33814 7046 33826 7098
rect 33878 7046 38570 7098
rect 38622 7046 38634 7098
rect 38686 7046 38698 7098
rect 38750 7046 38762 7098
rect 38814 7046 38826 7098
rect 38878 7046 43570 7098
rect 43622 7046 43634 7098
rect 43686 7046 43698 7098
rect 43750 7046 43762 7098
rect 43814 7046 43826 7098
rect 43878 7046 45540 7098
rect 460 7024 45540 7046
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7650 6984 7656 6996
rect 7055 6956 7656 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10137 6987 10195 6993
rect 10137 6984 10149 6987
rect 10100 6956 10149 6984
rect 10100 6944 10106 6956
rect 10137 6953 10149 6956
rect 10183 6953 10195 6987
rect 10137 6947 10195 6953
rect 10594 6944 10600 6996
rect 10652 6944 10658 6996
rect 11057 6987 11115 6993
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11333 6987 11391 6993
rect 11333 6984 11345 6987
rect 11103 6956 11345 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11333 6953 11345 6956
rect 11379 6984 11391 6987
rect 11882 6984 11888 6996
rect 11379 6956 11888 6984
rect 11379 6953 11391 6956
rect 11333 6947 11391 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 15102 6993 15108 6996
rect 15092 6987 15108 6993
rect 15092 6953 15104 6987
rect 15092 6947 15108 6953
rect 15102 6944 15108 6947
rect 15160 6944 15166 6996
rect 16574 6944 16580 6996
rect 16632 6944 16638 6996
rect 17034 6944 17040 6996
rect 17092 6944 17098 6996
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 17954 6984 17960 6996
rect 17368 6956 17960 6984
rect 17368 6944 17374 6956
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 18414 6944 18420 6996
rect 18472 6984 18478 6996
rect 19521 6987 19579 6993
rect 19521 6984 19533 6987
rect 18472 6956 19533 6984
rect 18472 6944 18478 6956
rect 19521 6953 19533 6956
rect 19567 6953 19579 6987
rect 19521 6947 19579 6953
rect 20622 6944 20628 6996
rect 20680 6944 20686 6996
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 20956 6956 22784 6984
rect 20956 6944 20962 6956
rect 8113 6919 8171 6925
rect 8113 6885 8125 6919
rect 8159 6916 8171 6919
rect 8938 6916 8944 6928
rect 8159 6888 8944 6916
rect 8159 6885 8171 6888
rect 8113 6879 8171 6885
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6848 7343 6851
rect 8128 6848 8156 6879
rect 8938 6876 8944 6888
rect 8996 6916 9002 6928
rect 9217 6919 9275 6925
rect 9217 6916 9229 6919
rect 8996 6888 9229 6916
rect 8996 6876 9002 6888
rect 9217 6885 9229 6888
rect 9263 6916 9275 6919
rect 9582 6916 9588 6928
rect 9263 6888 9588 6916
rect 9263 6885 9275 6888
rect 9217 6879 9275 6885
rect 9582 6876 9588 6888
rect 9640 6916 9646 6928
rect 9640 6876 9674 6916
rect 7331 6820 8156 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 9456 6820 9505 6848
rect 9456 6808 9462 6820
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9646 6848 9674 6876
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9646 6820 9965 6848
rect 9493 6811 9551 6817
rect 9953 6817 9965 6820
rect 9999 6848 10011 6851
rect 10321 6851 10379 6857
rect 9999 6820 10272 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8478 6780 8484 6792
rect 7791 6752 8484 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10244 6780 10272 6820
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10612 6848 10640 6944
rect 16669 6919 16727 6925
rect 16669 6885 16681 6919
rect 16715 6916 16727 6919
rect 17862 6916 17868 6928
rect 16715 6888 17868 6916
rect 16715 6885 16727 6888
rect 16669 6879 16727 6885
rect 10367 6820 10640 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16684 6848 16712 6879
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 17972 6916 18000 6944
rect 19153 6919 19211 6925
rect 19153 6916 19165 6919
rect 17972 6888 19165 6916
rect 19153 6885 19165 6888
rect 19199 6885 19211 6919
rect 20530 6916 20536 6928
rect 19153 6879 19211 6885
rect 19536 6888 20536 6916
rect 19536 6860 19564 6888
rect 20530 6876 20536 6888
rect 20588 6916 20594 6928
rect 20588 6888 21036 6916
rect 20588 6876 20594 6888
rect 15804 6820 16712 6848
rect 15804 6808 15810 6820
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 17678 6848 17684 6860
rect 16816 6820 17684 6848
rect 16816 6808 16822 6820
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 18340 6820 19472 6848
rect 18340 6792 18368 6820
rect 14829 6783 14887 6789
rect 10244 6752 10640 6780
rect 10045 6743 10103 6749
rect 10060 6712 10088 6743
rect 10410 6712 10416 6724
rect 10060 6684 10416 6712
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10612 6656 10640 6752
rect 14829 6749 14841 6783
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 12526 6712 12532 6724
rect 12084 6684 12532 6712
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 7708 6616 8769 6644
rect 7708 6604 7714 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 10284 6616 10333 6644
rect 10284 6604 10290 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 12084 6653 12112 6684
rect 12526 6672 12532 6684
rect 12584 6712 12590 6724
rect 12805 6715 12863 6721
rect 12805 6712 12817 6715
rect 12584 6684 12817 6712
rect 12584 6672 12590 6684
rect 12805 6681 12817 6684
rect 12851 6712 12863 6715
rect 13909 6715 13967 6721
rect 13909 6712 13921 6715
rect 12851 6684 13921 6712
rect 12851 6681 12863 6684
rect 12805 6675 12863 6681
rect 13909 6681 13921 6684
rect 13955 6712 13967 6715
rect 14277 6715 14335 6721
rect 14277 6712 14289 6715
rect 13955 6684 14289 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 14277 6681 14289 6684
rect 14323 6712 14335 6715
rect 14642 6712 14648 6724
rect 14323 6684 14648 6712
rect 14323 6681 14335 6684
rect 14277 6675 14335 6681
rect 14642 6672 14648 6684
rect 14700 6712 14706 6724
rect 14844 6712 14872 6743
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 17497 6783 17555 6789
rect 16540 6752 17448 6780
rect 16540 6740 16546 6752
rect 15378 6712 15384 6724
rect 14700 6684 15384 6712
rect 14700 6672 14706 6684
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 15654 6672 15660 6724
rect 15712 6672 15718 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 17037 6715 17095 6721
rect 17037 6712 17049 6715
rect 16816 6684 17049 6712
rect 16816 6672 16822 6684
rect 17037 6681 17049 6684
rect 17083 6681 17095 6715
rect 17313 6715 17371 6721
rect 17313 6712 17325 6715
rect 17037 6675 17095 6681
rect 17144 6684 17325 6712
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 10652 6616 11713 6644
rect 10652 6604 10658 6616
rect 11701 6613 11713 6616
rect 11747 6644 11759 6647
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 11747 6616 12081 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12618 6644 12624 6656
rect 12483 6616 12624 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12618 6604 12624 6616
rect 12676 6644 12682 6656
rect 13078 6644 13084 6656
rect 12676 6616 13084 6644
rect 12676 6604 12682 6616
rect 13078 6604 13084 6616
rect 13136 6644 13142 6656
rect 13173 6647 13231 6653
rect 13173 6644 13185 6647
rect 13136 6616 13185 6644
rect 13136 6604 13142 6616
rect 13173 6613 13185 6616
rect 13219 6613 13231 6647
rect 13173 6607 13231 6613
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 17144 6644 17172 6684
rect 17313 6681 17325 6684
rect 17359 6681 17371 6715
rect 17420 6712 17448 6752
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17586 6780 17592 6792
rect 17543 6752 17592 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 19334 6740 19340 6792
rect 19392 6740 19398 6792
rect 19444 6789 19472 6820
rect 19518 6808 19524 6860
rect 19576 6808 19582 6860
rect 20438 6848 20444 6860
rect 20088 6820 20444 6848
rect 20088 6789 20116 6820
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 21008 6857 21036 6888
rect 22370 6876 22376 6928
rect 22428 6876 22434 6928
rect 22756 6916 22784 6956
rect 22830 6944 22836 6996
rect 22888 6944 22894 6996
rect 24210 6984 24216 6996
rect 23124 6956 24216 6984
rect 23124 6916 23152 6956
rect 24210 6944 24216 6956
rect 24268 6944 24274 6996
rect 24302 6944 24308 6996
rect 24360 6944 24366 6996
rect 26418 6944 26424 6996
rect 26476 6984 26482 6996
rect 26789 6987 26847 6993
rect 26789 6984 26801 6987
rect 26476 6956 26801 6984
rect 26476 6944 26482 6956
rect 26789 6953 26801 6956
rect 26835 6953 26847 6987
rect 26789 6947 26847 6953
rect 27706 6944 27712 6996
rect 27764 6984 27770 6996
rect 27982 6984 27988 6996
rect 27764 6956 27988 6984
rect 27764 6944 27770 6956
rect 27982 6944 27988 6956
rect 28040 6984 28046 6996
rect 28718 6984 28724 6996
rect 28040 6956 28724 6984
rect 28040 6944 28046 6956
rect 28718 6944 28724 6956
rect 28776 6944 28782 6996
rect 33689 6987 33747 6993
rect 28966 6956 30236 6984
rect 22756 6888 23152 6916
rect 23198 6876 23204 6928
rect 23256 6916 23262 6928
rect 24320 6916 24348 6944
rect 25314 6916 25320 6928
rect 23256 6888 24348 6916
rect 25056 6888 25320 6916
rect 23256 6876 23262 6888
rect 20993 6851 21051 6857
rect 20772 6820 20852 6848
rect 20772 6808 20778 6820
rect 20824 6789 20852 6820
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 22002 6848 22008 6860
rect 21039 6820 22008 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 22388 6848 22416 6876
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22388 6820 22753 6848
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 22741 6811 22799 6817
rect 19430 6783 19488 6789
rect 19430 6749 19442 6783
rect 19476 6749 19488 6783
rect 19430 6743 19488 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 20809 6783 20867 6789
rect 20303 6752 20484 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 18414 6712 18420 6724
rect 17420 6684 18420 6712
rect 17313 6675 17371 6681
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 19812 6712 19840 6743
rect 19260 6684 19840 6712
rect 19996 6712 20024 6743
rect 20456 6712 20484 6752
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 22370 6740 22376 6792
rect 22428 6740 22434 6792
rect 22646 6740 22652 6792
rect 22704 6782 22710 6792
rect 23216 6789 23244 6876
rect 23290 6808 23296 6860
rect 23348 6808 23354 6860
rect 23385 6851 23443 6857
rect 23385 6817 23397 6851
rect 23431 6817 23443 6851
rect 23385 6811 23443 6817
rect 23201 6783 23259 6789
rect 22704 6754 22784 6782
rect 22704 6740 22710 6754
rect 20990 6712 20996 6724
rect 19996 6684 20392 6712
rect 20456 6684 20996 6712
rect 19260 6656 19288 6684
rect 20364 6656 20392 6684
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 21269 6715 21327 6721
rect 21269 6681 21281 6715
rect 21315 6712 21327 6715
rect 21542 6712 21548 6724
rect 21315 6684 21548 6712
rect 21315 6681 21327 6684
rect 21269 6675 21327 6681
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 22756 6712 22784 6754
rect 23201 6749 23213 6783
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 23400 6712 23428 6811
rect 24670 6808 24676 6860
rect 24728 6808 24734 6860
rect 24305 6715 24363 6721
rect 24305 6712 24317 6715
rect 22756 6684 23428 6712
rect 23952 6684 24317 6712
rect 15896 6616 17172 6644
rect 15896 6604 15902 6616
rect 17218 6604 17224 6656
rect 17276 6604 17282 6656
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 18325 6647 18383 6653
rect 18325 6644 18337 6647
rect 17460 6616 18337 6644
rect 17460 6604 17466 6616
rect 18325 6613 18337 6616
rect 18371 6644 18383 6647
rect 18506 6644 18512 6656
rect 18371 6616 18512 6644
rect 18371 6613 18383 6616
rect 18325 6607 18383 6613
rect 18506 6604 18512 6616
rect 18564 6644 18570 6656
rect 18785 6647 18843 6653
rect 18785 6644 18797 6647
rect 18564 6616 18797 6644
rect 18564 6604 18570 6616
rect 18785 6613 18797 6616
rect 18831 6644 18843 6647
rect 19150 6644 19156 6656
rect 18831 6616 19156 6644
rect 18831 6613 18843 6616
rect 18785 6607 18843 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19242 6604 19248 6656
rect 19300 6604 19306 6656
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 19886 6644 19892 6656
rect 19484 6616 19892 6644
rect 19484 6604 19490 6616
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 19978 6604 19984 6656
rect 20036 6604 20042 6656
rect 20162 6604 20168 6656
rect 20220 6604 20226 6656
rect 20346 6604 20352 6656
rect 20404 6604 20410 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 23952 6653 23980 6684
rect 24305 6681 24317 6684
rect 24351 6712 24363 6715
rect 25056 6712 25084 6888
rect 25314 6876 25320 6888
rect 25372 6916 25378 6928
rect 25372 6888 26556 6916
rect 25372 6876 25378 6888
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6848 25191 6851
rect 25590 6848 25596 6860
rect 25179 6820 25596 6848
rect 25179 6817 25191 6820
rect 25133 6811 25191 6817
rect 25590 6808 25596 6820
rect 25648 6848 25654 6860
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 25648 6820 26433 6848
rect 25648 6808 25654 6820
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26528 6848 26556 6888
rect 26602 6876 26608 6928
rect 26660 6916 26666 6928
rect 27724 6916 27752 6944
rect 28966 6916 28994 6956
rect 26660 6888 27752 6916
rect 28092 6888 28994 6916
rect 26660 6876 26666 6888
rect 27157 6851 27215 6857
rect 27157 6848 27169 6851
rect 26528 6820 27169 6848
rect 26421 6811 26479 6817
rect 27157 6817 27169 6820
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 25958 6740 25964 6792
rect 26016 6740 26022 6792
rect 27430 6740 27436 6792
rect 27488 6740 27494 6792
rect 28092 6780 28120 6888
rect 28169 6851 28227 6857
rect 28169 6817 28181 6851
rect 28215 6848 28227 6851
rect 29181 6851 29239 6857
rect 29181 6848 29193 6851
rect 28215 6820 29193 6848
rect 28215 6817 28227 6820
rect 28169 6811 28227 6817
rect 29181 6817 29193 6820
rect 29227 6817 29239 6851
rect 30208 6848 30236 6956
rect 31588 6956 32168 6984
rect 30282 6876 30288 6928
rect 30340 6916 30346 6928
rect 31478 6916 31484 6928
rect 30340 6888 31484 6916
rect 30340 6876 30346 6888
rect 31128 6857 31156 6888
rect 31478 6876 31484 6888
rect 31536 6876 31542 6928
rect 31021 6851 31079 6857
rect 31021 6848 31033 6851
rect 30208 6820 30512 6848
rect 29181 6811 29239 6817
rect 30484 6792 30512 6820
rect 30852 6820 31033 6848
rect 30852 6792 30880 6820
rect 31021 6817 31033 6820
rect 31067 6817 31079 6851
rect 31021 6811 31079 6817
rect 31113 6851 31171 6857
rect 31113 6817 31125 6851
rect 31159 6817 31171 6851
rect 31113 6811 31171 6817
rect 31205 6851 31263 6857
rect 31205 6817 31217 6851
rect 31251 6848 31263 6851
rect 31588 6848 31616 6956
rect 31251 6820 31616 6848
rect 31680 6888 31984 6916
rect 31251 6817 31263 6820
rect 31205 6811 31263 6817
rect 28353 6783 28411 6789
rect 28353 6780 28365 6783
rect 28092 6752 28365 6780
rect 28353 6749 28365 6752
rect 28399 6749 28411 6783
rect 28353 6743 28411 6749
rect 28445 6783 28503 6789
rect 28445 6749 28457 6783
rect 28491 6749 28503 6783
rect 28445 6743 28503 6749
rect 25409 6715 25467 6721
rect 25409 6712 25421 6715
rect 24351 6684 25421 6712
rect 24351 6681 24363 6684
rect 24305 6675 24363 6681
rect 25409 6681 25421 6684
rect 25455 6681 25467 6715
rect 25409 6675 25467 6681
rect 25685 6715 25743 6721
rect 25685 6681 25697 6715
rect 25731 6712 25743 6715
rect 27798 6712 27804 6724
rect 25731 6684 27804 6712
rect 25731 6681 25743 6684
rect 25685 6675 25743 6681
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 22244 6616 23949 6644
rect 22244 6604 22250 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 24210 6604 24216 6656
rect 24268 6644 24274 6656
rect 25038 6644 25044 6656
rect 24268 6616 25044 6644
rect 24268 6604 24274 6616
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 25648 6616 25789 6644
rect 25648 6604 25654 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 26142 6604 26148 6656
rect 26200 6604 26206 6656
rect 27430 6604 27436 6656
rect 27488 6644 27494 6656
rect 27617 6647 27675 6653
rect 27617 6644 27629 6647
rect 27488 6616 27629 6644
rect 27488 6604 27494 6616
rect 27617 6613 27629 6616
rect 27663 6613 27675 6647
rect 28460 6644 28488 6743
rect 28534 6740 28540 6792
rect 28592 6740 28598 6792
rect 28629 6783 28687 6789
rect 28629 6749 28641 6783
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 28644 6712 28672 6743
rect 28718 6740 28724 6792
rect 28776 6780 28782 6792
rect 28905 6783 28963 6789
rect 28905 6780 28917 6783
rect 28776 6752 28917 6780
rect 28776 6740 28782 6752
rect 28905 6749 28917 6752
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 30282 6740 30288 6792
rect 30340 6740 30346 6792
rect 30466 6740 30472 6792
rect 30524 6740 30530 6792
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 30834 6740 30840 6792
rect 30892 6740 30898 6792
rect 30929 6783 30987 6789
rect 30929 6749 30941 6783
rect 30975 6749 30987 6783
rect 31680 6780 31708 6888
rect 31757 6851 31815 6857
rect 31757 6817 31769 6851
rect 31803 6848 31815 6851
rect 31956 6848 31984 6888
rect 32033 6851 32091 6857
rect 32033 6848 32045 6851
rect 31803 6820 31892 6848
rect 31956 6820 32045 6848
rect 31803 6817 31815 6820
rect 31757 6811 31815 6817
rect 30929 6743 30987 6749
rect 31036 6752 31708 6780
rect 29454 6712 29460 6724
rect 28644 6684 29460 6712
rect 29454 6672 29460 6684
rect 29512 6672 29518 6724
rect 30484 6712 30512 6740
rect 30760 6712 30788 6740
rect 30944 6712 30972 6743
rect 31036 6724 31064 6752
rect 30484 6684 30972 6712
rect 31018 6672 31024 6724
rect 31076 6672 31082 6724
rect 31386 6672 31392 6724
rect 31444 6672 31450 6724
rect 31864 6712 31892 6820
rect 32033 6817 32045 6820
rect 32079 6817 32091 6851
rect 32140 6848 32168 6956
rect 33689 6953 33701 6987
rect 33735 6984 33747 6987
rect 33962 6984 33968 6996
rect 33735 6956 33968 6984
rect 33735 6953 33747 6956
rect 33689 6947 33747 6953
rect 33962 6944 33968 6956
rect 34020 6984 34026 6996
rect 34241 6987 34299 6993
rect 34241 6984 34253 6987
rect 34020 6956 34253 6984
rect 34020 6944 34026 6956
rect 34241 6953 34253 6956
rect 34287 6953 34299 6987
rect 34241 6947 34299 6953
rect 34422 6944 34428 6996
rect 34480 6944 34486 6996
rect 34882 6944 34888 6996
rect 34940 6984 34946 6996
rect 39472 6987 39530 6993
rect 34940 6956 39344 6984
rect 34940 6944 34946 6956
rect 32784 6888 33824 6916
rect 32784 6848 32812 6888
rect 32140 6820 32812 6848
rect 32033 6811 32091 6817
rect 32858 6808 32864 6860
rect 32916 6848 32922 6860
rect 33137 6851 33195 6857
rect 33137 6848 33149 6851
rect 32916 6820 33149 6848
rect 32916 6808 32922 6820
rect 33137 6817 33149 6820
rect 33183 6817 33195 6851
rect 33137 6811 33195 6817
rect 33321 6851 33379 6857
rect 33321 6817 33333 6851
rect 33367 6848 33379 6851
rect 33686 6848 33692 6860
rect 33367 6820 33692 6848
rect 33367 6817 33379 6820
rect 33321 6811 33379 6817
rect 33686 6808 33692 6820
rect 33744 6808 33750 6860
rect 33796 6848 33824 6888
rect 34974 6876 34980 6928
rect 35032 6876 35038 6928
rect 35360 6888 37044 6916
rect 34992 6848 35020 6876
rect 35360 6857 35388 6888
rect 33796 6820 35020 6848
rect 35345 6851 35403 6857
rect 35345 6817 35357 6851
rect 35391 6817 35403 6851
rect 35345 6811 35403 6817
rect 36173 6851 36231 6857
rect 36173 6817 36185 6851
rect 36219 6817 36231 6851
rect 36173 6811 36231 6817
rect 31938 6740 31944 6792
rect 31996 6780 32002 6792
rect 35897 6783 35955 6789
rect 31996 6755 33778 6780
rect 31996 6752 33793 6755
rect 31996 6740 32002 6752
rect 33735 6749 33793 6752
rect 31864 6684 32720 6712
rect 29546 6644 29552 6656
rect 28460 6616 29552 6644
rect 27617 6607 27675 6613
rect 29546 6604 29552 6616
rect 29604 6644 29610 6656
rect 30653 6647 30711 6653
rect 30653 6644 30665 6647
rect 29604 6616 30665 6644
rect 29604 6604 29610 6616
rect 30653 6613 30665 6616
rect 30699 6613 30711 6647
rect 30653 6607 30711 6613
rect 30742 6604 30748 6656
rect 30800 6604 30806 6656
rect 31404 6644 31432 6672
rect 31570 6644 31576 6656
rect 31404 6616 31576 6644
rect 31570 6604 31576 6616
rect 31628 6604 31634 6656
rect 31665 6647 31723 6653
rect 31665 6613 31677 6647
rect 31711 6644 31723 6647
rect 32490 6644 32496 6656
rect 31711 6616 32496 6644
rect 31711 6613 31723 6616
rect 31665 6607 31723 6613
rect 32490 6604 32496 6616
rect 32548 6604 32554 6656
rect 32692 6653 32720 6684
rect 33410 6672 33416 6724
rect 33468 6712 33474 6724
rect 33505 6715 33563 6721
rect 33505 6712 33517 6715
rect 33468 6684 33517 6712
rect 33468 6672 33474 6684
rect 33505 6681 33517 6684
rect 33551 6681 33563 6715
rect 33735 6715 33747 6749
rect 33781 6715 33793 6749
rect 35897 6749 35909 6783
rect 35943 6780 35955 6783
rect 35986 6780 35992 6792
rect 35943 6752 35992 6780
rect 35943 6749 35955 6752
rect 35897 6743 35955 6749
rect 35986 6740 35992 6752
rect 36044 6740 36050 6792
rect 36188 6724 36216 6811
rect 36906 6808 36912 6860
rect 36964 6808 36970 6860
rect 37016 6848 37044 6888
rect 37734 6876 37740 6928
rect 37792 6916 37798 6928
rect 37792 6888 38240 6916
rect 37792 6876 37798 6888
rect 37918 6848 37924 6860
rect 37016 6820 37924 6848
rect 37918 6808 37924 6820
rect 37976 6808 37982 6860
rect 38212 6848 38240 6888
rect 38657 6851 38715 6857
rect 38657 6848 38669 6851
rect 38212 6820 38669 6848
rect 38657 6817 38669 6820
rect 38703 6817 38715 6851
rect 38657 6811 38715 6817
rect 39206 6808 39212 6860
rect 39264 6808 39270 6860
rect 39316 6848 39344 6956
rect 39472 6953 39484 6987
rect 39518 6984 39530 6987
rect 39850 6984 39856 6996
rect 39518 6956 39856 6984
rect 39518 6953 39530 6956
rect 39472 6947 39530 6953
rect 39850 6944 39856 6956
rect 39908 6944 39914 6996
rect 40494 6944 40500 6996
rect 40552 6984 40558 6996
rect 41322 6993 41328 6996
rect 40957 6987 41015 6993
rect 40957 6984 40969 6987
rect 40552 6956 40969 6984
rect 40552 6944 40558 6956
rect 40957 6953 40969 6956
rect 41003 6953 41015 6987
rect 40957 6947 41015 6953
rect 41312 6987 41328 6993
rect 41312 6953 41324 6987
rect 41312 6947 41328 6953
rect 41322 6944 41328 6947
rect 41380 6944 41386 6996
rect 43438 6944 43444 6996
rect 43496 6984 43502 6996
rect 43901 6987 43959 6993
rect 43901 6984 43913 6987
rect 43496 6956 43913 6984
rect 43496 6944 43502 6956
rect 43901 6953 43913 6956
rect 43947 6984 43959 6987
rect 44545 6987 44603 6993
rect 44545 6984 44557 6987
rect 43947 6956 44557 6984
rect 43947 6953 43959 6956
rect 43901 6947 43959 6953
rect 44545 6953 44557 6956
rect 44591 6953 44603 6987
rect 44545 6947 44603 6953
rect 44910 6944 44916 6996
rect 44968 6944 44974 6996
rect 40678 6848 40684 6860
rect 39316 6820 40684 6848
rect 40678 6808 40684 6820
rect 40736 6808 40742 6860
rect 41049 6851 41107 6857
rect 41049 6848 41061 6851
rect 40880 6820 41061 6848
rect 40880 6792 40908 6820
rect 41049 6817 41061 6820
rect 41095 6848 41107 6851
rect 41874 6848 41880 6860
rect 41095 6820 41880 6848
rect 41095 6817 41107 6820
rect 41049 6811 41107 6817
rect 41874 6808 41880 6820
rect 41932 6808 41938 6860
rect 42518 6848 42524 6860
rect 42444 6820 42524 6848
rect 36722 6740 36728 6792
rect 36780 6740 36786 6792
rect 37461 6783 37519 6789
rect 37461 6749 37473 6783
rect 37507 6780 37519 6783
rect 38473 6783 38531 6789
rect 37507 6752 38148 6780
rect 37507 6749 37519 6752
rect 37461 6743 37519 6749
rect 33735 6709 33793 6715
rect 33505 6675 33563 6681
rect 34054 6672 34060 6724
rect 34112 6672 34118 6724
rect 34273 6715 34331 6721
rect 34273 6681 34285 6715
rect 34319 6712 34331 6715
rect 34606 6712 34612 6724
rect 34319 6684 34612 6712
rect 34319 6681 34331 6684
rect 34273 6675 34331 6681
rect 34606 6672 34612 6684
rect 34664 6672 34670 6724
rect 35161 6715 35219 6721
rect 35161 6681 35173 6715
rect 35207 6712 35219 6715
rect 35250 6712 35256 6724
rect 35207 6684 35256 6712
rect 35207 6681 35219 6684
rect 35161 6675 35219 6681
rect 35250 6672 35256 6684
rect 35308 6712 35314 6724
rect 35308 6684 35756 6712
rect 35308 6672 35314 6684
rect 32677 6647 32735 6653
rect 32677 6613 32689 6647
rect 32723 6613 32735 6647
rect 32677 6607 32735 6613
rect 33045 6647 33103 6653
rect 33045 6613 33057 6647
rect 33091 6644 33103 6647
rect 33778 6644 33784 6656
rect 33091 6616 33784 6644
rect 33091 6613 33103 6616
rect 33045 6607 33103 6613
rect 33778 6604 33784 6616
rect 33836 6604 33842 6656
rect 33873 6647 33931 6653
rect 33873 6613 33885 6647
rect 33919 6644 33931 6647
rect 33962 6644 33968 6656
rect 33919 6616 33968 6644
rect 33919 6613 33931 6616
rect 33873 6607 33931 6613
rect 33962 6604 33968 6616
rect 34020 6604 34026 6656
rect 34698 6604 34704 6656
rect 34756 6604 34762 6656
rect 34882 6604 34888 6656
rect 34940 6644 34946 6656
rect 35069 6647 35127 6653
rect 35069 6644 35081 6647
rect 34940 6616 35081 6644
rect 34940 6604 34946 6616
rect 35069 6613 35081 6616
rect 35115 6613 35127 6647
rect 35069 6607 35127 6613
rect 35526 6604 35532 6656
rect 35584 6604 35590 6656
rect 35728 6644 35756 6684
rect 36170 6672 36176 6724
rect 36228 6672 36234 6724
rect 37645 6715 37703 6721
rect 37645 6681 37657 6715
rect 37691 6712 37703 6715
rect 38010 6712 38016 6724
rect 37691 6684 38016 6712
rect 37691 6681 37703 6684
rect 37645 6675 37703 6681
rect 38010 6672 38016 6684
rect 38068 6672 38074 6724
rect 35989 6647 36047 6653
rect 35989 6644 36001 6647
rect 35728 6616 36001 6644
rect 35989 6613 36001 6616
rect 36035 6613 36047 6647
rect 35989 6607 36047 6613
rect 36357 6647 36415 6653
rect 36357 6613 36369 6647
rect 36403 6644 36415 6647
rect 36446 6644 36452 6656
rect 36403 6616 36452 6644
rect 36403 6613 36415 6616
rect 36357 6607 36415 6613
rect 36446 6604 36452 6616
rect 36504 6604 36510 6656
rect 36814 6604 36820 6656
rect 36872 6604 36878 6656
rect 37274 6604 37280 6656
rect 37332 6604 37338 6656
rect 38120 6653 38148 6752
rect 38473 6749 38485 6783
rect 38519 6780 38531 6783
rect 39114 6780 39120 6792
rect 38519 6752 39120 6780
rect 38519 6749 38531 6752
rect 38473 6743 38531 6749
rect 39114 6740 39120 6752
rect 39172 6740 39178 6792
rect 40862 6740 40868 6792
rect 40920 6740 40926 6792
rect 40710 6684 41000 6712
rect 38105 6647 38163 6653
rect 38105 6613 38117 6647
rect 38151 6613 38163 6647
rect 38105 6607 38163 6613
rect 38565 6647 38623 6653
rect 38565 6613 38577 6647
rect 38611 6644 38623 6647
rect 38838 6644 38844 6656
rect 38611 6616 38844 6644
rect 38611 6613 38623 6616
rect 38565 6607 38623 6613
rect 38838 6604 38844 6616
rect 38896 6604 38902 6656
rect 40310 6604 40316 6656
rect 40368 6644 40374 6656
rect 40972 6644 41000 6684
rect 42444 6644 42472 6820
rect 42518 6808 42524 6820
rect 42576 6808 42582 6860
rect 42794 6808 42800 6860
rect 42852 6848 42858 6860
rect 43349 6851 43407 6857
rect 43349 6848 43361 6851
rect 42852 6820 43361 6848
rect 42852 6808 42858 6820
rect 43349 6817 43361 6820
rect 43395 6817 43407 6851
rect 43349 6811 43407 6817
rect 43533 6851 43591 6857
rect 43533 6817 43545 6851
rect 43579 6848 43591 6851
rect 44174 6848 44180 6860
rect 43579 6820 44180 6848
rect 43579 6817 43591 6820
rect 43533 6811 43591 6817
rect 44174 6808 44180 6820
rect 44232 6808 44238 6860
rect 42886 6740 42892 6792
rect 42944 6740 42950 6792
rect 42904 6653 42932 6740
rect 40368 6616 42472 6644
rect 42889 6647 42947 6653
rect 40368 6604 40374 6616
rect 42889 6613 42901 6647
rect 42935 6613 42947 6647
rect 42889 6607 42947 6613
rect 43254 6604 43260 6656
rect 43312 6604 43318 6656
rect 460 6554 45540 6576
rect 460 6502 6070 6554
rect 6122 6502 6134 6554
rect 6186 6502 6198 6554
rect 6250 6502 6262 6554
rect 6314 6502 6326 6554
rect 6378 6502 11070 6554
rect 11122 6502 11134 6554
rect 11186 6502 11198 6554
rect 11250 6502 11262 6554
rect 11314 6502 11326 6554
rect 11378 6502 16070 6554
rect 16122 6502 16134 6554
rect 16186 6502 16198 6554
rect 16250 6502 16262 6554
rect 16314 6502 16326 6554
rect 16378 6502 21070 6554
rect 21122 6502 21134 6554
rect 21186 6502 21198 6554
rect 21250 6502 21262 6554
rect 21314 6502 21326 6554
rect 21378 6502 26070 6554
rect 26122 6502 26134 6554
rect 26186 6502 26198 6554
rect 26250 6502 26262 6554
rect 26314 6502 26326 6554
rect 26378 6502 31070 6554
rect 31122 6502 31134 6554
rect 31186 6502 31198 6554
rect 31250 6502 31262 6554
rect 31314 6502 31326 6554
rect 31378 6502 36070 6554
rect 36122 6502 36134 6554
rect 36186 6502 36198 6554
rect 36250 6502 36262 6554
rect 36314 6502 36326 6554
rect 36378 6502 41070 6554
rect 41122 6502 41134 6554
rect 41186 6502 41198 6554
rect 41250 6502 41262 6554
rect 41314 6502 41326 6554
rect 41378 6502 45540 6554
rect 460 6480 45540 6502
rect 15010 6440 15016 6452
rect 2746 6412 15016 6440
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 2746 6304 2774 6412
rect 15010 6400 15016 6412
rect 15068 6400 15074 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15988 6412 16405 6440
rect 15988 6400 15994 6412
rect 16393 6409 16405 6412
rect 16439 6440 16451 6443
rect 16574 6440 16580 6452
rect 16439 6412 16580 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17954 6440 17960 6452
rect 17000 6412 17172 6440
rect 17000 6400 17006 6412
rect 7650 6332 7656 6384
rect 7708 6332 7714 6384
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 9398 6372 9404 6384
rect 8159 6344 9404 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 9398 6332 9404 6344
rect 9456 6372 9462 6384
rect 9493 6375 9551 6381
rect 9493 6372 9505 6375
rect 9456 6344 9505 6372
rect 9456 6332 9462 6344
rect 9493 6341 9505 6344
rect 9539 6341 9551 6375
rect 9493 6335 9551 6341
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 17144 6381 17172 6412
rect 17788 6412 17960 6440
rect 10597 6375 10655 6381
rect 10597 6372 10609 6375
rect 10560 6344 10609 6372
rect 10560 6332 10566 6344
rect 10597 6341 10609 6344
rect 10643 6341 10655 6375
rect 10597 6335 10655 6341
rect 17129 6375 17187 6381
rect 17129 6341 17141 6375
rect 17175 6341 17187 6375
rect 17129 6335 17187 6341
rect 1360 6276 2774 6304
rect 7009 6307 7067 6313
rect 1360 6264 1366 6276
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 8478 6304 8484 6316
rect 7055 6276 8484 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 9180 6276 9229 6304
rect 9180 6264 9186 6276
rect 9217 6273 9229 6276
rect 9263 6304 9275 6307
rect 15654 6304 15660 6316
rect 9263 6276 10364 6304
rect 15502 6276 15660 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5040 6208 5273 6236
rect 5040 6196 5046 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 5307 6208 6653 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 6641 6205 6653 6208
rect 6687 6236 6699 6239
rect 9140 6236 9168 6264
rect 6687 6208 9168 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 8389 6171 8447 6177
rect 8389 6168 8401 6171
rect 7708 6140 8401 6168
rect 7708 6128 7714 6140
rect 8389 6137 8401 6140
rect 8435 6168 8447 6171
rect 8757 6171 8815 6177
rect 8757 6168 8769 6171
rect 8435 6140 8769 6168
rect 8435 6137 8447 6140
rect 8389 6131 8447 6137
rect 8757 6137 8769 6140
rect 8803 6168 8815 6171
rect 9861 6171 9919 6177
rect 9861 6168 9873 6171
rect 8803 6140 9873 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 9861 6137 9873 6140
rect 9907 6137 9919 6171
rect 9861 6131 9919 6137
rect 10336 6112 10364 6276
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16632 6276 16681 6304
rect 16632 6264 16638 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16758 6264 16764 6316
rect 16816 6264 16822 6316
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17678 6304 17684 6316
rect 17267 6276 17684 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 17788 6304 17816 6412
rect 17954 6400 17960 6412
rect 18012 6440 18018 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 18012 6412 18061 6440
rect 18012 6400 18018 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18506 6400 18512 6452
rect 18564 6400 18570 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 20990 6440 20996 6452
rect 19208 6412 20996 6440
rect 19208 6400 19214 6412
rect 20990 6400 20996 6412
rect 21048 6440 21054 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 21048 6412 21373 6440
rect 21048 6400 21054 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 21361 6403 21419 6409
rect 21542 6400 21548 6452
rect 21600 6400 21606 6452
rect 21910 6440 21916 6452
rect 21744 6412 21916 6440
rect 17862 6332 17868 6384
rect 17920 6372 17926 6384
rect 19168 6372 19196 6400
rect 17920 6344 19196 6372
rect 17920 6332 17926 6344
rect 19886 6332 19892 6384
rect 19944 6332 19950 6384
rect 17788 6276 18644 6304
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13188 6208 14105 6236
rect 13188 6180 13216 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 14415 6208 15424 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 12437 6171 12495 6177
rect 12437 6168 12449 6171
rect 11716 6140 12449 6168
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10594 6100 10600 6112
rect 10376 6072 10600 6100
rect 10376 6060 10382 6072
rect 10594 6060 10600 6072
rect 10652 6100 10658 6112
rect 11716 6109 11744 6140
rect 12437 6137 12449 6140
rect 12483 6168 12495 6171
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12483 6140 12817 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 12805 6137 12817 6140
rect 12851 6168 12863 6171
rect 13170 6168 13176 6180
rect 12851 6140 13176 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 13630 6128 13636 6180
rect 13688 6128 13694 6180
rect 15396 6168 15424 6208
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 16114 6236 16120 6248
rect 15620 6208 16120 6236
rect 15620 6196 15626 6208
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16298 6196 16304 6248
rect 16356 6236 16362 6248
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 16356 6208 17141 6236
rect 16356 6196 16362 6208
rect 17129 6205 17141 6208
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6236 17555 6239
rect 18046 6236 18052 6248
rect 17543 6208 18052 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18616 6245 18644 6276
rect 20438 6264 20444 6316
rect 20496 6264 20502 6316
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6304 20683 6307
rect 20898 6304 20904 6316
rect 20671 6276 20904 6304
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21450 6304 21456 6316
rect 21223 6276 21456 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 18877 6239 18935 6245
rect 18877 6205 18889 6239
rect 18923 6236 18935 6239
rect 18966 6236 18972 6248
rect 18923 6208 18972 6236
rect 18923 6205 18935 6208
rect 18877 6199 18935 6205
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 21192 6236 21220 6267
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 21744 6313 21772 6412
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 23382 6400 23388 6452
rect 23440 6440 23446 6452
rect 24121 6443 24179 6449
rect 24121 6440 24133 6443
rect 23440 6412 24133 6440
rect 23440 6400 23446 6412
rect 24121 6409 24133 6412
rect 24167 6409 24179 6443
rect 24121 6403 24179 6409
rect 25130 6400 25136 6452
rect 25188 6400 25194 6452
rect 25498 6400 25504 6452
rect 25556 6440 25562 6452
rect 25685 6443 25743 6449
rect 25685 6440 25697 6443
rect 25556 6412 25697 6440
rect 25556 6400 25562 6412
rect 25685 6409 25697 6412
rect 25731 6440 25743 6443
rect 25774 6440 25780 6452
rect 25731 6412 25780 6440
rect 25731 6409 25743 6412
rect 25685 6403 25743 6409
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 25958 6400 25964 6452
rect 26016 6440 26022 6452
rect 27709 6443 27767 6449
rect 27709 6440 27721 6443
rect 26016 6412 27721 6440
rect 26016 6400 26022 6412
rect 27709 6409 27721 6412
rect 27755 6409 27767 6443
rect 27709 6403 27767 6409
rect 27798 6400 27804 6452
rect 27856 6400 27862 6452
rect 28169 6443 28227 6449
rect 28169 6409 28181 6443
rect 28215 6440 28227 6443
rect 28350 6440 28356 6452
rect 28215 6412 28356 6440
rect 28215 6409 28227 6412
rect 28169 6403 28227 6409
rect 28350 6400 28356 6412
rect 28408 6400 28414 6452
rect 28537 6443 28595 6449
rect 28537 6409 28549 6443
rect 28583 6409 28595 6443
rect 28537 6403 28595 6409
rect 22002 6332 22008 6384
rect 22060 6372 22066 6384
rect 22554 6372 22560 6384
rect 22060 6344 22560 6372
rect 22060 6332 22066 6344
rect 22388 6313 22416 6344
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 22649 6375 22707 6381
rect 22649 6341 22661 6375
rect 22695 6372 22707 6375
rect 22738 6372 22744 6384
rect 22695 6344 22744 6372
rect 22695 6341 22707 6344
rect 22649 6335 22707 6341
rect 22738 6332 22744 6344
rect 22796 6332 22802 6384
rect 25314 6332 25320 6384
rect 25372 6332 25378 6384
rect 25406 6332 25412 6384
rect 25464 6372 25470 6384
rect 25593 6375 25651 6381
rect 25593 6372 25605 6375
rect 25464 6344 25605 6372
rect 25464 6332 25470 6344
rect 25593 6341 25605 6344
rect 25639 6372 25651 6375
rect 26421 6375 26479 6381
rect 25639 6344 26372 6372
rect 25639 6341 25651 6344
rect 25593 6335 25651 6341
rect 21729 6307 21787 6313
rect 21729 6273 21741 6307
rect 21775 6273 21787 6307
rect 21729 6267 21787 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 24118 6304 24124 6316
rect 23782 6276 24124 6304
rect 22373 6267 22431 6273
rect 24118 6264 24124 6276
rect 24176 6304 24182 6316
rect 24670 6304 24676 6316
rect 24176 6276 24676 6304
rect 24176 6264 24182 6276
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 24762 6264 24768 6316
rect 24820 6304 24826 6316
rect 25501 6307 25559 6313
rect 25501 6304 25513 6307
rect 24820 6276 25513 6304
rect 24820 6264 24826 6276
rect 25501 6273 25513 6276
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 19392 6208 21220 6236
rect 19392 6196 19398 6208
rect 23106 6196 23112 6248
rect 23164 6236 23170 6248
rect 25866 6236 25872 6248
rect 23164 6208 25872 6236
rect 23164 6196 23170 6208
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 15396 6140 16497 6168
rect 16485 6137 16497 6140
rect 16531 6137 16543 6171
rect 16485 6131 16543 6137
rect 16758 6128 16764 6180
rect 16816 6168 16822 6180
rect 17313 6171 17371 6177
rect 17313 6168 17325 6171
rect 16816 6140 17325 6168
rect 16816 6128 16822 6140
rect 17313 6137 17325 6140
rect 17359 6168 17371 6171
rect 17359 6140 17540 6168
rect 17359 6137 17371 6140
rect 17313 6131 17371 6137
rect 17512 6112 17540 6140
rect 20346 6128 20352 6180
rect 20404 6168 20410 6180
rect 20404 6140 21128 6168
rect 20404 6128 20410 6140
rect 21100 6112 21128 6140
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 21910 6168 21916 6180
rect 21692 6140 21916 6168
rect 21692 6128 21698 6140
rect 21910 6128 21916 6140
rect 21968 6128 21974 6180
rect 24026 6168 24032 6180
rect 23676 6140 24032 6168
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10652 6072 11345 6100
rect 10652 6060 10658 6072
rect 11333 6069 11345 6072
rect 11379 6100 11391 6103
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11379 6072 11713 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11701 6063 11759 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11848 6072 12081 6100
rect 11848 6060 11854 6072
rect 12069 6069 12081 6072
rect 12115 6100 12127 6103
rect 12618 6100 12624 6112
rect 12115 6072 12624 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12618 6060 12624 6072
rect 12676 6100 12682 6112
rect 13265 6103 13323 6109
rect 13265 6100 13277 6103
rect 12676 6072 13277 6100
rect 12676 6060 12682 6072
rect 13265 6069 13277 6072
rect 13311 6069 13323 6103
rect 13265 6063 13323 6069
rect 14001 6103 14059 6109
rect 14001 6069 14013 6103
rect 14047 6100 14059 6103
rect 14090 6100 14096 6112
rect 14047 6072 14096 6100
rect 14047 6069 14059 6072
rect 14001 6063 14059 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 15841 6103 15899 6109
rect 15841 6069 15853 6103
rect 15887 6100 15899 6103
rect 16206 6100 16212 6112
rect 15887 6072 16212 6100
rect 15887 6069 15899 6072
rect 15841 6063 15899 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 16724 6072 17417 6100
rect 16724 6060 16730 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 17494 6060 17500 6112
rect 17552 6060 17558 6112
rect 19242 6060 19248 6112
rect 19300 6100 19306 6112
rect 20809 6103 20867 6109
rect 20809 6100 20821 6103
rect 19300 6072 20821 6100
rect 19300 6060 19306 6072
rect 20809 6069 20821 6072
rect 20855 6069 20867 6103
rect 20809 6063 20867 6069
rect 21082 6060 21088 6112
rect 21140 6060 21146 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 22186 6100 22192 6112
rect 21232 6072 22192 6100
rect 21232 6060 21238 6072
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 22830 6060 22836 6112
rect 22888 6100 22894 6112
rect 23676 6100 23704 6140
rect 24026 6128 24032 6140
rect 24084 6168 24090 6180
rect 26344 6168 26372 6344
rect 26421 6341 26433 6375
rect 26467 6372 26479 6375
rect 27614 6372 27620 6384
rect 26467 6344 27620 6372
rect 26467 6341 26479 6344
rect 26421 6335 26479 6341
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 27816 6372 27844 6400
rect 28552 6372 28580 6403
rect 28902 6400 28908 6452
rect 28960 6440 28966 6452
rect 28997 6443 29055 6449
rect 28997 6440 29009 6443
rect 28960 6412 29009 6440
rect 28960 6400 28966 6412
rect 28997 6409 29009 6412
rect 29043 6409 29055 6443
rect 30742 6440 30748 6452
rect 28997 6403 29055 6409
rect 29840 6412 30748 6440
rect 29840 6381 29868 6412
rect 30742 6400 30748 6412
rect 30800 6400 30806 6452
rect 30834 6400 30840 6452
rect 30892 6440 30898 6452
rect 31297 6443 31355 6449
rect 31297 6440 31309 6443
rect 30892 6412 31309 6440
rect 30892 6400 30898 6412
rect 31297 6409 31309 6412
rect 31343 6409 31355 6443
rect 34698 6440 34704 6452
rect 31297 6403 31355 6409
rect 31726 6412 34704 6440
rect 29825 6375 29883 6381
rect 27816 6344 28580 6372
rect 28828 6344 29132 6372
rect 26605 6307 26663 6313
rect 26605 6273 26617 6307
rect 26651 6304 26663 6307
rect 26694 6304 26700 6316
rect 26651 6276 26700 6304
rect 26651 6273 26663 6276
rect 26605 6267 26663 6273
rect 26694 6264 26700 6276
rect 26752 6264 26758 6316
rect 26881 6307 26939 6313
rect 26881 6273 26893 6307
rect 26927 6304 26939 6307
rect 27890 6304 27896 6316
rect 26927 6276 27896 6304
rect 26927 6273 26939 6276
rect 26881 6267 26939 6273
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28828 6304 28856 6344
rect 28077 6267 28135 6273
rect 28368 6276 28856 6304
rect 28905 6307 28963 6313
rect 26418 6196 26424 6248
rect 26476 6236 26482 6248
rect 26789 6239 26847 6245
rect 26789 6236 26801 6239
rect 26476 6208 26801 6236
rect 26476 6196 26482 6208
rect 26789 6205 26801 6208
rect 26835 6205 26847 6239
rect 26789 6199 26847 6205
rect 27062 6196 27068 6248
rect 27120 6196 27126 6248
rect 27706 6236 27712 6248
rect 27172 6208 27712 6236
rect 26510 6168 26516 6180
rect 24084 6140 26004 6168
rect 26344 6140 26516 6168
rect 24084 6128 24090 6140
rect 22888 6072 23704 6100
rect 22888 6060 22894 6072
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 24394 6100 24400 6112
rect 23808 6072 24400 6100
rect 23808 6060 23814 6072
rect 24394 6060 24400 6072
rect 24452 6060 24458 6112
rect 24489 6103 24547 6109
rect 24489 6069 24501 6103
rect 24535 6100 24547 6103
rect 24857 6103 24915 6109
rect 24857 6100 24869 6103
rect 24535 6072 24869 6100
rect 24535 6069 24547 6072
rect 24489 6063 24547 6069
rect 24857 6069 24869 6072
rect 24903 6100 24915 6103
rect 25222 6100 25228 6112
rect 24903 6072 25228 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 25222 6060 25228 6072
rect 25280 6060 25286 6112
rect 25866 6060 25872 6112
rect 25924 6060 25930 6112
rect 25976 6100 26004 6140
rect 26510 6128 26516 6140
rect 26568 6128 26574 6180
rect 26602 6128 26608 6180
rect 26660 6168 26666 6180
rect 26697 6171 26755 6177
rect 26697 6168 26709 6171
rect 26660 6140 26709 6168
rect 26660 6128 26666 6140
rect 26697 6137 26709 6140
rect 26743 6137 26755 6171
rect 26697 6131 26755 6137
rect 27172 6100 27200 6208
rect 27706 6196 27712 6208
rect 27764 6196 27770 6248
rect 27341 6171 27399 6177
rect 27341 6137 27353 6171
rect 27387 6137 27399 6171
rect 28092 6168 28120 6267
rect 28368 6245 28396 6276
rect 28905 6273 28917 6307
rect 28951 6273 28963 6307
rect 28905 6267 28963 6273
rect 28353 6239 28411 6245
rect 28353 6205 28365 6239
rect 28399 6205 28411 6239
rect 28353 6199 28411 6205
rect 28920 6168 28948 6267
rect 29104 6245 29132 6344
rect 29825 6341 29837 6375
rect 29871 6341 29883 6375
rect 29825 6335 29883 6341
rect 30098 6332 30104 6384
rect 30156 6372 30162 6384
rect 30282 6372 30288 6384
rect 30156 6344 30288 6372
rect 30156 6332 30162 6344
rect 30282 6332 30288 6344
rect 30340 6332 30346 6384
rect 31726 6372 31754 6412
rect 34698 6400 34704 6412
rect 34756 6400 34762 6452
rect 35250 6400 35256 6452
rect 35308 6440 35314 6452
rect 36081 6443 36139 6449
rect 36081 6440 36093 6443
rect 35308 6412 36093 6440
rect 35308 6400 35314 6412
rect 36081 6409 36093 6412
rect 36127 6409 36139 6443
rect 36081 6403 36139 6409
rect 36446 6400 36452 6452
rect 36504 6400 36510 6452
rect 36906 6400 36912 6452
rect 36964 6440 36970 6452
rect 36964 6412 38516 6440
rect 36964 6400 36970 6412
rect 31128 6344 31754 6372
rect 29270 6264 29276 6316
rect 29328 6304 29334 6316
rect 29549 6307 29607 6313
rect 29549 6304 29561 6307
rect 29328 6276 29561 6304
rect 29328 6264 29334 6276
rect 29549 6273 29561 6276
rect 29595 6273 29607 6307
rect 29549 6267 29607 6273
rect 29089 6239 29147 6245
rect 29089 6205 29101 6239
rect 29135 6236 29147 6239
rect 29454 6236 29460 6248
rect 29135 6208 29460 6236
rect 29135 6205 29147 6208
rect 29089 6199 29147 6205
rect 29454 6196 29460 6208
rect 29512 6196 29518 6248
rect 31128 6236 31156 6344
rect 32950 6332 32956 6384
rect 33008 6332 33014 6384
rect 33597 6375 33655 6381
rect 33597 6341 33609 6375
rect 33643 6372 33655 6375
rect 34146 6372 34152 6384
rect 33643 6344 34152 6372
rect 33643 6341 33655 6344
rect 33597 6335 33655 6341
rect 34146 6332 34152 6344
rect 34204 6332 34210 6384
rect 31570 6264 31576 6316
rect 31628 6304 31634 6316
rect 31665 6307 31723 6313
rect 31665 6304 31677 6307
rect 31628 6276 31677 6304
rect 31628 6264 31634 6276
rect 31665 6273 31677 6276
rect 31711 6273 31723 6307
rect 35986 6304 35992 6316
rect 35742 6276 35992 6304
rect 31665 6267 31723 6273
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 36357 6307 36415 6313
rect 36357 6273 36369 6307
rect 36403 6304 36415 6307
rect 36464 6304 36492 6400
rect 37274 6332 37280 6384
rect 37332 6372 37338 6384
rect 37369 6375 37427 6381
rect 37369 6372 37381 6375
rect 37332 6344 37381 6372
rect 37332 6332 37338 6344
rect 37369 6341 37381 6344
rect 37415 6341 37427 6375
rect 37369 6335 37427 6341
rect 38488 6316 38516 6412
rect 38838 6400 38844 6452
rect 38896 6400 38902 6452
rect 39114 6400 39120 6452
rect 39172 6440 39178 6452
rect 40681 6443 40739 6449
rect 40681 6440 40693 6443
rect 39172 6412 40693 6440
rect 39172 6400 39178 6412
rect 40681 6409 40693 6412
rect 40727 6440 40739 6443
rect 41233 6443 41291 6449
rect 41233 6440 41245 6443
rect 40727 6412 41245 6440
rect 40727 6409 40739 6412
rect 40681 6403 40739 6409
rect 41233 6409 41245 6412
rect 41279 6409 41291 6443
rect 41233 6403 41291 6409
rect 41506 6400 41512 6452
rect 41564 6440 41570 6452
rect 41785 6443 41843 6449
rect 41785 6440 41797 6443
rect 41564 6412 41797 6440
rect 41564 6400 41570 6412
rect 41785 6409 41797 6412
rect 41831 6409 41843 6443
rect 41785 6403 41843 6409
rect 42245 6443 42303 6449
rect 42245 6409 42257 6443
rect 42291 6440 42303 6443
rect 42794 6440 42800 6452
rect 42291 6412 42800 6440
rect 42291 6409 42303 6412
rect 42245 6403 42303 6409
rect 42794 6400 42800 6412
rect 42852 6400 42858 6452
rect 43070 6400 43076 6452
rect 43128 6400 43134 6452
rect 43346 6400 43352 6452
rect 43404 6440 43410 6452
rect 43625 6443 43683 6449
rect 43625 6440 43637 6443
rect 43404 6412 43637 6440
rect 43404 6400 43410 6412
rect 43625 6409 43637 6412
rect 43671 6440 43683 6443
rect 44361 6443 44419 6449
rect 44361 6440 44373 6443
rect 43671 6412 44373 6440
rect 43671 6409 43683 6412
rect 43625 6403 43683 6409
rect 44361 6409 44373 6412
rect 44407 6409 44419 6443
rect 44361 6403 44419 6409
rect 44726 6400 44732 6452
rect 44784 6400 44790 6452
rect 39206 6372 39212 6384
rect 38948 6344 39212 6372
rect 36403 6276 36492 6304
rect 36403 6273 36415 6276
rect 36357 6267 36415 6273
rect 36998 6264 37004 6316
rect 37056 6264 37062 6316
rect 38470 6264 38476 6316
rect 38528 6264 38534 6316
rect 38654 6264 38660 6316
rect 38712 6304 38718 6316
rect 38948 6313 38976 6344
rect 39206 6332 39212 6344
rect 39264 6332 39270 6384
rect 40494 6332 40500 6384
rect 40552 6372 40558 6384
rect 42153 6375 42211 6381
rect 42153 6372 42165 6375
rect 40552 6344 42165 6372
rect 40552 6332 40558 6344
rect 42153 6341 42165 6344
rect 42199 6341 42211 6375
rect 42153 6335 42211 6341
rect 38933 6307 38991 6313
rect 38712 6276 38884 6304
rect 38712 6264 38718 6276
rect 29656 6208 31156 6236
rect 31941 6239 31999 6245
rect 29656 6168 29684 6208
rect 31941 6205 31953 6239
rect 31987 6236 31999 6239
rect 33226 6236 33232 6248
rect 31987 6208 33232 6236
rect 31987 6205 31999 6208
rect 31941 6199 31999 6205
rect 33226 6196 33232 6208
rect 33284 6196 33290 6248
rect 34238 6196 34244 6248
rect 34296 6236 34302 6248
rect 34333 6239 34391 6245
rect 34333 6236 34345 6239
rect 34296 6208 34345 6236
rect 34296 6196 34302 6208
rect 34333 6205 34345 6208
rect 34379 6205 34391 6239
rect 34333 6199 34391 6205
rect 34606 6196 34612 6248
rect 34664 6196 34670 6248
rect 35250 6196 35256 6248
rect 35308 6236 35314 6248
rect 37090 6236 37096 6248
rect 35308 6208 37096 6236
rect 35308 6196 35314 6208
rect 37090 6196 37096 6208
rect 37148 6196 37154 6248
rect 38856 6236 38884 6276
rect 38933 6273 38945 6307
rect 38979 6273 38991 6307
rect 38933 6267 38991 6273
rect 40310 6264 40316 6316
rect 40368 6264 40374 6316
rect 40586 6264 40592 6316
rect 40644 6304 40650 6316
rect 41141 6307 41199 6313
rect 41141 6304 41153 6307
rect 40644 6276 41153 6304
rect 40644 6264 40650 6276
rect 41141 6273 41153 6276
rect 41187 6273 41199 6307
rect 42981 6307 43039 6313
rect 41141 6267 41199 6273
rect 41248 6276 42656 6304
rect 39209 6239 39267 6245
rect 39209 6236 39221 6239
rect 37200 6208 38792 6236
rect 38856 6208 39221 6236
rect 28092 6140 28856 6168
rect 28920 6140 29684 6168
rect 31220 6140 31754 6168
rect 27341 6131 27399 6137
rect 25976 6072 27200 6100
rect 27356 6100 27384 6131
rect 27430 6100 27436 6112
rect 27356 6072 27436 6100
rect 27430 6060 27436 6072
rect 27488 6060 27494 6112
rect 27525 6103 27583 6109
rect 27525 6069 27537 6103
rect 27571 6100 27583 6103
rect 28350 6100 28356 6112
rect 27571 6072 28356 6100
rect 27571 6069 27583 6072
rect 27525 6063 27583 6069
rect 28350 6060 28356 6072
rect 28408 6060 28414 6112
rect 28828 6100 28856 6140
rect 31220 6100 31248 6140
rect 28828 6072 31248 6100
rect 31726 6100 31754 6140
rect 33336 6140 34468 6168
rect 33336 6100 33364 6140
rect 31726 6072 33364 6100
rect 33410 6060 33416 6112
rect 33468 6060 33474 6112
rect 33686 6060 33692 6112
rect 33744 6100 33750 6112
rect 34146 6100 34152 6112
rect 33744 6072 34152 6100
rect 33744 6060 33750 6072
rect 34146 6060 34152 6072
rect 34204 6060 34210 6112
rect 34440 6100 34468 6140
rect 35802 6128 35808 6180
rect 35860 6168 35866 6180
rect 35986 6168 35992 6180
rect 35860 6140 35992 6168
rect 35860 6128 35866 6140
rect 35986 6128 35992 6140
rect 36044 6128 36050 6180
rect 37200 6168 37228 6208
rect 38654 6168 38660 6180
rect 36096 6140 37228 6168
rect 38396 6140 38660 6168
rect 36096 6100 36124 6140
rect 34440 6072 36124 6100
rect 36170 6060 36176 6112
rect 36228 6060 36234 6112
rect 36817 6103 36875 6109
rect 36817 6069 36829 6103
rect 36863 6100 36875 6103
rect 38396 6100 38424 6140
rect 38654 6128 38660 6140
rect 38712 6128 38718 6180
rect 36863 6072 38424 6100
rect 38764 6100 38792 6208
rect 39209 6205 39221 6208
rect 39255 6205 39267 6239
rect 39209 6199 39267 6205
rect 40678 6196 40684 6248
rect 40736 6236 40742 6248
rect 41248 6236 41276 6276
rect 40736 6208 41276 6236
rect 41325 6239 41383 6245
rect 40736 6196 40742 6208
rect 41325 6205 41337 6239
rect 41371 6205 41383 6239
rect 41325 6199 41383 6205
rect 40770 6128 40776 6180
rect 40828 6128 40834 6180
rect 39298 6100 39304 6112
rect 38764 6072 39304 6100
rect 36863 6069 36875 6072
rect 36817 6063 36875 6069
rect 39298 6060 39304 6072
rect 39356 6060 39362 6112
rect 39574 6060 39580 6112
rect 39632 6100 39638 6112
rect 41340 6100 41368 6199
rect 42058 6196 42064 6248
rect 42116 6236 42122 6248
rect 42337 6239 42395 6245
rect 42337 6236 42349 6239
rect 42116 6208 42349 6236
rect 42116 6196 42122 6208
rect 42337 6205 42349 6208
rect 42383 6205 42395 6239
rect 42337 6199 42395 6205
rect 39632 6072 41368 6100
rect 42352 6100 42380 6199
rect 42628 6177 42656 6276
rect 42981 6273 42993 6307
rect 43027 6304 43039 6307
rect 44358 6304 44364 6316
rect 43027 6276 44364 6304
rect 43027 6273 43039 6276
rect 42981 6267 43039 6273
rect 44358 6264 44364 6276
rect 44416 6264 44422 6316
rect 42702 6196 42708 6248
rect 42760 6236 42766 6248
rect 43257 6239 43315 6245
rect 43257 6236 43269 6239
rect 42760 6208 43269 6236
rect 42760 6196 42766 6208
rect 43257 6205 43269 6208
rect 43303 6236 43315 6239
rect 44174 6236 44180 6248
rect 43303 6208 44180 6236
rect 43303 6205 43315 6208
rect 43257 6199 43315 6205
rect 44174 6196 44180 6208
rect 44232 6196 44238 6248
rect 42613 6171 42671 6177
rect 42613 6137 42625 6171
rect 42659 6137 42671 6171
rect 42613 6131 42671 6137
rect 42978 6100 42984 6112
rect 42352 6072 42984 6100
rect 39632 6060 39638 6072
rect 42978 6060 42984 6072
rect 43036 6060 43042 6112
rect 43990 6060 43996 6112
rect 44048 6100 44054 6112
rect 45097 6103 45155 6109
rect 45097 6100 45109 6103
rect 44048 6072 45109 6100
rect 44048 6060 44054 6072
rect 45097 6069 45109 6072
rect 45143 6069 45155 6103
rect 45097 6063 45155 6069
rect 460 6010 45540 6032
rect 460 5958 3570 6010
rect 3622 5958 3634 6010
rect 3686 5958 3698 6010
rect 3750 5958 3762 6010
rect 3814 5958 3826 6010
rect 3878 5958 8570 6010
rect 8622 5958 8634 6010
rect 8686 5958 8698 6010
rect 8750 5958 8762 6010
rect 8814 5958 8826 6010
rect 8878 5958 13570 6010
rect 13622 5958 13634 6010
rect 13686 5958 13698 6010
rect 13750 5958 13762 6010
rect 13814 5958 13826 6010
rect 13878 5958 18570 6010
rect 18622 5958 18634 6010
rect 18686 5958 18698 6010
rect 18750 5958 18762 6010
rect 18814 5958 18826 6010
rect 18878 5958 23570 6010
rect 23622 5958 23634 6010
rect 23686 5958 23698 6010
rect 23750 5958 23762 6010
rect 23814 5958 23826 6010
rect 23878 5958 28570 6010
rect 28622 5958 28634 6010
rect 28686 5958 28698 6010
rect 28750 5958 28762 6010
rect 28814 5958 28826 6010
rect 28878 5958 33570 6010
rect 33622 5958 33634 6010
rect 33686 5958 33698 6010
rect 33750 5958 33762 6010
rect 33814 5958 33826 6010
rect 33878 5958 38570 6010
rect 38622 5958 38634 6010
rect 38686 5958 38698 6010
rect 38750 5958 38762 6010
rect 38814 5958 38826 6010
rect 38878 5958 43570 6010
rect 43622 5958 43634 6010
rect 43686 5958 43698 6010
rect 43750 5958 43762 6010
rect 43814 5958 43826 6010
rect 43878 5958 45540 6010
rect 460 5936 45540 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2498 5896 2504 5908
rect 1719 5868 2504 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2498 5856 2504 5868
rect 2556 5896 2562 5908
rect 3050 5896 3056 5908
rect 2556 5868 3056 5896
rect 2556 5856 2562 5868
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4304 5868 4537 5896
rect 4304 5856 4310 5868
rect 4525 5865 4537 5868
rect 4571 5896 4583 5899
rect 5442 5896 5448 5908
rect 4571 5868 5448 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7190 5896 7196 5908
rect 6779 5868 7196 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8352 5868 8769 5896
rect 8352 5856 8358 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 10502 5896 10508 5908
rect 9272 5868 10508 5896
rect 9272 5856 9278 5868
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 13170 5856 13176 5908
rect 13228 5856 13234 5908
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14424 5868 14841 5896
rect 14424 5856 14430 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 15194 5896 15200 5908
rect 14829 5859 14887 5865
rect 14936 5868 15200 5896
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 6365 5831 6423 5837
rect 6365 5828 6377 5831
rect 5776 5800 6377 5828
rect 5776 5788 5782 5800
rect 6365 5797 6377 5800
rect 6411 5828 6423 5831
rect 7668 5828 7696 5856
rect 6411 5800 7696 5828
rect 10689 5831 10747 5837
rect 6411 5797 6423 5800
rect 6365 5791 6423 5797
rect 10689 5797 10701 5831
rect 10735 5828 10747 5831
rect 12802 5828 12808 5840
rect 10735 5800 12808 5828
rect 10735 5797 10747 5800
rect 10689 5791 10747 5797
rect 12802 5788 12808 5800
rect 12860 5828 12866 5840
rect 13354 5828 13360 5840
rect 12860 5800 13360 5828
rect 12860 5788 12866 5800
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 14093 5831 14151 5837
rect 14093 5797 14105 5831
rect 14139 5828 14151 5831
rect 14458 5828 14464 5840
rect 14139 5800 14464 5828
rect 14139 5797 14151 5800
rect 14093 5791 14151 5797
rect 14458 5788 14464 5800
rect 14516 5788 14522 5840
rect 14936 5828 14964 5868
rect 15194 5856 15200 5868
rect 15252 5896 15258 5908
rect 16022 5896 16028 5908
rect 15252 5868 16028 5896
rect 15252 5856 15258 5868
rect 16022 5856 16028 5868
rect 16080 5896 16086 5908
rect 16942 5896 16948 5908
rect 16080 5868 16948 5896
rect 16080 5856 16086 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17126 5856 17132 5908
rect 17184 5896 17190 5908
rect 17678 5896 17684 5908
rect 17184 5868 17684 5896
rect 17184 5856 17190 5868
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 19794 5896 19800 5908
rect 17828 5868 19800 5896
rect 17828 5856 17834 5868
rect 19794 5856 19800 5868
rect 19852 5896 19858 5908
rect 20254 5896 20260 5908
rect 19852 5868 20260 5896
rect 19852 5856 19858 5868
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20496 5868 21281 5896
rect 20496 5856 20502 5868
rect 21269 5865 21281 5868
rect 21315 5896 21327 5899
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 21315 5868 21373 5896
rect 21315 5865 21327 5868
rect 21269 5859 21327 5865
rect 21361 5865 21373 5868
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 21508 5868 23980 5896
rect 21508 5856 21514 5868
rect 17865 5831 17923 5837
rect 17865 5828 17877 5831
rect 14568 5800 14964 5828
rect 16316 5800 17877 5828
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5123 5732 5825 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5813 5729 5825 5732
rect 5859 5760 5871 5763
rect 7282 5760 7288 5772
rect 5859 5732 7288 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 4982 5692 4988 5704
rect 3007 5664 4988 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 14568 5701 14596 5800
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15562 5760 15568 5772
rect 14691 5732 14964 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 12897 5695 12955 5701
rect 10376 5664 11100 5692
rect 10376 5652 10382 5664
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 9585 5627 9643 5633
rect 7515 5596 8156 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 1305 5559 1363 5565
rect 1305 5525 1317 5559
rect 1351 5556 1363 5559
rect 2590 5556 2596 5568
rect 1351 5528 2596 5556
rect 1351 5525 1363 5528
rect 1305 5519 1363 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3329 5559 3387 5565
rect 3329 5556 3341 5559
rect 2924 5528 3341 5556
rect 2924 5516 2930 5528
rect 3329 5525 3341 5528
rect 3375 5525 3387 5559
rect 3329 5519 3387 5525
rect 3970 5516 3976 5568
rect 4028 5516 4034 5568
rect 5442 5516 5448 5568
rect 5500 5516 5506 5568
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5556 7159 5559
rect 7742 5556 7748 5568
rect 7147 5528 7748 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8128 5565 8156 5596
rect 9585 5593 9597 5627
rect 9631 5624 9643 5627
rect 9631 5596 10456 5624
rect 9631 5593 9643 5596
rect 9585 5587 9643 5593
rect 10428 5568 10456 5596
rect 8113 5559 8171 5565
rect 8113 5525 8125 5559
rect 8159 5556 8171 5559
rect 9122 5556 9128 5568
rect 8159 5528 9128 5556
rect 8159 5525 8171 5528
rect 8113 5519 8171 5525
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9950 5516 9956 5568
rect 10008 5516 10014 5568
rect 10410 5516 10416 5568
rect 10468 5516 10474 5568
rect 11072 5565 11100 5664
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 14553 5695 14611 5701
rect 12943 5664 14412 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 11103 5528 11437 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11425 5525 11437 5528
rect 11471 5556 11483 5559
rect 11514 5556 11520 5568
rect 11471 5528 11520 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11848 5528 12173 5556
rect 11848 5516 11854 5528
rect 12161 5525 12173 5528
rect 12207 5556 12219 5559
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 12207 5528 12541 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 12529 5525 12541 5528
rect 12575 5556 12587 5559
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 12575 5528 13737 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 13725 5525 13737 5528
rect 13771 5556 13783 5559
rect 14182 5556 14188 5568
rect 13771 5528 14188 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 14384 5556 14412 5664
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 14553 5655 14611 5661
rect 14660 5664 14749 5692
rect 14660 5636 14688 5664
rect 14737 5661 14749 5664
rect 14783 5661 14795 5695
rect 14936 5692 14964 5732
rect 15396 5732 15568 5760
rect 15105 5705 15163 5711
rect 15105 5694 15117 5705
rect 15104 5692 15117 5694
rect 14936 5671 15117 5692
rect 15151 5671 15163 5705
rect 15396 5701 15424 5732
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 14936 5665 15163 5671
rect 15381 5695 15439 5701
rect 14936 5664 15132 5665
rect 14737 5655 14795 5661
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 14458 5584 14464 5636
rect 14516 5584 14522 5636
rect 14642 5584 14648 5636
rect 14700 5584 14706 5636
rect 14829 5627 14887 5633
rect 14829 5593 14841 5627
rect 14875 5624 14887 5627
rect 15102 5624 15108 5636
rect 14875 5596 15108 5624
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15194 5584 15200 5636
rect 15252 5633 15258 5636
rect 15252 5627 15273 5633
rect 15261 5593 15273 5627
rect 15252 5587 15273 5593
rect 15657 5627 15715 5633
rect 15657 5593 15669 5627
rect 15703 5593 15715 5627
rect 15657 5587 15715 5593
rect 15252 5584 15258 5587
rect 14918 5556 14924 5568
rect 14384 5528 14924 5556
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15013 5559 15071 5565
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 15059 5528 15577 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15672 5556 15700 5587
rect 15838 5584 15844 5636
rect 15896 5584 15902 5636
rect 16316 5556 16344 5800
rect 16758 5760 16764 5772
rect 16408 5732 16764 5760
rect 16408 5701 16436 5732
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5661 16635 5695
rect 16577 5655 16635 5661
rect 16592 5568 16620 5655
rect 16666 5652 16672 5704
rect 16724 5652 16730 5704
rect 16869 5701 16897 5800
rect 17865 5797 17877 5800
rect 17911 5797 17923 5831
rect 17865 5791 17923 5797
rect 17954 5788 17960 5840
rect 18012 5788 18018 5840
rect 18601 5831 18659 5837
rect 18601 5797 18613 5831
rect 18647 5828 18659 5831
rect 18647 5800 19380 5828
rect 18647 5797 18659 5800
rect 18601 5791 18659 5797
rect 18414 5760 18420 5772
rect 17052 5732 17448 5760
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 16761 5627 16819 5633
rect 16761 5593 16773 5627
rect 16807 5624 16819 5627
rect 17052 5624 17080 5732
rect 17420 5701 17448 5732
rect 17604 5732 18420 5760
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 16807 5596 17080 5624
rect 17144 5624 17172 5655
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 17604 5692 17632 5732
rect 18414 5720 18420 5732
rect 18472 5720 18478 5772
rect 19242 5760 19248 5772
rect 18800 5732 19248 5760
rect 17552 5664 17632 5692
rect 17681 5695 17739 5701
rect 17552 5652 17558 5664
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 18046 5692 18052 5704
rect 17727 5664 18052 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18800 5701 18828 5732
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 19352 5704 19380 5800
rect 20824 5800 23888 5828
rect 19518 5720 19524 5772
rect 19576 5720 19582 5772
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 20162 5760 20168 5772
rect 19843 5732 20168 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 20254 5720 20260 5772
rect 20312 5760 20318 5772
rect 20824 5760 20852 5800
rect 20312 5732 20852 5760
rect 20312 5720 20318 5732
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 21048 5732 21465 5760
rect 21048 5720 21054 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 21634 5720 21640 5772
rect 21692 5760 21698 5772
rect 23014 5760 23020 5772
rect 21692 5732 23020 5760
rect 21692 5720 21698 5732
rect 23014 5720 23020 5732
rect 23072 5720 23078 5772
rect 23860 5769 23888 5800
rect 23845 5763 23903 5769
rect 23845 5729 23857 5763
rect 23891 5729 23903 5763
rect 23845 5723 23903 5729
rect 23952 5760 23980 5868
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 24578 5856 24584 5908
rect 24636 5856 24642 5908
rect 25130 5856 25136 5908
rect 25188 5856 25194 5908
rect 25240 5868 26740 5896
rect 24596 5760 24624 5856
rect 25240 5828 25268 5868
rect 24964 5800 25268 5828
rect 24964 5760 24992 5800
rect 23952 5732 24624 5760
rect 24872 5732 24992 5760
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18785 5695 18843 5701
rect 18279 5664 18736 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18708 5636 18736 5664
rect 18785 5661 18797 5695
rect 18831 5661 18843 5695
rect 18785 5655 18843 5661
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 17862 5624 17868 5636
rect 17144 5596 17868 5624
rect 16807 5593 16819 5596
rect 16761 5587 16819 5593
rect 17862 5584 17868 5596
rect 17920 5624 17926 5636
rect 17957 5627 18015 5633
rect 17957 5624 17969 5627
rect 17920 5596 17969 5624
rect 17920 5584 17926 5596
rect 17957 5593 17969 5596
rect 18003 5593 18015 5627
rect 18322 5624 18328 5636
rect 17957 5587 18015 5593
rect 18064 5596 18328 5624
rect 16390 5556 16396 5568
rect 15672 5528 16396 5556
rect 15565 5519 15623 5525
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 16482 5516 16488 5568
rect 16540 5516 16546 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16850 5556 16856 5568
rect 16632 5528 16856 5556
rect 16632 5516 16638 5528
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 16942 5516 16948 5568
rect 17000 5516 17006 5568
rect 17313 5559 17371 5565
rect 17313 5525 17325 5559
rect 17359 5556 17371 5559
rect 18064 5556 18092 5596
rect 18322 5584 18328 5596
rect 18380 5624 18386 5636
rect 18380 5596 18460 5624
rect 18380 5584 18386 5596
rect 17359 5528 18092 5556
rect 17359 5525 17371 5528
rect 17313 5519 17371 5525
rect 18138 5516 18144 5568
rect 18196 5516 18202 5568
rect 18432 5556 18460 5596
rect 18506 5584 18512 5636
rect 18564 5624 18570 5636
rect 18601 5627 18659 5633
rect 18601 5624 18613 5627
rect 18564 5596 18613 5624
rect 18564 5584 18570 5596
rect 18601 5593 18613 5596
rect 18647 5593 18659 5627
rect 18601 5587 18659 5593
rect 18690 5584 18696 5636
rect 18748 5584 18754 5636
rect 18892 5624 18920 5655
rect 18966 5652 18972 5704
rect 19024 5652 19030 5704
rect 19150 5652 19156 5704
rect 19208 5652 19214 5704
rect 19334 5652 19340 5704
rect 19392 5652 19398 5704
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 19475 5664 19564 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19536 5624 19564 5664
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 21140 5664 21373 5692
rect 21140 5652 21146 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21818 5692 21824 5704
rect 21361 5655 21419 5661
rect 21468 5664 21824 5692
rect 21468 5624 21496 5664
rect 21818 5652 21824 5664
rect 21876 5692 21882 5704
rect 22370 5692 22376 5704
rect 21876 5664 22376 5692
rect 21876 5652 21882 5664
rect 22370 5652 22376 5664
rect 22428 5652 22434 5704
rect 22646 5652 22652 5704
rect 22704 5652 22710 5704
rect 22830 5652 22836 5704
rect 22888 5692 22894 5704
rect 23032 5692 23060 5720
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22888 5664 22968 5692
rect 23032 5664 23213 5692
rect 22888 5652 22894 5664
rect 18892 5596 19472 5624
rect 19536 5596 19748 5624
rect 21022 5596 21496 5624
rect 19337 5559 19395 5565
rect 19337 5556 19349 5559
rect 18432 5528 19349 5556
rect 19337 5525 19349 5528
rect 19383 5525 19395 5559
rect 19444 5556 19472 5596
rect 19720 5568 19748 5596
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 22940 5624 22968 5664
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 23201 5655 23259 5661
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23017 5627 23075 5633
rect 23017 5624 23029 5627
rect 21600 5596 22600 5624
rect 22940 5596 23029 5624
rect 21600 5584 21606 5596
rect 19518 5556 19524 5568
rect 19444 5528 19524 5556
rect 19337 5519 19395 5525
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 19702 5516 19708 5568
rect 19760 5516 19766 5568
rect 19794 5516 19800 5568
rect 19852 5556 19858 5568
rect 21729 5559 21787 5565
rect 21729 5556 21741 5559
rect 19852 5528 21741 5556
rect 19852 5516 19858 5528
rect 21729 5525 21741 5528
rect 21775 5525 21787 5559
rect 21729 5519 21787 5525
rect 22370 5516 22376 5568
rect 22428 5556 22434 5568
rect 22465 5559 22523 5565
rect 22465 5556 22477 5559
rect 22428 5528 22477 5556
rect 22428 5516 22434 5528
rect 22465 5525 22477 5528
rect 22511 5525 22523 5559
rect 22572 5556 22600 5596
rect 23017 5593 23029 5596
rect 23063 5593 23075 5627
rect 23860 5624 23888 5723
rect 23952 5701 23980 5732
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5661 23995 5695
rect 23937 5655 23995 5661
rect 24302 5652 24308 5704
rect 24360 5652 24366 5704
rect 24394 5652 24400 5704
rect 24452 5692 24458 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24452 5664 24685 5692
rect 24452 5652 24458 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 24872 5624 24900 5732
rect 25222 5720 25228 5772
rect 25280 5760 25286 5772
rect 25409 5763 25467 5769
rect 25409 5760 25421 5763
rect 25280 5732 25421 5760
rect 25280 5720 25286 5732
rect 25409 5729 25421 5732
rect 25455 5760 25467 5763
rect 26050 5760 26056 5772
rect 25455 5732 26056 5760
rect 25455 5729 25467 5732
rect 25409 5723 25467 5729
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 26712 5760 26740 5868
rect 27062 5856 27068 5908
rect 27120 5896 27126 5908
rect 27157 5899 27215 5905
rect 27157 5896 27169 5899
rect 27120 5868 27169 5896
rect 27120 5856 27126 5868
rect 27157 5865 27169 5868
rect 27203 5865 27215 5899
rect 27157 5859 27215 5865
rect 28074 5856 28080 5908
rect 28132 5856 28138 5908
rect 28902 5856 28908 5908
rect 28960 5896 28966 5908
rect 28960 5868 30236 5896
rect 28960 5856 28966 5868
rect 27982 5788 27988 5840
rect 28040 5828 28046 5840
rect 28040 5800 29040 5828
rect 28040 5788 28046 5800
rect 26712 5732 28120 5760
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 23860 5596 24900 5624
rect 24964 5624 24992 5655
rect 25038 5652 25044 5704
rect 25096 5692 25102 5704
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 25096 5664 25145 5692
rect 25096 5652 25102 5664
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 26786 5652 26792 5704
rect 26844 5652 26850 5704
rect 27062 5652 27068 5704
rect 27120 5692 27126 5704
rect 27341 5695 27399 5701
rect 27341 5692 27353 5695
rect 27120 5664 27353 5692
rect 27120 5652 27126 5664
rect 27341 5661 27353 5664
rect 27387 5661 27399 5695
rect 27341 5655 27399 5661
rect 27430 5652 27436 5704
rect 27488 5692 27494 5704
rect 27617 5695 27675 5701
rect 27617 5692 27629 5695
rect 27488 5664 27629 5692
rect 27488 5652 27494 5664
rect 27617 5661 27629 5664
rect 27663 5661 27675 5695
rect 27617 5655 27675 5661
rect 25590 5624 25596 5636
rect 24964 5596 25596 5624
rect 23017 5587 23075 5593
rect 25590 5584 25596 5596
rect 25648 5584 25654 5636
rect 25685 5627 25743 5633
rect 25685 5593 25697 5627
rect 25731 5593 25743 5627
rect 25685 5587 25743 5593
rect 22922 5556 22928 5568
rect 22572 5528 22928 5556
rect 22465 5519 22523 5525
rect 22922 5516 22928 5528
rect 22980 5556 22986 5568
rect 23293 5559 23351 5565
rect 23293 5556 23305 5559
rect 22980 5528 23305 5556
rect 22980 5516 22986 5528
rect 23293 5525 23305 5528
rect 23339 5525 23351 5559
rect 23293 5519 23351 5525
rect 23569 5559 23627 5565
rect 23569 5525 23581 5559
rect 23615 5556 23627 5559
rect 24394 5556 24400 5568
rect 23615 5528 24400 5556
rect 23615 5525 23627 5528
rect 23569 5519 23627 5525
rect 24394 5516 24400 5528
rect 24452 5516 24458 5568
rect 24489 5559 24547 5565
rect 24489 5525 24501 5559
rect 24535 5556 24547 5559
rect 24854 5556 24860 5568
rect 24535 5528 24860 5556
rect 24535 5525 24547 5528
rect 24489 5519 24547 5525
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 25317 5559 25375 5565
rect 25317 5525 25329 5559
rect 25363 5556 25375 5559
rect 25406 5556 25412 5568
rect 25363 5528 25412 5556
rect 25363 5525 25375 5528
rect 25317 5519 25375 5525
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 25700 5556 25728 5587
rect 27246 5584 27252 5636
rect 27304 5624 27310 5636
rect 27525 5627 27583 5633
rect 27525 5624 27537 5627
rect 27304 5596 27537 5624
rect 27304 5584 27310 5596
rect 27525 5593 27537 5596
rect 27571 5593 27583 5627
rect 27525 5587 27583 5593
rect 27632 5556 27660 5655
rect 27893 5627 27951 5633
rect 27893 5593 27905 5627
rect 27939 5624 27951 5627
rect 27982 5624 27988 5636
rect 27939 5596 27988 5624
rect 27939 5593 27951 5596
rect 27893 5587 27951 5593
rect 27982 5584 27988 5596
rect 28040 5584 28046 5636
rect 28092 5633 28120 5732
rect 28902 5720 28908 5772
rect 28960 5720 28966 5772
rect 29012 5760 29040 5800
rect 29270 5760 29276 5772
rect 29012 5732 29276 5760
rect 29270 5720 29276 5732
rect 29328 5720 29334 5772
rect 30208 5760 30236 5868
rect 30558 5856 30564 5908
rect 30616 5896 30622 5908
rect 30616 5868 30880 5896
rect 30616 5856 30622 5868
rect 30374 5788 30380 5840
rect 30432 5828 30438 5840
rect 30653 5831 30711 5837
rect 30653 5828 30665 5831
rect 30432 5800 30665 5828
rect 30432 5788 30438 5800
rect 30653 5797 30665 5800
rect 30699 5797 30711 5831
rect 30653 5791 30711 5797
rect 30745 5763 30803 5769
rect 30745 5760 30757 5763
rect 30208 5732 30757 5760
rect 30745 5729 30757 5732
rect 30791 5729 30803 5763
rect 30852 5760 30880 5868
rect 31018 5856 31024 5908
rect 31076 5896 31082 5908
rect 31754 5896 31760 5908
rect 31076 5868 31760 5896
rect 31076 5856 31082 5868
rect 31754 5856 31760 5868
rect 31812 5896 31818 5908
rect 32493 5899 32551 5905
rect 32493 5896 32505 5899
rect 31812 5868 32505 5896
rect 31812 5856 31818 5868
rect 32493 5865 32505 5868
rect 32539 5865 32551 5899
rect 32493 5859 32551 5865
rect 33226 5856 33232 5908
rect 33284 5856 33290 5908
rect 34606 5856 34612 5908
rect 34664 5896 34670 5908
rect 34885 5899 34943 5905
rect 34885 5896 34897 5899
rect 34664 5868 34897 5896
rect 34664 5856 34670 5868
rect 34885 5865 34897 5868
rect 34931 5865 34943 5899
rect 35526 5896 35532 5908
rect 34885 5859 34943 5865
rect 35084 5868 35532 5896
rect 32416 5800 34192 5828
rect 32416 5772 32444 5800
rect 31021 5763 31079 5769
rect 31021 5760 31033 5763
rect 30852 5732 31033 5760
rect 30745 5723 30803 5729
rect 31021 5729 31033 5732
rect 31067 5729 31079 5763
rect 31021 5723 31079 5729
rect 32398 5720 32404 5772
rect 32456 5720 32462 5772
rect 32674 5720 32680 5772
rect 32732 5760 32738 5772
rect 33045 5763 33103 5769
rect 33045 5760 33057 5763
rect 32732 5732 33057 5760
rect 32732 5720 32738 5732
rect 33045 5729 33057 5732
rect 33091 5729 33103 5763
rect 33045 5723 33103 5729
rect 33134 5720 33140 5772
rect 33192 5720 33198 5772
rect 33428 5769 33456 5800
rect 33409 5763 33467 5769
rect 33409 5729 33421 5763
rect 33455 5729 33467 5763
rect 33409 5723 33467 5729
rect 33962 5720 33968 5772
rect 34020 5720 34026 5772
rect 34054 5720 34060 5772
rect 34112 5720 34118 5772
rect 30282 5652 30288 5704
rect 30340 5652 30346 5704
rect 32416 5692 32444 5720
rect 32769 5695 32827 5701
rect 32769 5692 32781 5695
rect 32416 5664 32781 5692
rect 32769 5661 32781 5664
rect 32815 5661 32827 5695
rect 32769 5655 32827 5661
rect 32861 5695 32919 5701
rect 32861 5661 32873 5695
rect 32907 5661 32919 5695
rect 32861 5655 32919 5661
rect 32953 5695 33011 5701
rect 32953 5661 32965 5695
rect 32999 5692 33011 5695
rect 33152 5692 33180 5720
rect 32999 5664 33180 5692
rect 32999 5661 33011 5664
rect 32953 5655 33011 5661
rect 28092 5627 28156 5633
rect 28092 5596 28110 5627
rect 28098 5593 28110 5596
rect 28144 5624 28156 5627
rect 28537 5627 28595 5633
rect 28144 5596 28488 5624
rect 28144 5593 28156 5596
rect 28098 5587 28156 5593
rect 28460 5568 28488 5596
rect 28537 5593 28549 5627
rect 28583 5624 28595 5627
rect 29086 5624 29092 5636
rect 28583 5596 29092 5624
rect 28583 5593 28595 5596
rect 28537 5587 28595 5593
rect 29086 5584 29092 5596
rect 29144 5584 29150 5636
rect 29178 5584 29184 5636
rect 29236 5584 29242 5636
rect 25700 5528 27660 5556
rect 28258 5516 28264 5568
rect 28316 5516 28322 5568
rect 28442 5516 28448 5568
rect 28500 5556 28506 5568
rect 28629 5559 28687 5565
rect 28629 5556 28641 5559
rect 28500 5528 28641 5556
rect 28500 5516 28506 5528
rect 28629 5525 28641 5528
rect 28675 5525 28687 5559
rect 30300 5556 30328 5652
rect 32674 5624 32680 5636
rect 32246 5596 32680 5624
rect 32324 5556 32352 5596
rect 32674 5584 32680 5596
rect 32732 5584 32738 5636
rect 32876 5624 32904 5655
rect 32784 5596 32904 5624
rect 33152 5624 33180 5664
rect 33318 5652 33324 5704
rect 33376 5692 33382 5704
rect 33494 5695 33552 5701
rect 33494 5692 33506 5695
rect 33376 5664 33506 5692
rect 33376 5652 33382 5664
rect 33494 5661 33506 5664
rect 33540 5661 33552 5695
rect 33597 5695 33655 5701
rect 33597 5692 33609 5695
rect 33494 5655 33552 5661
rect 33594 5661 33609 5692
rect 33643 5661 33655 5695
rect 33594 5655 33655 5661
rect 33689 5695 33747 5701
rect 33689 5661 33701 5695
rect 33735 5692 33747 5695
rect 33980 5692 34008 5720
rect 33735 5664 34008 5692
rect 34164 5692 34192 5800
rect 34514 5720 34520 5772
rect 34572 5720 34578 5772
rect 34241 5695 34299 5701
rect 34241 5692 34253 5695
rect 34164 5664 34253 5692
rect 33735 5661 33747 5664
rect 33689 5655 33747 5661
rect 34241 5661 34253 5664
rect 34287 5661 34299 5695
rect 34241 5655 34299 5661
rect 33594 5624 33622 5655
rect 34330 5652 34336 5704
rect 34388 5652 34394 5704
rect 34425 5695 34483 5701
rect 34425 5661 34437 5695
rect 34471 5661 34483 5695
rect 34425 5655 34483 5661
rect 34440 5624 34468 5655
rect 34698 5652 34704 5704
rect 34756 5652 34762 5704
rect 35084 5701 35112 5868
rect 35526 5856 35532 5868
rect 35584 5856 35590 5908
rect 36814 5856 36820 5908
rect 36872 5896 36878 5908
rect 37001 5899 37059 5905
rect 37001 5896 37013 5899
rect 36872 5868 37013 5896
rect 36872 5856 36878 5868
rect 37001 5865 37013 5868
rect 37047 5865 37059 5899
rect 37001 5859 37059 5865
rect 37090 5856 37096 5908
rect 37148 5896 37154 5908
rect 37274 5896 37280 5908
rect 37148 5868 37280 5896
rect 37148 5856 37154 5868
rect 37274 5856 37280 5868
rect 37332 5856 37338 5908
rect 38102 5856 38108 5908
rect 38160 5856 38166 5908
rect 38470 5856 38476 5908
rect 38528 5896 38534 5908
rect 39022 5896 39028 5908
rect 38528 5868 39028 5896
rect 38528 5856 38534 5868
rect 39022 5856 39028 5868
rect 39080 5856 39086 5908
rect 42797 5899 42855 5905
rect 42797 5865 42809 5899
rect 42843 5896 42855 5899
rect 43070 5896 43076 5908
rect 42843 5868 43076 5896
rect 42843 5865 42855 5868
rect 42797 5859 42855 5865
rect 43070 5856 43076 5868
rect 43128 5856 43134 5908
rect 43346 5856 43352 5908
rect 43404 5896 43410 5908
rect 43441 5899 43499 5905
rect 43441 5896 43453 5899
rect 43404 5868 43453 5896
rect 43404 5856 43410 5868
rect 43441 5865 43453 5868
rect 43487 5896 43499 5899
rect 43809 5899 43867 5905
rect 43809 5896 43821 5899
rect 43487 5868 43821 5896
rect 43487 5865 43499 5868
rect 43441 5859 43499 5865
rect 43809 5865 43821 5868
rect 43855 5896 43867 5899
rect 44545 5899 44603 5905
rect 44545 5896 44557 5899
rect 43855 5868 44557 5896
rect 43855 5865 43867 5868
rect 43809 5859 43867 5865
rect 44545 5865 44557 5868
rect 44591 5896 44603 5899
rect 44910 5896 44916 5908
rect 44591 5868 44916 5896
rect 44591 5865 44603 5868
rect 44545 5859 44603 5865
rect 44910 5856 44916 5868
rect 44968 5856 44974 5908
rect 40954 5788 40960 5840
rect 41012 5788 41018 5840
rect 35529 5763 35587 5769
rect 35529 5729 35541 5763
rect 35575 5760 35587 5763
rect 36170 5760 36176 5772
rect 35575 5732 36176 5760
rect 35575 5729 35587 5732
rect 35529 5723 35587 5729
rect 36170 5720 36176 5732
rect 36228 5720 36234 5772
rect 36814 5720 36820 5772
rect 36872 5760 36878 5772
rect 37737 5763 37795 5769
rect 36872 5732 37504 5760
rect 36872 5720 36878 5732
rect 37200 5704 37228 5732
rect 35069 5695 35127 5701
rect 35069 5661 35081 5695
rect 35115 5661 35127 5695
rect 35069 5655 35127 5661
rect 35250 5652 35256 5704
rect 35308 5652 35314 5704
rect 36630 5652 36636 5704
rect 36688 5692 36694 5704
rect 36906 5692 36912 5704
rect 36688 5664 36912 5692
rect 36688 5652 36694 5664
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 37182 5652 37188 5704
rect 37240 5652 37246 5704
rect 37476 5701 37504 5732
rect 37737 5729 37749 5763
rect 37783 5729 37795 5763
rect 37737 5723 37795 5729
rect 37461 5695 37519 5701
rect 37461 5661 37473 5695
rect 37507 5661 37519 5695
rect 37752 5692 37780 5723
rect 37918 5720 37924 5772
rect 37976 5760 37982 5772
rect 38657 5763 38715 5769
rect 38657 5760 38669 5763
rect 37976 5732 38669 5760
rect 37976 5720 37982 5732
rect 38657 5729 38669 5732
rect 38703 5729 38715 5763
rect 39850 5760 39856 5772
rect 38657 5723 38715 5729
rect 39132 5732 39856 5760
rect 38194 5692 38200 5704
rect 37752 5664 38200 5692
rect 37461 5655 37519 5661
rect 38194 5652 38200 5664
rect 38252 5692 38258 5704
rect 39132 5692 39160 5732
rect 39850 5720 39856 5732
rect 39908 5720 39914 5772
rect 40972 5760 41000 5788
rect 41325 5763 41383 5769
rect 41325 5760 41337 5763
rect 40972 5732 41337 5760
rect 41325 5729 41337 5732
rect 41371 5729 41383 5763
rect 42518 5760 42524 5772
rect 41325 5723 41383 5729
rect 42444 5732 42524 5760
rect 38252 5664 39160 5692
rect 39209 5695 39267 5701
rect 38252 5652 38258 5664
rect 39209 5661 39221 5695
rect 39255 5661 39267 5695
rect 40862 5692 40868 5704
rect 39209 5655 39267 5661
rect 40788 5664 40868 5692
rect 33152 5596 34468 5624
rect 34716 5624 34744 5652
rect 35268 5624 35296 5652
rect 34716 5596 35296 5624
rect 32784 5568 32812 5596
rect 36814 5584 36820 5636
rect 36872 5624 36878 5636
rect 37553 5627 37611 5633
rect 37553 5624 37565 5627
rect 36872 5596 37565 5624
rect 36872 5584 36878 5596
rect 37553 5593 37565 5596
rect 37599 5593 37611 5627
rect 39114 5624 39120 5636
rect 37553 5587 37611 5593
rect 37660 5596 39120 5624
rect 30300 5528 32352 5556
rect 28629 5519 28687 5525
rect 32582 5516 32588 5568
rect 32640 5516 32646 5568
rect 32766 5516 32772 5568
rect 32824 5516 32830 5568
rect 32858 5516 32864 5568
rect 32916 5556 32922 5568
rect 36446 5556 36452 5568
rect 32916 5528 36452 5556
rect 32916 5516 32922 5528
rect 36446 5516 36452 5528
rect 36504 5516 36510 5568
rect 37090 5516 37096 5568
rect 37148 5516 37154 5568
rect 37274 5516 37280 5568
rect 37332 5556 37338 5568
rect 37660 5556 37688 5596
rect 39114 5584 39120 5596
rect 39172 5624 39178 5636
rect 39224 5624 39252 5655
rect 39172 5596 39252 5624
rect 39172 5584 39178 5596
rect 37332 5528 37688 5556
rect 37332 5516 37338 5528
rect 38470 5516 38476 5568
rect 38528 5516 38534 5568
rect 38565 5559 38623 5565
rect 38565 5525 38577 5559
rect 38611 5556 38623 5559
rect 38930 5556 38936 5568
rect 38611 5528 38936 5556
rect 38611 5525 38623 5528
rect 38565 5519 38623 5525
rect 38930 5516 38936 5528
rect 38988 5516 38994 5568
rect 39224 5556 39252 5596
rect 39482 5584 39488 5636
rect 39540 5584 39546 5636
rect 40218 5584 40224 5636
rect 40276 5584 40282 5636
rect 40788 5556 40816 5664
rect 40862 5652 40868 5664
rect 40920 5692 40926 5704
rect 41049 5695 41107 5701
rect 41049 5692 41061 5695
rect 40920 5664 41061 5692
rect 40920 5652 40926 5664
rect 41049 5661 41061 5664
rect 41095 5661 41107 5695
rect 42444 5678 42472 5732
rect 42518 5720 42524 5732
rect 42576 5720 42582 5772
rect 41049 5655 41107 5661
rect 39224 5528 40816 5556
rect 40862 5516 40868 5568
rect 40920 5556 40926 5568
rect 40957 5559 41015 5565
rect 40957 5556 40969 5559
rect 40920 5528 40969 5556
rect 40920 5516 40926 5528
rect 40957 5525 40969 5528
rect 41003 5525 41015 5559
rect 40957 5519 41015 5525
rect 43070 5516 43076 5568
rect 43128 5516 43134 5568
rect 460 5466 45540 5488
rect 460 5414 6070 5466
rect 6122 5414 6134 5466
rect 6186 5414 6198 5466
rect 6250 5414 6262 5466
rect 6314 5414 6326 5466
rect 6378 5414 11070 5466
rect 11122 5414 11134 5466
rect 11186 5414 11198 5466
rect 11250 5414 11262 5466
rect 11314 5414 11326 5466
rect 11378 5414 16070 5466
rect 16122 5414 16134 5466
rect 16186 5414 16198 5466
rect 16250 5414 16262 5466
rect 16314 5414 16326 5466
rect 16378 5414 21070 5466
rect 21122 5414 21134 5466
rect 21186 5414 21198 5466
rect 21250 5414 21262 5466
rect 21314 5414 21326 5466
rect 21378 5414 26070 5466
rect 26122 5414 26134 5466
rect 26186 5414 26198 5466
rect 26250 5414 26262 5466
rect 26314 5414 26326 5466
rect 26378 5414 31070 5466
rect 31122 5414 31134 5466
rect 31186 5414 31198 5466
rect 31250 5414 31262 5466
rect 31314 5414 31326 5466
rect 31378 5414 36070 5466
rect 36122 5414 36134 5466
rect 36186 5414 36198 5466
rect 36250 5414 36262 5466
rect 36314 5414 36326 5466
rect 36378 5414 41070 5466
rect 41122 5414 41134 5466
rect 41186 5414 41198 5466
rect 41250 5414 41262 5466
rect 41314 5414 41326 5466
rect 41378 5414 45540 5466
rect 460 5392 45540 5414
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 3418 5352 3424 5364
rect 2363 5324 3424 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4614 5352 4620 5364
rect 4295 5324 4620 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5321 4767 5355
rect 4709 5315 4767 5321
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5442 5352 5448 5364
rect 5123 5324 5448 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 4525 5219 4583 5225
rect 1903 5188 1992 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 1964 5089 1992 5188
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4724 5216 4752 5315
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6454 5352 6460 5364
rect 6319 5324 6460 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6454 5312 6460 5324
rect 6512 5352 6518 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6512 5324 7297 5352
rect 6512 5312 6518 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 7285 5315 7343 5321
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 7800 5324 8033 5352
rect 7800 5312 7806 5324
rect 8021 5321 8033 5324
rect 8067 5352 8079 5355
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8067 5324 8769 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8757 5321 8769 5324
rect 8803 5352 8815 5355
rect 9950 5352 9956 5364
rect 8803 5324 9956 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 9950 5312 9956 5324
rect 10008 5352 10014 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10008 5324 10701 5352
rect 10008 5312 10014 5324
rect 10689 5321 10701 5324
rect 10735 5352 10747 5355
rect 11790 5352 11796 5364
rect 10735 5324 11796 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13228 5324 14136 5352
rect 13228 5312 13234 5324
rect 8386 5244 8392 5296
rect 8444 5244 8450 5296
rect 9122 5244 9128 5296
rect 9180 5244 9186 5296
rect 11514 5244 11520 5296
rect 11572 5284 11578 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11572 5256 11897 5284
rect 11572 5244 11578 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 12176 5256 14044 5284
rect 4571 5188 4752 5216
rect 5169 5219 5227 5225
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5350 5216 5356 5228
rect 5215 5188 5356 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 8404 5216 8432 5244
rect 12176 5216 12204 5256
rect 6411 5188 6776 5216
rect 8404 5188 12204 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 6748 5160 6776 5188
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 13262 5216 13268 5228
rect 12943 5188 13268 5216
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 13722 5216 13728 5228
rect 13679 5188 13728 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 1949 5083 2007 5089
rect 1949 5049 1961 5083
rect 1995 5049 2007 5083
rect 1949 5043 2007 5049
rect 1121 5015 1179 5021
rect 1121 4981 1133 5015
rect 1167 5012 1179 5015
rect 1486 5012 1492 5024
rect 1167 4984 1492 5012
rect 1167 4981 1179 4984
rect 1121 4975 1179 4981
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1578 4972 1584 5024
rect 1636 5012 1642 5024
rect 1673 5015 1731 5021
rect 1673 5012 1685 5015
rect 1636 4984 1685 5012
rect 1636 4972 1642 4984
rect 1673 4981 1685 4984
rect 1719 4981 1731 5015
rect 1673 4975 1731 4981
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2424 5012 2452 5111
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 2648 5120 2774 5148
rect 2648 5108 2654 5120
rect 2372 4984 2452 5012
rect 2746 5012 2774 5120
rect 5258 5108 5264 5160
rect 5316 5148 5322 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 5316 5120 6561 5148
rect 5316 5108 5322 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6564 5080 6592 5111
rect 6730 5108 6736 5160
rect 6788 5108 6794 5160
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 10686 5148 10692 5160
rect 10367 5120 10692 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 12526 5148 12532 5160
rect 10744 5120 12532 5148
rect 10744 5108 10750 5120
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 13648 5148 13676 5179
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 12676 5120 13676 5148
rect 12676 5108 12682 5120
rect 14016 5092 14044 5256
rect 14108 5225 14136 5324
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 16482 5352 16488 5364
rect 15160 5324 15792 5352
rect 15160 5312 15166 5324
rect 15764 5296 15792 5324
rect 16316 5324 16488 5352
rect 14366 5244 14372 5296
rect 14424 5244 14430 5296
rect 15746 5244 15752 5296
rect 15804 5284 15810 5296
rect 16022 5284 16028 5296
rect 15804 5256 16028 5284
rect 15804 5244 15810 5256
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5185 14151 5219
rect 15654 5216 15660 5228
rect 15502 5188 15660 5216
rect 14093 5179 14151 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16316 5225 16344 5324
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 17052 5324 17264 5352
rect 17052 5296 17080 5324
rect 16574 5284 16580 5296
rect 16535 5256 16580 5284
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 16758 5244 16764 5296
rect 16816 5244 16822 5296
rect 17034 5244 17040 5296
rect 17092 5244 17098 5296
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 17236 5284 17264 5324
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 18196 5324 18613 5352
rect 18196 5312 18202 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 19794 5352 19800 5364
rect 18601 5315 18659 5321
rect 19260 5324 19800 5352
rect 18616 5284 18644 5315
rect 18877 5287 18935 5293
rect 18877 5284 18889 5287
rect 17236 5256 17618 5284
rect 18616 5256 18889 5284
rect 18877 5253 18889 5256
rect 18923 5253 18935 5287
rect 19260 5284 19288 5324
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 20070 5312 20076 5364
rect 20128 5352 20134 5364
rect 25593 5355 25651 5361
rect 20128 5324 24992 5352
rect 20128 5312 20134 5324
rect 18877 5247 18935 5253
rect 19168 5256 19288 5284
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16393 5219 16451 5225
rect 16393 5185 16405 5219
rect 16439 5216 16451 5219
rect 16776 5216 16804 5244
rect 16439 5188 16804 5216
rect 16439 5185 16451 5188
rect 16393 5179 16451 5185
rect 14734 5108 14740 5160
rect 14792 5148 14798 5160
rect 15562 5148 15568 5160
rect 14792 5120 15568 5148
rect 14792 5108 14798 5120
rect 15562 5108 15568 5120
rect 15620 5148 15626 5160
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 15620 5120 15853 5148
rect 15620 5108 15626 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 16224 5148 16252 5179
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 19168 5216 19196 5256
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 19429 5287 19487 5293
rect 19429 5284 19441 5287
rect 19392 5256 19441 5284
rect 19392 5244 19398 5256
rect 19429 5253 19441 5256
rect 19475 5253 19487 5287
rect 21818 5284 21824 5296
rect 20654 5256 21824 5284
rect 19429 5247 19487 5253
rect 21818 5244 21824 5256
rect 21876 5244 21882 5296
rect 22097 5287 22155 5293
rect 22097 5253 22109 5287
rect 22143 5284 22155 5287
rect 22554 5284 22560 5296
rect 22143 5256 22560 5284
rect 22143 5253 22155 5256
rect 22097 5247 22155 5253
rect 22554 5244 22560 5256
rect 22612 5244 22618 5296
rect 24581 5287 24639 5293
rect 24581 5284 24593 5287
rect 22756 5256 24593 5284
rect 22756 5228 22784 5256
rect 18748 5188 19196 5216
rect 21729 5219 21787 5225
rect 18748 5176 18754 5188
rect 21729 5185 21741 5219
rect 21775 5216 21787 5219
rect 21910 5216 21916 5228
rect 21775 5188 21916 5216
rect 21775 5185 21787 5188
rect 21729 5179 21787 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 22738 5176 22744 5228
rect 22796 5176 22802 5228
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 23290 5176 23296 5228
rect 23348 5176 23354 5228
rect 23768 5225 23796 5256
rect 24581 5253 24593 5256
rect 24627 5253 24639 5287
rect 24581 5247 24639 5253
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23753 5219 23811 5225
rect 23753 5185 23765 5219
rect 23799 5185 23811 5219
rect 23753 5179 23811 5185
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16224 5120 16773 5148
rect 15841 5111 15899 5117
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 19153 5151 19211 5157
rect 19153 5148 19165 5151
rect 16908 5120 19165 5148
rect 16908 5108 16914 5120
rect 19153 5117 19165 5120
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 20864 5120 21680 5148
rect 20864 5108 20870 5120
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6564 5052 7021 5080
rect 7009 5049 7021 5052
rect 7055 5080 7067 5083
rect 7282 5080 7288 5092
rect 7055 5052 7288 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 7282 5040 7288 5052
rect 7340 5080 7346 5092
rect 11241 5083 11299 5089
rect 7340 5052 8524 5080
rect 7340 5040 7346 5052
rect 8496 5024 8524 5052
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 11287 5052 13277 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 13265 5049 13277 5052
rect 13311 5080 13323 5083
rect 13311 5052 13860 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2746 4984 3065 5012
rect 2372 4972 2378 4984
rect 3053 4981 3065 4984
rect 3099 5012 3111 5015
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3099 4984 3893 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3881 4981 3893 4984
rect 3927 5012 3939 5015
rect 4062 5012 4068 5024
rect 3927 4984 4068 5012
rect 3927 4981 3939 4984
rect 3881 4975 3939 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4338 4972 4344 5024
rect 4396 4972 4402 5024
rect 5902 4972 5908 5024
rect 5960 4972 5966 5024
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 8294 5012 8300 5024
rect 7791 4984 8300 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8478 4972 8484 5024
rect 8536 4972 8542 5024
rect 9493 5015 9551 5021
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 11606 5012 11612 5024
rect 9539 4984 11612 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12066 4972 12072 5024
rect 12124 4972 12130 5024
rect 13832 5012 13860 5052
rect 13998 5040 14004 5092
rect 14056 5040 14062 5092
rect 21542 5080 21548 5092
rect 15948 5052 16804 5080
rect 15948 5012 15976 5052
rect 13832 4984 15976 5012
rect 16025 5015 16083 5021
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 16666 5012 16672 5024
rect 16071 4984 16672 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16776 5012 16804 5052
rect 20824 5052 21548 5080
rect 17218 5012 17224 5024
rect 16776 4984 17224 5012
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 19058 4972 19064 5024
rect 19116 4972 19122 5024
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 20824 5012 20852 5052
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 19484 4984 20852 5012
rect 19484 4972 19490 4984
rect 20898 4972 20904 5024
rect 20956 4972 20962 5024
rect 21652 5012 21680 5120
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 22833 5151 22891 5157
rect 22833 5148 22845 5151
rect 22520 5120 22845 5148
rect 22520 5108 22526 5120
rect 22833 5117 22845 5120
rect 22879 5148 22891 5151
rect 23124 5148 23152 5176
rect 22879 5120 23152 5148
rect 22879 5117 22891 5120
rect 22833 5111 22891 5117
rect 23676 5080 23704 5179
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 24964 5225 24992 5324
rect 25593 5321 25605 5355
rect 25639 5321 25651 5355
rect 25593 5315 25651 5321
rect 25608 5284 25636 5315
rect 25774 5312 25780 5364
rect 25832 5352 25838 5364
rect 26142 5352 26148 5364
rect 25832 5324 26148 5352
rect 25832 5312 25838 5324
rect 26142 5312 26148 5324
rect 26200 5312 26206 5364
rect 26786 5312 26792 5364
rect 26844 5352 26850 5364
rect 26844 5324 27016 5352
rect 26844 5312 26850 5324
rect 26988 5284 27016 5324
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27672 5324 28304 5352
rect 27672 5312 27678 5324
rect 25608 5256 26464 5284
rect 26988 5256 27094 5284
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5216 25007 5219
rect 25317 5219 25375 5225
rect 24995 5188 25176 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 24857 5151 24915 5157
rect 24857 5117 24869 5151
rect 24903 5148 24915 5151
rect 25038 5148 25044 5160
rect 24903 5120 25044 5148
rect 24903 5117 24915 5120
rect 24857 5111 24915 5117
rect 25038 5108 25044 5120
rect 25096 5108 25102 5160
rect 25148 5080 25176 5188
rect 25317 5185 25329 5219
rect 25363 5185 25375 5219
rect 25682 5216 25688 5228
rect 25317 5179 25375 5185
rect 25608 5188 25688 5216
rect 25332 5148 25360 5179
rect 25608 5148 25636 5188
rect 25682 5176 25688 5188
rect 25740 5176 25746 5228
rect 25774 5176 25780 5228
rect 25832 5176 25838 5228
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26326 5216 26332 5228
rect 26016 5188 26332 5216
rect 26016 5176 26022 5188
rect 26326 5176 26332 5188
rect 26384 5176 26390 5228
rect 26436 5216 26464 5256
rect 27890 5244 27896 5296
rect 27948 5284 27954 5296
rect 28123 5287 28181 5293
rect 28123 5284 28135 5287
rect 27948 5256 28135 5284
rect 27948 5244 27954 5256
rect 28123 5253 28135 5256
rect 28169 5253 28181 5287
rect 28123 5247 28181 5253
rect 28276 5225 28304 5324
rect 29086 5312 29092 5364
rect 29144 5312 29150 5364
rect 29546 5312 29552 5364
rect 29604 5312 29610 5364
rect 29917 5355 29975 5361
rect 29917 5321 29929 5355
rect 29963 5321 29975 5355
rect 29917 5315 29975 5321
rect 28813 5287 28871 5293
rect 28813 5253 28825 5287
rect 28859 5284 28871 5287
rect 29932 5284 29960 5315
rect 30374 5312 30380 5364
rect 30432 5312 30438 5364
rect 30742 5312 30748 5364
rect 30800 5312 30806 5364
rect 31570 5312 31576 5364
rect 31628 5312 31634 5364
rect 32582 5352 32588 5364
rect 31772 5324 32588 5352
rect 28859 5256 29960 5284
rect 28859 5253 28871 5256
rect 28813 5247 28871 5253
rect 26697 5219 26755 5225
rect 26697 5216 26709 5219
rect 26436 5188 26709 5216
rect 26697 5185 26709 5188
rect 26743 5185 26755 5219
rect 26697 5179 26755 5185
rect 28261 5219 28319 5225
rect 28261 5185 28273 5219
rect 28307 5185 28319 5219
rect 28261 5179 28319 5185
rect 28350 5176 28356 5228
rect 28408 5176 28414 5228
rect 29457 5219 29515 5225
rect 29457 5185 29469 5219
rect 29503 5185 29515 5219
rect 29457 5179 29515 5185
rect 28997 5151 29055 5157
rect 28997 5148 29009 5151
rect 25332 5120 25636 5148
rect 26344 5120 29009 5148
rect 26344 5080 26372 5120
rect 28997 5117 29009 5120
rect 29043 5117 29055 5151
rect 28997 5111 29055 5117
rect 28629 5083 28687 5089
rect 28629 5080 28641 5083
rect 22480 5052 23704 5080
rect 24136 5052 24532 5080
rect 25148 5052 26372 5080
rect 27448 5052 28641 5080
rect 22002 5012 22008 5024
rect 21652 4984 22008 5012
rect 22002 4972 22008 4984
rect 22060 5012 22066 5024
rect 22480 5012 22508 5052
rect 22060 4984 22508 5012
rect 22060 4972 22066 4984
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 23474 4972 23480 5024
rect 23532 4972 23538 5024
rect 24136 5021 24164 5052
rect 24504 5024 24532 5052
rect 24121 5015 24179 5021
rect 24121 4981 24133 5015
rect 24167 4981 24179 5015
rect 24121 4975 24179 4981
rect 24302 4972 24308 5024
rect 24360 4972 24366 5024
rect 24486 4972 24492 5024
rect 24544 4972 24550 5024
rect 25222 4972 25228 5024
rect 25280 4972 25286 5024
rect 25501 5015 25559 5021
rect 25501 4981 25513 5015
rect 25547 5012 25559 5015
rect 25774 5012 25780 5024
rect 25547 4984 25780 5012
rect 25547 4981 25559 4984
rect 25501 4975 25559 4981
rect 25774 4972 25780 4984
rect 25832 4972 25838 5024
rect 26050 4972 26056 5024
rect 26108 4972 26114 5024
rect 26142 4972 26148 5024
rect 26200 5012 26206 5024
rect 27448 5012 27476 5052
rect 28629 5049 28641 5052
rect 28675 5049 28687 5083
rect 29472 5080 29500 5179
rect 30282 5176 30288 5228
rect 30340 5176 30346 5228
rect 30392 5216 30420 5312
rect 30760 5284 30788 5312
rect 31588 5284 31616 5312
rect 31772 5293 31800 5324
rect 32582 5312 32588 5324
rect 32640 5312 32646 5364
rect 32674 5312 32680 5364
rect 32732 5352 32738 5364
rect 33781 5355 33839 5361
rect 32732 5324 32904 5352
rect 32732 5312 32738 5324
rect 30760 5256 31248 5284
rect 31220 5225 31248 5256
rect 31496 5256 31616 5284
rect 31757 5287 31815 5293
rect 31496 5225 31524 5256
rect 31757 5253 31769 5287
rect 31803 5253 31815 5287
rect 31757 5247 31815 5253
rect 32876 5228 32904 5324
rect 33781 5321 33793 5355
rect 33827 5352 33839 5355
rect 34330 5352 34336 5364
rect 33827 5324 34336 5352
rect 33827 5321 33839 5324
rect 33781 5315 33839 5321
rect 34330 5312 34336 5324
rect 34388 5312 34394 5364
rect 35360 5324 36308 5352
rect 33689 5287 33747 5293
rect 33689 5253 33701 5287
rect 33735 5284 33747 5287
rect 35360 5284 35388 5324
rect 33735 5256 35388 5284
rect 36280 5284 36308 5324
rect 36354 5312 36360 5364
rect 36412 5352 36418 5364
rect 36449 5355 36507 5361
rect 36449 5352 36461 5355
rect 36412 5324 36461 5352
rect 36412 5312 36418 5324
rect 36449 5321 36461 5324
rect 36495 5352 36507 5355
rect 36814 5352 36820 5364
rect 36495 5324 36820 5352
rect 36495 5321 36507 5324
rect 36449 5315 36507 5321
rect 36814 5312 36820 5324
rect 36872 5312 36878 5364
rect 39485 5355 39543 5361
rect 38396 5324 39436 5352
rect 38396 5284 38424 5324
rect 36280 5256 38424 5284
rect 39408 5284 39436 5324
rect 39485 5321 39497 5355
rect 39531 5352 39543 5355
rect 40034 5352 40040 5364
rect 39531 5324 40040 5352
rect 39531 5321 39543 5324
rect 39485 5315 39543 5321
rect 40034 5312 40040 5324
rect 40092 5352 40098 5364
rect 40586 5352 40592 5364
rect 40092 5324 40592 5352
rect 40092 5312 40098 5324
rect 40586 5312 40592 5324
rect 40644 5312 40650 5364
rect 40954 5312 40960 5364
rect 41012 5352 41018 5364
rect 41417 5355 41475 5361
rect 41417 5352 41429 5355
rect 41012 5324 41429 5352
rect 41012 5312 41018 5324
rect 41417 5321 41429 5324
rect 41463 5352 41475 5355
rect 41782 5352 41788 5364
rect 41463 5324 41788 5352
rect 41463 5321 41475 5324
rect 41417 5315 41475 5321
rect 41782 5312 41788 5324
rect 41840 5352 41846 5364
rect 42337 5355 42395 5361
rect 42337 5352 42349 5355
rect 41840 5324 42349 5352
rect 41840 5312 41846 5324
rect 42337 5321 42349 5324
rect 42383 5352 42395 5355
rect 43070 5352 43076 5364
rect 42383 5324 43076 5352
rect 42383 5321 42395 5324
rect 42337 5315 42395 5321
rect 43070 5312 43076 5324
rect 43128 5352 43134 5364
rect 43441 5355 43499 5361
rect 43441 5352 43453 5355
rect 43128 5324 43453 5352
rect 43128 5312 43134 5324
rect 43441 5321 43453 5324
rect 43487 5352 43499 5355
rect 43809 5355 43867 5361
rect 43809 5352 43821 5355
rect 43487 5324 43821 5352
rect 43487 5321 43499 5324
rect 43441 5315 43499 5321
rect 43809 5321 43821 5324
rect 43855 5352 43867 5355
rect 43990 5352 43996 5364
rect 43855 5324 43996 5352
rect 43855 5321 43867 5324
rect 43809 5315 43867 5321
rect 43990 5312 43996 5324
rect 44048 5312 44054 5364
rect 44542 5312 44548 5364
rect 44600 5312 44606 5364
rect 40126 5284 40132 5296
rect 39408 5256 40132 5284
rect 33735 5253 33747 5256
rect 33689 5247 33747 5253
rect 40126 5244 40132 5256
rect 40184 5244 40190 5296
rect 42797 5287 42855 5293
rect 42797 5253 42809 5287
rect 42843 5284 42855 5287
rect 42886 5284 42892 5296
rect 42843 5256 42892 5284
rect 42843 5253 42855 5256
rect 42797 5247 42855 5253
rect 42886 5244 42892 5256
rect 42944 5284 42950 5296
rect 43346 5284 43352 5296
rect 42944 5256 43352 5284
rect 42944 5244 42950 5256
rect 43346 5244 43352 5256
rect 43404 5244 43410 5296
rect 31021 5219 31079 5225
rect 31021 5216 31033 5219
rect 30392 5188 31033 5216
rect 31021 5185 31033 5188
rect 31067 5185 31079 5219
rect 31021 5179 31079 5185
rect 31205 5219 31263 5225
rect 31205 5185 31217 5219
rect 31251 5185 31263 5219
rect 31205 5179 31263 5185
rect 31481 5219 31539 5225
rect 31481 5185 31493 5219
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 32858 5176 32864 5228
rect 32916 5176 32922 5228
rect 34514 5176 34520 5228
rect 34572 5216 34578 5228
rect 34609 5219 34667 5225
rect 34609 5216 34621 5219
rect 34572 5188 34621 5216
rect 34572 5176 34578 5188
rect 34609 5185 34621 5188
rect 34655 5185 34667 5219
rect 34609 5179 34667 5185
rect 36078 5176 36084 5228
rect 36136 5216 36142 5228
rect 36630 5216 36636 5228
rect 36136 5188 36636 5216
rect 36136 5176 36142 5188
rect 36630 5176 36636 5188
rect 36688 5176 36694 5228
rect 36817 5219 36875 5225
rect 36817 5185 36829 5219
rect 36863 5216 36875 5219
rect 37090 5216 37096 5228
rect 36863 5188 37096 5216
rect 36863 5185 36875 5188
rect 36817 5179 36875 5185
rect 37090 5176 37096 5188
rect 37148 5176 37154 5228
rect 37274 5176 37280 5228
rect 37332 5216 37338 5228
rect 37737 5219 37795 5225
rect 37737 5216 37749 5219
rect 37332 5188 37749 5216
rect 37332 5176 37338 5188
rect 37737 5185 37749 5188
rect 37783 5185 37795 5219
rect 37737 5179 37795 5185
rect 39022 5176 39028 5228
rect 39080 5216 39086 5228
rect 39390 5216 39396 5228
rect 39080 5188 39396 5216
rect 39080 5176 39086 5188
rect 39390 5176 39396 5188
rect 39448 5176 39454 5228
rect 39942 5176 39948 5228
rect 40000 5176 40006 5228
rect 40773 5219 40831 5225
rect 40773 5185 40785 5219
rect 40819 5216 40831 5219
rect 42058 5216 42064 5228
rect 40819 5188 42064 5216
rect 40819 5185 40831 5188
rect 40773 5179 40831 5185
rect 42058 5176 42064 5188
rect 42116 5176 42122 5228
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 29641 5151 29699 5157
rect 29641 5148 29653 5151
rect 29604 5120 29653 5148
rect 29604 5108 29610 5120
rect 29641 5117 29653 5120
rect 29687 5148 29699 5151
rect 30190 5148 30196 5160
rect 29687 5120 30196 5148
rect 29687 5117 29699 5120
rect 29641 5111 29699 5117
rect 30190 5108 30196 5120
rect 30248 5148 30254 5160
rect 30469 5151 30527 5157
rect 30469 5148 30481 5151
rect 30248 5120 30481 5148
rect 30248 5108 30254 5120
rect 30469 5117 30481 5120
rect 30515 5117 30527 5151
rect 30469 5111 30527 5117
rect 30558 5108 30564 5160
rect 30616 5148 30622 5160
rect 30929 5151 30987 5157
rect 30929 5148 30941 5151
rect 30616 5120 30941 5148
rect 30616 5108 30622 5120
rect 30929 5117 30941 5120
rect 30975 5117 30987 5151
rect 30929 5111 30987 5117
rect 31113 5151 31171 5157
rect 31113 5117 31125 5151
rect 31159 5148 31171 5151
rect 31386 5148 31392 5160
rect 31159 5120 31392 5148
rect 31159 5117 31171 5120
rect 31113 5111 31171 5117
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 33965 5151 34023 5157
rect 31588 5120 33824 5148
rect 31588 5080 31616 5120
rect 33796 5080 33824 5120
rect 33965 5117 33977 5151
rect 34011 5148 34023 5151
rect 34146 5148 34152 5160
rect 34011 5120 34152 5148
rect 34011 5117 34023 5120
rect 33965 5111 34023 5117
rect 34146 5108 34152 5120
rect 34204 5108 34210 5160
rect 34238 5108 34244 5160
rect 34296 5148 34302 5160
rect 34698 5148 34704 5160
rect 34296 5120 34704 5148
rect 34296 5108 34302 5120
rect 34698 5108 34704 5120
rect 34756 5108 34762 5160
rect 34977 5151 35035 5157
rect 34977 5117 34989 5151
rect 35023 5148 35035 5151
rect 35023 5120 36676 5148
rect 35023 5117 35035 5120
rect 34977 5111 35035 5117
rect 36648 5089 36676 5120
rect 36722 5108 36728 5160
rect 36780 5148 36786 5160
rect 37461 5151 37519 5157
rect 37461 5148 37473 5151
rect 36780 5120 37473 5148
rect 36780 5108 36786 5120
rect 37461 5117 37473 5120
rect 37507 5117 37519 5151
rect 37461 5111 37519 5117
rect 38010 5108 38016 5160
rect 38068 5108 38074 5160
rect 39298 5108 39304 5160
rect 39356 5108 39362 5160
rect 39574 5108 39580 5160
rect 39632 5148 39638 5160
rect 40129 5151 40187 5157
rect 40129 5148 40141 5151
rect 39632 5120 40141 5148
rect 39632 5108 39638 5120
rect 40129 5117 40141 5120
rect 40175 5117 40187 5151
rect 40129 5111 40187 5117
rect 40862 5108 40868 5160
rect 40920 5108 40926 5160
rect 40954 5108 40960 5160
rect 41012 5108 41018 5160
rect 36633 5083 36691 5089
rect 29472 5052 31616 5080
rect 32784 5052 33456 5080
rect 33796 5052 34836 5080
rect 28629 5043 28687 5049
rect 26200 4984 27476 5012
rect 26200 4972 26206 4984
rect 28258 4972 28264 5024
rect 28316 4972 28322 5024
rect 29178 4972 29184 5024
rect 29236 5012 29242 5024
rect 30745 5015 30803 5021
rect 30745 5012 30757 5015
rect 29236 4984 30757 5012
rect 29236 4972 29242 4984
rect 30745 4981 30757 4984
rect 30791 4981 30803 5015
rect 30745 4975 30803 4981
rect 31386 4972 31392 5024
rect 31444 5012 31450 5024
rect 32784 5012 32812 5052
rect 31444 4984 32812 5012
rect 31444 4972 31450 4984
rect 32858 4972 32864 5024
rect 32916 5012 32922 5024
rect 33229 5015 33287 5021
rect 33229 5012 33241 5015
rect 32916 4984 33241 5012
rect 32916 4972 32922 4984
rect 33229 4981 33241 4984
rect 33275 4981 33287 5015
rect 33229 4975 33287 4981
rect 33318 4972 33324 5024
rect 33376 4972 33382 5024
rect 33428 5012 33456 5052
rect 34146 5012 34152 5024
rect 33428 4984 34152 5012
rect 34146 4972 34152 4984
rect 34204 4972 34210 5024
rect 34422 4972 34428 5024
rect 34480 4972 34486 5024
rect 34808 5012 34836 5052
rect 36633 5049 36645 5083
rect 36679 5049 36691 5083
rect 39316 5080 39344 5108
rect 40405 5083 40463 5089
rect 40405 5080 40417 5083
rect 39316 5052 40417 5080
rect 36633 5043 36691 5049
rect 40405 5049 40417 5052
rect 40451 5049 40463 5083
rect 44913 5083 44971 5089
rect 44913 5080 44925 5083
rect 40405 5043 40463 5049
rect 44100 5052 44925 5080
rect 44100 5024 44128 5052
rect 44913 5049 44925 5052
rect 44959 5049 44971 5083
rect 44913 5043 44971 5049
rect 35342 5012 35348 5024
rect 34808 4984 35348 5012
rect 35342 4972 35348 4984
rect 35400 4972 35406 5024
rect 36446 4972 36452 5024
rect 36504 5012 36510 5024
rect 37093 5015 37151 5021
rect 37093 5012 37105 5015
rect 36504 4984 37105 5012
rect 36504 4972 36510 4984
rect 37093 4981 37105 4984
rect 37139 4981 37151 5015
rect 37093 4975 37151 4981
rect 39206 4972 39212 5024
rect 39264 5012 39270 5024
rect 39577 5015 39635 5021
rect 39577 5012 39589 5015
rect 39264 4984 39589 5012
rect 39264 4972 39270 4984
rect 39577 4981 39589 4984
rect 39623 4981 39635 5015
rect 39577 4975 39635 4981
rect 41966 4972 41972 5024
rect 42024 4972 42030 5024
rect 44082 4972 44088 5024
rect 44140 4972 44146 5024
rect 44174 4972 44180 5024
rect 44232 4972 44238 5024
rect 460 4922 45540 4944
rect 460 4870 3570 4922
rect 3622 4870 3634 4922
rect 3686 4870 3698 4922
rect 3750 4870 3762 4922
rect 3814 4870 3826 4922
rect 3878 4870 8570 4922
rect 8622 4870 8634 4922
rect 8686 4870 8698 4922
rect 8750 4870 8762 4922
rect 8814 4870 8826 4922
rect 8878 4870 13570 4922
rect 13622 4870 13634 4922
rect 13686 4870 13698 4922
rect 13750 4870 13762 4922
rect 13814 4870 13826 4922
rect 13878 4870 18570 4922
rect 18622 4870 18634 4922
rect 18686 4870 18698 4922
rect 18750 4870 18762 4922
rect 18814 4870 18826 4922
rect 18878 4870 23570 4922
rect 23622 4870 23634 4922
rect 23686 4870 23698 4922
rect 23750 4870 23762 4922
rect 23814 4870 23826 4922
rect 23878 4870 28570 4922
rect 28622 4870 28634 4922
rect 28686 4870 28698 4922
rect 28750 4870 28762 4922
rect 28814 4870 28826 4922
rect 28878 4870 33570 4922
rect 33622 4870 33634 4922
rect 33686 4870 33698 4922
rect 33750 4870 33762 4922
rect 33814 4870 33826 4922
rect 33878 4870 38570 4922
rect 38622 4870 38634 4922
rect 38686 4870 38698 4922
rect 38750 4870 38762 4922
rect 38814 4870 38826 4922
rect 38878 4870 43570 4922
rect 43622 4870 43634 4922
rect 43686 4870 43698 4922
rect 43750 4870 43762 4922
rect 43814 4870 43826 4922
rect 43878 4870 45540 4922
rect 460 4848 45540 4870
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 1228 4780 3157 4808
rect 1228 4672 1256 4780
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 11609 4811 11667 4817
rect 3145 4771 3203 4777
rect 9508 4780 10916 4808
rect 9508 4749 9536 4780
rect 9493 4743 9551 4749
rect 9493 4709 9505 4743
rect 9539 4709 9551 4743
rect 9493 4703 9551 4709
rect 10045 4743 10103 4749
rect 10045 4709 10057 4743
rect 10091 4709 10103 4743
rect 10888 4740 10916 4780
rect 11609 4777 11621 4811
rect 11655 4808 11667 4811
rect 11790 4808 11796 4820
rect 11655 4780 11796 4808
rect 11655 4777 11667 4780
rect 11609 4771 11667 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 12308 4780 12541 4808
rect 12308 4768 12314 4780
rect 12529 4777 12541 4780
rect 12575 4777 12587 4811
rect 12529 4771 12587 4777
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14090 4808 14096 4820
rect 14047 4780 14096 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14090 4768 14096 4780
rect 14148 4808 14154 4820
rect 14148 4780 15792 4808
rect 14148 4768 14154 4780
rect 13906 4740 13912 4752
rect 10888 4712 13912 4740
rect 10045 4703 10103 4709
rect 1136 4644 1256 4672
rect 1489 4675 1547 4681
rect 1136 4613 1164 4644
rect 1489 4641 1501 4675
rect 1535 4672 1547 4675
rect 1578 4672 1584 4684
rect 1535 4644 1584 4672
rect 1535 4641 1547 4644
rect 1489 4635 1547 4641
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4672 3847 4675
rect 4062 4672 4068 4684
rect 3835 4644 4068 4672
rect 3835 4641 3847 4644
rect 3789 4635 3847 4641
rect 4062 4632 4068 4644
rect 4120 4672 4126 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4120 4644 4813 4672
rect 4120 4632 4126 4644
rect 4801 4641 4813 4644
rect 4847 4672 4859 4675
rect 5258 4672 5264 4684
rect 4847 4644 5264 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 8113 4675 8171 4681
rect 8113 4641 8125 4675
rect 8159 4672 8171 4675
rect 8294 4672 8300 4684
rect 8159 4644 8300 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8536 4644 8953 4672
rect 8536 4632 8542 4644
rect 8941 4641 8953 4644
rect 8987 4672 8999 4675
rect 9306 4672 9312 4684
rect 8987 4644 9312 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 1121 4607 1179 4613
rect 1121 4573 1133 4607
rect 1167 4573 1179 4607
rect 1121 4567 1179 4573
rect 1213 4607 1271 4613
rect 1213 4573 1225 4607
rect 1259 4573 1271 4607
rect 1213 4567 1271 4573
rect 1228 4536 1256 4567
rect 2590 4564 2596 4616
rect 2648 4564 2654 4616
rect 3510 4564 3516 4616
rect 3568 4604 3574 4616
rect 3970 4604 3976 4616
rect 3568 4576 3976 4604
rect 3568 4564 3574 4576
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 4614 4604 4620 4616
rect 4571 4576 4620 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7331 4576 8340 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 1486 4536 1492 4548
rect 1228 4508 1492 4536
rect 1486 4496 1492 4508
rect 1544 4496 1550 4548
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3605 4539 3663 4545
rect 3605 4536 3617 4539
rect 2832 4508 3617 4536
rect 2832 4496 2838 4508
rect 3605 4505 3617 4508
rect 3651 4505 3663 4539
rect 3605 4499 3663 4505
rect 4706 4496 4712 4548
rect 4764 4496 4770 4548
rect 5261 4539 5319 4545
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5534 4536 5540 4548
rect 5307 4508 5540 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 5644 4508 5750 4536
rect 934 4428 940 4480
rect 992 4428 998 4480
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2372 4440 2973 4468
rect 2372 4428 2378 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 4154 4428 4160 4480
rect 4212 4428 4218 4480
rect 4614 4428 4620 4480
rect 4672 4428 4678 4480
rect 4724 4468 4752 4496
rect 5644 4468 5672 4508
rect 4724 4440 5672 4468
rect 6730 4428 6736 4480
rect 6788 4428 6794 4480
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 6972 4440 7113 4468
rect 6972 4428 6978 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 7926 4468 7932 4480
rect 7791 4440 7932 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8312 4477 8340 4576
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8665 4607 8723 4613
rect 8665 4604 8677 4607
rect 8444 4576 8677 4604
rect 8444 4564 8450 4576
rect 8665 4573 8677 4576
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 10060 4604 10088 4703
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 10652 4644 12265 4672
rect 10652 4632 10658 4644
rect 12253 4641 12265 4644
rect 12299 4672 12311 4675
rect 13081 4675 13139 4681
rect 13081 4672 13093 4675
rect 12299 4644 13093 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 13081 4641 13093 4644
rect 13127 4672 13139 4675
rect 13998 4672 14004 4684
rect 13127 4644 14004 4672
rect 13127 4641 13139 4644
rect 13081 4635 13139 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 15764 4616 15792 4780
rect 15838 4768 15844 4820
rect 15896 4768 15902 4820
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 17126 4768 17132 4820
rect 17184 4808 17190 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 17184 4780 18337 4808
rect 17184 4768 17190 4780
rect 18325 4777 18337 4780
rect 18371 4777 18383 4811
rect 18325 4771 18383 4777
rect 19426 4768 19432 4820
rect 19484 4768 19490 4820
rect 19702 4768 19708 4820
rect 19760 4768 19766 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 20990 4808 20996 4820
rect 20763 4780 20996 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 21453 4811 21511 4817
rect 21453 4777 21465 4811
rect 21499 4808 21511 4811
rect 21818 4808 21824 4820
rect 21499 4780 21824 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 22554 4808 22560 4820
rect 21928 4780 22560 4808
rect 9815 4576 10088 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13228 4576 14105 4604
rect 13228 4564 13234 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 15746 4564 15752 4616
rect 15804 4564 15810 4616
rect 15856 4604 15884 4768
rect 15930 4700 15936 4752
rect 15988 4700 15994 4752
rect 16408 4672 16436 4768
rect 17954 4700 17960 4752
rect 18012 4700 18018 4752
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18141 4743 18199 4749
rect 18141 4740 18153 4743
rect 18104 4712 18153 4740
rect 18104 4700 18110 4712
rect 18141 4709 18153 4712
rect 18187 4709 18199 4743
rect 18141 4703 18199 4709
rect 19518 4700 19524 4752
rect 19576 4740 19582 4752
rect 19981 4743 20039 4749
rect 19981 4740 19993 4743
rect 19576 4712 19993 4740
rect 19576 4700 19582 4712
rect 19981 4709 19993 4712
rect 20027 4709 20039 4743
rect 19981 4703 20039 4709
rect 16224 4644 16436 4672
rect 16224 4613 16252 4644
rect 16117 4607 16175 4613
rect 16117 4604 16129 4607
rect 15856 4576 16129 4604
rect 16117 4573 16129 4576
rect 16163 4573 16175 4607
rect 16117 4567 16175 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4573 16267 4607
rect 16209 4567 16267 4573
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 17972 4604 18000 4700
rect 20438 4672 20444 4684
rect 19996 4644 20444 4672
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 17972 4576 18245 4604
rect 16393 4567 16451 4573
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 8757 4539 8815 4545
rect 8757 4536 8769 4539
rect 8404 4508 8769 4536
rect 8404 4480 8432 4508
rect 8757 4505 8769 4508
rect 8803 4505 8815 4539
rect 8757 4499 8815 4505
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 11664 4508 14320 4536
rect 11664 4496 11670 4508
rect 8297 4471 8355 4477
rect 8297 4437 8309 4471
rect 8343 4437 8355 4471
rect 8297 4431 8355 4437
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 9582 4428 9588 4480
rect 9640 4428 9646 4480
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 10505 4471 10563 4477
rect 10505 4437 10517 4471
rect 10551 4468 10563 4471
rect 10686 4468 10692 4480
rect 10551 4440 10692 4468
rect 10551 4437 10563 4440
rect 10505 4431 10563 4437
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 11514 4468 11520 4480
rect 11287 4440 11520 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 11698 4428 11704 4480
rect 11756 4428 11762 4480
rect 12084 4477 12112 4508
rect 12069 4471 12127 4477
rect 12069 4437 12081 4471
rect 12115 4437 12127 4471
rect 12069 4431 12127 4437
rect 12158 4428 12164 4480
rect 12216 4428 12222 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 12860 4440 12909 4468
rect 12860 4428 12866 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 12986 4428 12992 4480
rect 13044 4428 13050 4480
rect 14292 4468 14320 4508
rect 14366 4496 14372 4548
rect 14424 4496 14430 4548
rect 15654 4536 15660 4548
rect 15594 4508 15660 4536
rect 15654 4496 15660 4508
rect 15712 4536 15718 4548
rect 15838 4536 15844 4548
rect 15712 4508 15844 4536
rect 15712 4496 15718 4508
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 15933 4539 15991 4545
rect 15933 4505 15945 4539
rect 15979 4536 15991 4539
rect 16022 4536 16028 4548
rect 15979 4508 16028 4536
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 16408 4536 16436 4567
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 19058 4604 19064 4616
rect 18472 4576 19064 4604
rect 18472 4564 18478 4576
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 16574 4536 16580 4548
rect 16408 4508 16580 4536
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16669 4539 16727 4545
rect 16669 4505 16681 4539
rect 16715 4536 16727 4539
rect 16942 4536 16948 4548
rect 16715 4508 16948 4536
rect 16715 4505 16727 4508
rect 16669 4499 16727 4505
rect 16942 4496 16948 4508
rect 17000 4496 17006 4548
rect 17126 4496 17132 4548
rect 17184 4496 17190 4548
rect 19628 4536 19656 4567
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 19996 4604 20024 4644
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 20990 4632 20996 4684
rect 21048 4672 21054 4684
rect 21085 4675 21143 4681
rect 21085 4672 21097 4675
rect 21048 4644 21097 4672
rect 21048 4632 21054 4644
rect 21085 4641 21097 4644
rect 21131 4672 21143 4675
rect 21928 4672 21956 4780
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 22646 4768 22652 4820
rect 22704 4808 22710 4820
rect 23753 4811 23811 4817
rect 23753 4808 23765 4811
rect 22704 4780 23765 4808
rect 22704 4768 22710 4780
rect 23753 4777 23765 4780
rect 23799 4777 23811 4811
rect 23753 4771 23811 4777
rect 23842 4768 23848 4820
rect 23900 4808 23906 4820
rect 24578 4808 24584 4820
rect 23900 4780 24584 4808
rect 23900 4768 23906 4780
rect 24578 4768 24584 4780
rect 24636 4808 24642 4820
rect 25409 4811 25467 4817
rect 25409 4808 25421 4811
rect 24636 4780 25421 4808
rect 24636 4768 24642 4780
rect 25409 4777 25421 4780
rect 25455 4777 25467 4811
rect 25409 4771 25467 4777
rect 25792 4780 30236 4808
rect 24670 4740 24676 4752
rect 23216 4712 24676 4740
rect 21131 4644 21956 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 19935 4576 20024 4604
rect 20073 4607 20131 4613
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20898 4604 20904 4616
rect 20119 4576 20904 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21836 4613 21864 4644
rect 22094 4632 22100 4684
rect 22152 4632 22158 4684
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4573 21787 4607
rect 21729 4567 21787 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4573 21879 4607
rect 21821 4567 21879 4573
rect 19978 4536 19984 4548
rect 19076 4508 19564 4536
rect 19628 4508 19984 4536
rect 19076 4477 19104 4508
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 14292 4440 19073 4468
rect 19061 4437 19073 4440
rect 19107 4437 19119 4471
rect 19536 4468 19564 4508
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 21634 4536 21640 4548
rect 20916 4508 21640 4536
rect 20916 4468 20944 4508
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 21744 4536 21772 4567
rect 23106 4564 23112 4616
rect 23164 4604 23170 4616
rect 23216 4604 23244 4712
rect 24670 4700 24676 4712
rect 24728 4740 24734 4752
rect 24765 4743 24823 4749
rect 24765 4740 24777 4743
rect 24728 4712 24777 4740
rect 24728 4700 24734 4712
rect 24765 4709 24777 4712
rect 24811 4709 24823 4743
rect 24765 4703 24823 4709
rect 25130 4700 25136 4752
rect 25188 4700 25194 4752
rect 23290 4632 23296 4684
rect 23348 4632 23354 4684
rect 23934 4632 23940 4684
rect 23992 4672 23998 4684
rect 24305 4675 24363 4681
rect 24305 4672 24317 4675
rect 23992 4644 24317 4672
rect 23992 4632 23998 4644
rect 24305 4641 24317 4644
rect 24351 4641 24363 4675
rect 24305 4635 24363 4641
rect 24946 4632 24952 4684
rect 25004 4672 25010 4684
rect 25041 4675 25099 4681
rect 25041 4672 25053 4675
rect 25004 4644 25053 4672
rect 25004 4632 25010 4644
rect 25041 4641 25053 4644
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 23164 4590 23244 4604
rect 23308 4604 23336 4632
rect 25148 4613 25176 4700
rect 25792 4672 25820 4780
rect 27430 4700 27436 4752
rect 27488 4740 27494 4752
rect 30006 4740 30012 4752
rect 27488 4712 30012 4740
rect 27488 4700 27494 4712
rect 30006 4700 30012 4712
rect 30064 4700 30070 4752
rect 30208 4740 30236 4780
rect 30282 4768 30288 4820
rect 30340 4808 30346 4820
rect 32950 4808 32956 4820
rect 30340 4780 32956 4808
rect 30340 4768 30346 4780
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 33781 4811 33839 4817
rect 33781 4777 33793 4811
rect 33827 4808 33839 4811
rect 34330 4808 34336 4820
rect 33827 4780 34336 4808
rect 33827 4777 33839 4780
rect 33781 4771 33839 4777
rect 34330 4768 34336 4780
rect 34388 4768 34394 4820
rect 34514 4768 34520 4820
rect 34572 4808 34578 4820
rect 36725 4811 36783 4817
rect 36725 4808 36737 4811
rect 34572 4780 36737 4808
rect 34572 4768 34578 4780
rect 36725 4777 36737 4780
rect 36771 4777 36783 4811
rect 36725 4771 36783 4777
rect 38010 4768 38016 4820
rect 38068 4808 38074 4820
rect 38197 4811 38255 4817
rect 38197 4808 38209 4811
rect 38068 4780 38209 4808
rect 38068 4768 38074 4780
rect 38197 4777 38209 4780
rect 38243 4777 38255 4811
rect 38197 4771 38255 4777
rect 38378 4768 38384 4820
rect 38436 4808 38442 4820
rect 38657 4811 38715 4817
rect 38657 4808 38669 4811
rect 38436 4780 38669 4808
rect 38436 4768 38442 4780
rect 38657 4777 38669 4780
rect 38703 4777 38715 4811
rect 38657 4771 38715 4777
rect 38841 4811 38899 4817
rect 38841 4777 38853 4811
rect 38887 4808 38899 4811
rect 39482 4808 39488 4820
rect 38887 4780 39488 4808
rect 38887 4777 38899 4780
rect 38841 4771 38899 4777
rect 39482 4768 39488 4780
rect 39540 4768 39546 4820
rect 40586 4808 40592 4820
rect 39592 4780 40592 4808
rect 31846 4740 31852 4752
rect 30208 4712 31852 4740
rect 31846 4700 31852 4712
rect 31904 4700 31910 4752
rect 34054 4700 34060 4752
rect 34112 4700 34118 4752
rect 35342 4700 35348 4752
rect 35400 4740 35406 4752
rect 35897 4743 35955 4749
rect 35897 4740 35909 4743
rect 35400 4712 35909 4740
rect 35400 4700 35406 4712
rect 35897 4709 35909 4712
rect 35943 4709 35955 4743
rect 35897 4703 35955 4709
rect 35986 4700 35992 4752
rect 36044 4740 36050 4752
rect 36446 4740 36452 4752
rect 36044 4712 36452 4740
rect 36044 4700 36050 4712
rect 36446 4700 36452 4712
rect 36504 4700 36510 4752
rect 37918 4740 37924 4752
rect 36556 4712 37924 4740
rect 25516 4644 25820 4672
rect 25516 4613 25544 4644
rect 26786 4632 26792 4684
rect 26844 4672 26850 4684
rect 27525 4675 27583 4681
rect 26844 4644 27200 4672
rect 26844 4632 26850 4644
rect 25133 4607 25191 4613
rect 23164 4576 23230 4590
rect 23308 4576 25084 4604
rect 23164 4564 23170 4576
rect 22370 4536 22376 4548
rect 21744 4508 22376 4536
rect 22370 4496 22376 4508
rect 22428 4496 22434 4548
rect 24213 4539 24271 4545
rect 24213 4536 24225 4539
rect 23584 4508 24225 4536
rect 19536 4440 20944 4468
rect 19061 4431 19119 4437
rect 21542 4428 21548 4480
rect 21600 4428 21606 4480
rect 22462 4428 22468 4480
rect 22520 4468 22526 4480
rect 23584 4477 23612 4508
rect 24213 4505 24225 4508
rect 24259 4505 24271 4539
rect 24762 4536 24768 4548
rect 24213 4499 24271 4505
rect 24596 4508 24768 4536
rect 23569 4471 23627 4477
rect 23569 4468 23581 4471
rect 22520 4440 23581 4468
rect 22520 4428 22526 4440
rect 23569 4437 23581 4440
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 24118 4428 24124 4480
rect 24176 4468 24182 4480
rect 24596 4468 24624 4508
rect 24762 4496 24768 4508
rect 24820 4496 24826 4548
rect 25056 4536 25084 4576
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 25501 4607 25559 4613
rect 25501 4573 25513 4607
rect 25547 4573 25559 4607
rect 25777 4607 25835 4613
rect 25777 4600 25789 4607
rect 25501 4567 25559 4573
rect 25700 4573 25789 4600
rect 25823 4573 25835 4607
rect 27172 4590 27200 4644
rect 27525 4641 27537 4675
rect 27571 4672 27583 4675
rect 27982 4672 27988 4684
rect 27571 4644 27988 4672
rect 27571 4641 27583 4644
rect 27525 4635 27583 4641
rect 25700 4572 25835 4573
rect 25516 4536 25544 4567
rect 25056 4508 25544 4536
rect 25590 4496 25596 4548
rect 25648 4536 25654 4548
rect 25700 4536 25728 4572
rect 25777 4567 25835 4572
rect 27706 4564 27712 4616
rect 27764 4564 27770 4616
rect 27816 4613 27844 4644
rect 27982 4632 27988 4644
rect 28040 4632 28046 4684
rect 28261 4675 28319 4681
rect 28261 4641 28273 4675
rect 28307 4672 28319 4675
rect 28442 4672 28448 4684
rect 28307 4644 28448 4672
rect 28307 4641 28319 4644
rect 28261 4635 28319 4641
rect 28442 4632 28448 4644
rect 28500 4632 28506 4684
rect 28718 4632 28724 4684
rect 28776 4672 28782 4684
rect 28776 4644 30144 4672
rect 28776 4632 28782 4644
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4604 27859 4607
rect 28123 4607 28181 4613
rect 27847 4576 27881 4604
rect 27847 4573 27859 4576
rect 27801 4567 27859 4573
rect 28123 4573 28135 4607
rect 28169 4604 28181 4607
rect 28350 4604 28356 4616
rect 28169 4576 28356 4604
rect 28169 4573 28181 4576
rect 28123 4567 28181 4573
rect 28350 4564 28356 4576
rect 28408 4604 28414 4616
rect 28905 4607 28963 4613
rect 28905 4604 28917 4607
rect 28408 4576 28917 4604
rect 28408 4564 28414 4576
rect 28905 4573 28917 4576
rect 28951 4573 28963 4607
rect 28905 4567 28963 4573
rect 29089 4607 29147 4613
rect 29089 4573 29101 4607
rect 29135 4573 29147 4607
rect 29089 4567 29147 4573
rect 25648 4508 25912 4536
rect 25648 4496 25654 4508
rect 24176 4440 24624 4468
rect 24176 4428 24182 4440
rect 25682 4428 25688 4480
rect 25740 4428 25746 4480
rect 25884 4468 25912 4508
rect 25958 4496 25964 4548
rect 26016 4536 26022 4548
rect 26053 4539 26111 4545
rect 26053 4536 26065 4539
rect 26016 4508 26065 4536
rect 26016 4496 26022 4508
rect 26053 4505 26065 4508
rect 26099 4505 26111 4539
rect 26053 4499 26111 4505
rect 26326 4496 26332 4548
rect 26384 4496 26390 4548
rect 27614 4496 27620 4548
rect 27672 4536 27678 4548
rect 28997 4539 29055 4545
rect 28997 4536 29009 4539
rect 27672 4508 29009 4536
rect 27672 4496 27678 4508
rect 28997 4505 29009 4508
rect 29043 4505 29055 4539
rect 28997 4499 29055 4505
rect 26344 4468 26372 4496
rect 29104 4480 29132 4567
rect 29270 4564 29276 4616
rect 29328 4564 29334 4616
rect 30116 4604 30144 4644
rect 30190 4632 30196 4684
rect 30248 4672 30254 4684
rect 30653 4675 30711 4681
rect 30653 4672 30665 4675
rect 30248 4644 30665 4672
rect 30248 4632 30254 4644
rect 30653 4641 30665 4644
rect 30699 4672 30711 4675
rect 31386 4672 31392 4684
rect 30699 4644 31392 4672
rect 30699 4641 30711 4644
rect 30653 4635 30711 4641
rect 31386 4632 31392 4644
rect 31444 4672 31450 4684
rect 31481 4675 31539 4681
rect 31481 4672 31493 4675
rect 31444 4644 31493 4672
rect 31444 4632 31450 4644
rect 31481 4641 31493 4644
rect 31527 4641 31539 4675
rect 31481 4635 31539 4641
rect 31570 4632 31576 4684
rect 31628 4672 31634 4684
rect 32033 4675 32091 4681
rect 32033 4672 32045 4675
rect 31628 4644 32045 4672
rect 31628 4632 31634 4644
rect 32033 4641 32045 4644
rect 32079 4641 32091 4675
rect 32033 4635 32091 4641
rect 32309 4675 32367 4681
rect 32309 4641 32321 4675
rect 32355 4672 32367 4675
rect 34072 4672 34100 4700
rect 36556 4684 36584 4712
rect 37918 4700 37924 4712
rect 37976 4700 37982 4752
rect 39592 4740 39620 4780
rect 40586 4768 40592 4780
rect 40644 4768 40650 4820
rect 41782 4768 41788 4820
rect 41840 4768 41846 4820
rect 42242 4768 42248 4820
rect 42300 4808 42306 4820
rect 42886 4808 42892 4820
rect 42300 4780 42892 4808
rect 42300 4768 42306 4780
rect 42886 4768 42892 4780
rect 42944 4768 42950 4820
rect 42978 4768 42984 4820
rect 43036 4808 43042 4820
rect 44082 4808 44088 4820
rect 43036 4780 44088 4808
rect 43036 4768 43042 4780
rect 44082 4768 44088 4780
rect 44140 4808 44146 4820
rect 44545 4811 44603 4817
rect 44545 4808 44557 4811
rect 44140 4780 44557 4808
rect 44140 4768 44146 4780
rect 44545 4777 44557 4780
rect 44591 4777 44603 4811
rect 44545 4771 44603 4777
rect 39850 4740 39856 4752
rect 38028 4712 39620 4740
rect 39776 4712 39856 4740
rect 32355 4644 34100 4672
rect 34333 4675 34391 4681
rect 32355 4641 32367 4644
rect 32309 4635 32367 4641
rect 34333 4641 34345 4675
rect 34379 4672 34391 4675
rect 34422 4672 34428 4684
rect 34379 4644 34428 4672
rect 34379 4641 34391 4644
rect 34333 4635 34391 4641
rect 34422 4632 34428 4644
rect 34480 4632 34486 4684
rect 36354 4632 36360 4684
rect 36412 4632 36418 4684
rect 36538 4632 36544 4684
rect 36596 4632 36602 4684
rect 36998 4632 37004 4684
rect 37056 4672 37062 4684
rect 37277 4675 37335 4681
rect 37277 4672 37289 4675
rect 37056 4644 37289 4672
rect 37056 4632 37062 4644
rect 37277 4641 37289 4644
rect 37323 4641 37335 4675
rect 37277 4635 37335 4641
rect 30116 4576 30236 4604
rect 29825 4539 29883 4545
rect 29825 4505 29837 4539
rect 29871 4536 29883 4539
rect 29871 4508 30144 4536
rect 29871 4505 29883 4508
rect 29825 4499 29883 4505
rect 25884 4440 26372 4468
rect 26786 4428 26792 4480
rect 26844 4468 26850 4480
rect 28537 4471 28595 4477
rect 28537 4468 28549 4471
rect 26844 4440 28549 4468
rect 26844 4428 26850 4440
rect 28537 4437 28549 4440
rect 28583 4437 28595 4471
rect 28537 4431 28595 4437
rect 29086 4428 29092 4480
rect 29144 4468 29150 4480
rect 30116 4477 30144 4508
rect 29365 4471 29423 4477
rect 29365 4468 29377 4471
rect 29144 4440 29377 4468
rect 29144 4428 29150 4440
rect 29365 4437 29377 4440
rect 29411 4437 29423 4471
rect 29365 4431 29423 4437
rect 30101 4471 30159 4477
rect 30101 4437 30113 4471
rect 30147 4437 30159 4471
rect 30208 4468 30236 4576
rect 30484 4576 31754 4604
rect 30484 4545 30512 4576
rect 30469 4539 30527 4545
rect 30469 4505 30481 4539
rect 30515 4505 30527 4539
rect 30469 4499 30527 4505
rect 30561 4539 30619 4545
rect 30561 4505 30573 4539
rect 30607 4536 30619 4539
rect 30834 4536 30840 4548
rect 30607 4508 30840 4536
rect 30607 4505 30619 4508
rect 30561 4499 30619 4505
rect 30834 4496 30840 4508
rect 30892 4496 30898 4548
rect 31726 4536 31754 4576
rect 34054 4564 34060 4616
rect 34112 4564 34118 4616
rect 36078 4604 36084 4616
rect 35466 4576 36084 4604
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 36265 4607 36323 4613
rect 36265 4573 36277 4607
rect 36311 4604 36323 4607
rect 36906 4604 36912 4616
rect 36311 4576 36912 4604
rect 36311 4573 36323 4576
rect 36265 4567 36323 4573
rect 36906 4564 36912 4576
rect 36964 4564 36970 4616
rect 37093 4607 37151 4613
rect 37093 4573 37105 4607
rect 37139 4604 37151 4607
rect 37182 4604 37188 4616
rect 37139 4576 37188 4604
rect 37139 4573 37151 4576
rect 37093 4567 37151 4573
rect 37182 4564 37188 4576
rect 37240 4564 37246 4616
rect 38028 4604 38056 4712
rect 39206 4672 39212 4684
rect 38396 4644 39212 4672
rect 38396 4613 38424 4644
rect 39206 4632 39212 4644
rect 39264 4632 39270 4684
rect 39776 4681 39804 4712
rect 39850 4700 39856 4712
rect 39908 4740 39914 4752
rect 40402 4740 40408 4752
rect 39908 4712 40408 4740
rect 39908 4700 39914 4712
rect 40402 4700 40408 4712
rect 40460 4740 40466 4752
rect 41141 4743 41199 4749
rect 40460 4712 40632 4740
rect 40460 4700 40466 4712
rect 39761 4675 39819 4681
rect 39761 4641 39773 4675
rect 39807 4641 39819 4675
rect 40034 4672 40040 4684
rect 39761 4635 39819 4641
rect 39868 4644 40040 4672
rect 37292 4576 38056 4604
rect 38381 4607 38439 4613
rect 31312 4508 31524 4536
rect 31726 4508 32720 4536
rect 30650 4468 30656 4480
rect 30208 4440 30656 4468
rect 30101 4431 30159 4437
rect 30650 4428 30656 4440
rect 30708 4428 30714 4480
rect 30926 4428 30932 4480
rect 30984 4428 30990 4480
rect 31312 4477 31340 4508
rect 31297 4471 31355 4477
rect 31297 4437 31309 4471
rect 31343 4437 31355 4471
rect 31297 4431 31355 4437
rect 31386 4428 31392 4480
rect 31444 4428 31450 4480
rect 31496 4468 31524 4508
rect 32582 4468 32588 4480
rect 31496 4440 32588 4468
rect 32582 4428 32588 4440
rect 32640 4428 32646 4480
rect 32692 4468 32720 4508
rect 33042 4496 33048 4548
rect 33100 4496 33106 4548
rect 35710 4496 35716 4548
rect 35768 4536 35774 4548
rect 37292 4536 37320 4576
rect 38381 4573 38393 4607
rect 38427 4573 38439 4607
rect 38381 4567 38439 4573
rect 39025 4607 39083 4613
rect 39025 4573 39037 4607
rect 39071 4604 39083 4607
rect 39577 4607 39635 4613
rect 39071 4576 39252 4604
rect 39071 4573 39083 4576
rect 39025 4567 39083 4573
rect 35768 4508 37320 4536
rect 35768 4496 35774 4508
rect 37734 4496 37740 4548
rect 37792 4496 37798 4548
rect 35342 4468 35348 4480
rect 32692 4440 35348 4468
rect 35342 4428 35348 4440
rect 35400 4428 35406 4480
rect 35802 4428 35808 4480
rect 35860 4468 35866 4480
rect 39224 4477 39252 4576
rect 39577 4573 39589 4607
rect 39623 4604 39635 4607
rect 39868 4604 39896 4644
rect 40034 4632 40040 4644
rect 40092 4632 40098 4684
rect 40604 4681 40632 4712
rect 41141 4709 41153 4743
rect 41187 4740 41199 4743
rect 42260 4740 42288 4768
rect 41187 4712 42288 4740
rect 42904 4740 42932 4768
rect 43257 4743 43315 4749
rect 43257 4740 43269 4743
rect 42904 4712 43269 4740
rect 41187 4709 41199 4712
rect 41141 4703 41199 4709
rect 43257 4709 43269 4712
rect 43303 4740 43315 4743
rect 43625 4743 43683 4749
rect 43625 4740 43637 4743
rect 43303 4712 43637 4740
rect 43303 4709 43315 4712
rect 43257 4703 43315 4709
rect 43625 4709 43637 4712
rect 43671 4709 43683 4743
rect 43625 4703 43683 4709
rect 43990 4700 43996 4752
rect 44048 4700 44054 4752
rect 40589 4675 40647 4681
rect 40589 4641 40601 4675
rect 40635 4641 40647 4675
rect 40589 4635 40647 4641
rect 42518 4632 42524 4684
rect 42576 4672 42582 4684
rect 43438 4672 43444 4684
rect 42576 4644 43444 4672
rect 42576 4632 42582 4644
rect 43438 4632 43444 4644
rect 43496 4672 43502 4684
rect 44913 4675 44971 4681
rect 44913 4672 44925 4675
rect 43496 4644 44925 4672
rect 43496 4632 43502 4644
rect 44913 4641 44925 4644
rect 44959 4641 44971 4675
rect 44913 4635 44971 4641
rect 39623 4576 39896 4604
rect 39623 4573 39635 4576
rect 39577 4567 39635 4573
rect 39942 4564 39948 4616
rect 40000 4604 40006 4616
rect 40405 4607 40463 4613
rect 40405 4604 40417 4607
rect 40000 4576 40417 4604
rect 40000 4564 40006 4576
rect 40405 4573 40417 4576
rect 40451 4573 40463 4607
rect 40405 4567 40463 4573
rect 39669 4539 39727 4545
rect 39669 4505 39681 4539
rect 39715 4536 39727 4539
rect 40862 4536 40868 4548
rect 39715 4508 40868 4536
rect 39715 4505 39727 4508
rect 39669 4499 39727 4505
rect 40862 4496 40868 4508
rect 40920 4496 40926 4548
rect 41506 4496 41512 4548
rect 41564 4536 41570 4548
rect 42521 4539 42579 4545
rect 42521 4536 42533 4539
rect 41564 4508 42533 4536
rect 41564 4496 41570 4508
rect 42521 4505 42533 4508
rect 42567 4505 42579 4539
rect 42521 4499 42579 4505
rect 37185 4471 37243 4477
rect 37185 4468 37197 4471
rect 35860 4440 37197 4468
rect 35860 4428 35866 4440
rect 37185 4437 37197 4440
rect 37231 4437 37243 4471
rect 37185 4431 37243 4437
rect 39209 4471 39267 4477
rect 39209 4437 39221 4471
rect 39255 4437 39267 4471
rect 39209 4431 39267 4437
rect 40034 4428 40040 4480
rect 40092 4428 40098 4480
rect 40494 4428 40500 4480
rect 40552 4428 40558 4480
rect 460 4378 45540 4400
rect 460 4326 6070 4378
rect 6122 4326 6134 4378
rect 6186 4326 6198 4378
rect 6250 4326 6262 4378
rect 6314 4326 6326 4378
rect 6378 4326 11070 4378
rect 11122 4326 11134 4378
rect 11186 4326 11198 4378
rect 11250 4326 11262 4378
rect 11314 4326 11326 4378
rect 11378 4326 16070 4378
rect 16122 4326 16134 4378
rect 16186 4326 16198 4378
rect 16250 4326 16262 4378
rect 16314 4326 16326 4378
rect 16378 4326 21070 4378
rect 21122 4326 21134 4378
rect 21186 4326 21198 4378
rect 21250 4326 21262 4378
rect 21314 4326 21326 4378
rect 21378 4326 26070 4378
rect 26122 4326 26134 4378
rect 26186 4326 26198 4378
rect 26250 4326 26262 4378
rect 26314 4326 26326 4378
rect 26378 4326 31070 4378
rect 31122 4326 31134 4378
rect 31186 4326 31198 4378
rect 31250 4326 31262 4378
rect 31314 4326 31326 4378
rect 31378 4326 36070 4378
rect 36122 4326 36134 4378
rect 36186 4326 36198 4378
rect 36250 4326 36262 4378
rect 36314 4326 36326 4378
rect 36378 4326 41070 4378
rect 41122 4326 41134 4378
rect 41186 4326 41198 4378
rect 41250 4326 41262 4378
rect 41314 4326 41326 4378
rect 41378 4326 45540 4378
rect 460 4304 45540 4326
rect 4706 4264 4712 4276
rect 3804 4236 4712 4264
rect 1486 4196 1492 4208
rect 1228 4168 1492 4196
rect 1228 4137 1256 4168
rect 1486 4156 1492 4168
rect 1544 4156 1550 4208
rect 1213 4131 1271 4137
rect 1213 4097 1225 4131
rect 1259 4097 1271 4131
rect 1213 4091 1271 4097
rect 2590 4088 2596 4140
rect 2648 4088 2654 4140
rect 3804 4128 3832 4236
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 4338 4196 4344 4208
rect 4111 4168 4344 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 4448 4196 4476 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5592 4236 5733 4264
rect 5592 4224 5598 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 5902 4224 5908 4276
rect 5960 4224 5966 4276
rect 6932 4236 8340 4264
rect 4448 4168 4554 4196
rect 3620 4100 3832 4128
rect 1489 4063 1547 4069
rect 1489 4060 1501 4063
rect 1320 4032 1501 4060
rect 934 3952 940 4004
rect 992 3992 998 4004
rect 1320 3992 1348 4032
rect 1489 4029 1501 4032
rect 1535 4029 1547 4063
rect 1489 4023 1547 4029
rect 2608 4060 2636 4088
rect 3620 4069 3648 4100
rect 5074 4088 5080 4140
rect 5132 4088 5138 4140
rect 5920 4137 5948 4224
rect 6932 4196 6960 4236
rect 8312 4208 8340 4236
rect 9122 4224 9128 4276
rect 9180 4224 9186 4276
rect 9582 4224 9588 4276
rect 9640 4224 9646 4276
rect 11698 4224 11704 4276
rect 11756 4224 11762 4276
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 12584 4236 14105 4264
rect 12584 4224 12590 4236
rect 14093 4233 14105 4236
rect 14139 4264 14151 4267
rect 14274 4264 14280 4276
rect 14139 4236 14280 4264
rect 14139 4233 14151 4236
rect 14093 4227 14151 4233
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14424 4236 15025 4264
rect 14424 4224 14430 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 22278 4264 22284 4276
rect 15804 4236 22284 4264
rect 15804 4224 15810 4236
rect 22278 4224 22284 4236
rect 22336 4224 22342 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 23109 4267 23167 4273
rect 23109 4264 23121 4267
rect 22428 4236 23121 4264
rect 22428 4224 22434 4236
rect 23109 4233 23121 4236
rect 23155 4233 23167 4267
rect 23109 4227 23167 4233
rect 23474 4224 23480 4276
rect 23532 4224 23538 4276
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24305 4267 24363 4273
rect 24305 4264 24317 4267
rect 24176 4236 24317 4264
rect 24176 4224 24182 4236
rect 24305 4233 24317 4236
rect 24351 4264 24363 4267
rect 25590 4264 25596 4276
rect 24351 4236 25596 4264
rect 24351 4233 24363 4236
rect 24305 4227 24363 4233
rect 25590 4224 25596 4236
rect 25648 4224 25654 4276
rect 26418 4224 26424 4276
rect 26476 4224 26482 4276
rect 26694 4224 26700 4276
rect 26752 4264 26758 4276
rect 27614 4264 27620 4276
rect 26752 4236 27620 4264
rect 26752 4224 26758 4236
rect 6564 4168 6960 4196
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 6564 4137 6592 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9140 4196 9168 4224
rect 8352 4168 9168 4196
rect 9217 4199 9275 4205
rect 8352 4156 8358 4168
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6512 4100 6561 4128
rect 6512 4088 6518 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 7926 4088 7932 4140
rect 7984 4088 7990 4140
rect 8956 4137 8984 4168
rect 9217 4165 9229 4199
rect 9263 4196 9275 4199
rect 9600 4196 9628 4224
rect 11716 4196 11744 4224
rect 9263 4168 9628 4196
rect 11440 4168 11744 4196
rect 11793 4199 11851 4205
rect 9263 4165 9275 4168
rect 9217 4159 9275 4165
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 3605 4063 3663 4069
rect 3605 4060 3617 4063
rect 2608 4032 3617 4060
rect 992 3964 1348 3992
rect 992 3952 998 3964
rect 1121 3927 1179 3933
rect 1121 3893 1133 3927
rect 1167 3924 1179 3927
rect 2608 3924 2636 4032
rect 3605 4029 3617 4032
rect 3651 4029 3663 4063
rect 3605 4023 3663 4029
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 5092 4060 5120 4088
rect 3835 4032 5120 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 3804 3992 3832 4023
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5408 4032 5549 4060
rect 5408 4020 5414 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 3384 3964 3832 3992
rect 3384 3952 3390 3964
rect 1167 3896 2636 3924
rect 1167 3893 1179 3896
rect 1121 3887 1179 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2832 3896 2973 3924
rect 2832 3884 2838 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 7944 3924 7972 4088
rect 8864 3992 8892 4091
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 11440 4137 11468 4168
rect 11793 4165 11805 4199
rect 11839 4196 11851 4199
rect 12066 4196 12072 4208
rect 11839 4168 12072 4196
rect 11839 4165 11851 4168
rect 11793 4159 11851 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 15930 4196 15936 4208
rect 15028 4168 15936 4196
rect 11425 4131 11483 4137
rect 10284 4100 10350 4128
rect 10284 4088 10290 4100
rect 11425 4097 11437 4131
rect 11471 4097 11483 4131
rect 11425 4091 11483 4097
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 13541 4131 13599 4137
rect 12952 4100 13492 4128
rect 12952 4088 12958 4100
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 11164 3992 11192 4023
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 13262 4060 13268 4072
rect 11624 4032 13268 4060
rect 11624 3992 11652 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 8864 3964 9076 3992
rect 11164 3964 11652 3992
rect 9048 3936 9076 3964
rect 6696 3896 7972 3924
rect 8297 3927 8355 3933
rect 6696 3884 6702 3896
rect 8297 3893 8309 3927
rect 8343 3924 8355 3927
rect 8386 3924 8392 3936
rect 8343 3896 8392 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 8938 3924 8944 3936
rect 8711 3896 8944 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9030 3884 9036 3936
rect 9088 3884 9094 3936
rect 10686 3884 10692 3936
rect 10744 3884 10750 3936
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 12986 3924 12992 3936
rect 12584 3896 12992 3924
rect 12584 3884 12590 3896
rect 12986 3884 12992 3896
rect 13044 3924 13050 3936
rect 13265 3927 13323 3933
rect 13265 3924 13277 3927
rect 13044 3896 13277 3924
rect 13044 3884 13050 3896
rect 13265 3893 13277 3896
rect 13311 3893 13323 3927
rect 13265 3887 13323 3893
rect 13354 3884 13360 3936
rect 13412 3884 13418 3936
rect 13464 3924 13492 4100
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 14185 4131 14243 4137
rect 13587 4100 13768 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13740 4001 13768 4100
rect 14185 4097 14197 4131
rect 14231 4128 14243 4131
rect 14458 4128 14464 4140
rect 14231 4100 14464 4128
rect 14231 4097 14243 4100
rect 14185 4091 14243 4097
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15028 4128 15056 4168
rect 15930 4156 15936 4168
rect 15988 4156 15994 4208
rect 16574 4196 16580 4208
rect 16408 4168 16580 4196
rect 14967 4100 15056 4128
rect 15105 4131 15163 4137
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15105 4097 15117 4131
rect 15151 4128 15163 4131
rect 15194 4128 15200 4140
rect 15151 4100 15200 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16206 4128 16212 4140
rect 15887 4100 16212 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 16408 4137 16436 4168
rect 16574 4156 16580 4168
rect 16632 4196 16638 4208
rect 16758 4196 16764 4208
rect 16632 4168 16764 4196
rect 16632 4156 16638 4168
rect 16758 4156 16764 4168
rect 16816 4156 16822 4208
rect 17126 4156 17132 4208
rect 17184 4156 17190 4208
rect 19058 4156 19064 4208
rect 19116 4196 19122 4208
rect 20165 4199 20223 4205
rect 19116 4168 19932 4196
rect 19116 4156 19122 4168
rect 16393 4131 16451 4137
rect 16393 4097 16405 4131
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19904 4128 19932 4168
rect 20165 4165 20177 4199
rect 20211 4196 20223 4199
rect 20346 4196 20352 4208
rect 20211 4168 20352 4196
rect 20211 4165 20223 4168
rect 20165 4159 20223 4165
rect 20346 4156 20352 4168
rect 20404 4156 20410 4208
rect 23492 4196 23520 4224
rect 23492 4168 24716 4196
rect 20070 4128 20076 4140
rect 19904 4100 20076 4128
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20438 4128 20444 4140
rect 20303 4100 20444 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 20990 4128 20996 4140
rect 20588 4100 20996 4128
rect 20588 4088 20594 4100
rect 20990 4088 20996 4100
rect 21048 4128 21054 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 21048 4100 21281 4128
rect 21048 4088 21054 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 23106 4128 23112 4140
rect 22678 4100 23112 4128
rect 21269 4091 21327 4097
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4128 23535 4131
rect 23842 4128 23848 4140
rect 23523 4100 23848 4128
rect 23523 4097 23535 4100
rect 23477 4091 23535 4097
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 24302 4088 24308 4140
rect 24360 4088 24366 4140
rect 24394 4088 24400 4140
rect 24452 4128 24458 4140
rect 24581 4131 24639 4137
rect 24581 4128 24593 4131
rect 24452 4100 24593 4128
rect 24452 4088 24458 4100
rect 24581 4097 24593 4100
rect 24627 4097 24639 4131
rect 24688 4128 24716 4168
rect 25130 4156 25136 4208
rect 25188 4156 25194 4208
rect 25317 4199 25375 4205
rect 25317 4165 25329 4199
rect 25363 4196 25375 4199
rect 25866 4196 25872 4208
rect 25363 4168 25872 4196
rect 25363 4165 25375 4168
rect 25317 4159 25375 4165
rect 25866 4156 25872 4168
rect 25924 4156 25930 4208
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 24688 4100 25053 4128
rect 24581 4091 24639 4097
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25041 4091 25099 4097
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14056 4032 14289 4060
rect 14056 4020 14062 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 16298 4020 16304 4072
rect 16356 4020 16362 4072
rect 16666 4020 16672 4072
rect 16724 4020 16730 4072
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17736 4032 18153 4060
rect 17736 4020 17742 4032
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18141 4023 18199 4029
rect 19061 4063 19119 4069
rect 19061 4029 19073 4063
rect 19107 4060 19119 4063
rect 19150 4060 19156 4072
rect 19107 4032 19156 4060
rect 19107 4029 19119 4032
rect 19061 4023 19119 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 19567 4032 20361 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 20349 4029 20361 4032
rect 20395 4060 20407 4063
rect 20714 4060 20720 4072
rect 20395 4032 20720 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 21542 4020 21548 4072
rect 21600 4020 21606 4072
rect 23569 4063 23627 4069
rect 23569 4060 23581 4063
rect 23032 4032 23581 4060
rect 13725 3995 13783 4001
rect 13725 3961 13737 3995
rect 13771 3961 13783 3995
rect 13725 3955 13783 3961
rect 13906 3952 13912 4004
rect 13964 3992 13970 4004
rect 18693 3995 18751 4001
rect 13964 3964 16344 3992
rect 13964 3952 13970 3964
rect 14090 3924 14096 3936
rect 13464 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3924 14154 3936
rect 14829 3927 14887 3933
rect 14829 3924 14841 3927
rect 14148 3896 14841 3924
rect 14148 3884 14154 3896
rect 14829 3893 14841 3896
rect 14875 3924 14887 3927
rect 15473 3927 15531 3933
rect 15473 3924 15485 3927
rect 14875 3896 15485 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15473 3893 15485 3896
rect 15519 3924 15531 3927
rect 15838 3924 15844 3936
rect 15519 3896 15844 3924
rect 15519 3893 15531 3896
rect 15473 3887 15531 3893
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 16316 3924 16344 3964
rect 18693 3961 18705 3995
rect 18739 3992 18751 3995
rect 18739 3964 21036 3992
rect 18739 3961 18751 3964
rect 18693 3955 18751 3961
rect 18708 3924 18736 3955
rect 16316 3896 18736 3924
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 19797 3927 19855 3933
rect 19797 3924 19809 3927
rect 19760 3896 19809 3924
rect 19760 3884 19766 3896
rect 19797 3893 19809 3896
rect 19843 3893 19855 3927
rect 21008 3924 21036 3964
rect 22186 3924 22192 3936
rect 21008 3896 22192 3924
rect 19797 3887 19855 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 23032 3933 23060 4032
rect 23569 4029 23581 4032
rect 23615 4029 23627 4063
rect 23569 4023 23627 4029
rect 23753 4063 23811 4069
rect 23753 4029 23765 4063
rect 23799 4060 23811 4063
rect 23934 4060 23940 4072
rect 23799 4032 23940 4060
rect 23799 4029 23811 4032
rect 23753 4023 23811 4029
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 24320 4060 24348 4088
rect 24857 4063 24915 4069
rect 24857 4060 24869 4063
rect 24320 4032 24869 4060
rect 24857 4029 24869 4032
rect 24903 4029 24915 4063
rect 24857 4023 24915 4029
rect 23106 3952 23112 4004
rect 23164 3992 23170 4004
rect 25148 3992 25176 4156
rect 25682 4088 25688 4140
rect 25740 4088 25746 4140
rect 25774 4088 25780 4140
rect 25832 4088 25838 4140
rect 25958 4020 25964 4072
rect 26016 4060 26022 4072
rect 26329 4063 26387 4069
rect 26329 4060 26341 4063
rect 26016 4032 26341 4060
rect 26016 4020 26022 4032
rect 26329 4029 26341 4032
rect 26375 4029 26387 4063
rect 26329 4023 26387 4029
rect 23164 3964 25176 3992
rect 25225 3995 25283 4001
rect 23164 3952 23170 3964
rect 25225 3961 25237 3995
rect 25271 3992 25283 3995
rect 25866 3992 25872 4004
rect 25271 3964 25872 3992
rect 25271 3961 25283 3964
rect 25225 3955 25283 3961
rect 25866 3952 25872 3964
rect 25924 3992 25930 4004
rect 26436 3992 26464 4224
rect 27474 4205 27502 4236
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 28258 4224 28264 4276
rect 28316 4264 28322 4276
rect 28316 4236 29040 4264
rect 28316 4224 28322 4236
rect 27459 4199 27517 4205
rect 27459 4165 27471 4199
rect 27505 4165 27517 4199
rect 27459 4159 27517 4165
rect 27706 4156 27712 4208
rect 27764 4156 27770 4208
rect 27925 4199 27983 4205
rect 27925 4165 27937 4199
rect 27971 4196 27983 4199
rect 28074 4196 28080 4208
rect 27971 4168 28080 4196
rect 27971 4165 27983 4168
rect 27925 4159 27983 4165
rect 28074 4156 28080 4168
rect 28132 4196 28138 4208
rect 28718 4196 28724 4208
rect 28132 4168 28724 4196
rect 28132 4156 28138 4168
rect 26513 4131 26571 4137
rect 26513 4097 26525 4131
rect 26559 4097 26571 4131
rect 26513 4091 26571 4097
rect 26528 4060 26556 4091
rect 26694 4088 26700 4140
rect 26752 4088 26758 4140
rect 26789 4131 26847 4137
rect 26789 4097 26801 4131
rect 26835 4128 26847 4131
rect 27157 4131 27215 4137
rect 26835 4100 27108 4128
rect 26835 4097 26847 4100
rect 26789 4091 26847 4097
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26528 4032 26985 4060
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 25924 3964 26464 3992
rect 25924 3952 25930 3964
rect 26602 3952 26608 4004
rect 26660 3952 26666 4004
rect 27080 3992 27108 4100
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27172 4060 27200 4091
rect 27246 4088 27252 4140
rect 27304 4088 27310 4140
rect 27338 4088 27344 4140
rect 27396 4088 27402 4140
rect 27724 4128 27752 4156
rect 28166 4128 28172 4140
rect 27724 4100 28172 4128
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 28460 4137 28488 4168
rect 28718 4156 28724 4168
rect 28776 4156 28782 4208
rect 29012 4205 29040 4236
rect 29178 4224 29184 4276
rect 29236 4264 29242 4276
rect 29638 4264 29644 4276
rect 29236 4236 29644 4264
rect 29236 4224 29242 4236
rect 29638 4224 29644 4236
rect 29696 4224 29702 4276
rect 30926 4264 30932 4276
rect 30760 4236 30932 4264
rect 30760 4205 30788 4236
rect 30926 4224 30932 4236
rect 30984 4224 30990 4276
rect 31018 4224 31024 4276
rect 31076 4224 31082 4276
rect 33318 4224 33324 4276
rect 33376 4264 33382 4276
rect 39853 4267 39911 4273
rect 33376 4236 33824 4264
rect 33376 4224 33382 4236
rect 28997 4199 29055 4205
rect 28997 4196 29009 4199
rect 28920 4168 29009 4196
rect 28445 4131 28503 4137
rect 28445 4097 28457 4131
rect 28491 4097 28503 4131
rect 28445 4091 28503 4097
rect 28626 4088 28632 4140
rect 28684 4128 28690 4140
rect 28813 4131 28871 4137
rect 28813 4128 28825 4131
rect 28684 4100 28825 4128
rect 28684 4088 28690 4100
rect 28813 4097 28825 4100
rect 28859 4097 28871 4131
rect 28813 4091 28871 4097
rect 27522 4060 27528 4072
rect 27172 4032 27528 4060
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 27617 4063 27675 4069
rect 27617 4029 27629 4063
rect 27663 4060 27675 4063
rect 27982 4060 27988 4072
rect 27663 4032 27988 4060
rect 27663 4029 27675 4032
rect 27617 4023 27675 4029
rect 27982 4020 27988 4032
rect 28040 4020 28046 4072
rect 28721 4063 28779 4069
rect 28721 4029 28733 4063
rect 28767 4060 28779 4063
rect 28920 4060 28948 4168
rect 28997 4165 29009 4168
rect 29043 4165 29055 4199
rect 30745 4199 30803 4205
rect 28997 4159 29055 4165
rect 29656 4168 29960 4196
rect 29270 4088 29276 4140
rect 29328 4128 29334 4140
rect 29656 4128 29684 4168
rect 29328 4100 29684 4128
rect 29328 4088 29334 4100
rect 29730 4088 29736 4140
rect 29788 4088 29794 4140
rect 29825 4131 29883 4137
rect 29825 4097 29837 4131
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 28767 4032 28948 4060
rect 29181 4063 29239 4069
rect 28767 4029 28779 4032
rect 28721 4023 28779 4029
rect 29181 4029 29193 4063
rect 29227 4060 29239 4063
rect 29362 4060 29368 4072
rect 29227 4032 29368 4060
rect 29227 4029 29239 4032
rect 29181 4023 29239 4029
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 28077 3995 28135 4001
rect 28077 3992 28089 3995
rect 27080 3964 28089 3992
rect 28077 3961 28089 3964
rect 28123 3961 28135 3995
rect 28077 3955 28135 3961
rect 28261 3995 28319 4001
rect 28261 3961 28273 3995
rect 28307 3992 28319 3995
rect 29840 3992 29868 4091
rect 29932 4060 29960 4168
rect 30745 4165 30757 4199
rect 30791 4165 30803 4199
rect 30745 4159 30803 4165
rect 31665 4199 31723 4205
rect 31665 4165 31677 4199
rect 31711 4196 31723 4199
rect 32398 4196 32404 4208
rect 31711 4168 32404 4196
rect 31711 4165 31723 4168
rect 31665 4159 31723 4165
rect 32398 4156 32404 4168
rect 32456 4156 32462 4208
rect 33796 4205 33824 4236
rect 33888 4236 39712 4264
rect 33229 4199 33287 4205
rect 33229 4165 33241 4199
rect 33275 4196 33287 4199
rect 33781 4199 33839 4205
rect 33275 4168 33732 4196
rect 33275 4165 33287 4168
rect 33229 4159 33287 4165
rect 30101 4131 30159 4137
rect 30101 4097 30113 4131
rect 30147 4097 30159 4131
rect 30101 4091 30159 4097
rect 30116 4060 30144 4091
rect 30190 4088 30196 4140
rect 30248 4088 30254 4140
rect 30834 4128 30840 4140
rect 30300 4100 30840 4128
rect 30300 4069 30328 4100
rect 30834 4088 30840 4100
rect 30892 4088 30898 4140
rect 30926 4088 30932 4140
rect 30984 4128 30990 4140
rect 31205 4131 31263 4137
rect 31205 4128 31217 4131
rect 30984 4100 31217 4128
rect 30984 4088 30990 4100
rect 31205 4097 31217 4100
rect 31251 4097 31263 4131
rect 31205 4091 31263 4097
rect 32214 4088 32220 4140
rect 32272 4088 32278 4140
rect 33321 4131 33379 4137
rect 33321 4097 33333 4131
rect 33367 4128 33379 4131
rect 33410 4128 33416 4140
rect 33367 4100 33416 4128
rect 33367 4097 33379 4100
rect 33321 4091 33379 4097
rect 33410 4088 33416 4100
rect 33468 4088 33474 4140
rect 33704 4128 33732 4168
rect 33781 4165 33793 4199
rect 33827 4165 33839 4199
rect 33781 4159 33839 4165
rect 33888 4128 33916 4236
rect 34146 4156 34152 4208
rect 34204 4156 34210 4208
rect 35986 4196 35992 4208
rect 35650 4168 35992 4196
rect 35986 4156 35992 4168
rect 36044 4196 36050 4208
rect 36044 4168 37228 4196
rect 36044 4156 36050 4168
rect 34164 4128 34192 4156
rect 33704 4100 33916 4128
rect 33980 4100 34192 4128
rect 30285 4063 30343 4069
rect 30285 4060 30297 4063
rect 29932 4032 30297 4060
rect 30285 4029 30297 4032
rect 30331 4029 30343 4063
rect 30285 4023 30343 4029
rect 30650 4020 30656 4072
rect 30708 4060 30714 4072
rect 31941 4063 31999 4069
rect 30708 4032 31340 4060
rect 30708 4020 30714 4032
rect 31202 3992 31208 4004
rect 28307 3964 31208 3992
rect 28307 3961 28319 3964
rect 28261 3955 28319 3961
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 23017 3927 23075 3933
rect 23017 3924 23029 3927
rect 22336 3896 23029 3924
rect 22336 3884 22342 3896
rect 23017 3893 23029 3896
rect 23063 3893 23075 3927
rect 23017 3887 23075 3893
rect 24854 3884 24860 3936
rect 24912 3884 24918 3936
rect 25406 3884 25412 3936
rect 25464 3884 25470 3936
rect 25961 3927 26019 3933
rect 25961 3893 25973 3927
rect 26007 3924 26019 3927
rect 26418 3924 26424 3936
rect 26007 3896 26424 3924
rect 26007 3893 26019 3896
rect 25961 3887 26019 3893
rect 26418 3884 26424 3896
rect 26476 3924 26482 3936
rect 26620 3924 26648 3952
rect 26476 3896 26648 3924
rect 26476 3884 26482 3896
rect 27890 3884 27896 3936
rect 27948 3884 27954 3936
rect 28442 3884 28448 3936
rect 28500 3924 28506 3936
rect 28626 3924 28632 3936
rect 28500 3896 28632 3924
rect 28500 3884 28506 3896
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 29365 3927 29423 3933
rect 29365 3893 29377 3927
rect 29411 3924 29423 3927
rect 29454 3924 29460 3936
rect 29411 3896 29460 3924
rect 29411 3893 29423 3896
rect 29365 3887 29423 3893
rect 29454 3884 29460 3896
rect 29512 3884 29518 3936
rect 29546 3884 29552 3936
rect 29604 3884 29610 3936
rect 30006 3884 30012 3936
rect 30064 3884 30070 3936
rect 30377 3927 30435 3933
rect 30377 3893 30389 3927
rect 30423 3924 30435 3927
rect 30466 3924 30472 3936
rect 30423 3896 30472 3924
rect 30423 3893 30435 3896
rect 30377 3887 30435 3893
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 30558 3884 30564 3936
rect 30616 3884 30622 3936
rect 30837 3927 30895 3933
rect 30837 3893 30849 3927
rect 30883 3924 30895 3927
rect 31312 3924 31340 4032
rect 31941 4029 31953 4063
rect 31987 4029 31999 4063
rect 31941 4023 31999 4029
rect 31846 3952 31852 4004
rect 31904 3952 31910 4004
rect 31956 3992 31984 4023
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 33505 4063 33563 4069
rect 33505 4060 33517 4063
rect 33192 4032 33517 4060
rect 33192 4020 33198 4032
rect 33505 4029 33517 4032
rect 33551 4060 33563 4063
rect 33980 4060 34008 4100
rect 35894 4088 35900 4140
rect 35952 4128 35958 4140
rect 36173 4131 36231 4137
rect 36173 4128 36185 4131
rect 35952 4100 36185 4128
rect 35952 4088 35958 4100
rect 36173 4097 36185 4100
rect 36219 4097 36231 4131
rect 37200 4128 37228 4168
rect 37274 4156 37280 4208
rect 37332 4196 37338 4208
rect 38286 4196 38292 4208
rect 37332 4168 38292 4196
rect 37332 4156 37338 4168
rect 37458 4128 37464 4140
rect 37200 4100 37464 4128
rect 36173 4091 36231 4097
rect 37458 4088 37464 4100
rect 37516 4088 37522 4140
rect 38120 4137 38148 4168
rect 38286 4156 38292 4168
rect 38344 4156 38350 4208
rect 39684 4196 39712 4236
rect 39853 4233 39865 4267
rect 39899 4264 39911 4267
rect 39942 4264 39948 4276
rect 39899 4236 39948 4264
rect 39899 4233 39911 4236
rect 39853 4227 39911 4233
rect 39942 4224 39948 4236
rect 40000 4264 40006 4276
rect 40405 4267 40463 4273
rect 40405 4264 40417 4267
rect 40000 4236 40417 4264
rect 40000 4224 40006 4236
rect 40405 4233 40417 4236
rect 40451 4233 40463 4267
rect 40405 4227 40463 4233
rect 40494 4224 40500 4276
rect 40552 4264 40558 4276
rect 40954 4264 40960 4276
rect 40552 4236 40960 4264
rect 40552 4224 40558 4236
rect 40954 4224 40960 4236
rect 41012 4264 41018 4276
rect 41233 4267 41291 4273
rect 41233 4264 41245 4267
rect 41012 4236 41245 4264
rect 41012 4224 41018 4236
rect 41233 4233 41245 4236
rect 41279 4233 41291 4267
rect 41233 4227 41291 4233
rect 41874 4224 41880 4276
rect 41932 4224 41938 4276
rect 41966 4224 41972 4276
rect 42024 4224 42030 4276
rect 42978 4224 42984 4276
rect 43036 4264 43042 4276
rect 43073 4267 43131 4273
rect 43073 4264 43085 4267
rect 43036 4236 43085 4264
rect 43036 4224 43042 4236
rect 43073 4233 43085 4236
rect 43119 4233 43131 4267
rect 43073 4227 43131 4233
rect 43438 4224 43444 4276
rect 43496 4224 43502 4276
rect 43901 4267 43959 4273
rect 43901 4233 43913 4267
rect 43947 4264 43959 4267
rect 43990 4264 43996 4276
rect 43947 4236 43996 4264
rect 43947 4233 43959 4236
rect 43901 4227 43959 4233
rect 43990 4224 43996 4236
rect 44048 4264 44054 4276
rect 44545 4267 44603 4273
rect 44545 4264 44557 4267
rect 44048 4236 44557 4264
rect 44048 4224 44054 4236
rect 44545 4233 44557 4236
rect 44591 4264 44603 4267
rect 44726 4264 44732 4276
rect 44591 4236 44732 4264
rect 44591 4233 44603 4236
rect 44545 4227 44603 4233
rect 44726 4224 44732 4236
rect 44784 4264 44790 4276
rect 44913 4267 44971 4273
rect 44913 4264 44925 4267
rect 44784 4236 44925 4264
rect 44784 4224 44790 4236
rect 44913 4233 44925 4236
rect 44959 4233 44971 4267
rect 44913 4227 44971 4233
rect 41141 4199 41199 4205
rect 39684 4168 40448 4196
rect 38105 4131 38163 4137
rect 38105 4097 38117 4131
rect 38151 4097 38163 4131
rect 38105 4091 38163 4097
rect 39390 4088 39396 4140
rect 39448 4128 39454 4140
rect 40218 4128 40224 4140
rect 39448 4100 40224 4128
rect 39448 4088 39454 4100
rect 40218 4088 40224 4100
rect 40276 4088 40282 4140
rect 40310 4088 40316 4140
rect 40368 4088 40374 4140
rect 40420 4128 40448 4168
rect 41141 4165 41153 4199
rect 41187 4196 41199 4199
rect 41782 4196 41788 4208
rect 41187 4168 41788 4196
rect 41187 4165 41199 4168
rect 41141 4159 41199 4165
rect 41782 4156 41788 4168
rect 41840 4156 41846 4208
rect 41892 4196 41920 4224
rect 42337 4199 42395 4205
rect 42337 4196 42349 4199
rect 41892 4168 42349 4196
rect 42337 4165 42349 4168
rect 42383 4196 42395 4199
rect 42705 4199 42763 4205
rect 42705 4196 42717 4199
rect 42383 4168 42717 4196
rect 42383 4165 42395 4168
rect 42337 4159 42395 4165
rect 42705 4165 42717 4168
rect 42751 4165 42763 4199
rect 43456 4196 43484 4224
rect 44177 4199 44235 4205
rect 44177 4196 44189 4199
rect 43456 4168 44189 4196
rect 42705 4159 42763 4165
rect 44177 4165 44189 4168
rect 44223 4165 44235 4199
rect 44177 4159 44235 4165
rect 40420 4100 40632 4128
rect 33551 4032 34008 4060
rect 33551 4029 33563 4032
rect 33505 4023 33563 4029
rect 34146 4020 34152 4072
rect 34204 4020 34210 4072
rect 34422 4020 34428 4072
rect 34480 4020 34486 4072
rect 36446 4020 36452 4072
rect 36504 4060 36510 4072
rect 37185 4063 37243 4069
rect 37185 4060 37197 4063
rect 36504 4032 37197 4060
rect 36504 4020 36510 4032
rect 37185 4029 37197 4032
rect 37231 4029 37243 4063
rect 37185 4023 37243 4029
rect 38378 4020 38384 4072
rect 38436 4020 38442 4072
rect 39758 4020 39764 4072
rect 39816 4060 39822 4072
rect 40497 4063 40555 4069
rect 40497 4060 40509 4063
rect 39816 4032 40509 4060
rect 39816 4020 39822 4032
rect 40497 4029 40509 4032
rect 40543 4029 40555 4063
rect 40497 4023 40555 4029
rect 32861 3995 32919 4001
rect 32861 3992 32873 3995
rect 31956 3964 32873 3992
rect 32861 3961 32873 3964
rect 32907 3961 32919 3995
rect 32861 3955 32919 3961
rect 33962 3952 33968 4004
rect 34020 3952 34026 4004
rect 35452 3964 36032 3992
rect 35452 3924 35480 3964
rect 30883 3896 35480 3924
rect 30883 3893 30895 3896
rect 30837 3887 30895 3893
rect 35894 3884 35900 3936
rect 35952 3884 35958 3936
rect 36004 3924 36032 3964
rect 36814 3952 36820 4004
rect 36872 3952 36878 4004
rect 40604 3992 40632 4100
rect 41325 4063 41383 4069
rect 41325 4060 41337 4063
rect 40880 4032 41337 4060
rect 40773 3995 40831 4001
rect 40773 3992 40785 3995
rect 39868 3964 40080 3992
rect 40604 3964 40785 3992
rect 37553 3927 37611 3933
rect 37553 3924 37565 3927
rect 36004 3896 37565 3924
rect 37553 3893 37565 3896
rect 37599 3893 37611 3927
rect 37553 3887 37611 3893
rect 37918 3884 37924 3936
rect 37976 3884 37982 3936
rect 38194 3884 38200 3936
rect 38252 3924 38258 3936
rect 39868 3924 39896 3964
rect 38252 3896 39896 3924
rect 38252 3884 38258 3896
rect 39942 3884 39948 3936
rect 40000 3884 40006 3936
rect 40052 3924 40080 3964
rect 40773 3961 40785 3964
rect 40819 3961 40831 3995
rect 40773 3955 40831 3961
rect 40880 3936 40908 4032
rect 41325 4029 41337 4032
rect 41371 4029 41383 4063
rect 41325 4023 41383 4029
rect 40862 3924 40868 3936
rect 40052 3896 40868 3924
rect 40862 3884 40868 3896
rect 40920 3884 40926 3936
rect 460 3834 45540 3856
rect 460 3782 3570 3834
rect 3622 3782 3634 3834
rect 3686 3782 3698 3834
rect 3750 3782 3762 3834
rect 3814 3782 3826 3834
rect 3878 3782 8570 3834
rect 8622 3782 8634 3834
rect 8686 3782 8698 3834
rect 8750 3782 8762 3834
rect 8814 3782 8826 3834
rect 8878 3782 13570 3834
rect 13622 3782 13634 3834
rect 13686 3782 13698 3834
rect 13750 3782 13762 3834
rect 13814 3782 13826 3834
rect 13878 3782 18570 3834
rect 18622 3782 18634 3834
rect 18686 3782 18698 3834
rect 18750 3782 18762 3834
rect 18814 3782 18826 3834
rect 18878 3782 23570 3834
rect 23622 3782 23634 3834
rect 23686 3782 23698 3834
rect 23750 3782 23762 3834
rect 23814 3782 23826 3834
rect 23878 3782 28570 3834
rect 28622 3782 28634 3834
rect 28686 3782 28698 3834
rect 28750 3782 28762 3834
rect 28814 3782 28826 3834
rect 28878 3782 33570 3834
rect 33622 3782 33634 3834
rect 33686 3782 33698 3834
rect 33750 3782 33762 3834
rect 33814 3782 33826 3834
rect 33878 3782 38570 3834
rect 38622 3782 38634 3834
rect 38686 3782 38698 3834
rect 38750 3782 38762 3834
rect 38814 3782 38826 3834
rect 38878 3782 43570 3834
rect 43622 3782 43634 3834
rect 43686 3782 43698 3834
rect 43750 3782 43762 3834
rect 43814 3782 43826 3834
rect 43878 3782 45540 3834
rect 460 3760 45540 3782
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4672 3692 5089 3720
rect 4672 3680 4678 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5718 3720 5724 3732
rect 5583 3692 5724 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6454 3720 6460 3732
rect 5960 3692 6460 3720
rect 5960 3680 5966 3692
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 8021 3723 8079 3729
rect 8021 3720 8033 3723
rect 7984 3692 8033 3720
rect 7984 3680 7990 3692
rect 8021 3689 8033 3692
rect 8067 3689 8079 3723
rect 8021 3683 8079 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 9088 3692 10149 3720
rect 9088 3680 9094 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10137 3683 10195 3689
rect 11238 3680 11244 3732
rect 11296 3680 11302 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12216 3692 13093 3720
rect 12216 3680 12222 3692
rect 13081 3689 13093 3692
rect 13127 3689 13139 3723
rect 13081 3683 13139 3689
rect 13262 3680 13268 3732
rect 13320 3680 13326 3732
rect 14826 3680 14832 3732
rect 14884 3680 14890 3732
rect 19058 3720 19064 3732
rect 14936 3692 19064 3720
rect 1489 3655 1547 3661
rect 1489 3621 1501 3655
rect 1535 3652 1547 3655
rect 1578 3652 1584 3664
rect 1535 3624 1584 3652
rect 1535 3621 1547 3624
rect 1489 3615 1547 3621
rect 1578 3612 1584 3624
rect 1636 3652 1642 3664
rect 2593 3655 2651 3661
rect 2593 3652 2605 3655
rect 1636 3624 2605 3652
rect 1636 3612 1642 3624
rect 2593 3621 2605 3624
rect 2639 3621 2651 3655
rect 2593 3615 2651 3621
rect 2608 3584 2636 3615
rect 9674 3612 9680 3664
rect 9732 3612 9738 3664
rect 2961 3587 3019 3593
rect 2961 3584 2973 3587
rect 2608 3556 2973 3584
rect 2961 3553 2973 3556
rect 3007 3584 3019 3587
rect 3326 3584 3332 3596
rect 3007 3556 3332 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3584 7435 3587
rect 9306 3584 9312 3596
rect 7423 3556 9312 3584
rect 7423 3553 7435 3556
rect 7377 3547 7435 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9692 3584 9720 3612
rect 10594 3584 10600 3596
rect 9692 3556 10600 3584
rect 10594 3544 10600 3556
rect 10652 3584 10658 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10652 3556 10701 3584
rect 10652 3544 10658 3556
rect 10689 3553 10701 3556
rect 10735 3584 10747 3587
rect 10962 3584 10968 3596
rect 10735 3556 10968 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11256 3584 11284 3680
rect 13280 3652 13308 3680
rect 14936 3652 14964 3692
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19242 3680 19248 3732
rect 19300 3720 19306 3732
rect 21726 3720 21732 3732
rect 19300 3692 21732 3720
rect 19300 3680 19306 3692
rect 21726 3680 21732 3692
rect 21784 3680 21790 3732
rect 21818 3680 21824 3732
rect 21876 3680 21882 3732
rect 23382 3680 23388 3732
rect 23440 3720 23446 3732
rect 23440 3692 25636 3720
rect 23440 3680 23446 3692
rect 13280 3624 14964 3652
rect 16298 3612 16304 3664
rect 16356 3652 16362 3664
rect 16356 3624 18276 3652
rect 16356 3612 16362 3624
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 11256 3556 11621 3584
rect 11609 3553 11621 3556
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 14056 3556 14105 3584
rect 14056 3544 14062 3556
rect 14093 3553 14105 3556
rect 14139 3584 14151 3587
rect 16666 3584 16672 3596
rect 14139 3556 16672 3584
rect 14139 3553 14151 3556
rect 14093 3547 14151 3553
rect 16666 3544 16672 3556
rect 16724 3584 16730 3596
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 16724 3556 17417 3584
rect 16724 3544 16730 3556
rect 17405 3553 17417 3556
rect 17451 3584 17463 3587
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17451 3556 18061 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18248 3584 18276 3624
rect 18322 3612 18328 3664
rect 18380 3652 18386 3664
rect 19260 3652 19288 3680
rect 18380 3624 19288 3652
rect 18380 3612 18386 3624
rect 18248 3556 19196 3584
rect 18049 3547 18107 3553
rect 1121 3519 1179 3525
rect 1121 3485 1133 3519
rect 1167 3516 1179 3519
rect 1486 3516 1492 3528
rect 1167 3488 1492 3516
rect 1167 3485 1179 3488
rect 1121 3479 1179 3485
rect 1486 3476 1492 3488
rect 1544 3516 1550 3528
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1544 3488 1869 3516
rect 1544 3476 1550 3488
rect 1857 3485 1869 3488
rect 1903 3516 1915 3519
rect 2590 3516 2596 3528
rect 1903 3488 2596 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 4764 3488 6193 3516
rect 4764 3476 4770 3488
rect 6181 3485 6193 3488
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 7101 3519 7159 3525
rect 6595 3488 6776 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 3605 3451 3663 3457
rect 3605 3417 3617 3451
rect 3651 3417 3663 3451
rect 6196 3448 6224 3479
rect 6638 3448 6644 3460
rect 6196 3420 6644 3448
rect 3605 3411 3663 3417
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 3620 3380 3648 3411
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 4430 3380 4436 3392
rect 3620 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6454 3380 6460 3392
rect 6411 3352 6460 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6748 3389 6776 3488
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7190 3516 7196 3528
rect 7147 3488 7196 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 10502 3476 10508 3528
rect 10560 3476 10566 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 12894 3516 12900 3528
rect 12742 3488 12900 3516
rect 11333 3479 11391 3485
rect 8570 3408 8576 3460
rect 8628 3408 8634 3460
rect 10134 3448 10140 3460
rect 9798 3420 10140 3448
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 11348 3448 11376 3479
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13906 3476 13912 3528
rect 13964 3476 13970 3528
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14976 3488 15025 3516
rect 14976 3476 14982 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 17034 3516 17040 3528
rect 16422 3488 17040 3516
rect 15013 3479 15071 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 17218 3476 17224 3528
rect 17276 3476 17282 3528
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18322 3516 18328 3528
rect 17819 3488 18328 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18463 3488 18736 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 11514 3448 11520 3460
rect 11348 3420 11520 3448
rect 11514 3408 11520 3420
rect 11572 3448 11578 3460
rect 11882 3448 11888 3460
rect 11572 3420 11888 3448
rect 11572 3408 11578 3420
rect 11882 3408 11888 3420
rect 11940 3408 11946 3460
rect 13096 3420 15240 3448
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3349 6791 3383
rect 6733 3343 6791 3349
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 10042 3340 10048 3392
rect 10100 3340 10106 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 11241 3383 11299 3389
rect 11241 3349 11253 3383
rect 11287 3380 11299 3383
rect 13096 3380 13124 3420
rect 11287 3352 13124 3380
rect 11287 3349 11299 3352
rect 11241 3343 11299 3349
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 13541 3383 13599 3389
rect 13541 3380 13553 3383
rect 13228 3352 13553 3380
rect 13228 3340 13234 3352
rect 13541 3349 13553 3352
rect 13587 3349 13599 3383
rect 13541 3343 13599 3349
rect 13998 3340 14004 3392
rect 14056 3340 14062 3392
rect 15212 3380 15240 3420
rect 15286 3408 15292 3460
rect 15344 3408 15350 3460
rect 17313 3451 17371 3457
rect 17313 3448 17325 3451
rect 16776 3420 17325 3448
rect 16298 3380 16304 3392
rect 15212 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 16574 3340 16580 3392
rect 16632 3380 16638 3392
rect 16776 3389 16804 3420
rect 17313 3417 17325 3420
rect 17359 3417 17371 3451
rect 17313 3411 17371 3417
rect 16761 3383 16819 3389
rect 16761 3380 16773 3383
rect 16632 3352 16773 3380
rect 16632 3340 16638 3352
rect 16761 3349 16773 3352
rect 16807 3349 16819 3383
rect 16761 3343 16819 3349
rect 16850 3340 16856 3392
rect 16908 3340 16914 3392
rect 18230 3340 18236 3392
rect 18288 3340 18294 3392
rect 18708 3389 18736 3488
rect 19058 3476 19064 3528
rect 19116 3476 19122 3528
rect 19168 3516 19196 3556
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 19300 3556 19349 3584
rect 19300 3544 19306 3556
rect 19337 3553 19349 3556
rect 19383 3584 19395 3587
rect 20165 3587 20223 3593
rect 20165 3584 20177 3587
rect 19383 3556 20177 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 20165 3553 20177 3556
rect 20211 3584 20223 3587
rect 20714 3584 20720 3596
rect 20211 3556 20720 3584
rect 20211 3553 20223 3556
rect 20165 3547 20223 3553
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 19886 3516 19892 3528
rect 19168 3488 19892 3516
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3485 20407 3519
rect 21836 3516 21864 3680
rect 22002 3544 22008 3596
rect 22060 3584 22066 3596
rect 22649 3587 22707 3593
rect 22649 3584 22661 3587
rect 22060 3556 22661 3584
rect 22060 3544 22066 3556
rect 22649 3553 22661 3556
rect 22695 3553 22707 3587
rect 22649 3547 22707 3553
rect 22738 3544 22744 3596
rect 22796 3544 22802 3596
rect 23934 3584 23940 3596
rect 23492 3556 23940 3584
rect 21910 3516 21916 3528
rect 21758 3488 21916 3516
rect 20349 3479 20407 3485
rect 18782 3408 18788 3460
rect 18840 3408 18846 3460
rect 19150 3408 19156 3460
rect 19208 3408 19214 3460
rect 20364 3448 20392 3479
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 23106 3516 23112 3528
rect 22572 3488 23112 3516
rect 20530 3448 20536 3460
rect 19306 3420 20536 3448
rect 18693 3383 18751 3389
rect 18693 3349 18705 3383
rect 18739 3349 18751 3383
rect 18800 3380 18828 3408
rect 19306 3380 19334 3420
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 20622 3408 20628 3460
rect 20680 3408 20686 3460
rect 22370 3408 22376 3460
rect 22428 3448 22434 3460
rect 22572 3457 22600 3488
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 22557 3451 22615 3457
rect 22557 3448 22569 3451
rect 22428 3420 22569 3448
rect 22428 3408 22434 3420
rect 22557 3417 22569 3420
rect 22603 3417 22615 3451
rect 23216 3448 23244 3479
rect 22557 3411 22615 3417
rect 22940 3420 23244 3448
rect 18800 3352 19334 3380
rect 19521 3383 19579 3389
rect 18693 3343 18751 3349
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 19886 3380 19892 3392
rect 19567 3352 19892 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3380 20039 3383
rect 20990 3380 20996 3392
rect 20027 3352 20996 3380
rect 20027 3349 20039 3352
rect 19981 3343 20039 3349
rect 20990 3340 20996 3352
rect 21048 3380 21054 3392
rect 22097 3383 22155 3389
rect 22097 3380 22109 3383
rect 21048 3352 22109 3380
rect 21048 3340 21054 3352
rect 22097 3349 22109 3352
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 22189 3383 22247 3389
rect 22189 3349 22201 3383
rect 22235 3380 22247 3383
rect 22940 3380 22968 3420
rect 23492 3392 23520 3556
rect 23934 3544 23940 3556
rect 23992 3584 23998 3596
rect 24305 3587 24363 3593
rect 24305 3584 24317 3587
rect 23992 3556 24317 3584
rect 23992 3544 23998 3556
rect 24305 3553 24317 3556
rect 24351 3553 24363 3587
rect 24946 3584 24952 3596
rect 24305 3547 24363 3553
rect 24780 3556 24952 3584
rect 23566 3476 23572 3528
rect 23624 3516 23630 3528
rect 24026 3516 24032 3528
rect 23624 3488 24032 3516
rect 23624 3476 23630 3488
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 24121 3519 24179 3525
rect 24121 3485 24133 3519
rect 24167 3516 24179 3519
rect 24780 3516 24808 3556
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 25608 3593 25636 3692
rect 27246 3680 27252 3732
rect 27304 3720 27310 3732
rect 27433 3723 27491 3729
rect 27433 3720 27445 3723
rect 27304 3692 27445 3720
rect 27304 3680 27310 3692
rect 27433 3689 27445 3692
rect 27479 3689 27491 3723
rect 27433 3683 27491 3689
rect 28077 3723 28135 3729
rect 28077 3689 28089 3723
rect 28123 3720 28135 3723
rect 28442 3720 28448 3732
rect 28123 3692 28448 3720
rect 28123 3689 28135 3692
rect 28077 3683 28135 3689
rect 27448 3652 27476 3683
rect 28442 3680 28448 3692
rect 28500 3680 28506 3732
rect 29638 3720 29644 3732
rect 29196 3692 29644 3720
rect 28534 3652 28540 3664
rect 27448 3624 28120 3652
rect 28092 3596 28120 3624
rect 28195 3624 28540 3652
rect 28195 3596 28223 3624
rect 28534 3612 28540 3624
rect 28592 3652 28598 3664
rect 29086 3652 29092 3664
rect 28592 3624 29092 3652
rect 28592 3612 28598 3624
rect 29086 3612 29092 3624
rect 29144 3612 29150 3664
rect 25593 3587 25651 3593
rect 25593 3553 25605 3587
rect 25639 3584 25651 3587
rect 26421 3587 26479 3593
rect 26421 3584 26433 3587
rect 25639 3556 26433 3584
rect 25639 3553 25651 3556
rect 25593 3547 25651 3553
rect 26421 3553 26433 3556
rect 26467 3584 26479 3587
rect 26786 3584 26792 3596
rect 26467 3556 26792 3584
rect 26467 3553 26479 3556
rect 26421 3547 26479 3553
rect 24167 3488 24808 3516
rect 24857 3519 24915 3525
rect 24167 3485 24179 3488
rect 24121 3479 24179 3485
rect 24857 3485 24869 3519
rect 24903 3516 24915 3519
rect 26237 3519 26295 3525
rect 24903 3488 25084 3516
rect 24903 3485 24915 3488
rect 24857 3479 24915 3485
rect 22235 3352 22968 3380
rect 22235 3349 22247 3352
rect 22189 3343 22247 3349
rect 23014 3340 23020 3392
rect 23072 3340 23078 3392
rect 23474 3340 23480 3392
rect 23532 3340 23538 3392
rect 23750 3340 23756 3392
rect 23808 3340 23814 3392
rect 24210 3340 24216 3392
rect 24268 3340 24274 3392
rect 24670 3340 24676 3392
rect 24728 3340 24734 3392
rect 25056 3389 25084 3488
rect 26237 3485 26249 3519
rect 26283 3516 26295 3519
rect 26326 3516 26332 3528
rect 26283 3488 26332 3516
rect 26283 3485 26295 3488
rect 26237 3479 26295 3485
rect 26326 3476 26332 3488
rect 26384 3476 26390 3528
rect 26712 3525 26740 3556
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27338 3544 27344 3596
rect 27396 3584 27402 3596
rect 27396 3556 28028 3584
rect 27396 3544 27402 3556
rect 26697 3519 26755 3525
rect 26697 3485 26709 3519
rect 26743 3485 26755 3519
rect 26697 3479 26755 3485
rect 26988 3488 27614 3516
rect 25130 3408 25136 3460
rect 25188 3448 25194 3460
rect 26988 3457 27016 3488
rect 26973 3451 27031 3457
rect 26973 3448 26985 3451
rect 25188 3420 26985 3448
rect 25188 3408 25194 3420
rect 26973 3417 26985 3420
rect 27019 3417 27031 3451
rect 26973 3411 27031 3417
rect 27249 3451 27307 3457
rect 27249 3417 27261 3451
rect 27295 3448 27307 3451
rect 27338 3448 27344 3460
rect 27295 3420 27344 3448
rect 27295 3417 27307 3420
rect 27249 3411 27307 3417
rect 27338 3408 27344 3420
rect 27396 3408 27402 3460
rect 27430 3408 27436 3460
rect 27488 3457 27494 3460
rect 27488 3451 27523 3457
rect 27511 3417 27523 3451
rect 27586 3448 27614 3488
rect 27890 3476 27896 3528
rect 27948 3476 27954 3528
rect 28000 3525 28028 3556
rect 28074 3544 28080 3596
rect 28132 3544 28138 3596
rect 28166 3544 28172 3596
rect 28224 3544 28230 3596
rect 29196 3593 29224 3692
rect 29638 3680 29644 3692
rect 29696 3680 29702 3732
rect 30006 3680 30012 3732
rect 30064 3720 30070 3732
rect 31113 3723 31171 3729
rect 31113 3720 31125 3723
rect 30064 3692 31125 3720
rect 30064 3680 30070 3692
rect 31113 3689 31125 3692
rect 31159 3689 31171 3723
rect 31113 3683 31171 3689
rect 31202 3680 31208 3732
rect 31260 3720 31266 3732
rect 31938 3720 31944 3732
rect 31260 3692 31944 3720
rect 31260 3680 31266 3692
rect 30834 3612 30840 3664
rect 30892 3652 30898 3664
rect 30929 3655 30987 3661
rect 30929 3652 30941 3655
rect 30892 3624 30941 3652
rect 30892 3612 30898 3624
rect 30929 3621 30941 3624
rect 30975 3621 30987 3655
rect 30929 3615 30987 3621
rect 29181 3587 29239 3593
rect 28552 3556 29040 3584
rect 27985 3519 28043 3525
rect 27985 3485 27997 3519
rect 28031 3516 28043 3519
rect 28350 3516 28356 3528
rect 28031 3488 28356 3516
rect 28031 3485 28043 3488
rect 27985 3479 28043 3485
rect 28350 3476 28356 3488
rect 28408 3476 28414 3528
rect 28442 3476 28448 3528
rect 28500 3476 28506 3528
rect 28552 3525 28580 3556
rect 29012 3528 29040 3556
rect 29181 3553 29193 3587
rect 29227 3553 29239 3587
rect 29181 3547 29239 3553
rect 29457 3587 29515 3593
rect 29457 3553 29469 3587
rect 29503 3584 29515 3587
rect 29546 3584 29552 3596
rect 29503 3556 29552 3584
rect 29503 3553 29515 3556
rect 29457 3547 29515 3553
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 30650 3544 30656 3596
rect 30708 3584 30714 3596
rect 31018 3584 31024 3596
rect 30708 3556 31024 3584
rect 30708 3544 30714 3556
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 28537 3519 28595 3525
rect 28537 3485 28549 3519
rect 28583 3485 28595 3519
rect 28537 3479 28595 3485
rect 28721 3519 28779 3525
rect 28721 3485 28733 3519
rect 28767 3516 28779 3519
rect 28905 3519 28963 3525
rect 28905 3516 28917 3519
rect 28767 3488 28917 3516
rect 28767 3485 28779 3488
rect 28721 3479 28779 3485
rect 28905 3485 28917 3488
rect 28951 3485 28963 3519
rect 28905 3479 28963 3485
rect 27706 3448 27712 3460
rect 27586 3420 27712 3448
rect 27488 3411 27523 3417
rect 27488 3408 27494 3411
rect 27706 3408 27712 3420
rect 27764 3408 27770 3460
rect 28920 3448 28948 3479
rect 28994 3476 29000 3528
rect 29052 3476 29058 3528
rect 29086 3476 29092 3528
rect 29144 3476 29150 3528
rect 30834 3476 30840 3528
rect 30892 3516 30898 3528
rect 31312 3525 31340 3692
rect 31938 3680 31944 3692
rect 31996 3680 32002 3732
rect 32398 3680 32404 3732
rect 32456 3680 32462 3732
rect 32950 3680 32956 3732
rect 33008 3680 33014 3732
rect 33226 3680 33232 3732
rect 33284 3720 33290 3732
rect 34241 3723 34299 3729
rect 34241 3720 34253 3723
rect 33284 3692 34253 3720
rect 33284 3680 33290 3692
rect 34241 3689 34253 3692
rect 34287 3689 34299 3723
rect 34241 3683 34299 3689
rect 34422 3680 34428 3732
rect 34480 3720 34486 3732
rect 34701 3723 34759 3729
rect 34701 3720 34713 3723
rect 34480 3692 34713 3720
rect 34480 3680 34486 3692
rect 34701 3689 34713 3692
rect 34747 3689 34759 3723
rect 34701 3683 34759 3689
rect 35894 3680 35900 3732
rect 35952 3680 35958 3732
rect 38378 3680 38384 3732
rect 38436 3720 38442 3732
rect 38473 3723 38531 3729
rect 38473 3720 38485 3723
rect 38436 3692 38485 3720
rect 38436 3680 38442 3692
rect 38473 3689 38485 3692
rect 38519 3689 38531 3723
rect 39942 3720 39948 3732
rect 38473 3683 38531 3689
rect 38948 3692 39948 3720
rect 32968 3652 32996 3680
rect 35912 3652 35940 3680
rect 32968 3624 33824 3652
rect 32674 3584 32680 3596
rect 31726 3556 32680 3584
rect 31119 3519 31177 3525
rect 31119 3516 31131 3519
rect 30892 3488 31131 3516
rect 30892 3476 30898 3488
rect 31119 3485 31131 3488
rect 31165 3485 31177 3519
rect 31119 3479 31177 3485
rect 31297 3519 31355 3525
rect 31297 3485 31309 3519
rect 31343 3485 31355 3519
rect 31297 3479 31355 3485
rect 31527 3519 31585 3525
rect 31527 3485 31539 3519
rect 31573 3516 31585 3519
rect 31726 3516 31754 3556
rect 32674 3544 32680 3556
rect 32732 3544 32738 3596
rect 32858 3544 32864 3596
rect 32916 3544 32922 3596
rect 33045 3587 33103 3593
rect 33045 3553 33057 3587
rect 33091 3584 33103 3587
rect 33134 3584 33140 3596
rect 33091 3556 33140 3584
rect 33091 3553 33103 3556
rect 33045 3547 33103 3553
rect 33134 3544 33140 3556
rect 33192 3544 33198 3596
rect 33796 3584 33824 3624
rect 35544 3624 35940 3652
rect 35544 3593 35572 3624
rect 35529 3587 35587 3593
rect 33796 3556 35204 3584
rect 31573 3488 31754 3516
rect 31849 3519 31907 3525
rect 31573 3485 31585 3488
rect 31527 3479 31585 3485
rect 31849 3485 31861 3519
rect 31895 3512 31907 3519
rect 31938 3512 31944 3528
rect 31895 3485 31944 3512
rect 31849 3484 31944 3485
rect 31849 3479 31907 3484
rect 31938 3476 31944 3484
rect 31996 3476 32002 3528
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 29362 3448 29368 3460
rect 28920 3420 29368 3448
rect 29362 3408 29368 3420
rect 29420 3408 29426 3460
rect 29546 3408 29552 3460
rect 29604 3448 29610 3460
rect 29604 3420 29946 3448
rect 30852 3420 31064 3448
rect 29604 3408 29610 3420
rect 25041 3383 25099 3389
rect 25041 3349 25053 3383
rect 25087 3349 25099 3383
rect 25041 3343 25099 3349
rect 25222 3340 25228 3392
rect 25280 3380 25286 3392
rect 25406 3380 25412 3392
rect 25280 3352 25412 3380
rect 25280 3340 25286 3352
rect 25406 3340 25412 3352
rect 25464 3340 25470 3392
rect 25501 3383 25559 3389
rect 25501 3349 25513 3383
rect 25547 3380 25559 3383
rect 25682 3380 25688 3392
rect 25547 3352 25688 3380
rect 25547 3349 25559 3352
rect 25501 3343 25559 3349
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 25869 3383 25927 3389
rect 25869 3349 25881 3383
rect 25915 3380 25927 3383
rect 25958 3380 25964 3392
rect 25915 3352 25964 3380
rect 25915 3349 25927 3352
rect 25869 3343 25927 3349
rect 25958 3340 25964 3352
rect 26016 3340 26022 3392
rect 26329 3383 26387 3389
rect 26329 3349 26341 3383
rect 26375 3380 26387 3383
rect 27062 3380 27068 3392
rect 26375 3352 27068 3380
rect 26375 3349 26387 3352
rect 26329 3343 26387 3349
rect 27062 3340 27068 3352
rect 27120 3340 27126 3392
rect 27614 3340 27620 3392
rect 27672 3340 27678 3392
rect 28258 3340 28264 3392
rect 28316 3340 28322 3392
rect 28629 3383 28687 3389
rect 28629 3349 28641 3383
rect 28675 3380 28687 3383
rect 28902 3380 28908 3392
rect 28675 3352 28908 3380
rect 28675 3349 28687 3352
rect 28629 3343 28687 3349
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 28997 3383 29055 3389
rect 28997 3349 29009 3383
rect 29043 3380 29055 3383
rect 29270 3380 29276 3392
rect 29043 3352 29276 3380
rect 29043 3349 29055 3352
rect 28997 3343 29055 3349
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 29454 3340 29460 3392
rect 29512 3380 29518 3392
rect 30852 3380 30880 3420
rect 29512 3352 30880 3380
rect 31036 3380 31064 3420
rect 31386 3408 31392 3460
rect 31444 3448 31450 3460
rect 31665 3451 31723 3457
rect 31665 3448 31677 3451
rect 31444 3420 31677 3448
rect 31444 3408 31450 3420
rect 31665 3417 31677 3420
rect 31711 3417 31723 3451
rect 31665 3411 31723 3417
rect 31754 3408 31760 3460
rect 31812 3408 31818 3460
rect 32140 3448 32168 3479
rect 32306 3476 32312 3528
rect 32364 3476 32370 3528
rect 33410 3476 33416 3528
rect 33468 3476 33474 3528
rect 34606 3476 34612 3528
rect 34664 3476 34670 3528
rect 34885 3519 34943 3525
rect 34885 3485 34897 3519
rect 34931 3516 34943 3519
rect 34931 3488 35112 3516
rect 34931 3485 34943 3488
rect 34885 3479 34943 3485
rect 33134 3448 33140 3460
rect 31956 3420 32168 3448
rect 32324 3420 33140 3448
rect 31956 3380 31984 3420
rect 31036 3352 31984 3380
rect 29512 3340 29518 3352
rect 32030 3340 32036 3392
rect 32088 3340 32094 3392
rect 32324 3389 32352 3420
rect 33134 3408 33140 3420
rect 33192 3408 33198 3460
rect 33686 3408 33692 3460
rect 33744 3408 33750 3460
rect 32309 3383 32367 3389
rect 32309 3349 32321 3383
rect 32355 3349 32367 3383
rect 32309 3343 32367 3349
rect 32766 3340 32772 3392
rect 32824 3340 32830 3392
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 33229 3383 33287 3389
rect 33229 3380 33241 3383
rect 33100 3352 33241 3380
rect 33100 3340 33106 3352
rect 33229 3349 33241 3352
rect 33275 3349 33287 3383
rect 33229 3343 33287 3349
rect 34422 3340 34428 3392
rect 34480 3340 34486 3392
rect 35084 3389 35112 3488
rect 35069 3383 35127 3389
rect 35069 3349 35081 3383
rect 35115 3349 35127 3383
rect 35176 3380 35204 3556
rect 35529 3553 35541 3587
rect 35575 3553 35587 3587
rect 35529 3547 35587 3553
rect 35710 3544 35716 3596
rect 35768 3544 35774 3596
rect 35912 3584 35940 3624
rect 36556 3624 38240 3652
rect 36556 3596 36584 3624
rect 38212 3596 38240 3624
rect 36357 3587 36415 3593
rect 36357 3584 36369 3587
rect 35912 3556 36369 3584
rect 36357 3553 36369 3556
rect 36403 3553 36415 3587
rect 36357 3547 36415 3553
rect 36538 3544 36544 3596
rect 36596 3544 36602 3596
rect 37369 3587 37427 3593
rect 37369 3584 37381 3587
rect 37200 3556 37381 3584
rect 35802 3516 35808 3528
rect 35544 3488 35808 3516
rect 35437 3451 35495 3457
rect 35437 3417 35449 3451
rect 35483 3448 35495 3451
rect 35544 3448 35572 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36998 3516 37004 3528
rect 35952 3488 37004 3516
rect 35952 3476 35958 3488
rect 36998 3476 37004 3488
rect 37056 3516 37062 3528
rect 37200 3516 37228 3556
rect 37369 3553 37381 3556
rect 37415 3553 37427 3587
rect 37369 3547 37427 3553
rect 38194 3544 38200 3596
rect 38252 3544 38258 3596
rect 37056 3488 37228 3516
rect 38657 3519 38715 3525
rect 37056 3476 37062 3488
rect 38657 3485 38669 3519
rect 38703 3516 38715 3519
rect 38948 3516 38976 3692
rect 39942 3680 39948 3692
rect 40000 3680 40006 3732
rect 40954 3680 40960 3732
rect 41012 3680 41018 3732
rect 41693 3723 41751 3729
rect 41693 3689 41705 3723
rect 41739 3720 41751 3723
rect 41874 3720 41880 3732
rect 41739 3692 41880 3720
rect 41739 3689 41751 3692
rect 41693 3683 41751 3689
rect 41874 3680 41880 3692
rect 41932 3720 41938 3732
rect 42705 3723 42763 3729
rect 42705 3720 42717 3723
rect 41932 3692 42717 3720
rect 41932 3680 41938 3692
rect 42705 3689 42717 3692
rect 42751 3720 42763 3723
rect 43073 3723 43131 3729
rect 43073 3720 43085 3723
rect 42751 3692 43085 3720
rect 42751 3689 42763 3692
rect 42705 3683 42763 3689
rect 43073 3689 43085 3692
rect 43119 3689 43131 3723
rect 43073 3683 43131 3689
rect 43901 3723 43959 3729
rect 43901 3689 43913 3723
rect 43947 3720 43959 3723
rect 44542 3720 44548 3732
rect 43947 3692 44548 3720
rect 43947 3689 43959 3692
rect 43901 3683 43959 3689
rect 44542 3680 44548 3692
rect 44600 3720 44606 3732
rect 44818 3720 44824 3732
rect 44600 3692 44824 3720
rect 44600 3680 44606 3692
rect 44818 3680 44824 3692
rect 44876 3680 44882 3732
rect 44910 3680 44916 3732
rect 44968 3680 44974 3732
rect 40586 3612 40592 3664
rect 40644 3652 40650 3664
rect 41233 3655 41291 3661
rect 41233 3652 41245 3655
rect 40644 3624 41245 3652
rect 40644 3612 40650 3624
rect 41233 3621 41245 3624
rect 41279 3621 41291 3655
rect 41233 3615 41291 3621
rect 42061 3655 42119 3661
rect 42061 3621 42073 3655
rect 42107 3652 42119 3655
rect 42242 3652 42248 3664
rect 42107 3624 42248 3652
rect 42107 3621 42119 3624
rect 42061 3615 42119 3621
rect 42242 3612 42248 3624
rect 42300 3612 42306 3664
rect 42429 3655 42487 3661
rect 42429 3621 42441 3655
rect 42475 3652 42487 3655
rect 42518 3652 42524 3664
rect 42475 3624 42524 3652
rect 42475 3621 42487 3624
rect 42429 3615 42487 3621
rect 40034 3584 40040 3596
rect 39040 3556 40040 3584
rect 39040 3525 39068 3556
rect 40034 3544 40040 3556
rect 40092 3544 40098 3596
rect 40218 3544 40224 3596
rect 40276 3584 40282 3596
rect 40276 3556 40632 3584
rect 40276 3544 40282 3556
rect 38703 3488 38976 3516
rect 39025 3519 39083 3525
rect 38703 3485 38715 3488
rect 38657 3479 38715 3485
rect 39025 3485 39037 3519
rect 39071 3485 39083 3519
rect 39025 3479 39083 3485
rect 39209 3519 39267 3525
rect 39209 3485 39221 3519
rect 39255 3485 39267 3519
rect 40604 3516 40632 3556
rect 42444 3516 42472 3615
rect 42518 3612 42524 3624
rect 42576 3652 42582 3664
rect 43346 3652 43352 3664
rect 42576 3624 43352 3652
rect 42576 3612 42582 3624
rect 43346 3612 43352 3624
rect 43404 3652 43410 3664
rect 43441 3655 43499 3661
rect 43441 3652 43453 3655
rect 43404 3624 43453 3652
rect 43404 3612 43410 3624
rect 43441 3621 43453 3624
rect 43487 3621 43499 3655
rect 43441 3615 43499 3621
rect 44637 3655 44695 3661
rect 44637 3621 44649 3655
rect 44683 3652 44695 3655
rect 44726 3652 44732 3664
rect 44683 3624 44732 3652
rect 44683 3621 44695 3624
rect 44637 3615 44695 3621
rect 44726 3612 44732 3624
rect 44784 3612 44790 3664
rect 40604 3502 42472 3516
rect 40618 3488 42472 3502
rect 39209 3479 39267 3485
rect 37182 3448 37188 3460
rect 35483 3420 35572 3448
rect 36004 3420 37188 3448
rect 35483 3417 35495 3420
rect 35437 3411 35495 3417
rect 36004 3392 36032 3420
rect 37182 3408 37188 3420
rect 37240 3408 37246 3460
rect 38746 3408 38752 3460
rect 38804 3448 38810 3460
rect 39224 3448 39252 3479
rect 38804 3420 39252 3448
rect 39485 3451 39543 3457
rect 38804 3408 38810 3420
rect 39485 3417 39497 3451
rect 39531 3417 39543 3451
rect 39485 3411 39543 3417
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35176 3352 35909 3380
rect 35069 3343 35127 3349
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 35986 3340 35992 3392
rect 36044 3340 36050 3392
rect 36265 3383 36323 3389
rect 36265 3349 36277 3383
rect 36311 3380 36323 3383
rect 36722 3380 36728 3392
rect 36311 3352 36728 3380
rect 36311 3349 36323 3352
rect 36265 3343 36323 3349
rect 36722 3340 36728 3352
rect 36780 3340 36786 3392
rect 36814 3340 36820 3392
rect 36872 3340 36878 3392
rect 37274 3340 37280 3392
rect 37332 3340 37338 3392
rect 37642 3340 37648 3392
rect 37700 3340 37706 3392
rect 38010 3340 38016 3392
rect 38068 3340 38074 3392
rect 38102 3340 38108 3392
rect 38160 3340 38166 3392
rect 38841 3383 38899 3389
rect 38841 3349 38853 3383
rect 38887 3380 38899 3383
rect 39500 3380 39528 3411
rect 38887 3352 39528 3380
rect 38887 3349 38899 3352
rect 38841 3343 38899 3349
rect 460 3290 45540 3312
rect 460 3238 6070 3290
rect 6122 3238 6134 3290
rect 6186 3238 6198 3290
rect 6250 3238 6262 3290
rect 6314 3238 6326 3290
rect 6378 3238 11070 3290
rect 11122 3238 11134 3290
rect 11186 3238 11198 3290
rect 11250 3238 11262 3290
rect 11314 3238 11326 3290
rect 11378 3238 16070 3290
rect 16122 3238 16134 3290
rect 16186 3238 16198 3290
rect 16250 3238 16262 3290
rect 16314 3238 16326 3290
rect 16378 3238 21070 3290
rect 21122 3238 21134 3290
rect 21186 3238 21198 3290
rect 21250 3238 21262 3290
rect 21314 3238 21326 3290
rect 21378 3238 26070 3290
rect 26122 3238 26134 3290
rect 26186 3238 26198 3290
rect 26250 3238 26262 3290
rect 26314 3238 26326 3290
rect 26378 3238 31070 3290
rect 31122 3238 31134 3290
rect 31186 3238 31198 3290
rect 31250 3238 31262 3290
rect 31314 3238 31326 3290
rect 31378 3238 36070 3290
rect 36122 3238 36134 3290
rect 36186 3238 36198 3290
rect 36250 3238 36262 3290
rect 36314 3238 36326 3290
rect 36378 3238 41070 3290
rect 41122 3238 41134 3290
rect 41186 3238 41198 3290
rect 41250 3238 41262 3290
rect 41314 3238 41326 3290
rect 41378 3238 45540 3290
rect 460 3216 45540 3238
rect 937 3179 995 3185
rect 937 3145 949 3179
rect 983 3176 995 3179
rect 1302 3176 1308 3188
rect 983 3148 1308 3176
rect 983 3145 995 3148
rect 937 3139 995 3145
rect 1302 3136 1308 3148
rect 1360 3136 1366 3188
rect 1578 3136 1584 3188
rect 1636 3136 1642 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 2648 3148 2912 3176
rect 2648 3136 2654 3148
rect 1596 3108 1624 3136
rect 1504 3080 1624 3108
rect 750 3000 756 3052
rect 808 3000 814 3052
rect 1504 3049 1532 3080
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3009 1547 3043
rect 2884 3026 2912 3148
rect 4154 3136 4160 3188
rect 4212 3136 4218 3188
rect 4430 3136 4436 3188
rect 4488 3136 4494 3188
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5718 3176 5724 3188
rect 5583 3148 5724 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 6454 3136 6460 3188
rect 6512 3136 6518 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7248 3148 7665 3176
rect 7248 3136 7254 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8570 3176 8576 3188
rect 8435 3148 8576 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 10413 3179 10471 3185
rect 10413 3145 10425 3179
rect 10459 3176 10471 3179
rect 10594 3176 10600 3188
rect 10459 3148 10600 3176
rect 10459 3145 10471 3148
rect 10413 3139 10471 3145
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 13170 3136 13176 3188
rect 13228 3136 13234 3188
rect 14458 3136 14464 3188
rect 14516 3136 14522 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15657 3179 15715 3185
rect 15657 3176 15669 3179
rect 15344 3148 15669 3176
rect 15344 3136 15350 3148
rect 15657 3145 15669 3148
rect 15703 3145 15715 3179
rect 15657 3139 15715 3145
rect 16850 3136 16856 3188
rect 16908 3136 16914 3188
rect 18230 3176 18236 3188
rect 17328 3148 18236 3176
rect 3973 3111 4031 3117
rect 3973 3077 3985 3111
rect 4019 3108 4031 3111
rect 4062 3108 4068 3120
rect 4019 3080 4068 3108
rect 4019 3077 4031 3080
rect 3973 3071 4031 3077
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4172 3040 4200 3136
rect 6181 3111 6239 3117
rect 6181 3077 6193 3111
rect 6227 3108 6239 3111
rect 6472 3108 6500 3136
rect 6227 3080 6500 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 6638 3068 6644 3120
rect 6696 3068 6702 3120
rect 11425 3111 11483 3117
rect 11425 3077 11437 3111
rect 11471 3108 11483 3111
rect 11790 3108 11796 3120
rect 11471 3080 11796 3108
rect 11471 3077 11483 3080
rect 11425 3071 11483 3077
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 13188 3108 13216 3136
rect 16868 3108 16896 3136
rect 17328 3117 17356 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 19334 3176 19340 3188
rect 18380 3148 19340 3176
rect 18380 3136 18386 3148
rect 19334 3136 19340 3148
rect 19392 3176 19398 3188
rect 19392 3148 19564 3176
rect 19392 3136 19398 3148
rect 12636 3080 13216 3108
rect 15856 3080 16896 3108
rect 17313 3111 17371 3117
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4172 3012 4629 3040
rect 1489 3003 1547 3009
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5902 3040 5908 3052
rect 5215 3012 5908 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 8570 3000 8576 3052
rect 8628 3000 8634 3052
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10008 3012 10074 3040
rect 10008 3000 10014 3012
rect 11330 3000 11336 3052
rect 11388 3000 11394 3052
rect 12636 3049 12664 3080
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 14090 3000 14096 3052
rect 14148 3000 14154 3052
rect 15856 3049 15884 3080
rect 17313 3077 17325 3111
rect 17359 3077 17371 3111
rect 17313 3071 17371 3077
rect 17770 3068 17776 3120
rect 17828 3068 17834 3120
rect 19153 3111 19211 3117
rect 19153 3077 19165 3111
rect 19199 3108 19211 3111
rect 19426 3108 19432 3120
rect 19199 3080 19432 3108
rect 19199 3077 19211 3080
rect 19153 3071 19211 3077
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 19536 3108 19564 3148
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 20530 3176 20536 3188
rect 19944 3148 20536 3176
rect 19944 3136 19950 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 20622 3136 20628 3188
rect 20680 3176 20686 3188
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 20680 3148 20821 3176
rect 20680 3136 20686 3148
rect 20809 3145 20821 3148
rect 20855 3145 20867 3179
rect 23014 3176 23020 3188
rect 20809 3139 20867 3145
rect 21468 3148 23020 3176
rect 21468 3117 21496 3148
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 24670 3176 24676 3188
rect 24412 3148 24676 3176
rect 21453 3111 21511 3117
rect 19536 3080 19642 3108
rect 21453 3077 21465 3111
rect 21499 3077 21511 3111
rect 21453 3071 21511 3077
rect 21542 3068 21548 3120
rect 21600 3108 21606 3120
rect 21910 3108 21916 3120
rect 21600 3080 21916 3108
rect 21600 3068 21606 3080
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 23474 3108 23480 3120
rect 22756 3080 23480 3108
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3009 15071 3043
rect 15013 3003 15071 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 1762 2932 1768 2984
rect 1820 2932 1826 2984
rect 3970 2932 3976 2984
rect 4028 2932 4034 2984
rect 4062 2932 4068 2984
rect 4120 2932 4126 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2941 4215 2975
rect 8312 2972 8340 3000
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8312 2944 8677 2972
rect 4157 2935 4215 2941
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 3988 2904 4016 2932
rect 4172 2904 4200 2935
rect 8938 2932 8944 2984
rect 8996 2932 9002 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9364 2944 9996 2972
rect 9364 2932 9370 2944
rect 2884 2876 4200 2904
rect 1397 2839 1455 2845
rect 1397 2805 1409 2839
rect 1443 2836 1455 2839
rect 2406 2836 2412 2848
rect 1443 2808 2412 2836
rect 1443 2805 1455 2808
rect 1397 2799 1455 2805
rect 2406 2796 2412 2808
rect 2464 2836 2470 2848
rect 2884 2836 2912 2876
rect 8294 2864 8300 2916
rect 8352 2864 8358 2916
rect 9968 2904 9996 2944
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 11020 2944 11529 2972
rect 11020 2932 11026 2944
rect 11517 2941 11529 2944
rect 11563 2941 11575 2975
rect 11517 2935 11575 2941
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12342 2972 12348 2984
rect 11940 2944 12348 2972
rect 11940 2932 11946 2944
rect 12342 2932 12348 2944
rect 12400 2972 12406 2984
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 12400 2944 12725 2972
rect 12400 2932 12406 2944
rect 12713 2941 12725 2944
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13354 2972 13360 2984
rect 13035 2944 13360 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 15028 2972 15056 3003
rect 16390 3000 16396 3052
rect 16448 3000 16454 3052
rect 16666 3000 16672 3052
rect 16724 3000 16730 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16816 3012 17049 3040
rect 16816 3000 16822 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 15028 2944 16068 2972
rect 16040 2913 16068 2944
rect 16482 2932 16488 2984
rect 16540 2932 16546 2984
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2972 16635 2975
rect 16684 2972 16712 3000
rect 16623 2944 16712 2972
rect 17052 2972 17080 3003
rect 18782 3000 18788 3052
rect 18840 3000 18846 3052
rect 20530 3000 20536 3052
rect 20588 3040 20594 3052
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20588 3012 21005 3040
rect 20588 3000 20594 3012
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 20993 3003 21051 3009
rect 18800 2972 18828 3000
rect 22756 2984 22784 3080
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 23753 3111 23811 3117
rect 23753 3077 23765 3111
rect 23799 3108 23811 3111
rect 24302 3108 24308 3120
rect 23799 3080 24308 3108
rect 23799 3077 23811 3080
rect 23753 3071 23811 3077
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 24412 3117 24440 3148
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 24762 3136 24768 3188
rect 24820 3136 24826 3188
rect 25682 3136 25688 3188
rect 25740 3176 25746 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 25740 3148 25881 3176
rect 25740 3136 25746 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 25958 3136 25964 3188
rect 26016 3136 26022 3188
rect 26053 3179 26111 3185
rect 26053 3145 26065 3179
rect 26099 3176 26111 3179
rect 26602 3176 26608 3188
rect 26099 3148 26608 3176
rect 26099 3145 26111 3148
rect 26053 3139 26111 3145
rect 26602 3136 26608 3148
rect 26660 3136 26666 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 29641 3179 29699 3185
rect 29641 3176 29653 3179
rect 27580 3148 29653 3176
rect 27580 3136 27586 3148
rect 29641 3145 29653 3148
rect 29687 3145 29699 3179
rect 29641 3139 29699 3145
rect 29730 3136 29736 3188
rect 29788 3136 29794 3188
rect 30558 3176 30564 3188
rect 30116 3148 30564 3176
rect 24397 3111 24455 3117
rect 24397 3077 24409 3111
rect 24443 3077 24455 3111
rect 24780 3108 24808 3136
rect 25976 3108 26004 3136
rect 24780 3080 24886 3108
rect 25976 3080 26556 3108
rect 24397 3071 24455 3077
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3040 23259 3043
rect 23247 3012 23336 3040
rect 23247 3009 23259 3012
rect 23201 3003 23259 3009
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 17052 2944 18889 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 19150 2972 19156 2984
rect 18877 2935 18935 2941
rect 18984 2944 19156 2972
rect 16025 2907 16083 2913
rect 9968 2876 12848 2904
rect 2464 2808 2912 2836
rect 2464 2796 2470 2808
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3237 2839 3295 2845
rect 3237 2836 3249 2839
rect 3016 2808 3249 2836
rect 3016 2796 3022 2808
rect 3237 2805 3249 2808
rect 3283 2805 3295 2839
rect 3237 2799 3295 2805
rect 3326 2796 3332 2848
rect 3384 2836 3390 2848
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3384 2808 3617 2836
rect 3384 2796 3390 2808
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 3605 2799 3663 2805
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2836 11023 2839
rect 11422 2836 11428 2848
rect 11011 2808 11428 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 12342 2796 12348 2848
rect 12400 2796 12406 2848
rect 12434 2796 12440 2848
rect 12492 2796 12498 2848
rect 12820 2836 12848 2876
rect 14016 2876 15976 2904
rect 14016 2836 14044 2876
rect 12820 2808 14044 2836
rect 14826 2796 14832 2848
rect 14884 2796 14890 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15381 2839 15439 2845
rect 15381 2836 15393 2839
rect 14976 2808 15393 2836
rect 14976 2796 14982 2808
rect 15381 2805 15393 2808
rect 15427 2805 15439 2839
rect 15948 2836 15976 2876
rect 16025 2873 16037 2907
rect 16071 2873 16083 2907
rect 16025 2867 16083 2873
rect 18785 2907 18843 2913
rect 18785 2873 18797 2907
rect 18831 2904 18843 2907
rect 18984 2904 19012 2944
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19886 2932 19892 2984
rect 19944 2972 19950 2984
rect 20438 2972 20444 2984
rect 19944 2944 20444 2972
rect 19944 2932 19950 2944
rect 20438 2932 20444 2944
rect 20496 2972 20502 2984
rect 20625 2975 20683 2981
rect 20625 2972 20637 2975
rect 20496 2944 20637 2972
rect 20496 2932 20502 2944
rect 20625 2941 20637 2944
rect 20671 2941 20683 2975
rect 20625 2935 20683 2941
rect 21082 2932 21088 2984
rect 21140 2972 21146 2984
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 21140 2944 21189 2972
rect 21140 2932 21146 2944
rect 21177 2941 21189 2944
rect 21223 2941 21235 2975
rect 22738 2972 22744 2984
rect 21177 2935 21235 2941
rect 21284 2944 22744 2972
rect 18831 2876 19012 2904
rect 18831 2873 18843 2876
rect 18785 2867 18843 2873
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 21284 2904 21312 2944
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 23308 2913 23336 3012
rect 23492 2972 23520 3068
rect 23661 3043 23719 3049
rect 23661 3009 23673 3043
rect 23707 3040 23719 3043
rect 23707 3012 24072 3040
rect 23707 3009 23719 3012
rect 23661 3003 23719 3009
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23492 2944 23857 2972
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 24044 2972 24072 3012
rect 24118 3000 24124 3052
rect 24176 3000 24182 3052
rect 25406 3000 25412 3052
rect 25464 3000 25470 3052
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25924 3012 25973 3040
rect 25924 3000 25930 3012
rect 25961 3009 25973 3012
rect 26007 3009 26019 3043
rect 25961 3003 26019 3009
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26418 3040 26424 3052
rect 26191 3012 26424 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 26528 3049 26556 3080
rect 26878 3068 26884 3120
rect 26936 3108 26942 3120
rect 28905 3111 28963 3117
rect 26936 3080 27370 3108
rect 26936 3068 26942 3080
rect 28905 3077 28917 3111
rect 28951 3108 28963 3111
rect 30116 3108 30144 3148
rect 30558 3136 30564 3148
rect 30616 3136 30622 3188
rect 32030 3176 32036 3188
rect 31956 3148 32036 3176
rect 31956 3117 31984 3148
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 32674 3136 32680 3188
rect 32732 3176 32738 3188
rect 33597 3179 33655 3185
rect 33597 3176 33609 3179
rect 32732 3148 33609 3176
rect 32732 3136 32738 3148
rect 33597 3145 33609 3148
rect 33643 3145 33655 3179
rect 33597 3139 33655 3145
rect 34606 3136 34612 3188
rect 34664 3176 34670 3188
rect 34977 3179 35035 3185
rect 34977 3176 34989 3179
rect 34664 3148 34989 3176
rect 34664 3136 34670 3148
rect 34977 3145 34989 3148
rect 35023 3145 35035 3179
rect 34977 3139 35035 3145
rect 35345 3179 35403 3185
rect 35345 3145 35357 3179
rect 35391 3176 35403 3179
rect 35802 3176 35808 3188
rect 35391 3148 35808 3176
rect 35391 3145 35403 3148
rect 35345 3139 35403 3145
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 35986 3176 35992 3188
rect 35912 3148 35992 3176
rect 28951 3080 30144 3108
rect 31941 3111 31999 3117
rect 28951 3077 28963 3080
rect 28905 3071 28963 3077
rect 31941 3077 31953 3111
rect 31987 3077 31999 3111
rect 31941 3071 31999 3077
rect 32950 3068 32956 3120
rect 33008 3068 33014 3120
rect 34517 3111 34575 3117
rect 34517 3077 34529 3111
rect 34563 3108 34575 3111
rect 35250 3108 35256 3120
rect 34563 3080 35256 3108
rect 34563 3077 34575 3080
rect 34517 3071 34575 3077
rect 35250 3068 35256 3080
rect 35308 3108 35314 3120
rect 35437 3111 35495 3117
rect 35437 3108 35449 3111
rect 35308 3080 35449 3108
rect 35308 3068 35314 3080
rect 35437 3077 35449 3080
rect 35483 3077 35495 3111
rect 35437 3071 35495 3077
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 28166 3000 28172 3052
rect 28224 3040 28230 3052
rect 28721 3043 28779 3049
rect 28721 3040 28733 3043
rect 28224 3012 28733 3040
rect 28224 3000 28230 3012
rect 28721 3009 28733 3012
rect 28767 3009 28779 3043
rect 28721 3003 28779 3009
rect 29270 3000 29276 3052
rect 29328 3040 29334 3052
rect 29328 3012 29500 3040
rect 29328 3000 29334 3012
rect 25424 2972 25452 3000
rect 24044 2944 25452 2972
rect 23845 2935 23903 2941
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 26605 2975 26663 2981
rect 26605 2972 26617 2975
rect 25648 2944 26617 2972
rect 25648 2932 25654 2944
rect 26605 2941 26617 2944
rect 26651 2941 26663 2975
rect 26605 2935 26663 2941
rect 26881 2975 26939 2981
rect 26881 2941 26893 2975
rect 26927 2972 26939 2975
rect 27430 2972 27436 2984
rect 26927 2944 27436 2972
rect 26927 2941 26939 2944
rect 26881 2935 26939 2941
rect 20772 2876 21312 2904
rect 20772 2864 20778 2876
rect 21174 2836 21180 2848
rect 15948 2808 21180 2836
rect 15381 2799 15439 2805
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21284 2836 21312 2876
rect 23293 2907 23351 2913
rect 23293 2873 23305 2907
rect 23339 2873 23351 2907
rect 23293 2867 23351 2873
rect 21910 2836 21916 2848
rect 21284 2808 21916 2836
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 22925 2839 22983 2845
rect 22925 2836 22937 2839
rect 22060 2808 22937 2836
rect 22060 2796 22066 2808
rect 22925 2805 22937 2808
rect 22971 2805 22983 2839
rect 22925 2799 22983 2805
rect 23014 2796 23020 2848
rect 23072 2796 23078 2848
rect 26326 2796 26332 2848
rect 26384 2796 26390 2848
rect 26620 2836 26648 2935
rect 27430 2932 27436 2944
rect 27488 2932 27494 2984
rect 28258 2932 28264 2984
rect 28316 2972 28322 2984
rect 28534 2972 28540 2984
rect 28316 2944 28540 2972
rect 28316 2932 28322 2944
rect 28534 2932 28540 2944
rect 28592 2972 28598 2984
rect 29472 2981 29500 3012
rect 29546 3000 29552 3052
rect 29604 3040 29610 3052
rect 30009 3043 30067 3049
rect 30009 3040 30021 3043
rect 29604 3012 30021 3040
rect 29604 3000 29610 3012
rect 30009 3009 30021 3012
rect 30055 3009 30067 3043
rect 30009 3003 30067 3009
rect 30098 3000 30104 3052
rect 30156 3000 30162 3052
rect 30193 3043 30251 3049
rect 30193 3009 30205 3043
rect 30239 3040 30251 3043
rect 30282 3040 30288 3052
rect 30239 3012 30288 3040
rect 30239 3009 30251 3012
rect 30193 3003 30251 3009
rect 30282 3000 30288 3012
rect 30340 3000 30346 3052
rect 30374 3000 30380 3052
rect 30432 3000 30438 3052
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30653 3043 30711 3049
rect 30653 3040 30665 3043
rect 30524 3012 30665 3040
rect 30524 3000 30530 3012
rect 30653 3009 30665 3012
rect 30699 3040 30711 3043
rect 31478 3040 31484 3052
rect 30699 3012 31484 3040
rect 30699 3009 30711 3012
rect 30653 3003 30711 3009
rect 31478 3000 31484 3012
rect 31536 3000 31542 3052
rect 33502 3000 33508 3052
rect 33560 3000 33566 3052
rect 33689 3043 33747 3049
rect 33689 3009 33701 3043
rect 33735 3009 33747 3043
rect 33689 3003 33747 3009
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3009 34115 3043
rect 34057 3003 34115 3009
rect 34609 3043 34667 3049
rect 34609 3009 34621 3043
rect 34655 3040 34667 3043
rect 35912 3040 35940 3148
rect 35986 3136 35992 3148
rect 36044 3136 36050 3188
rect 36814 3136 36820 3188
rect 36872 3136 36878 3188
rect 36998 3136 37004 3188
rect 37056 3176 37062 3188
rect 40221 3179 40279 3185
rect 37056 3148 40080 3176
rect 37056 3136 37062 3148
rect 36832 3108 36860 3136
rect 36464 3080 36860 3108
rect 36464 3049 36492 3080
rect 37458 3068 37464 3120
rect 37516 3068 37522 3120
rect 38746 3108 38752 3120
rect 38488 3080 38752 3108
rect 34655 3012 35940 3040
rect 35989 3043 36047 3049
rect 34655 3009 34667 3012
rect 34609 3003 34667 3009
rect 35989 3009 36001 3043
rect 36035 3009 36047 3043
rect 35989 3003 36047 3009
rect 36449 3043 36507 3049
rect 36449 3009 36461 3043
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 28592 2944 29377 2972
rect 28592 2932 28598 2944
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 29457 2975 29515 2981
rect 29457 2941 29469 2975
rect 29503 2972 29515 2975
rect 30745 2975 30803 2981
rect 30745 2972 30757 2975
rect 29503 2944 30757 2972
rect 29503 2941 29515 2944
rect 29457 2935 29515 2941
rect 30745 2941 30757 2944
rect 30791 2972 30803 2975
rect 30791 2944 30880 2972
rect 30791 2941 30803 2944
rect 30745 2935 30803 2941
rect 27890 2864 27896 2916
rect 27948 2904 27954 2916
rect 28905 2907 28963 2913
rect 27948 2876 28580 2904
rect 27948 2864 27954 2876
rect 27982 2836 27988 2848
rect 26620 2808 27988 2836
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 28350 2796 28356 2848
rect 28408 2796 28414 2848
rect 28552 2845 28580 2876
rect 28905 2873 28917 2907
rect 28951 2904 28963 2907
rect 28951 2876 29776 2904
rect 28951 2873 28963 2876
rect 28905 2867 28963 2873
rect 28537 2839 28595 2845
rect 28537 2805 28549 2839
rect 28583 2805 28595 2839
rect 28537 2799 28595 2805
rect 29178 2796 29184 2848
rect 29236 2836 29242 2848
rect 29454 2836 29460 2848
rect 29236 2808 29460 2836
rect 29236 2796 29242 2808
rect 29454 2796 29460 2808
rect 29512 2796 29518 2848
rect 29638 2796 29644 2848
rect 29696 2836 29702 2848
rect 29748 2836 29776 2876
rect 30098 2864 30104 2916
rect 30156 2904 30162 2916
rect 30852 2904 30880 2944
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 31665 2975 31723 2981
rect 31665 2972 31677 2975
rect 31352 2944 31677 2972
rect 31352 2932 31358 2944
rect 31665 2941 31677 2944
rect 31711 2941 31723 2975
rect 33704 2972 33732 3003
rect 31665 2935 31723 2941
rect 31772 2944 33732 2972
rect 34072 2972 34100 3003
rect 34514 2972 34520 2984
rect 34072 2944 34520 2972
rect 31478 2904 31484 2916
rect 30156 2876 30788 2904
rect 30852 2876 31484 2904
rect 30156 2864 30162 2876
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 29696 2808 30665 2836
rect 29696 2796 29702 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30760 2836 30788 2876
rect 31478 2864 31484 2876
rect 31536 2864 31542 2916
rect 31772 2904 31800 2944
rect 34514 2932 34520 2944
rect 34572 2932 34578 2984
rect 34793 2975 34851 2981
rect 34793 2941 34805 2975
rect 34839 2972 34851 2975
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 34839 2944 35541 2972
rect 34839 2941 34851 2944
rect 34793 2935 34851 2941
rect 35529 2941 35541 2944
rect 35575 2972 35587 2975
rect 35894 2972 35900 2984
rect 35575 2944 35900 2972
rect 35575 2941 35587 2944
rect 35529 2935 35587 2941
rect 35894 2932 35900 2944
rect 35952 2932 35958 2984
rect 33778 2904 33784 2916
rect 31588 2876 31800 2904
rect 33428 2876 33784 2904
rect 30834 2836 30840 2848
rect 30760 2808 30840 2836
rect 30653 2799 30711 2805
rect 30834 2796 30840 2808
rect 30892 2836 30898 2848
rect 31021 2839 31079 2845
rect 31021 2836 31033 2839
rect 30892 2808 31033 2836
rect 30892 2796 30898 2808
rect 31021 2805 31033 2808
rect 31067 2836 31079 2839
rect 31588 2836 31616 2876
rect 31067 2808 31616 2836
rect 31067 2805 31079 2808
rect 31021 2799 31079 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 33428 2845 33456 2876
rect 33778 2864 33784 2876
rect 33836 2864 33842 2916
rect 34149 2907 34207 2913
rect 34149 2873 34161 2907
rect 34195 2904 34207 2907
rect 36004 2904 36032 3003
rect 38286 3000 38292 3052
rect 38344 3040 38350 3052
rect 38488 3049 38516 3080
rect 38746 3068 38752 3080
rect 38804 3108 38810 3120
rect 39022 3108 39028 3120
rect 38804 3080 39028 3108
rect 38804 3068 38810 3080
rect 39022 3068 39028 3080
rect 39080 3068 39086 3120
rect 39390 3068 39396 3120
rect 39448 3068 39454 3120
rect 40052 3108 40080 3148
rect 40221 3145 40233 3179
rect 40267 3176 40279 3179
rect 40310 3176 40316 3188
rect 40267 3148 40316 3176
rect 40267 3145 40279 3148
rect 40221 3139 40279 3145
rect 40310 3136 40316 3148
rect 40368 3136 40374 3188
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 41969 3179 42027 3185
rect 41969 3176 41981 3179
rect 41932 3148 41981 3176
rect 41932 3136 41938 3148
rect 41969 3145 41981 3148
rect 42015 3176 42027 3179
rect 42705 3179 42763 3185
rect 42705 3176 42717 3179
rect 42015 3148 42717 3176
rect 42015 3145 42027 3148
rect 41969 3139 42027 3145
rect 42705 3145 42717 3148
rect 42751 3176 42763 3179
rect 43073 3179 43131 3185
rect 43073 3176 43085 3179
rect 42751 3148 43085 3176
rect 42751 3145 42763 3148
rect 42705 3139 42763 3145
rect 43073 3145 43085 3148
rect 43119 3145 43131 3179
rect 43073 3139 43131 3145
rect 44726 3136 44732 3188
rect 44784 3136 44790 3188
rect 40586 3108 40592 3120
rect 40052 3080 40592 3108
rect 40586 3068 40592 3080
rect 40644 3068 40650 3120
rect 41325 3111 41383 3117
rect 41325 3077 41337 3111
rect 41371 3108 41383 3111
rect 42242 3108 42248 3120
rect 41371 3080 42248 3108
rect 41371 3077 41383 3080
rect 41325 3071 41383 3077
rect 42242 3068 42248 3080
rect 42300 3108 42306 3120
rect 42337 3111 42395 3117
rect 42337 3108 42349 3111
rect 42300 3080 42349 3108
rect 42300 3068 42306 3080
rect 42337 3077 42349 3080
rect 42383 3077 42395 3111
rect 42337 3071 42395 3077
rect 38473 3043 38531 3049
rect 38473 3040 38485 3043
rect 38344 3012 38485 3040
rect 38344 3000 38350 3012
rect 38473 3009 38485 3012
rect 38519 3009 38531 3043
rect 38473 3003 38531 3009
rect 40126 3000 40132 3052
rect 40184 3000 40190 3052
rect 40681 3043 40739 3049
rect 40681 3009 40693 3043
rect 40727 3040 40739 3043
rect 41414 3040 41420 3052
rect 40727 3012 41420 3040
rect 40727 3009 40739 3012
rect 40681 3003 40739 3009
rect 41414 3000 41420 3012
rect 41472 3000 41478 3052
rect 43441 3043 43499 3049
rect 43441 3009 43453 3043
rect 43487 3040 43499 3043
rect 44634 3040 44640 3052
rect 43487 3012 44640 3040
rect 43487 3009 43499 3012
rect 43441 3003 43499 3009
rect 44634 3000 44640 3012
rect 44692 3000 44698 3052
rect 36354 2932 36360 2984
rect 36412 2972 36418 2984
rect 36633 2975 36691 2981
rect 36633 2972 36645 2975
rect 36412 2944 36645 2972
rect 36412 2932 36418 2944
rect 36633 2941 36645 2944
rect 36679 2941 36691 2975
rect 36909 2975 36967 2981
rect 36909 2972 36921 2975
rect 36633 2935 36691 2941
rect 36740 2944 36921 2972
rect 34195 2876 36032 2904
rect 36265 2907 36323 2913
rect 34195 2873 34207 2876
rect 34149 2867 34207 2873
rect 36265 2873 36277 2907
rect 36311 2904 36323 2907
rect 36740 2904 36768 2944
rect 36909 2941 36921 2944
rect 36955 2941 36967 2975
rect 36909 2935 36967 2941
rect 37274 2932 37280 2984
rect 37332 2972 37338 2984
rect 37332 2944 38148 2972
rect 37332 2932 37338 2944
rect 36311 2876 36768 2904
rect 38120 2904 38148 2944
rect 38746 2932 38752 2984
rect 38804 2932 38810 2984
rect 38381 2907 38439 2913
rect 38381 2904 38393 2907
rect 38120 2876 38393 2904
rect 36311 2873 36323 2876
rect 36265 2867 36323 2873
rect 38381 2873 38393 2876
rect 38427 2873 38439 2907
rect 40144 2904 40172 3000
rect 40494 2932 40500 2984
rect 40552 2972 40558 2984
rect 40773 2975 40831 2981
rect 40773 2972 40785 2975
rect 40552 2944 40785 2972
rect 40552 2932 40558 2944
rect 40773 2941 40785 2944
rect 40819 2941 40831 2975
rect 40773 2935 40831 2941
rect 40862 2932 40868 2984
rect 40920 2932 40926 2984
rect 40313 2907 40371 2913
rect 40313 2904 40325 2907
rect 40144 2876 40325 2904
rect 38381 2867 38439 2873
rect 40313 2873 40325 2876
rect 40359 2873 40371 2907
rect 40313 2867 40371 2873
rect 33413 2839 33471 2845
rect 33413 2836 33425 2839
rect 31720 2808 33425 2836
rect 31720 2796 31726 2808
rect 33413 2805 33425 2808
rect 33459 2805 33471 2839
rect 33413 2799 33471 2805
rect 33873 2839 33931 2845
rect 33873 2805 33885 2839
rect 33919 2836 33931 2839
rect 34054 2836 34060 2848
rect 33919 2808 34060 2836
rect 33919 2805 33931 2808
rect 33873 2799 33931 2805
rect 34054 2796 34060 2808
rect 34112 2796 34118 2848
rect 35802 2796 35808 2848
rect 35860 2796 35866 2848
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38286 2836 38292 2848
rect 36044 2808 38292 2836
rect 36044 2796 36050 2808
rect 38286 2796 38292 2808
rect 38344 2796 38350 2848
rect 38396 2836 38424 2867
rect 39390 2836 39396 2848
rect 38396 2808 39396 2836
rect 39390 2796 39396 2808
rect 39448 2796 39454 2848
rect 460 2746 45540 2768
rect 460 2694 3570 2746
rect 3622 2694 3634 2746
rect 3686 2694 3698 2746
rect 3750 2694 3762 2746
rect 3814 2694 3826 2746
rect 3878 2694 8570 2746
rect 8622 2694 8634 2746
rect 8686 2694 8698 2746
rect 8750 2694 8762 2746
rect 8814 2694 8826 2746
rect 8878 2694 13570 2746
rect 13622 2694 13634 2746
rect 13686 2694 13698 2746
rect 13750 2694 13762 2746
rect 13814 2694 13826 2746
rect 13878 2694 18570 2746
rect 18622 2694 18634 2746
rect 18686 2694 18698 2746
rect 18750 2694 18762 2746
rect 18814 2694 18826 2746
rect 18878 2694 23570 2746
rect 23622 2694 23634 2746
rect 23686 2694 23698 2746
rect 23750 2694 23762 2746
rect 23814 2694 23826 2746
rect 23878 2694 28570 2746
rect 28622 2694 28634 2746
rect 28686 2694 28698 2746
rect 28750 2694 28762 2746
rect 28814 2694 28826 2746
rect 28878 2694 33570 2746
rect 33622 2694 33634 2746
rect 33686 2694 33698 2746
rect 33750 2694 33762 2746
rect 33814 2694 33826 2746
rect 33878 2694 38570 2746
rect 38622 2694 38634 2746
rect 38686 2694 38698 2746
rect 38750 2694 38762 2746
rect 38814 2694 38826 2746
rect 38878 2694 43570 2746
rect 43622 2694 43634 2746
rect 43686 2694 43698 2746
rect 43750 2694 43762 2746
rect 43814 2694 43826 2746
rect 43878 2694 45540 2746
rect 460 2672 45540 2694
rect 1486 2592 1492 2644
rect 1544 2592 1550 2644
rect 1762 2592 1768 2644
rect 1820 2632 1826 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1820 2604 1961 2632
rect 1820 2592 1826 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 2774 2632 2780 2644
rect 1949 2595 2007 2601
rect 2746 2592 2780 2632
rect 2832 2592 2838 2644
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8536 2604 9137 2632
rect 8536 2592 8542 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 9508 2604 11376 2632
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 1581 2567 1639 2573
rect 1581 2564 1593 2567
rect 1360 2536 1593 2564
rect 1360 2524 1366 2536
rect 1581 2533 1593 2536
rect 1627 2533 1639 2567
rect 2746 2564 2774 2592
rect 1581 2527 1639 2533
rect 1780 2536 2774 2564
rect 1780 2437 1808 2536
rect 7006 2524 7012 2576
rect 7064 2524 7070 2576
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2464 2468 2789 2496
rect 2464 2456 2470 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 3142 2456 3148 2508
rect 3200 2456 3206 2508
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 9508 2496 9536 2604
rect 11348 2564 11376 2604
rect 11790 2592 11796 2644
rect 11848 2592 11854 2644
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 11940 2604 12173 2632
rect 11940 2592 11946 2604
rect 12161 2601 12173 2604
rect 12207 2632 12219 2635
rect 13265 2635 13323 2641
rect 12207 2604 12940 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 12618 2564 12624 2576
rect 11348 2536 12624 2564
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 12912 2573 12940 2604
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13311 2604 15884 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 14090 2564 14096 2576
rect 12943 2536 14096 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 15856 2564 15884 2604
rect 15930 2592 15936 2644
rect 15988 2632 15994 2644
rect 16025 2635 16083 2641
rect 16025 2632 16037 2635
rect 15988 2604 16037 2632
rect 15988 2592 15994 2604
rect 16025 2601 16037 2604
rect 16071 2632 16083 2635
rect 16482 2632 16488 2644
rect 16071 2604 16488 2632
rect 16071 2601 16083 2604
rect 16025 2595 16083 2601
rect 16482 2592 16488 2604
rect 16540 2592 16546 2644
rect 19426 2592 19432 2644
rect 19484 2592 19490 2644
rect 20346 2632 20352 2644
rect 19996 2604 20352 2632
rect 19996 2564 20024 2604
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 22554 2632 22560 2644
rect 22336 2604 22560 2632
rect 22336 2592 22342 2604
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 23569 2635 23627 2641
rect 23569 2601 23581 2635
rect 23615 2632 23627 2635
rect 24210 2632 24216 2644
rect 23615 2604 24216 2632
rect 23615 2601 23627 2604
rect 23569 2595 23627 2601
rect 24210 2592 24216 2604
rect 24268 2592 24274 2644
rect 25682 2592 25688 2644
rect 25740 2632 25746 2644
rect 25740 2604 27108 2632
rect 25740 2592 25746 2604
rect 15856 2536 16804 2564
rect 5491 2468 9536 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2179 2400 2268 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 1121 2295 1179 2301
rect 1121 2261 1133 2295
rect 1167 2292 1179 2295
rect 1670 2292 1676 2304
rect 1167 2264 1676 2292
rect 1167 2261 1179 2264
rect 1121 2255 1179 2261
rect 1670 2252 1676 2264
rect 1728 2252 1734 2304
rect 2240 2301 2268 2400
rect 2498 2388 2504 2440
rect 2556 2428 2562 2440
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2556 2400 2605 2428
rect 2556 2388 2562 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2958 2428 2964 2440
rect 2731 2400 2964 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 4706 2428 4712 2440
rect 4554 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 9508 2437 9536 2468
rect 9674 2456 9680 2508
rect 9732 2456 9738 2508
rect 9858 2456 9864 2508
rect 9916 2456 9922 2508
rect 14182 2496 14188 2508
rect 9968 2468 14188 2496
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9876 2428 9904 2456
rect 9631 2400 9904 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 3418 2320 3424 2372
rect 3476 2320 3482 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 9033 2363 9091 2369
rect 6963 2332 8984 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 2225 2295 2283 2301
rect 2225 2261 2237 2295
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4120 2264 4905 2292
rect 4120 2252 4126 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 5718 2252 5724 2304
rect 5776 2252 5782 2304
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6089 2295 6147 2301
rect 6089 2292 6101 2295
rect 6052 2264 6101 2292
rect 6052 2252 6058 2264
rect 6089 2261 6101 2264
rect 6135 2261 6147 2295
rect 6089 2255 6147 2261
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 6595 2264 7757 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 7745 2261 7757 2264
rect 7791 2292 7803 2295
rect 8110 2292 8116 2304
rect 7791 2264 8116 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 8570 2252 8576 2304
rect 8628 2252 8634 2304
rect 8956 2292 8984 2332
rect 9033 2329 9045 2363
rect 9079 2360 9091 2363
rect 9968 2360 9996 2468
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14918 2496 14924 2508
rect 14323 2468 14924 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14918 2456 14924 2468
rect 14976 2496 14982 2508
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 14976 2468 16497 2496
rect 14976 2456 14982 2468
rect 16485 2465 16497 2468
rect 16531 2496 16543 2499
rect 16666 2496 16672 2508
rect 16531 2468 16672 2496
rect 16531 2465 16543 2468
rect 16485 2459 16543 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 16776 2496 16804 2536
rect 17972 2536 20024 2564
rect 17972 2496 18000 2536
rect 16776 2468 18000 2496
rect 18417 2499 18475 2505
rect 18417 2465 18429 2499
rect 18463 2496 18475 2499
rect 18506 2496 18512 2508
rect 18463 2468 18512 2496
rect 18463 2465 18475 2468
rect 18417 2459 18475 2465
rect 18506 2456 18512 2468
rect 18564 2496 18570 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18564 2468 19073 2496
rect 18564 2456 18570 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 19242 2456 19248 2508
rect 19300 2456 19306 2508
rect 19702 2456 19708 2508
rect 19760 2456 19766 2508
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19852 2468 19901 2496
rect 19852 2456 19858 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 21174 2496 21180 2508
rect 19935 2468 21180 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21232 2468 21833 2496
rect 21232 2456 21238 2468
rect 21821 2465 21833 2468
rect 21867 2496 21879 2499
rect 24118 2496 24124 2508
rect 21867 2468 24124 2496
rect 21867 2465 21879 2468
rect 21821 2459 21879 2465
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 11882 2428 11888 2440
rect 11454 2400 11888 2428
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2428 13967 2431
rect 13998 2428 14004 2440
rect 13955 2400 14004 2428
rect 13955 2397 13967 2400
rect 13909 2391 13967 2397
rect 13998 2388 14004 2400
rect 14056 2428 14062 2440
rect 19613 2431 19671 2437
rect 14056 2400 14320 2428
rect 14056 2388 14062 2400
rect 14292 2372 14320 2400
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 19720 2428 19748 2456
rect 23768 2440 23796 2468
rect 24118 2456 24124 2468
rect 24176 2456 24182 2508
rect 25590 2456 25596 2508
rect 25648 2456 25654 2508
rect 25869 2499 25927 2505
rect 25869 2465 25881 2499
rect 25915 2496 25927 2499
rect 26326 2496 26332 2508
rect 25915 2468 26332 2496
rect 25915 2465 25927 2468
rect 25869 2459 25927 2465
rect 26326 2456 26332 2468
rect 26384 2456 26390 2508
rect 27080 2496 27108 2604
rect 27246 2592 27252 2644
rect 27304 2632 27310 2644
rect 27341 2635 27399 2641
rect 27341 2632 27353 2635
rect 27304 2604 27353 2632
rect 27304 2592 27310 2604
rect 27341 2601 27353 2604
rect 27387 2601 27399 2635
rect 27341 2595 27399 2601
rect 27522 2592 27528 2644
rect 27580 2592 27586 2644
rect 28261 2635 28319 2641
rect 28261 2601 28273 2635
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 27154 2524 27160 2576
rect 27212 2564 27218 2576
rect 27801 2567 27859 2573
rect 27801 2564 27813 2567
rect 27212 2536 27813 2564
rect 27212 2524 27218 2536
rect 27801 2533 27813 2536
rect 27847 2533 27859 2567
rect 28276 2564 28304 2595
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 29052 2604 29745 2632
rect 29052 2592 29058 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 29733 2595 29791 2601
rect 30745 2635 30803 2641
rect 30745 2601 30757 2635
rect 30791 2632 30803 2635
rect 33226 2632 33232 2644
rect 30791 2604 33232 2632
rect 30791 2601 30803 2604
rect 30745 2595 30803 2601
rect 33226 2592 33232 2604
rect 33284 2592 33290 2644
rect 34146 2632 34152 2644
rect 34072 2604 34152 2632
rect 28276 2536 28580 2564
rect 27801 2527 27859 2533
rect 27080 2468 27568 2496
rect 21542 2428 21548 2440
rect 19659 2400 19748 2428
rect 21298 2400 21548 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 23750 2388 23756 2440
rect 23808 2388 23814 2440
rect 26878 2388 26884 2440
rect 26936 2428 26942 2440
rect 26936 2400 27002 2428
rect 26936 2388 26942 2400
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 27540 2428 27568 2468
rect 27706 2456 27712 2508
rect 27764 2456 27770 2508
rect 28552 2440 28580 2536
rect 29362 2524 29368 2576
rect 29420 2524 29426 2576
rect 29457 2567 29515 2573
rect 29457 2533 29469 2567
rect 29503 2564 29515 2567
rect 30098 2564 30104 2576
rect 29503 2536 30104 2564
rect 29503 2533 29515 2536
rect 29457 2527 29515 2533
rect 30098 2524 30104 2536
rect 30156 2524 30162 2576
rect 30190 2524 30196 2576
rect 30248 2524 30254 2576
rect 31294 2564 31300 2576
rect 30576 2536 31300 2564
rect 28718 2456 28724 2508
rect 28776 2456 28782 2508
rect 30009 2499 30067 2505
rect 29472 2468 29960 2496
rect 29472 2440 29500 2468
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 27540 2400 27997 2428
rect 27985 2397 27997 2400
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 28442 2428 28448 2440
rect 28132 2400 28448 2428
rect 28132 2388 28138 2400
rect 28442 2388 28448 2400
rect 28500 2388 28506 2440
rect 28534 2388 28540 2440
rect 28592 2388 28598 2440
rect 28629 2431 28687 2437
rect 28629 2397 28641 2431
rect 28675 2428 28687 2431
rect 29089 2431 29147 2437
rect 29089 2428 29101 2431
rect 28675 2400 29101 2428
rect 28675 2397 28687 2400
rect 28629 2391 28687 2397
rect 29089 2397 29101 2400
rect 29135 2397 29147 2431
rect 29089 2391 29147 2397
rect 29273 2431 29331 2437
rect 29273 2397 29285 2431
rect 29319 2428 29331 2431
rect 29454 2428 29460 2440
rect 29319 2400 29460 2428
rect 29319 2397 29331 2400
rect 29273 2391 29331 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 29932 2437 29960 2468
rect 30009 2465 30021 2499
rect 30055 2496 30067 2499
rect 30208 2496 30236 2524
rect 30576 2508 30604 2536
rect 31294 2524 31300 2536
rect 31352 2564 31358 2576
rect 31352 2536 31616 2564
rect 31352 2524 31358 2536
rect 30055 2468 30236 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 29549 2431 29607 2437
rect 29549 2397 29561 2431
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 29917 2431 29975 2437
rect 29917 2397 29929 2431
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 9079 2332 9996 2360
rect 9079 2329 9091 2332
rect 9033 2323 9091 2329
rect 10318 2320 10324 2372
rect 10376 2320 10382 2372
rect 12437 2363 12495 2369
rect 12437 2360 12449 2363
rect 12360 2332 12449 2360
rect 12360 2304 12388 2332
rect 12437 2329 12449 2332
rect 12483 2329 12495 2363
rect 12437 2323 12495 2329
rect 14182 2320 14188 2372
rect 14240 2320 14246 2372
rect 14274 2320 14280 2372
rect 14332 2320 14338 2372
rect 14550 2320 14556 2372
rect 14608 2320 14614 2372
rect 15838 2360 15844 2372
rect 15778 2332 15844 2360
rect 15838 2320 15844 2332
rect 15896 2320 15902 2372
rect 16942 2320 16948 2372
rect 17000 2320 17006 2372
rect 17678 2320 17684 2372
rect 17736 2320 17742 2372
rect 18969 2363 19027 2369
rect 18969 2360 18981 2363
rect 18248 2332 18981 2360
rect 11330 2292 11336 2304
rect 8956 2264 11336 2292
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 12342 2252 12348 2304
rect 12400 2252 12406 2304
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13504 2264 13737 2292
rect 13504 2252 13510 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 14200 2292 14228 2320
rect 18248 2292 18276 2332
rect 18969 2329 18981 2332
rect 19015 2360 19027 2363
rect 19058 2360 19064 2372
rect 19015 2332 19064 2360
rect 19015 2329 19027 2332
rect 18969 2323 19027 2329
rect 19058 2320 19064 2332
rect 19116 2320 19122 2372
rect 20162 2320 20168 2372
rect 20220 2320 20226 2372
rect 21560 2360 21588 2388
rect 21560 2332 22048 2360
rect 14200 2264 18276 2292
rect 13725 2255 13783 2261
rect 18598 2252 18604 2304
rect 18656 2252 18662 2304
rect 21634 2252 21640 2304
rect 21692 2252 21698 2304
rect 22020 2292 22048 2332
rect 22094 2320 22100 2372
rect 22152 2320 22158 2372
rect 22480 2332 22586 2360
rect 22480 2292 22508 2332
rect 24026 2320 24032 2372
rect 24084 2320 24090 2372
rect 24762 2320 24768 2372
rect 24820 2320 24826 2372
rect 27522 2320 27528 2372
rect 27580 2360 27586 2372
rect 27709 2363 27767 2369
rect 27709 2360 27721 2363
rect 27580 2332 27721 2360
rect 27580 2320 27586 2332
rect 27709 2329 27721 2332
rect 27755 2329 27767 2363
rect 29564 2360 29592 2391
rect 30024 2372 30052 2459
rect 30558 2456 30564 2508
rect 30616 2456 30622 2508
rect 31202 2456 31208 2508
rect 31260 2456 31266 2508
rect 31389 2499 31447 2505
rect 31389 2465 31401 2499
rect 31435 2496 31447 2499
rect 31435 2468 31524 2496
rect 31435 2465 31447 2468
rect 31389 2459 31447 2465
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2428 30251 2431
rect 30282 2428 30288 2440
rect 30239 2400 30288 2428
rect 30239 2397 30251 2400
rect 30193 2391 30251 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30377 2431 30435 2437
rect 30377 2397 30389 2431
rect 30423 2428 30435 2431
rect 30650 2428 30656 2440
rect 30423 2400 30656 2428
rect 30423 2397 30435 2400
rect 30377 2391 30435 2397
rect 30650 2388 30656 2400
rect 30708 2388 30714 2440
rect 30006 2360 30012 2372
rect 29564 2332 30012 2360
rect 27709 2323 27767 2329
rect 30006 2320 30012 2332
rect 30064 2320 30070 2372
rect 31113 2363 31171 2369
rect 31113 2329 31125 2363
rect 31159 2360 31171 2363
rect 31386 2360 31392 2372
rect 31159 2332 31392 2360
rect 31159 2329 31171 2332
rect 31113 2323 31171 2329
rect 31386 2320 31392 2332
rect 31444 2320 31450 2372
rect 31496 2304 31524 2468
rect 31588 2437 31616 2536
rect 31849 2499 31907 2505
rect 31849 2465 31861 2499
rect 31895 2496 31907 2499
rect 32858 2496 32864 2508
rect 31895 2468 32864 2496
rect 31895 2465 31907 2468
rect 31849 2459 31907 2465
rect 32858 2456 32864 2468
rect 32916 2456 32922 2508
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2397 31631 2431
rect 31573 2391 31631 2397
rect 31588 2360 31616 2391
rect 32950 2388 32956 2440
rect 33008 2388 33014 2440
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33192 2400 33701 2428
rect 33192 2388 33198 2400
rect 33689 2397 33701 2400
rect 33735 2397 33747 2431
rect 33689 2391 33747 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34072 2437 34100 2604
rect 34146 2592 34152 2604
rect 34204 2632 34210 2644
rect 35805 2635 35863 2641
rect 34204 2604 35756 2632
rect 34204 2592 34210 2604
rect 34330 2456 34336 2508
rect 34388 2456 34394 2508
rect 34057 2431 34115 2437
rect 34057 2428 34069 2431
rect 33836 2400 34069 2428
rect 33836 2388 33842 2400
rect 34057 2397 34069 2400
rect 34103 2397 34115 2431
rect 35728 2428 35756 2604
rect 35805 2601 35817 2635
rect 35851 2632 35863 2635
rect 35894 2632 35900 2644
rect 35851 2604 35900 2632
rect 35851 2601 35863 2604
rect 35805 2595 35863 2601
rect 35894 2592 35900 2604
rect 35952 2592 35958 2644
rect 37274 2592 37280 2644
rect 37332 2632 37338 2644
rect 37642 2632 37648 2644
rect 37332 2604 37648 2632
rect 37332 2592 37338 2604
rect 37642 2592 37648 2604
rect 37700 2592 37706 2644
rect 38841 2635 38899 2641
rect 38841 2601 38853 2635
rect 38887 2632 38899 2635
rect 38930 2632 38936 2644
rect 38887 2604 38936 2632
rect 38887 2601 38899 2604
rect 38841 2595 38899 2601
rect 38930 2592 38936 2604
rect 38988 2592 38994 2644
rect 40402 2632 40408 2644
rect 39316 2604 40408 2632
rect 38565 2567 38623 2573
rect 38565 2564 38577 2567
rect 37660 2536 38577 2564
rect 35802 2456 35808 2508
rect 35860 2496 35866 2508
rect 36173 2499 36231 2505
rect 36173 2496 36185 2499
rect 35860 2468 36185 2496
rect 35860 2456 35866 2468
rect 36173 2465 36185 2468
rect 36219 2465 36231 2499
rect 36173 2459 36231 2465
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 37660 2496 37688 2536
rect 38565 2533 38577 2536
rect 38611 2533 38623 2567
rect 38565 2527 38623 2533
rect 39209 2567 39267 2573
rect 39209 2533 39221 2567
rect 39255 2533 39267 2567
rect 39209 2527 39267 2533
rect 36964 2468 37688 2496
rect 36964 2456 36970 2468
rect 38102 2456 38108 2508
rect 38160 2496 38166 2508
rect 38197 2499 38255 2505
rect 38197 2496 38209 2499
rect 38160 2468 38209 2496
rect 38160 2456 38166 2468
rect 38197 2465 38209 2468
rect 38243 2465 38255 2499
rect 38197 2459 38255 2465
rect 38286 2456 38292 2508
rect 38344 2456 38350 2508
rect 35897 2431 35955 2437
rect 35897 2428 35909 2431
rect 35728 2400 35909 2428
rect 34057 2391 34115 2397
rect 35897 2397 35909 2400
rect 35943 2397 35955 2431
rect 35897 2391 35955 2397
rect 31938 2360 31944 2372
rect 31588 2332 31944 2360
rect 31938 2320 31944 2332
rect 31996 2320 32002 2372
rect 35912 2360 35940 2391
rect 36446 2360 36452 2372
rect 35558 2332 35848 2360
rect 35912 2332 36452 2360
rect 22020 2264 22508 2292
rect 25406 2252 25412 2304
rect 25464 2292 25470 2304
rect 25501 2295 25559 2301
rect 25501 2292 25513 2295
rect 25464 2264 25513 2292
rect 25464 2252 25470 2264
rect 25501 2261 25513 2264
rect 25547 2261 25559 2295
rect 25501 2255 25559 2261
rect 27430 2252 27436 2304
rect 27488 2292 27494 2304
rect 29086 2292 29092 2304
rect 27488 2264 29092 2292
rect 27488 2252 27494 2264
rect 29086 2252 29092 2264
rect 29144 2252 29150 2304
rect 29178 2252 29184 2304
rect 29236 2292 29242 2304
rect 30561 2295 30619 2301
rect 30561 2292 30573 2295
rect 29236 2264 30573 2292
rect 29236 2252 29242 2264
rect 30561 2261 30573 2264
rect 30607 2261 30619 2295
rect 30561 2255 30619 2261
rect 31478 2252 31484 2304
rect 31536 2292 31542 2304
rect 33226 2292 33232 2304
rect 31536 2264 33232 2292
rect 31536 2252 31542 2264
rect 33226 2252 33232 2264
rect 33284 2292 33290 2304
rect 33321 2295 33379 2301
rect 33321 2292 33333 2295
rect 33284 2264 33333 2292
rect 33284 2252 33290 2264
rect 33321 2261 33333 2264
rect 33367 2261 33379 2295
rect 33321 2255 33379 2261
rect 33502 2252 33508 2304
rect 33560 2252 33566 2304
rect 35250 2252 35256 2304
rect 35308 2292 35314 2304
rect 35710 2292 35716 2304
rect 35308 2264 35716 2292
rect 35308 2252 35314 2264
rect 35710 2252 35716 2264
rect 35768 2252 35774 2304
rect 35820 2292 35848 2332
rect 36446 2320 36452 2332
rect 36504 2320 36510 2372
rect 37458 2360 37464 2372
rect 37398 2332 37464 2360
rect 37458 2320 37464 2332
rect 37516 2320 37522 2372
rect 37642 2320 37648 2372
rect 37700 2360 37706 2372
rect 38105 2363 38163 2369
rect 38105 2360 38117 2363
rect 37700 2332 38117 2360
rect 37700 2320 37706 2332
rect 38105 2329 38117 2332
rect 38151 2329 38163 2363
rect 38304 2360 38332 2456
rect 38378 2388 38384 2440
rect 38436 2428 38442 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38436 2400 38761 2428
rect 38436 2388 38442 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 39025 2431 39083 2437
rect 39025 2397 39037 2431
rect 39071 2428 39083 2431
rect 39224 2428 39252 2527
rect 39071 2400 39252 2428
rect 39071 2397 39083 2400
rect 39025 2391 39083 2397
rect 39316 2360 39344 2604
rect 40402 2592 40408 2604
rect 40460 2592 40466 2644
rect 41874 2592 41880 2644
rect 41932 2632 41938 2644
rect 42337 2635 42395 2641
rect 42337 2632 42349 2635
rect 41932 2604 42349 2632
rect 41932 2592 41938 2604
rect 42337 2601 42349 2604
rect 42383 2632 42395 2635
rect 42426 2632 42432 2644
rect 42383 2604 42432 2632
rect 42383 2601 42395 2604
rect 42337 2595 42395 2601
rect 42426 2592 42432 2604
rect 42484 2632 42490 2644
rect 43073 2635 43131 2641
rect 43073 2632 43085 2635
rect 42484 2604 43085 2632
rect 42484 2592 42490 2604
rect 43073 2601 43085 2604
rect 43119 2601 43131 2635
rect 43073 2595 43131 2601
rect 43346 2592 43352 2644
rect 43404 2632 43410 2644
rect 43717 2635 43775 2641
rect 43717 2632 43729 2635
rect 43404 2604 43729 2632
rect 43404 2592 43410 2604
rect 43717 2601 43729 2604
rect 43763 2601 43775 2635
rect 43717 2595 43775 2601
rect 39574 2524 39580 2576
rect 39632 2564 39638 2576
rect 39632 2536 40356 2564
rect 39632 2524 39638 2536
rect 39684 2505 39712 2536
rect 40328 2508 40356 2536
rect 39669 2499 39727 2505
rect 39669 2465 39681 2499
rect 39715 2465 39727 2499
rect 39669 2459 39727 2465
rect 39758 2456 39764 2508
rect 39816 2456 39822 2508
rect 40310 2456 40316 2508
rect 40368 2456 40374 2508
rect 40420 2496 40448 2592
rect 41969 2567 42027 2573
rect 41969 2533 41981 2567
rect 42015 2564 42027 2567
rect 42242 2564 42248 2576
rect 42015 2536 42248 2564
rect 42015 2533 42027 2536
rect 41969 2527 42027 2533
rect 42242 2524 42248 2536
rect 42300 2564 42306 2576
rect 42613 2567 42671 2573
rect 42613 2564 42625 2567
rect 42300 2536 42625 2564
rect 42300 2524 42306 2536
rect 42613 2533 42625 2536
rect 42659 2533 42671 2567
rect 42613 2527 42671 2533
rect 40589 2499 40647 2505
rect 40589 2496 40601 2499
rect 40420 2468 40601 2496
rect 40589 2465 40601 2468
rect 40635 2465 40647 2499
rect 40589 2459 40647 2465
rect 40862 2456 40868 2508
rect 40920 2496 40926 2508
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 40920 2468 41429 2496
rect 40920 2456 40926 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 43732 2496 43760 2595
rect 44174 2592 44180 2644
rect 44232 2592 44238 2644
rect 44726 2592 44732 2644
rect 44784 2632 44790 2644
rect 45005 2635 45063 2641
rect 45005 2632 45017 2635
rect 44784 2604 45017 2632
rect 44784 2592 44790 2604
rect 45005 2601 45017 2604
rect 45051 2601 45063 2635
rect 45005 2595 45063 2601
rect 43806 2496 43812 2508
rect 43732 2468 43812 2496
rect 41417 2459 41475 2465
rect 43806 2456 43812 2468
rect 43864 2496 43870 2508
rect 44545 2499 44603 2505
rect 44545 2496 44557 2499
rect 43864 2468 44557 2496
rect 43864 2456 43870 2468
rect 44545 2465 44557 2468
rect 44591 2465 44603 2499
rect 44545 2459 44603 2465
rect 39390 2388 39396 2440
rect 39448 2428 39454 2440
rect 39577 2431 39635 2437
rect 39577 2428 39589 2431
rect 39448 2400 39589 2428
rect 39448 2388 39454 2400
rect 39577 2397 39589 2400
rect 39623 2428 39635 2431
rect 40405 2431 40463 2437
rect 40405 2428 40417 2431
rect 39623 2400 40417 2428
rect 39623 2397 39635 2400
rect 39577 2391 39635 2397
rect 40405 2397 40417 2400
rect 40451 2397 40463 2431
rect 40405 2391 40463 2397
rect 39758 2360 39764 2372
rect 38304 2332 39764 2360
rect 38105 2323 38163 2329
rect 39758 2320 39764 2332
rect 39816 2320 39822 2372
rect 40126 2320 40132 2372
rect 40184 2360 40190 2372
rect 40497 2363 40555 2369
rect 40497 2360 40509 2363
rect 40184 2332 40509 2360
rect 40184 2320 40190 2332
rect 40497 2329 40509 2332
rect 40543 2360 40555 2363
rect 41325 2363 41383 2369
rect 41325 2360 41337 2363
rect 40543 2332 41337 2360
rect 40543 2329 40555 2332
rect 40497 2323 40555 2329
rect 41325 2329 41337 2332
rect 41371 2329 41383 2363
rect 41325 2323 41383 2329
rect 35894 2292 35900 2304
rect 35820 2264 35900 2292
rect 35894 2252 35900 2264
rect 35952 2292 35958 2304
rect 37476 2292 37504 2320
rect 35952 2264 37504 2292
rect 37737 2295 37795 2301
rect 35952 2252 35958 2264
rect 37737 2261 37749 2295
rect 37783 2292 37795 2295
rect 37826 2292 37832 2304
rect 37783 2264 37832 2292
rect 37783 2261 37795 2264
rect 37737 2255 37795 2261
rect 37826 2252 37832 2264
rect 37884 2252 37890 2304
rect 40037 2295 40095 2301
rect 40037 2261 40049 2295
rect 40083 2292 40095 2295
rect 40310 2292 40316 2304
rect 40083 2264 40316 2292
rect 40083 2261 40095 2264
rect 40037 2255 40095 2261
rect 40310 2252 40316 2264
rect 40368 2252 40374 2304
rect 40862 2252 40868 2304
rect 40920 2252 40926 2304
rect 40954 2252 40960 2304
rect 41012 2292 41018 2304
rect 41233 2295 41291 2301
rect 41233 2292 41245 2295
rect 41012 2264 41245 2292
rect 41012 2252 41018 2264
rect 41233 2261 41245 2264
rect 41279 2261 41291 2295
rect 41233 2255 41291 2261
rect 460 2202 45540 2224
rect 460 2150 6070 2202
rect 6122 2150 6134 2202
rect 6186 2150 6198 2202
rect 6250 2150 6262 2202
rect 6314 2150 6326 2202
rect 6378 2150 11070 2202
rect 11122 2150 11134 2202
rect 11186 2150 11198 2202
rect 11250 2150 11262 2202
rect 11314 2150 11326 2202
rect 11378 2150 16070 2202
rect 16122 2150 16134 2202
rect 16186 2150 16198 2202
rect 16250 2150 16262 2202
rect 16314 2150 16326 2202
rect 16378 2150 21070 2202
rect 21122 2150 21134 2202
rect 21186 2150 21198 2202
rect 21250 2150 21262 2202
rect 21314 2150 21326 2202
rect 21378 2150 26070 2202
rect 26122 2150 26134 2202
rect 26186 2150 26198 2202
rect 26250 2150 26262 2202
rect 26314 2150 26326 2202
rect 26378 2150 31070 2202
rect 31122 2150 31134 2202
rect 31186 2150 31198 2202
rect 31250 2150 31262 2202
rect 31314 2150 31326 2202
rect 31378 2150 36070 2202
rect 36122 2150 36134 2202
rect 36186 2150 36198 2202
rect 36250 2150 36262 2202
rect 36314 2150 36326 2202
rect 36378 2150 41070 2202
rect 41122 2150 41134 2202
rect 41186 2150 41198 2202
rect 41250 2150 41262 2202
rect 41314 2150 41326 2202
rect 41378 2150 45540 2202
rect 460 2128 45540 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 2041 2091 2099 2097
rect 2041 2088 2053 2091
rect 1728 2060 2053 2088
rect 1728 2048 1734 2060
rect 2041 2057 2053 2060
rect 2087 2088 2099 2091
rect 2222 2088 2228 2100
rect 2087 2060 2228 2088
rect 2087 2057 2099 2060
rect 2041 2051 2099 2057
rect 2222 2048 2228 2060
rect 2280 2048 2286 2100
rect 2958 2048 2964 2100
rect 3016 2048 3022 2100
rect 3329 2091 3387 2097
rect 3329 2057 3341 2091
rect 3375 2088 3387 2091
rect 3418 2088 3424 2100
rect 3375 2060 3424 2088
rect 3375 2057 3387 2060
rect 3329 2051 3387 2057
rect 3418 2048 3424 2060
rect 3476 2048 3482 2100
rect 4062 2048 4068 2100
rect 4120 2048 4126 2100
rect 4433 2091 4491 2097
rect 4433 2057 4445 2091
rect 4479 2088 4491 2091
rect 4706 2088 4712 2100
rect 4479 2060 4712 2088
rect 4479 2057 4491 2060
rect 4433 2051 4491 2057
rect 4706 2048 4712 2060
rect 4764 2048 4770 2100
rect 9858 2048 9864 2100
rect 9916 2048 9922 2100
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 10137 2091 10195 2097
rect 10137 2088 10149 2091
rect 10100 2060 10149 2088
rect 10100 2048 10106 2060
rect 10137 2057 10149 2060
rect 10183 2057 10195 2091
rect 10137 2051 10195 2057
rect 10318 2048 10324 2100
rect 10376 2088 10382 2100
rect 10873 2091 10931 2097
rect 10873 2088 10885 2091
rect 10376 2060 10885 2088
rect 10376 2048 10382 2060
rect 10873 2057 10885 2060
rect 10919 2057 10931 2091
rect 10873 2051 10931 2057
rect 11790 2048 11796 2100
rect 11848 2048 11854 2100
rect 11882 2048 11888 2100
rect 11940 2048 11946 2100
rect 12434 2048 12440 2100
rect 12492 2088 12498 2100
rect 12492 2060 12848 2088
rect 12492 2048 12498 2060
rect 2314 1912 2320 1964
rect 2372 1912 2378 1964
rect 2869 1955 2927 1961
rect 2869 1921 2881 1955
rect 2915 1952 2927 1955
rect 2976 1952 3004 2048
rect 2915 1924 3004 1952
rect 2915 1921 2927 1924
rect 2869 1915 2927 1921
rect 3510 1912 3516 1964
rect 3568 1912 3574 1964
rect 3973 1955 4031 1961
rect 3973 1921 3985 1955
rect 4019 1952 4031 1955
rect 4080 1952 4108 2048
rect 9876 2020 9904 2048
rect 11422 2020 11428 2032
rect 9140 1992 9904 2020
rect 11072 1992 11428 2020
rect 4019 1924 4108 1952
rect 4019 1921 4031 1924
rect 3973 1915 4031 1921
rect 4706 1912 4712 1964
rect 4764 1912 4770 1964
rect 5350 1912 5356 1964
rect 5408 1912 5414 1964
rect 6365 1955 6423 1961
rect 6365 1921 6377 1955
rect 6411 1952 6423 1955
rect 6730 1952 6736 1964
rect 6411 1924 6736 1952
rect 6411 1921 6423 1924
rect 6365 1915 6423 1921
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1952 7987 1955
rect 8294 1952 8300 1964
rect 7975 1924 8300 1952
rect 7975 1921 7987 1924
rect 7929 1915 7987 1921
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 9140 1961 9168 1992
rect 9125 1955 9183 1961
rect 9125 1921 9137 1955
rect 9171 1921 9183 1955
rect 9125 1915 9183 1921
rect 9861 1955 9919 1961
rect 9861 1921 9873 1955
rect 9907 1952 9919 1955
rect 10410 1952 10416 1964
rect 9907 1924 10416 1952
rect 9907 1921 9919 1924
rect 9861 1915 9919 1921
rect 10410 1912 10416 1924
rect 10468 1912 10474 1964
rect 10502 1912 10508 1964
rect 10560 1912 10566 1964
rect 11072 1961 11100 1992
rect 11422 1980 11428 1992
rect 11480 1980 11486 2032
rect 11057 1955 11115 1961
rect 11057 1921 11069 1955
rect 11103 1921 11115 1955
rect 11057 1915 11115 1921
rect 11333 1955 11391 1961
rect 11333 1921 11345 1955
rect 11379 1952 11391 1955
rect 11808 1952 11836 2048
rect 11379 1924 11836 1952
rect 11379 1921 11391 1924
rect 11333 1915 11391 1921
rect 3142 1844 3148 1896
rect 3200 1884 3206 1896
rect 3237 1887 3295 1893
rect 3237 1884 3249 1887
rect 3200 1856 3249 1884
rect 3200 1844 3206 1856
rect 3237 1853 3249 1856
rect 3283 1884 3295 1887
rect 5077 1887 5135 1893
rect 5077 1884 5089 1887
rect 3283 1856 5089 1884
rect 3283 1853 3295 1856
rect 3237 1847 3295 1853
rect 5077 1853 5089 1856
rect 5123 1884 5135 1887
rect 5994 1884 6000 1896
rect 5123 1856 6000 1884
rect 5123 1853 5135 1856
rect 5077 1847 5135 1853
rect 5994 1844 6000 1856
rect 6052 1884 6058 1896
rect 6089 1887 6147 1893
rect 6089 1884 6101 1887
rect 6052 1856 6101 1884
rect 6052 1844 6058 1856
rect 6089 1853 6101 1856
rect 6135 1884 6147 1887
rect 6917 1887 6975 1893
rect 6917 1884 6929 1887
rect 6135 1856 6929 1884
rect 6135 1853 6147 1856
rect 6089 1847 6147 1853
rect 6917 1853 6929 1856
rect 6963 1884 6975 1887
rect 7653 1887 7711 1893
rect 7653 1884 7665 1887
rect 6963 1856 7665 1884
rect 6963 1853 6975 1856
rect 6917 1847 6975 1853
rect 7653 1853 7665 1856
rect 7699 1884 7711 1887
rect 8481 1887 8539 1893
rect 8481 1884 8493 1887
rect 7699 1856 8493 1884
rect 7699 1853 7711 1856
rect 7653 1847 7711 1853
rect 8481 1853 8493 1856
rect 8527 1884 8539 1887
rect 8570 1884 8576 1896
rect 8527 1856 8576 1884
rect 8527 1853 8539 1856
rect 8481 1847 8539 1853
rect 8570 1844 8576 1856
rect 8628 1884 8634 1896
rect 8849 1887 8907 1893
rect 8849 1884 8861 1887
rect 8628 1856 8861 1884
rect 8628 1844 8634 1856
rect 8849 1853 8861 1856
rect 8895 1884 8907 1887
rect 9214 1884 9220 1896
rect 8895 1856 9220 1884
rect 8895 1853 8907 1856
rect 8849 1847 8907 1853
rect 9214 1844 9220 1856
rect 9272 1844 9278 1896
rect 7285 1819 7343 1825
rect 7285 1785 7297 1819
rect 7331 1816 7343 1819
rect 8110 1816 8116 1828
rect 7331 1788 8116 1816
rect 7331 1785 7343 1788
rect 7285 1779 7343 1785
rect 8110 1776 8116 1788
rect 8168 1816 8174 1828
rect 9585 1819 9643 1825
rect 9585 1816 9597 1819
rect 8168 1788 9597 1816
rect 8168 1776 8174 1788
rect 9585 1785 9597 1788
rect 9631 1816 9643 1819
rect 9950 1816 9956 1828
rect 9631 1788 9956 1816
rect 9631 1785 9643 1788
rect 9585 1779 9643 1785
rect 9950 1776 9956 1788
rect 10008 1816 10014 1828
rect 11900 1816 11928 2048
rect 12820 2029 12848 2060
rect 14274 2048 14280 2100
rect 14332 2048 14338 2100
rect 15930 2048 15936 2100
rect 15988 2048 15994 2100
rect 16942 2048 16948 2100
rect 17000 2088 17006 2100
rect 17773 2091 17831 2097
rect 17773 2088 17785 2091
rect 17000 2060 17785 2088
rect 17000 2048 17006 2060
rect 17773 2057 17785 2060
rect 17819 2057 17831 2091
rect 17773 2051 17831 2057
rect 18598 2048 18604 2100
rect 18656 2048 18662 2100
rect 19150 2048 19156 2100
rect 19208 2048 19214 2100
rect 19242 2048 19248 2100
rect 19300 2048 19306 2100
rect 19613 2091 19671 2097
rect 19613 2057 19625 2091
rect 19659 2088 19671 2091
rect 19794 2088 19800 2100
rect 19659 2060 19800 2088
rect 19659 2057 19671 2060
rect 19613 2051 19671 2057
rect 19794 2048 19800 2060
rect 19852 2048 19858 2100
rect 20162 2048 20168 2100
rect 20220 2088 20226 2100
rect 20441 2091 20499 2097
rect 20441 2088 20453 2091
rect 20220 2060 20453 2088
rect 20220 2048 20226 2060
rect 20441 2057 20453 2060
rect 20487 2057 20499 2091
rect 20441 2051 20499 2057
rect 21177 2091 21235 2097
rect 21177 2057 21189 2091
rect 21223 2057 21235 2091
rect 21177 2051 21235 2057
rect 12805 2023 12863 2029
rect 12360 1992 12572 2020
rect 12360 1964 12388 1992
rect 12158 1912 12164 1964
rect 12216 1912 12222 1964
rect 12342 1912 12348 1964
rect 12400 1912 12406 1964
rect 12434 1912 12440 1964
rect 12492 1912 12498 1964
rect 12544 1961 12572 1992
rect 12805 1989 12817 2023
rect 12851 1989 12863 2023
rect 14090 2020 14096 2032
rect 14030 1992 14096 2020
rect 12805 1983 12863 1989
rect 14090 1980 14096 1992
rect 14148 1980 14154 2032
rect 12529 1955 12587 1961
rect 12529 1921 12541 1955
rect 12575 1921 12587 1955
rect 12529 1915 12587 1921
rect 12544 1884 12572 1915
rect 14550 1912 14556 1964
rect 14608 1912 14614 1964
rect 15565 1955 15623 1961
rect 15565 1921 15577 1955
rect 15611 1952 15623 1955
rect 15948 1952 15976 2048
rect 16853 2023 16911 2029
rect 16853 1989 16865 2023
rect 16899 2020 16911 2023
rect 17034 2020 17040 2032
rect 16899 1992 17040 2020
rect 16899 1989 16911 1992
rect 16853 1983 16911 1989
rect 17034 1980 17040 1992
rect 17092 2020 17098 2032
rect 17678 2020 17684 2032
rect 17092 1992 17684 2020
rect 17092 1980 17098 1992
rect 17678 1980 17684 1992
rect 17736 1980 17742 2032
rect 18616 2020 18644 2048
rect 17972 1992 18644 2020
rect 15611 1924 15976 1952
rect 16393 1955 16451 1961
rect 15611 1921 15623 1924
rect 15565 1915 15623 1921
rect 16393 1921 16405 1955
rect 16439 1952 16451 1955
rect 16574 1952 16580 1964
rect 16439 1924 16580 1952
rect 16439 1921 16451 1924
rect 16393 1915 16451 1921
rect 16574 1912 16580 1924
rect 16632 1912 16638 1964
rect 16666 1912 16672 1964
rect 16724 1952 16730 1964
rect 17972 1961 18000 1992
rect 17221 1955 17279 1961
rect 17221 1952 17233 1955
rect 16724 1924 17233 1952
rect 16724 1912 16730 1924
rect 17221 1921 17233 1924
rect 17267 1921 17279 1955
rect 17221 1915 17279 1921
rect 17405 1955 17463 1961
rect 17405 1921 17417 1955
rect 17451 1921 17463 1955
rect 17405 1915 17463 1921
rect 17957 1955 18015 1961
rect 17957 1921 17969 1955
rect 18003 1921 18015 1955
rect 17957 1915 18015 1921
rect 14918 1884 14924 1896
rect 12544 1856 14924 1884
rect 14918 1844 14924 1856
rect 14976 1884 14982 1896
rect 15197 1887 15255 1893
rect 15197 1884 15209 1887
rect 14976 1856 15209 1884
rect 14976 1844 14982 1856
rect 15197 1853 15209 1856
rect 15243 1853 15255 1887
rect 17420 1884 17448 1915
rect 18506 1912 18512 1964
rect 18564 1912 18570 1964
rect 18877 1955 18935 1961
rect 18877 1921 18889 1955
rect 18923 1952 18935 1955
rect 19168 1952 19196 2048
rect 21192 2020 21220 2051
rect 21634 2048 21640 2100
rect 21692 2048 21698 2100
rect 22094 2048 22100 2100
rect 22152 2088 22158 2100
rect 22465 2091 22523 2097
rect 22465 2088 22477 2091
rect 22152 2060 22477 2088
rect 22152 2048 22158 2060
rect 22465 2057 22477 2060
rect 22511 2057 22523 2091
rect 23750 2088 23756 2100
rect 22465 2051 22523 2057
rect 22756 2060 23756 2088
rect 20640 1992 21220 2020
rect 18923 1924 19196 1952
rect 18923 1921 18935 1924
rect 18877 1915 18935 1921
rect 19886 1912 19892 1964
rect 19944 1912 19950 1964
rect 20640 1961 20668 1992
rect 20349 1955 20407 1961
rect 20349 1921 20361 1955
rect 20395 1921 20407 1955
rect 20349 1915 20407 1921
rect 20625 1955 20683 1961
rect 20625 1921 20637 1955
rect 20671 1921 20683 1955
rect 20625 1915 20683 1921
rect 18233 1887 18291 1893
rect 18233 1884 18245 1887
rect 17420 1856 18245 1884
rect 15197 1847 15255 1853
rect 18233 1853 18245 1856
rect 18279 1853 18291 1887
rect 20364 1884 20392 1915
rect 20990 1912 20996 1964
rect 21048 1912 21054 1964
rect 21542 1912 21548 1964
rect 21600 1912 21606 1964
rect 21652 1884 21680 2048
rect 22373 1955 22431 1961
rect 22373 1921 22385 1955
rect 22419 1952 22431 1955
rect 22554 1952 22560 1964
rect 22419 1924 22560 1952
rect 22419 1921 22431 1924
rect 22373 1915 22431 1921
rect 22554 1912 22560 1924
rect 22612 1912 22618 1964
rect 22756 1961 22784 2060
rect 23750 2048 23756 2060
rect 23808 2048 23814 2100
rect 24026 2048 24032 2100
rect 24084 2088 24090 2100
rect 25133 2091 25191 2097
rect 25133 2088 25145 2091
rect 24084 2060 25145 2088
rect 24084 2048 24090 2060
rect 25133 2057 25145 2060
rect 25179 2057 25191 2091
rect 27614 2088 27620 2100
rect 25133 2051 25191 2057
rect 25332 2060 27620 2088
rect 23014 1980 23020 2032
rect 23072 1980 23078 2032
rect 24762 2020 24768 2032
rect 24242 1992 24768 2020
rect 24762 1980 24768 1992
rect 24820 1980 24826 2032
rect 22649 1955 22707 1961
rect 22649 1921 22661 1955
rect 22695 1921 22707 1955
rect 22649 1915 22707 1921
rect 22741 1955 22799 1961
rect 22741 1921 22753 1955
rect 22787 1921 22799 1955
rect 22741 1915 22799 1921
rect 20364 1856 21680 1884
rect 21821 1887 21879 1893
rect 18233 1847 18291 1853
rect 21821 1853 21833 1887
rect 21867 1884 21879 1887
rect 21910 1884 21916 1896
rect 21867 1856 21916 1884
rect 21867 1853 21879 1856
rect 21821 1847 21879 1853
rect 21910 1844 21916 1856
rect 21968 1844 21974 1896
rect 22664 1884 22692 1915
rect 24486 1912 24492 1964
rect 24544 1952 24550 1964
rect 25332 1961 25360 2060
rect 27614 2048 27620 2060
rect 27672 2048 27678 2100
rect 28074 2048 28080 2100
rect 28132 2088 28138 2100
rect 29917 2091 29975 2097
rect 28132 2060 29592 2088
rect 28132 2048 28138 2060
rect 25682 1980 25688 2032
rect 25740 2020 25746 2032
rect 25740 1992 26372 2020
rect 25740 1980 25746 1992
rect 24673 1955 24731 1961
rect 24673 1952 24685 1955
rect 24544 1924 24685 1952
rect 24544 1912 24550 1924
rect 24673 1921 24685 1924
rect 24719 1921 24731 1955
rect 24673 1915 24731 1921
rect 25317 1955 25375 1961
rect 25317 1921 25329 1955
rect 25363 1921 25375 1955
rect 25317 1915 25375 1921
rect 25406 1912 25412 1964
rect 25464 1912 25470 1964
rect 25590 1912 25596 1964
rect 25648 1912 25654 1964
rect 26344 1961 26372 1992
rect 26878 1980 26884 2032
rect 26936 2020 26942 2032
rect 26936 1992 27094 2020
rect 26936 1980 26942 1992
rect 29564 1964 29592 2060
rect 29917 2057 29929 2091
rect 29963 2088 29975 2091
rect 30006 2088 30012 2100
rect 29963 2060 30012 2088
rect 29963 2057 29975 2060
rect 29917 2051 29975 2057
rect 30006 2048 30012 2060
rect 30064 2048 30070 2100
rect 30926 2048 30932 2100
rect 30984 2088 30990 2100
rect 31113 2091 31171 2097
rect 31113 2088 31125 2091
rect 30984 2060 31125 2088
rect 30984 2048 30990 2060
rect 31113 2057 31125 2060
rect 31159 2057 31171 2091
rect 31113 2051 31171 2057
rect 31846 2048 31852 2100
rect 31904 2088 31910 2100
rect 33502 2088 33508 2100
rect 31904 2060 33508 2088
rect 31904 2048 31910 2060
rect 33502 2048 33508 2060
rect 33560 2048 33566 2100
rect 34072 2060 35480 2088
rect 32306 2020 32312 2032
rect 30024 1992 32312 2020
rect 26053 1955 26111 1961
rect 26053 1952 26065 1955
rect 25700 1924 26065 1952
rect 23658 1884 23664 1896
rect 22664 1856 23664 1884
rect 23658 1844 23664 1856
rect 23716 1844 23722 1896
rect 25424 1884 25452 1912
rect 25148 1856 25452 1884
rect 25148 1828 25176 1856
rect 10008 1788 11928 1816
rect 14936 1788 20944 1816
rect 10008 1776 10014 1788
rect 1210 1708 1216 1760
rect 1268 1708 1274 1760
rect 2130 1708 2136 1760
rect 2188 1708 2194 1760
rect 2685 1751 2743 1757
rect 2685 1717 2697 1751
rect 2731 1748 2743 1751
rect 2958 1748 2964 1760
rect 2731 1720 2964 1748
rect 2731 1717 2743 1720
rect 2685 1711 2743 1717
rect 2958 1708 2964 1720
rect 3016 1708 3022 1760
rect 3789 1751 3847 1757
rect 3789 1717 3801 1751
rect 3835 1748 3847 1751
rect 3970 1748 3976 1760
rect 3835 1720 3976 1748
rect 3835 1717 3847 1720
rect 3789 1711 3847 1717
rect 3970 1708 3976 1720
rect 4028 1708 4034 1760
rect 4522 1708 4528 1760
rect 4580 1708 4586 1760
rect 5166 1708 5172 1760
rect 5224 1708 5230 1760
rect 6178 1708 6184 1760
rect 6236 1708 6242 1760
rect 7742 1708 7748 1760
rect 7800 1708 7806 1760
rect 8938 1708 8944 1760
rect 8996 1708 9002 1760
rect 9674 1708 9680 1760
rect 9732 1708 9738 1760
rect 10318 1708 10324 1760
rect 10376 1708 10382 1760
rect 11146 1708 11152 1760
rect 11204 1708 11210 1760
rect 11974 1708 11980 1760
rect 12032 1708 12038 1760
rect 12250 1708 12256 1760
rect 12308 1708 12314 1760
rect 14366 1708 14372 1760
rect 14424 1708 14430 1760
rect 14936 1757 14964 1788
rect 14921 1751 14979 1757
rect 14921 1717 14933 1751
rect 14967 1717 14979 1751
rect 14921 1711 14979 1717
rect 15378 1708 15384 1760
rect 15436 1708 15442 1760
rect 16206 1708 16212 1760
rect 16264 1708 16270 1760
rect 17586 1708 17592 1760
rect 17644 1708 17650 1760
rect 18322 1708 18328 1760
rect 18380 1708 18386 1760
rect 18414 1708 18420 1760
rect 18472 1748 18478 1760
rect 18693 1751 18751 1757
rect 18693 1748 18705 1751
rect 18472 1720 18705 1748
rect 18472 1708 18478 1720
rect 18693 1717 18705 1720
rect 18739 1717 18751 1751
rect 18693 1711 18751 1717
rect 19702 1708 19708 1760
rect 19760 1708 19766 1760
rect 20162 1708 20168 1760
rect 20220 1708 20226 1760
rect 20806 1708 20812 1760
rect 20864 1708 20870 1760
rect 20916 1748 20944 1788
rect 22066 1788 22416 1816
rect 22066 1748 22094 1788
rect 22388 1760 22416 1788
rect 24302 1776 24308 1828
rect 24360 1776 24366 1828
rect 24394 1776 24400 1828
rect 24452 1816 24458 1828
rect 24857 1819 24915 1825
rect 24857 1816 24869 1819
rect 24452 1788 24869 1816
rect 24452 1776 24458 1788
rect 24857 1785 24869 1788
rect 24903 1785 24915 1819
rect 24857 1779 24915 1785
rect 25130 1776 25136 1828
rect 25188 1776 25194 1828
rect 20916 1720 22094 1748
rect 22186 1708 22192 1760
rect 22244 1708 22250 1760
rect 22370 1708 22376 1760
rect 22428 1708 22434 1760
rect 24320 1748 24348 1776
rect 24489 1751 24547 1757
rect 24489 1748 24501 1751
rect 24320 1720 24501 1748
rect 24489 1717 24501 1720
rect 24535 1748 24547 1751
rect 25700 1748 25728 1924
rect 26053 1921 26065 1924
rect 26099 1921 26111 1955
rect 26053 1915 26111 1921
rect 26329 1955 26387 1961
rect 26329 1921 26341 1955
rect 26375 1921 26387 1955
rect 26329 1915 26387 1921
rect 27982 1912 27988 1964
rect 28040 1952 28046 1964
rect 28169 1955 28227 1961
rect 28169 1952 28181 1955
rect 28040 1924 28181 1952
rect 28040 1912 28046 1924
rect 28169 1921 28181 1924
rect 28215 1921 28227 1955
rect 28169 1915 28227 1921
rect 26605 1887 26663 1893
rect 26605 1853 26617 1887
rect 26651 1884 26663 1887
rect 27890 1884 27896 1896
rect 26651 1856 27896 1884
rect 26651 1853 26663 1856
rect 26605 1847 26663 1853
rect 27890 1844 27896 1856
rect 27948 1844 27954 1896
rect 28184 1884 28212 1915
rect 29546 1912 29552 1964
rect 29604 1912 29610 1964
rect 29730 1912 29736 1964
rect 29788 1952 29794 1964
rect 30024 1961 30052 1992
rect 30576 1961 30604 1992
rect 32306 1980 32312 1992
rect 32364 1980 32370 2032
rect 34072 2020 34100 2060
rect 33442 2006 34100 2020
rect 33428 1992 34100 2006
rect 30009 1955 30067 1961
rect 30009 1952 30021 1955
rect 29788 1924 30021 1952
rect 29788 1912 29794 1924
rect 30009 1921 30021 1924
rect 30055 1921 30067 1955
rect 30009 1915 30067 1921
rect 30561 1955 30619 1961
rect 30561 1921 30573 1955
rect 30607 1921 30619 1955
rect 31297 1955 31355 1961
rect 31297 1952 31309 1955
rect 30561 1915 30619 1921
rect 30668 1924 31309 1952
rect 28445 1887 28503 1893
rect 28184 1856 28304 1884
rect 25777 1819 25835 1825
rect 25777 1785 25789 1819
rect 25823 1816 25835 1819
rect 25823 1788 26464 1816
rect 25823 1785 25835 1788
rect 25777 1779 25835 1785
rect 24535 1720 25728 1748
rect 25869 1751 25927 1757
rect 24535 1717 24547 1720
rect 24489 1711 24547 1717
rect 25869 1717 25881 1751
rect 25915 1748 25927 1751
rect 26234 1748 26240 1760
rect 25915 1720 26240 1748
rect 25915 1717 25927 1720
rect 25869 1711 25927 1717
rect 26234 1708 26240 1720
rect 26292 1708 26298 1760
rect 26436 1748 26464 1788
rect 27632 1788 28212 1816
rect 27632 1748 27660 1788
rect 28184 1760 28212 1788
rect 26436 1720 27660 1748
rect 28074 1708 28080 1760
rect 28132 1708 28138 1760
rect 28166 1708 28172 1760
rect 28224 1708 28230 1760
rect 28276 1748 28304 1856
rect 28445 1853 28457 1887
rect 28491 1884 28503 1887
rect 28534 1884 28540 1896
rect 28491 1856 28540 1884
rect 28491 1853 28503 1856
rect 28445 1847 28503 1853
rect 28534 1844 28540 1856
rect 28592 1844 28598 1896
rect 29914 1844 29920 1896
rect 29972 1884 29978 1896
rect 30668 1884 30696 1924
rect 31297 1921 31309 1924
rect 31343 1921 31355 1955
rect 31297 1915 31355 1921
rect 31481 1955 31539 1961
rect 31481 1921 31493 1955
rect 31527 1952 31539 1955
rect 31846 1952 31852 1964
rect 31527 1924 31852 1952
rect 31527 1921 31539 1924
rect 31481 1915 31539 1921
rect 31846 1912 31852 1924
rect 31904 1912 31910 1964
rect 31938 1912 31944 1964
rect 31996 1912 32002 1964
rect 29972 1856 30696 1884
rect 31021 1887 31079 1893
rect 29972 1844 29978 1856
rect 31021 1853 31033 1887
rect 31067 1884 31079 1887
rect 31067 1856 31892 1884
rect 31067 1853 31079 1856
rect 31021 1847 31079 1853
rect 30558 1816 30564 1828
rect 29932 1788 30564 1816
rect 29932 1748 29960 1788
rect 30558 1776 30564 1788
rect 30616 1776 30622 1828
rect 31570 1816 31576 1828
rect 30760 1788 31576 1816
rect 28276 1720 29960 1748
rect 30006 1708 30012 1760
rect 30064 1748 30070 1760
rect 30101 1751 30159 1757
rect 30101 1748 30113 1751
rect 30064 1720 30113 1748
rect 30064 1708 30070 1720
rect 30101 1717 30113 1720
rect 30147 1717 30159 1751
rect 30101 1711 30159 1717
rect 30466 1708 30472 1760
rect 30524 1708 30530 1760
rect 30760 1757 30788 1788
rect 31570 1776 31576 1788
rect 31628 1776 31634 1828
rect 30745 1751 30803 1757
rect 30745 1717 30757 1751
rect 30791 1717 30803 1751
rect 30745 1711 30803 1717
rect 30834 1708 30840 1760
rect 30892 1748 30898 1760
rect 31665 1751 31723 1757
rect 31665 1748 31677 1751
rect 30892 1720 31677 1748
rect 30892 1708 30898 1720
rect 31665 1717 31677 1720
rect 31711 1717 31723 1751
rect 31864 1748 31892 1856
rect 32214 1844 32220 1896
rect 32272 1844 32278 1896
rect 32950 1844 32956 1896
rect 33008 1884 33014 1896
rect 33428 1884 33456 1992
rect 34146 1980 34152 2032
rect 34204 1980 34210 2032
rect 35452 2020 35480 2060
rect 35526 2048 35532 2100
rect 35584 2088 35590 2100
rect 35713 2091 35771 2097
rect 35713 2088 35725 2091
rect 35584 2060 35725 2088
rect 35584 2048 35590 2060
rect 35713 2057 35725 2060
rect 35759 2057 35771 2091
rect 35713 2051 35771 2057
rect 35894 2048 35900 2100
rect 35952 2048 35958 2100
rect 36081 2091 36139 2097
rect 36081 2057 36093 2091
rect 36127 2088 36139 2091
rect 36127 2060 38240 2088
rect 36127 2057 36139 2060
rect 36081 2051 36139 2057
rect 35912 2020 35940 2048
rect 35374 1992 35940 2020
rect 37458 1980 37464 2032
rect 37516 1980 37522 2032
rect 38212 2020 38240 2060
rect 39022 2048 39028 2100
rect 39080 2048 39086 2100
rect 39482 2048 39488 2100
rect 39540 2048 39546 2100
rect 40034 2048 40040 2100
rect 40092 2088 40098 2100
rect 40494 2088 40500 2100
rect 40092 2060 40500 2088
rect 40092 2048 40098 2060
rect 40494 2048 40500 2060
rect 40552 2088 40558 2100
rect 40589 2091 40647 2097
rect 40589 2088 40601 2091
rect 40552 2060 40601 2088
rect 40552 2048 40558 2060
rect 40589 2057 40601 2060
rect 40635 2057 40647 2091
rect 40589 2051 40647 2057
rect 40678 2048 40684 2100
rect 40736 2048 40742 2100
rect 42061 2091 42119 2097
rect 42061 2057 42073 2091
rect 42107 2088 42119 2091
rect 42242 2088 42248 2100
rect 42107 2060 42248 2088
rect 42107 2057 42119 2060
rect 42061 2051 42119 2057
rect 42242 2048 42248 2060
rect 42300 2088 42306 2100
rect 42705 2091 42763 2097
rect 42705 2088 42717 2091
rect 42300 2060 42717 2088
rect 42300 2048 42306 2060
rect 42705 2057 42717 2060
rect 42751 2088 42763 2091
rect 42978 2088 42984 2100
rect 42751 2060 42984 2088
rect 42751 2057 42763 2060
rect 42705 2051 42763 2057
rect 42978 2048 42984 2060
rect 43036 2048 43042 2100
rect 43806 2048 43812 2100
rect 43864 2088 43870 2100
rect 44177 2091 44235 2097
rect 44177 2088 44189 2091
rect 43864 2060 44189 2088
rect 43864 2048 43870 2060
rect 44177 2057 44189 2060
rect 44223 2057 44235 2091
rect 44177 2051 44235 2057
rect 44542 2048 44548 2100
rect 44600 2048 44606 2100
rect 44726 2048 44732 2100
rect 44784 2088 44790 2100
rect 44913 2091 44971 2097
rect 44913 2088 44925 2091
rect 44784 2060 44925 2088
rect 44784 2048 44790 2060
rect 44913 2057 44925 2060
rect 44959 2057 44971 2091
rect 44913 2051 44971 2057
rect 39040 2020 39068 2048
rect 38212 1992 38792 2020
rect 33778 1912 33784 1964
rect 33836 1912 33842 1964
rect 36446 1912 36452 1964
rect 36504 1952 36510 1964
rect 36633 1955 36691 1961
rect 36633 1952 36645 1955
rect 36504 1924 36645 1952
rect 36504 1912 36510 1924
rect 36633 1921 36645 1924
rect 36679 1921 36691 1955
rect 36633 1915 36691 1921
rect 38194 1912 38200 1964
rect 38252 1952 38258 1964
rect 38657 1955 38715 1961
rect 38657 1952 38669 1955
rect 38252 1924 38669 1952
rect 38252 1912 38258 1924
rect 38657 1921 38669 1924
rect 38703 1921 38715 1955
rect 38657 1915 38715 1921
rect 33008 1856 33456 1884
rect 33796 1884 33824 1912
rect 33873 1887 33931 1893
rect 33873 1884 33885 1887
rect 33796 1856 33885 1884
rect 33008 1844 33014 1856
rect 33873 1853 33885 1856
rect 33919 1853 33931 1887
rect 34238 1884 34244 1896
rect 33873 1847 33931 1853
rect 33980 1856 34244 1884
rect 33980 1816 34008 1856
rect 34238 1844 34244 1856
rect 34296 1844 34302 1896
rect 34882 1844 34888 1896
rect 34940 1884 34946 1896
rect 34940 1856 35572 1884
rect 34940 1844 34946 1856
rect 33244 1788 34008 1816
rect 35544 1816 35572 1856
rect 35618 1844 35624 1896
rect 35676 1884 35682 1896
rect 36173 1887 36231 1893
rect 36173 1884 36185 1887
rect 35676 1856 36185 1884
rect 35676 1844 35682 1856
rect 36173 1853 36185 1856
rect 36219 1853 36231 1887
rect 36173 1847 36231 1853
rect 36357 1887 36415 1893
rect 36357 1853 36369 1887
rect 36403 1884 36415 1887
rect 36538 1884 36544 1896
rect 36403 1856 36544 1884
rect 36403 1853 36415 1856
rect 36357 1847 36415 1853
rect 36538 1844 36544 1856
rect 36596 1844 36602 1896
rect 38764 1884 38792 1992
rect 38856 1992 39068 2020
rect 39500 2020 39528 2048
rect 39500 1992 39606 2020
rect 38856 1961 38884 1992
rect 40402 1980 40408 2032
rect 40460 2020 40466 2032
rect 40460 1992 41184 2020
rect 40460 1980 40466 1992
rect 38841 1955 38899 1961
rect 38841 1921 38853 1955
rect 38887 1921 38899 1955
rect 38841 1915 38899 1921
rect 40586 1912 40592 1964
rect 40644 1952 40650 1964
rect 41156 1961 41184 1992
rect 41506 1980 41512 2032
rect 41564 1980 41570 2032
rect 42426 1980 42432 2032
rect 42484 2020 42490 2032
rect 43073 2023 43131 2029
rect 43073 2020 43085 2023
rect 42484 1992 43085 2020
rect 42484 1980 42490 1992
rect 43073 1989 43085 1992
rect 43119 2020 43131 2023
rect 43441 2023 43499 2029
rect 43441 2020 43453 2023
rect 43119 1992 43453 2020
rect 43119 1989 43131 1992
rect 43073 1983 43131 1989
rect 43441 1989 43453 1992
rect 43487 1989 43499 2023
rect 43441 1983 43499 1989
rect 40865 1955 40923 1961
rect 40865 1952 40877 1955
rect 40644 1924 40877 1952
rect 40644 1912 40650 1924
rect 40865 1921 40877 1924
rect 40911 1921 40923 1955
rect 40865 1915 40923 1921
rect 41141 1955 41199 1961
rect 41141 1921 41153 1955
rect 41187 1921 41199 1955
rect 41141 1915 41199 1921
rect 39117 1887 39175 1893
rect 36740 1856 38516 1884
rect 38764 1856 38976 1884
rect 36740 1816 36768 1856
rect 35544 1788 36768 1816
rect 33244 1748 33272 1788
rect 38102 1776 38108 1828
rect 38160 1816 38166 1828
rect 38488 1825 38516 1856
rect 38381 1819 38439 1825
rect 38381 1816 38393 1819
rect 38160 1788 38393 1816
rect 38160 1776 38166 1788
rect 38381 1785 38393 1788
rect 38427 1785 38439 1819
rect 38381 1779 38439 1785
rect 38473 1819 38531 1825
rect 38473 1785 38485 1819
rect 38519 1785 38531 1819
rect 38473 1779 38531 1785
rect 31864 1720 33272 1748
rect 31665 1711 31723 1717
rect 33318 1708 33324 1760
rect 33376 1748 33382 1760
rect 33689 1751 33747 1757
rect 33689 1748 33701 1751
rect 33376 1720 33701 1748
rect 33376 1708 33382 1720
rect 33689 1717 33701 1720
rect 33735 1717 33747 1751
rect 33689 1711 33747 1717
rect 36896 1751 36954 1757
rect 36896 1717 36908 1751
rect 36942 1748 36954 1751
rect 38838 1748 38844 1760
rect 36942 1720 38844 1748
rect 36942 1717 36954 1720
rect 36896 1711 36954 1717
rect 38838 1708 38844 1720
rect 38896 1708 38902 1760
rect 38948 1748 38976 1856
rect 39117 1853 39129 1887
rect 39163 1884 39175 1887
rect 39163 1856 41000 1884
rect 39163 1853 39175 1856
rect 39117 1847 39175 1853
rect 40972 1825 41000 1856
rect 40957 1819 41015 1825
rect 40957 1785 40969 1819
rect 41003 1785 41015 1819
rect 40957 1779 41015 1785
rect 40218 1748 40224 1760
rect 38948 1720 40224 1748
rect 40218 1708 40224 1720
rect 40276 1708 40282 1760
rect 460 1658 45540 1680
rect 460 1606 3570 1658
rect 3622 1606 3634 1658
rect 3686 1606 3698 1658
rect 3750 1606 3762 1658
rect 3814 1606 3826 1658
rect 3878 1606 8570 1658
rect 8622 1606 8634 1658
rect 8686 1606 8698 1658
rect 8750 1606 8762 1658
rect 8814 1606 8826 1658
rect 8878 1606 13570 1658
rect 13622 1606 13634 1658
rect 13686 1606 13698 1658
rect 13750 1606 13762 1658
rect 13814 1606 13826 1658
rect 13878 1606 18570 1658
rect 18622 1606 18634 1658
rect 18686 1606 18698 1658
rect 18750 1606 18762 1658
rect 18814 1606 18826 1658
rect 18878 1606 23570 1658
rect 23622 1606 23634 1658
rect 23686 1606 23698 1658
rect 23750 1606 23762 1658
rect 23814 1606 23826 1658
rect 23878 1606 28570 1658
rect 28622 1606 28634 1658
rect 28686 1606 28698 1658
rect 28750 1606 28762 1658
rect 28814 1606 28826 1658
rect 28878 1606 33570 1658
rect 33622 1606 33634 1658
rect 33686 1606 33698 1658
rect 33750 1606 33762 1658
rect 33814 1606 33826 1658
rect 33878 1606 38570 1658
rect 38622 1606 38634 1658
rect 38686 1606 38698 1658
rect 38750 1606 38762 1658
rect 38814 1606 38826 1658
rect 38878 1606 43570 1658
rect 43622 1606 43634 1658
rect 43686 1606 43698 1658
rect 43750 1606 43762 1658
rect 43814 1606 43826 1658
rect 43878 1606 45540 1658
rect 460 1584 45540 1606
rect 2866 1504 2872 1556
rect 2924 1544 2930 1556
rect 3329 1547 3387 1553
rect 3329 1544 3341 1547
rect 2924 1516 3341 1544
rect 2924 1504 2930 1516
rect 3329 1513 3341 1516
rect 3375 1513 3387 1547
rect 3329 1507 3387 1513
rect 5169 1547 5227 1553
rect 5169 1513 5181 1547
rect 5215 1544 5227 1547
rect 5994 1544 6000 1556
rect 5215 1516 6000 1544
rect 5215 1513 5227 1516
rect 5169 1507 5227 1513
rect 5994 1504 6000 1516
rect 6052 1504 6058 1556
rect 6914 1504 6920 1556
rect 6972 1504 6978 1556
rect 7653 1547 7711 1553
rect 7653 1513 7665 1547
rect 7699 1544 7711 1547
rect 8110 1544 8116 1556
rect 7699 1516 8116 1544
rect 7699 1513 7711 1516
rect 7653 1507 7711 1513
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 9214 1504 9220 1556
rect 9272 1504 9278 1556
rect 10042 1504 10048 1556
rect 10100 1504 10106 1556
rect 11054 1504 11060 1556
rect 11112 1504 11118 1556
rect 15194 1504 15200 1556
rect 15252 1504 15258 1556
rect 16666 1504 16672 1556
rect 16724 1504 16730 1556
rect 17678 1504 17684 1556
rect 17736 1544 17742 1556
rect 17957 1547 18015 1553
rect 17957 1544 17969 1547
rect 17736 1516 17969 1544
rect 17736 1504 17742 1516
rect 17957 1513 17969 1516
rect 18003 1513 18015 1547
rect 17957 1507 18015 1513
rect 19334 1504 19340 1556
rect 19392 1504 19398 1556
rect 24210 1504 24216 1556
rect 24268 1504 24274 1556
rect 25590 1504 25596 1556
rect 25648 1544 25654 1556
rect 25961 1547 26019 1553
rect 25961 1544 25973 1547
rect 25648 1516 25973 1544
rect 25648 1504 25654 1516
rect 25961 1513 25973 1516
rect 26007 1513 26019 1547
rect 25961 1507 26019 1513
rect 26513 1547 26571 1553
rect 26513 1513 26525 1547
rect 26559 1513 26571 1547
rect 26513 1507 26571 1513
rect 27065 1547 27123 1553
rect 27065 1513 27077 1547
rect 27111 1513 27123 1547
rect 27065 1507 27123 1513
rect 1029 1479 1087 1485
rect 1029 1445 1041 1479
rect 1075 1476 1087 1479
rect 1210 1476 1216 1488
rect 1075 1448 1216 1476
rect 1075 1445 1087 1448
rect 1029 1439 1087 1445
rect 1210 1436 1216 1448
rect 1268 1476 1274 1488
rect 1857 1479 1915 1485
rect 1857 1476 1869 1479
rect 1268 1448 1869 1476
rect 1268 1436 1274 1448
rect 1857 1445 1869 1448
rect 1903 1476 1915 1479
rect 2961 1479 3019 1485
rect 2961 1476 2973 1479
rect 1903 1448 2973 1476
rect 1903 1445 1915 1448
rect 1857 1439 1915 1445
rect 2961 1445 2973 1448
rect 3007 1476 3019 1479
rect 3142 1476 3148 1488
rect 3007 1448 3148 1476
rect 3007 1445 3019 1448
rect 2961 1439 3019 1445
rect 3142 1436 3148 1448
rect 3200 1436 3206 1488
rect 10060 1476 10088 1504
rect 11701 1479 11759 1485
rect 11701 1476 11713 1479
rect 10060 1448 11713 1476
rect 11701 1445 11713 1448
rect 11747 1476 11759 1479
rect 12342 1476 12348 1488
rect 11747 1448 12348 1476
rect 11747 1445 11759 1448
rect 11701 1439 11759 1445
rect 12342 1436 12348 1448
rect 12400 1476 12406 1488
rect 12529 1479 12587 1485
rect 12529 1476 12541 1479
rect 12400 1448 12541 1476
rect 12400 1436 12406 1448
rect 12529 1445 12541 1448
rect 12575 1445 12587 1479
rect 12529 1439 12587 1445
rect 15838 1436 15844 1488
rect 15896 1476 15902 1488
rect 17696 1476 17724 1504
rect 15896 1448 17724 1476
rect 22066 1448 22784 1476
rect 15896 1436 15902 1448
rect 22066 1408 22094 1448
rect 21652 1380 22094 1408
rect 22204 1380 22692 1408
rect 1121 1343 1179 1349
rect 1121 1309 1133 1343
rect 1167 1340 1179 1343
rect 1302 1340 1308 1352
rect 1167 1312 1308 1340
rect 1167 1309 1179 1312
rect 1121 1303 1179 1309
rect 1302 1300 1308 1312
rect 1360 1300 1366 1352
rect 1949 1343 2007 1349
rect 1949 1309 1961 1343
rect 1995 1340 2007 1343
rect 2130 1340 2136 1352
rect 1995 1312 2136 1340
rect 1995 1309 2007 1312
rect 1949 1303 2007 1309
rect 2130 1300 2136 1312
rect 2188 1300 2194 1352
rect 2958 1300 2964 1352
rect 3016 1340 3022 1352
rect 3237 1343 3295 1349
rect 3237 1340 3249 1343
rect 3016 1312 3249 1340
rect 3016 1300 3022 1312
rect 3237 1309 3249 1312
rect 3283 1309 3295 1343
rect 3237 1303 3295 1309
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1340 3755 1343
rect 3970 1340 3976 1352
rect 3743 1312 3976 1340
rect 3743 1309 3755 1312
rect 3697 1303 3755 1309
rect 3970 1300 3976 1312
rect 4028 1300 4034 1352
rect 4433 1343 4491 1349
rect 4433 1309 4445 1343
rect 4479 1340 4491 1343
rect 4522 1340 4528 1352
rect 4479 1312 4528 1340
rect 4479 1309 4491 1312
rect 4433 1303 4491 1309
rect 4522 1300 4528 1312
rect 4580 1300 4586 1352
rect 5166 1300 5172 1352
rect 5224 1340 5230 1352
rect 5261 1343 5319 1349
rect 5261 1340 5273 1343
rect 5224 1312 5273 1340
rect 5224 1300 5230 1312
rect 5261 1309 5273 1312
rect 5307 1309 5319 1343
rect 5261 1303 5319 1309
rect 6089 1343 6147 1349
rect 6089 1309 6101 1343
rect 6135 1340 6147 1343
rect 6178 1340 6184 1352
rect 6135 1312 6184 1340
rect 6135 1309 6147 1312
rect 6089 1303 6147 1309
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1340 6883 1343
rect 7006 1340 7012 1352
rect 6871 1312 7012 1340
rect 6871 1309 6883 1312
rect 6825 1303 6883 1309
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7742 1300 7748 1352
rect 7800 1300 7806 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8938 1340 8944 1352
rect 8619 1312 8944 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8938 1300 8944 1312
rect 8996 1300 9002 1352
rect 9401 1343 9459 1349
rect 9401 1309 9413 1343
rect 9447 1340 9459 1343
rect 9674 1340 9680 1352
rect 9447 1312 9680 1340
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 9674 1300 9680 1312
rect 9732 1300 9738 1352
rect 10229 1343 10287 1349
rect 10229 1309 10241 1343
rect 10275 1340 10287 1343
rect 10318 1340 10324 1352
rect 10275 1312 10324 1340
rect 10275 1309 10287 1312
rect 10229 1303 10287 1309
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1340 11023 1343
rect 11146 1340 11152 1352
rect 11011 1312 11152 1340
rect 11011 1309 11023 1312
rect 10965 1303 11023 1309
rect 11146 1300 11152 1312
rect 11204 1300 11210 1352
rect 11885 1343 11943 1349
rect 11885 1309 11897 1343
rect 11931 1340 11943 1343
rect 11974 1340 11980 1352
rect 11931 1312 11980 1340
rect 11931 1309 11943 1312
rect 11885 1303 11943 1309
rect 11974 1300 11980 1312
rect 12032 1300 12038 1352
rect 12250 1300 12256 1352
rect 12308 1340 12314 1352
rect 12713 1343 12771 1349
rect 12713 1340 12725 1343
rect 12308 1312 12725 1340
rect 12308 1300 12314 1312
rect 12713 1309 12725 1312
rect 12759 1309 12771 1343
rect 12713 1303 12771 1309
rect 13446 1300 13452 1352
rect 13504 1340 13510 1352
rect 13541 1343 13599 1349
rect 13541 1340 13553 1343
rect 13504 1312 13553 1340
rect 13504 1300 13510 1312
rect 13541 1309 13553 1312
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 14366 1300 14372 1352
rect 14424 1300 14430 1352
rect 15105 1343 15163 1349
rect 15105 1309 15117 1343
rect 15151 1340 15163 1343
rect 15378 1340 15384 1352
rect 15151 1312 15384 1340
rect 15151 1309 15163 1312
rect 15105 1303 15163 1309
rect 15378 1300 15384 1312
rect 15436 1300 15442 1352
rect 16025 1343 16083 1349
rect 16025 1309 16037 1343
rect 16071 1340 16083 1343
rect 16206 1340 16212 1352
rect 16071 1312 16212 1340
rect 16071 1309 16083 1312
rect 16025 1303 16083 1309
rect 16206 1300 16212 1312
rect 16264 1300 16270 1352
rect 16853 1343 16911 1349
rect 16853 1309 16865 1343
rect 16899 1340 16911 1343
rect 18322 1340 18328 1352
rect 16899 1312 18328 1340
rect 16899 1309 16911 1312
rect 16853 1303 16911 1309
rect 18322 1300 18328 1312
rect 18380 1300 18386 1352
rect 18414 1300 18420 1352
rect 18472 1340 18478 1352
rect 18601 1343 18659 1349
rect 18601 1340 18613 1343
rect 18472 1312 18613 1340
rect 18472 1300 18478 1312
rect 18601 1309 18613 1312
rect 18647 1309 18659 1343
rect 18601 1303 18659 1309
rect 19245 1343 19303 1349
rect 19245 1309 19257 1343
rect 19291 1340 19303 1343
rect 19702 1340 19708 1352
rect 19291 1312 19708 1340
rect 19291 1309 19303 1312
rect 19245 1303 19303 1309
rect 19702 1300 19708 1312
rect 19760 1300 19766 1352
rect 20162 1300 20168 1352
rect 20220 1300 20226 1352
rect 20806 1300 20812 1352
rect 20864 1340 20870 1352
rect 21177 1343 21235 1349
rect 21177 1340 21189 1343
rect 20864 1312 21189 1340
rect 20864 1300 20870 1312
rect 21177 1309 21189 1312
rect 21223 1309 21235 1343
rect 21652 1340 21680 1380
rect 22204 1352 22232 1380
rect 21177 1303 21235 1309
rect 21468 1312 21680 1340
rect 2222 1232 2228 1284
rect 2280 1272 2286 1284
rect 2593 1275 2651 1281
rect 2593 1272 2605 1275
rect 2280 1244 2605 1272
rect 2280 1232 2286 1244
rect 2593 1241 2605 1244
rect 2639 1272 2651 1275
rect 4249 1275 4307 1281
rect 4249 1272 4261 1275
rect 2639 1244 4261 1272
rect 2639 1241 2651 1244
rect 2593 1235 2651 1241
rect 4249 1241 4261 1244
rect 4295 1272 4307 1275
rect 5718 1272 5724 1284
rect 4295 1244 5724 1272
rect 4295 1241 4307 1244
rect 4249 1235 4307 1241
rect 5718 1232 5724 1244
rect 5776 1232 5782 1284
rect 10137 1275 10195 1281
rect 10137 1241 10149 1275
rect 10183 1272 10195 1275
rect 14090 1272 14096 1284
rect 10183 1244 14096 1272
rect 10183 1241 10195 1244
rect 10137 1235 10195 1241
rect 14090 1232 14096 1244
rect 14148 1232 14154 1284
rect 19518 1272 19524 1284
rect 18340 1244 19524 1272
rect 1302 1164 1308 1216
rect 1360 1164 1366 1216
rect 1854 1164 1860 1216
rect 1912 1204 1918 1216
rect 2133 1207 2191 1213
rect 2133 1204 2145 1207
rect 1912 1176 2145 1204
rect 1912 1164 1918 1176
rect 2133 1173 2145 1176
rect 2179 1173 2191 1207
rect 2133 1167 2191 1173
rect 3510 1164 3516 1216
rect 3568 1204 3574 1216
rect 3881 1207 3939 1213
rect 3881 1204 3893 1207
rect 3568 1176 3893 1204
rect 3568 1164 3574 1176
rect 3881 1173 3893 1176
rect 3927 1173 3939 1207
rect 3881 1167 3939 1173
rect 4614 1164 4620 1216
rect 4672 1164 4678 1216
rect 5442 1164 5448 1216
rect 5500 1164 5506 1216
rect 5994 1164 6000 1216
rect 6052 1204 6058 1216
rect 6273 1207 6331 1213
rect 6273 1204 6285 1207
rect 6052 1176 6285 1204
rect 6052 1164 6058 1176
rect 6273 1173 6285 1176
rect 6319 1173 6331 1207
rect 6273 1167 6331 1173
rect 7926 1164 7932 1216
rect 7984 1164 7990 1216
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9582 1164 9588 1216
rect 9640 1164 9646 1216
rect 10410 1164 10416 1216
rect 10468 1164 10474 1216
rect 12066 1164 12072 1216
rect 12124 1164 12130 1216
rect 12894 1164 12900 1216
rect 12952 1164 12958 1216
rect 13722 1164 13728 1216
rect 13780 1164 13786 1216
rect 14182 1164 14188 1216
rect 14240 1164 14246 1216
rect 14274 1164 14280 1216
rect 14332 1204 14338 1216
rect 14553 1207 14611 1213
rect 14553 1204 14565 1207
rect 14332 1176 14565 1204
rect 14332 1164 14338 1176
rect 14553 1173 14565 1176
rect 14599 1173 14611 1207
rect 14553 1167 14611 1173
rect 15930 1164 15936 1216
rect 15988 1204 15994 1216
rect 16209 1207 16267 1213
rect 16209 1204 16221 1207
rect 15988 1176 16221 1204
rect 15988 1164 15994 1176
rect 16209 1173 16221 1176
rect 16255 1173 16267 1207
rect 16209 1167 16267 1173
rect 17034 1164 17040 1216
rect 17092 1164 17098 1216
rect 18340 1213 18368 1244
rect 19518 1232 19524 1244
rect 19576 1232 19582 1284
rect 20901 1275 20959 1281
rect 20901 1241 20913 1275
rect 20947 1272 20959 1275
rect 21468 1272 21496 1312
rect 21726 1300 21732 1352
rect 21784 1300 21790 1352
rect 21821 1343 21879 1349
rect 21821 1309 21833 1343
rect 21867 1309 21879 1343
rect 21821 1303 21879 1309
rect 21836 1272 21864 1303
rect 22186 1300 22192 1352
rect 22244 1300 22250 1352
rect 22554 1300 22560 1352
rect 22612 1300 22618 1352
rect 22664 1349 22692 1380
rect 22649 1343 22707 1349
rect 22649 1309 22661 1343
rect 22695 1309 22707 1343
rect 22756 1340 22784 1448
rect 24228 1408 24256 1504
rect 25498 1436 25504 1488
rect 25556 1476 25562 1488
rect 26528 1476 26556 1507
rect 25556 1448 26556 1476
rect 25556 1436 25562 1448
rect 23952 1380 24256 1408
rect 24489 1411 24547 1417
rect 23014 1340 23020 1352
rect 22756 1312 23020 1340
rect 22649 1303 22707 1309
rect 23014 1300 23020 1312
rect 23072 1300 23078 1352
rect 23952 1349 23980 1380
rect 24489 1377 24501 1411
rect 24535 1408 24547 1411
rect 25130 1408 25136 1420
rect 24535 1380 25136 1408
rect 24535 1377 24547 1380
rect 24489 1371 24547 1377
rect 25130 1368 25136 1380
rect 25188 1368 25194 1420
rect 26142 1368 26148 1420
rect 26200 1408 26206 1420
rect 27080 1408 27108 1507
rect 27614 1504 27620 1556
rect 27672 1544 27678 1556
rect 27801 1547 27859 1553
rect 27801 1544 27813 1547
rect 27672 1516 27813 1544
rect 27672 1504 27678 1516
rect 27801 1513 27813 1516
rect 27847 1513 27859 1547
rect 27801 1507 27859 1513
rect 28629 1547 28687 1553
rect 28629 1513 28641 1547
rect 28675 1544 28687 1547
rect 29086 1544 29092 1556
rect 28675 1516 29092 1544
rect 28675 1513 28687 1516
rect 28629 1507 28687 1513
rect 29086 1504 29092 1516
rect 29144 1504 29150 1556
rect 29181 1547 29239 1553
rect 29181 1513 29193 1547
rect 29227 1544 29239 1547
rect 29270 1544 29276 1556
rect 29227 1516 29276 1544
rect 29227 1513 29239 1516
rect 29181 1507 29239 1513
rect 29270 1504 29276 1516
rect 29328 1504 29334 1556
rect 29638 1504 29644 1556
rect 29696 1504 29702 1556
rect 29914 1504 29920 1556
rect 29972 1504 29978 1556
rect 30006 1504 30012 1556
rect 30064 1544 30070 1556
rect 30377 1547 30435 1553
rect 30377 1544 30389 1547
rect 30064 1516 30389 1544
rect 30064 1504 30070 1516
rect 30377 1513 30389 1516
rect 30423 1513 30435 1547
rect 30377 1507 30435 1513
rect 31036 1516 31524 1544
rect 28258 1436 28264 1488
rect 28316 1476 28322 1488
rect 29656 1476 29684 1504
rect 31036 1476 31064 1516
rect 28316 1448 28948 1476
rect 29656 1448 31064 1476
rect 31113 1479 31171 1485
rect 28316 1436 28322 1448
rect 26200 1380 27108 1408
rect 26200 1368 26206 1380
rect 28350 1368 28356 1420
rect 28408 1408 28414 1420
rect 28920 1408 28948 1448
rect 31113 1445 31125 1479
rect 31159 1445 31171 1479
rect 31113 1439 31171 1445
rect 29270 1408 29276 1420
rect 28408 1380 28764 1408
rect 28408 1368 28414 1380
rect 23937 1343 23995 1349
rect 23124 1312 23888 1340
rect 23124 1272 23152 1312
rect 20947 1244 21496 1272
rect 21560 1244 21864 1272
rect 22388 1244 23152 1272
rect 23201 1275 23259 1281
rect 20947 1241 20959 1244
rect 20901 1235 20959 1241
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1173 18383 1207
rect 18325 1167 18383 1173
rect 18414 1164 18420 1216
rect 18472 1204 18478 1216
rect 18785 1207 18843 1213
rect 18785 1204 18797 1207
rect 18472 1176 18797 1204
rect 18472 1164 18478 1176
rect 18785 1173 18797 1176
rect 18831 1173 18843 1207
rect 18785 1167 18843 1173
rect 20070 1164 20076 1216
rect 20128 1164 20134 1216
rect 20346 1164 20352 1216
rect 20404 1164 20410 1216
rect 20990 1164 20996 1216
rect 21048 1204 21054 1216
rect 21560 1213 21588 1244
rect 21361 1207 21419 1213
rect 21361 1204 21373 1207
rect 21048 1176 21373 1204
rect 21048 1164 21054 1176
rect 21361 1173 21373 1176
rect 21407 1173 21419 1207
rect 21361 1167 21419 1173
rect 21545 1207 21603 1213
rect 21545 1173 21557 1207
rect 21591 1173 21603 1207
rect 21545 1167 21603 1173
rect 21726 1164 21732 1216
rect 21784 1204 21790 1216
rect 22388 1213 22416 1244
rect 23201 1241 23213 1275
rect 23247 1272 23259 1275
rect 23860 1272 23888 1312
rect 23937 1309 23949 1343
rect 23983 1309 23995 1343
rect 23937 1303 23995 1309
rect 24118 1300 24124 1352
rect 24176 1340 24182 1352
rect 24213 1343 24271 1349
rect 24213 1340 24225 1343
rect 24176 1312 24225 1340
rect 24176 1300 24182 1312
rect 24213 1309 24225 1312
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 26234 1300 26240 1352
rect 26292 1340 26298 1352
rect 26421 1343 26479 1349
rect 26421 1340 26433 1343
rect 26292 1312 26433 1340
rect 26292 1300 26298 1312
rect 26421 1309 26433 1312
rect 26467 1309 26479 1343
rect 26421 1303 26479 1309
rect 26973 1343 27031 1349
rect 26973 1309 26985 1343
rect 27019 1340 27031 1343
rect 27154 1340 27160 1352
rect 27019 1312 27160 1340
rect 27019 1309 27031 1312
rect 26973 1303 27031 1309
rect 27154 1300 27160 1312
rect 27212 1300 27218 1352
rect 27709 1343 27767 1349
rect 27709 1309 27721 1343
rect 27755 1340 27767 1343
rect 28074 1340 28080 1352
rect 27755 1312 28080 1340
rect 27755 1309 27767 1312
rect 27709 1303 27767 1309
rect 28074 1300 28080 1312
rect 28132 1300 28138 1352
rect 28169 1343 28227 1349
rect 28169 1309 28181 1343
rect 28215 1309 28227 1343
rect 28169 1303 28227 1309
rect 24486 1272 24492 1284
rect 23247 1244 23796 1272
rect 23860 1244 24492 1272
rect 23247 1241 23259 1244
rect 23201 1235 23259 1241
rect 22005 1207 22063 1213
rect 22005 1204 22017 1207
rect 21784 1176 22017 1204
rect 21784 1164 21790 1176
rect 22005 1173 22017 1176
rect 22051 1173 22063 1207
rect 22005 1167 22063 1173
rect 22373 1207 22431 1213
rect 22373 1173 22385 1207
rect 22419 1173 22431 1207
rect 22373 1167 22431 1173
rect 22554 1164 22560 1216
rect 22612 1204 22618 1216
rect 22833 1207 22891 1213
rect 22833 1204 22845 1207
rect 22612 1176 22845 1204
rect 22612 1164 22618 1176
rect 22833 1173 22845 1176
rect 22879 1173 22891 1207
rect 22833 1167 22891 1173
rect 23290 1164 23296 1216
rect 23348 1164 23354 1216
rect 23768 1213 23796 1244
rect 24486 1232 24492 1244
rect 24544 1232 24550 1284
rect 24762 1232 24768 1284
rect 24820 1272 24826 1284
rect 28184 1272 28212 1303
rect 28442 1300 28448 1352
rect 28500 1340 28506 1352
rect 28736 1349 28764 1380
rect 28920 1380 29276 1408
rect 28920 1349 28948 1380
rect 29270 1368 29276 1380
rect 29328 1368 29334 1420
rect 31128 1408 31156 1439
rect 29380 1380 29592 1408
rect 28537 1343 28595 1349
rect 28537 1340 28549 1343
rect 28500 1312 28549 1340
rect 28500 1300 28506 1312
rect 28537 1309 28549 1312
rect 28583 1309 28595 1343
rect 28537 1303 28595 1309
rect 28721 1343 28779 1349
rect 28721 1309 28733 1343
rect 28767 1309 28779 1343
rect 28721 1303 28779 1309
rect 28905 1343 28963 1349
rect 28905 1309 28917 1343
rect 28951 1309 28963 1343
rect 29380 1340 29408 1380
rect 28905 1303 28963 1309
rect 29012 1312 29408 1340
rect 29457 1343 29515 1349
rect 24820 1244 24978 1272
rect 28184 1244 28764 1272
rect 24820 1232 24826 1244
rect 23753 1207 23811 1213
rect 23753 1173 23765 1207
rect 23799 1173 23811 1207
rect 23753 1167 23811 1173
rect 27062 1164 27068 1216
rect 27120 1204 27126 1216
rect 28353 1207 28411 1213
rect 28353 1204 28365 1207
rect 27120 1176 28365 1204
rect 27120 1164 27126 1176
rect 28353 1173 28365 1176
rect 28399 1173 28411 1207
rect 28736 1204 28764 1244
rect 29012 1204 29040 1312
rect 29457 1309 29469 1343
rect 29503 1309 29515 1343
rect 29564 1340 29592 1380
rect 30668 1380 31156 1408
rect 31496 1408 31524 1516
rect 31662 1504 31668 1556
rect 31720 1544 31726 1556
rect 31720 1516 32168 1544
rect 31720 1504 31726 1516
rect 32030 1436 32036 1488
rect 32088 1436 32094 1488
rect 32140 1476 32168 1516
rect 32214 1504 32220 1556
rect 32272 1544 32278 1556
rect 32677 1547 32735 1553
rect 32677 1544 32689 1547
rect 32272 1516 32689 1544
rect 32272 1504 32278 1516
rect 32677 1513 32689 1516
rect 32723 1513 32735 1547
rect 32677 1507 32735 1513
rect 34974 1504 34980 1556
rect 35032 1544 35038 1556
rect 38194 1544 38200 1556
rect 35032 1516 38200 1544
rect 35032 1504 35038 1516
rect 38194 1504 38200 1516
rect 38252 1504 38258 1556
rect 38930 1504 38936 1556
rect 38988 1544 38994 1556
rect 40037 1547 40095 1553
rect 40037 1544 40049 1547
rect 38988 1516 40049 1544
rect 38988 1504 38994 1516
rect 40037 1513 40049 1516
rect 40083 1513 40095 1547
rect 40037 1507 40095 1513
rect 40218 1504 40224 1556
rect 40276 1544 40282 1556
rect 40589 1547 40647 1553
rect 40589 1544 40601 1547
rect 40276 1516 40601 1544
rect 40276 1504 40282 1516
rect 40589 1513 40601 1516
rect 40635 1513 40647 1547
rect 40589 1507 40647 1513
rect 40954 1504 40960 1556
rect 41012 1544 41018 1556
rect 41141 1547 41199 1553
rect 41141 1544 41153 1547
rect 41012 1516 41153 1544
rect 41012 1504 41018 1516
rect 41141 1513 41153 1516
rect 41187 1513 41199 1547
rect 41141 1507 41199 1513
rect 42978 1504 42984 1556
rect 43036 1504 43042 1556
rect 43898 1504 43904 1556
rect 43956 1504 43962 1556
rect 33137 1479 33195 1485
rect 33137 1476 33149 1479
rect 32140 1448 33149 1476
rect 33137 1445 33149 1448
rect 33183 1445 33195 1479
rect 33137 1439 33195 1445
rect 33318 1436 33324 1488
rect 33376 1436 33382 1488
rect 35250 1436 35256 1488
rect 35308 1476 35314 1488
rect 36173 1479 36231 1485
rect 35308 1448 35388 1476
rect 35308 1436 35314 1448
rect 31573 1411 31631 1417
rect 31573 1408 31585 1411
rect 31496 1380 31585 1408
rect 30668 1340 30696 1380
rect 31573 1377 31585 1380
rect 31619 1408 31631 1411
rect 32306 1408 32312 1420
rect 31619 1380 32312 1408
rect 31619 1377 31631 1380
rect 31573 1371 31631 1377
rect 32306 1368 32312 1380
rect 32364 1368 32370 1420
rect 33336 1408 33364 1436
rect 33413 1411 33471 1417
rect 33413 1408 33425 1411
rect 32416 1380 32996 1408
rect 29564 1312 30696 1340
rect 30745 1343 30803 1349
rect 29457 1303 29515 1309
rect 30745 1309 30757 1343
rect 30791 1309 30803 1343
rect 30745 1303 30803 1309
rect 31297 1343 31355 1349
rect 31297 1309 31309 1343
rect 31343 1340 31355 1343
rect 31386 1340 31392 1352
rect 31343 1312 31392 1340
rect 31343 1309 31355 1312
rect 31297 1303 31355 1309
rect 29270 1232 29276 1284
rect 29328 1272 29334 1284
rect 29472 1272 29500 1303
rect 29730 1272 29736 1284
rect 29328 1244 29736 1272
rect 29328 1232 29334 1244
rect 29730 1232 29736 1244
rect 29788 1232 29794 1284
rect 30282 1232 30288 1284
rect 30340 1232 30346 1284
rect 30760 1272 30788 1303
rect 31386 1300 31392 1312
rect 31444 1300 31450 1352
rect 31478 1300 31484 1352
rect 31536 1340 31542 1352
rect 31665 1343 31723 1349
rect 31665 1340 31677 1343
rect 31536 1312 31677 1340
rect 31536 1300 31542 1312
rect 31665 1309 31677 1312
rect 31711 1309 31723 1343
rect 31665 1303 31723 1309
rect 32030 1300 32036 1352
rect 32088 1340 32094 1352
rect 32125 1343 32183 1349
rect 32125 1340 32137 1343
rect 32088 1312 32137 1340
rect 32088 1300 32094 1312
rect 32125 1309 32137 1312
rect 32171 1309 32183 1343
rect 32416 1340 32444 1380
rect 32125 1303 32183 1309
rect 32232 1312 32444 1340
rect 32232 1272 32260 1312
rect 32490 1300 32496 1352
rect 32548 1300 32554 1352
rect 30760 1244 32260 1272
rect 32309 1275 32367 1281
rect 32309 1241 32321 1275
rect 32355 1241 32367 1275
rect 32309 1235 32367 1241
rect 28736 1176 29040 1204
rect 28353 1167 28411 1173
rect 29086 1164 29092 1216
rect 29144 1204 29150 1216
rect 29365 1207 29423 1213
rect 29365 1204 29377 1207
rect 29144 1176 29377 1204
rect 29144 1164 29150 1176
rect 29365 1173 29377 1176
rect 29411 1173 29423 1207
rect 29365 1167 29423 1173
rect 30374 1164 30380 1216
rect 30432 1204 30438 1216
rect 30929 1207 30987 1213
rect 30929 1204 30941 1207
rect 30432 1176 30941 1204
rect 30432 1164 30438 1176
rect 30929 1173 30941 1176
rect 30975 1173 30987 1207
rect 30929 1167 30987 1173
rect 32122 1164 32128 1216
rect 32180 1204 32186 1216
rect 32324 1204 32352 1235
rect 32398 1232 32404 1284
rect 32456 1232 32462 1284
rect 32858 1281 32864 1284
rect 32843 1275 32864 1281
rect 32843 1241 32855 1275
rect 32843 1235 32864 1241
rect 32858 1232 32864 1235
rect 32916 1232 32922 1284
rect 32968 1272 32996 1380
rect 33060 1380 33425 1408
rect 33060 1352 33088 1380
rect 33413 1377 33425 1380
rect 33459 1377 33471 1411
rect 33413 1371 33471 1377
rect 33597 1411 33655 1417
rect 33597 1377 33609 1411
rect 33643 1408 33655 1411
rect 33962 1408 33968 1420
rect 33643 1380 33968 1408
rect 33643 1377 33655 1380
rect 33597 1371 33655 1377
rect 33962 1368 33968 1380
rect 34020 1368 34026 1420
rect 35360 1417 35388 1448
rect 36173 1445 36185 1479
rect 36219 1445 36231 1479
rect 36173 1439 36231 1445
rect 35345 1411 35403 1417
rect 35345 1377 35357 1411
rect 35391 1377 35403 1411
rect 35345 1371 35403 1377
rect 35618 1368 35624 1420
rect 35676 1368 35682 1420
rect 35728 1380 36032 1408
rect 33042 1300 33048 1352
rect 33100 1300 33106 1352
rect 33226 1300 33232 1352
rect 33284 1340 33290 1352
rect 33321 1343 33379 1349
rect 33321 1340 33333 1343
rect 33284 1312 33333 1340
rect 33284 1300 33290 1312
rect 33321 1309 33333 1312
rect 33367 1309 33379 1343
rect 33321 1303 33379 1309
rect 33870 1300 33876 1352
rect 33928 1300 33934 1352
rect 34238 1300 34244 1352
rect 34296 1300 34302 1352
rect 34517 1343 34575 1349
rect 34517 1309 34529 1343
rect 34563 1309 34575 1343
rect 34517 1303 34575 1309
rect 34532 1272 34560 1303
rect 34698 1300 34704 1352
rect 34756 1300 34762 1352
rect 35158 1300 35164 1352
rect 35216 1300 35222 1352
rect 35253 1343 35311 1349
rect 35253 1309 35265 1343
rect 35299 1340 35311 1343
rect 35636 1340 35664 1368
rect 35728 1352 35756 1380
rect 35299 1312 35664 1340
rect 35299 1309 35311 1312
rect 35253 1303 35311 1309
rect 35710 1300 35716 1352
rect 35768 1300 35774 1352
rect 35805 1343 35863 1349
rect 35805 1309 35817 1343
rect 35851 1340 35863 1343
rect 35851 1312 35940 1340
rect 35851 1309 35863 1312
rect 35805 1303 35863 1309
rect 32968 1244 33732 1272
rect 32180 1176 32352 1204
rect 32416 1204 32444 1232
rect 33042 1204 33048 1216
rect 32416 1176 33048 1204
rect 32180 1164 32186 1176
rect 33042 1164 33048 1176
rect 33100 1164 33106 1216
rect 33410 1164 33416 1216
rect 33468 1204 33474 1216
rect 33704 1213 33732 1244
rect 34072 1244 34560 1272
rect 34072 1213 34100 1244
rect 33597 1207 33655 1213
rect 33597 1204 33609 1207
rect 33468 1176 33609 1204
rect 33468 1164 33474 1176
rect 33597 1173 33609 1176
rect 33643 1173 33655 1207
rect 33597 1167 33655 1173
rect 33689 1207 33747 1213
rect 33689 1173 33701 1207
rect 33735 1173 33747 1207
rect 33689 1167 33747 1173
rect 34057 1207 34115 1213
rect 34057 1173 34069 1207
rect 34103 1173 34115 1207
rect 34057 1167 34115 1173
rect 34330 1164 34336 1216
rect 34388 1164 34394 1216
rect 34716 1204 34744 1300
rect 34793 1207 34851 1213
rect 34793 1204 34805 1207
rect 34716 1176 34805 1204
rect 34793 1173 34805 1176
rect 34839 1173 34851 1207
rect 34793 1167 34851 1173
rect 35618 1164 35624 1216
rect 35676 1164 35682 1216
rect 35912 1213 35940 1312
rect 36004 1272 36032 1380
rect 36188 1352 36216 1439
rect 36446 1436 36452 1488
rect 36504 1476 36510 1488
rect 40313 1479 40371 1485
rect 40313 1476 40325 1479
rect 36504 1448 37320 1476
rect 36504 1436 36510 1448
rect 37292 1417 37320 1448
rect 38948 1448 40325 1476
rect 37277 1411 37335 1417
rect 37277 1377 37289 1411
rect 37323 1377 37335 1411
rect 37277 1371 37335 1377
rect 37553 1411 37611 1417
rect 37553 1377 37565 1411
rect 37599 1408 37611 1411
rect 38948 1408 38976 1448
rect 40313 1445 40325 1448
rect 40359 1445 40371 1479
rect 40313 1439 40371 1445
rect 39853 1411 39911 1417
rect 39853 1408 39865 1411
rect 37599 1380 38976 1408
rect 39776 1380 39865 1408
rect 37599 1377 37611 1380
rect 37553 1371 37611 1377
rect 39776 1352 39804 1380
rect 39853 1377 39865 1380
rect 39899 1377 39911 1411
rect 39853 1371 39911 1377
rect 36078 1300 36084 1352
rect 36136 1300 36142 1352
rect 36170 1300 36176 1352
rect 36228 1300 36234 1352
rect 36354 1300 36360 1352
rect 36412 1300 36418 1352
rect 36814 1300 36820 1352
rect 36872 1300 36878 1352
rect 37090 1300 37096 1352
rect 37148 1300 37154 1352
rect 39482 1340 39488 1352
rect 38686 1312 39488 1340
rect 39482 1300 39488 1312
rect 39540 1300 39546 1352
rect 39574 1300 39580 1352
rect 39632 1300 39638 1352
rect 39666 1300 39672 1352
rect 39724 1300 39730 1352
rect 39758 1300 39764 1352
rect 39816 1300 39822 1352
rect 40221 1343 40279 1349
rect 40221 1340 40233 1343
rect 39868 1312 40233 1340
rect 36004 1244 36952 1272
rect 35897 1207 35955 1213
rect 35897 1173 35909 1207
rect 35943 1173 35955 1207
rect 35897 1167 35955 1173
rect 35986 1164 35992 1216
rect 36044 1204 36050 1216
rect 36924 1213 36952 1244
rect 37826 1232 37832 1284
rect 37884 1232 37890 1284
rect 39868 1272 39896 1312
rect 40221 1309 40233 1312
rect 40267 1309 40279 1343
rect 40221 1303 40279 1309
rect 40310 1300 40316 1352
rect 40368 1340 40374 1352
rect 40497 1343 40555 1349
rect 40497 1340 40509 1343
rect 40368 1312 40509 1340
rect 40368 1300 40374 1312
rect 40497 1309 40509 1312
rect 40543 1309 40555 1343
rect 40497 1303 40555 1309
rect 40770 1300 40776 1352
rect 40828 1300 40834 1352
rect 40862 1300 40868 1352
rect 40920 1340 40926 1352
rect 41049 1343 41107 1349
rect 41049 1340 41061 1343
rect 40920 1312 41061 1340
rect 40920 1300 40926 1312
rect 41049 1309 41061 1312
rect 41095 1309 41107 1343
rect 41049 1303 41107 1309
rect 41322 1300 41328 1352
rect 41380 1300 41386 1352
rect 41601 1343 41659 1349
rect 41601 1309 41613 1343
rect 41647 1309 41659 1343
rect 41601 1303 41659 1309
rect 38948 1244 39896 1272
rect 36633 1207 36691 1213
rect 36633 1204 36645 1207
rect 36044 1176 36645 1204
rect 36044 1164 36050 1176
rect 36633 1173 36645 1176
rect 36679 1173 36691 1207
rect 36633 1167 36691 1173
rect 36909 1207 36967 1213
rect 36909 1173 36921 1207
rect 36955 1173 36967 1207
rect 37844 1204 37872 1232
rect 38948 1204 38976 1244
rect 39942 1232 39948 1284
rect 40000 1272 40006 1284
rect 41616 1272 41644 1303
rect 41966 1300 41972 1352
rect 42024 1300 42030 1352
rect 42245 1343 42303 1349
rect 42245 1309 42257 1343
rect 42291 1309 42303 1343
rect 42245 1303 42303 1309
rect 40000 1244 41644 1272
rect 40000 1232 40006 1244
rect 41690 1232 41696 1284
rect 41748 1272 41754 1284
rect 42260 1272 42288 1303
rect 42702 1300 42708 1352
rect 42760 1300 42766 1352
rect 43254 1300 43260 1352
rect 43312 1300 43318 1352
rect 43530 1300 43536 1352
rect 43588 1300 43594 1352
rect 44358 1300 44364 1352
rect 44416 1300 44422 1352
rect 44542 1300 44548 1352
rect 44600 1300 44606 1352
rect 44818 1300 44824 1352
rect 44876 1300 44882 1352
rect 45002 1300 45008 1352
rect 45060 1300 45066 1352
rect 45186 1300 45192 1352
rect 45244 1300 45250 1352
rect 41748 1244 42288 1272
rect 41748 1232 41754 1244
rect 37844 1176 38976 1204
rect 36909 1167 36967 1173
rect 39022 1164 39028 1216
rect 39080 1164 39086 1216
rect 39209 1207 39267 1213
rect 39209 1173 39221 1207
rect 39255 1204 39267 1207
rect 40402 1204 40408 1216
rect 39255 1176 40408 1204
rect 39255 1173 39267 1176
rect 39209 1167 39267 1173
rect 40402 1164 40408 1176
rect 40460 1164 40466 1216
rect 40678 1164 40684 1216
rect 40736 1204 40742 1216
rect 40865 1207 40923 1213
rect 40865 1204 40877 1207
rect 40736 1176 40877 1204
rect 40736 1164 40742 1176
rect 40865 1173 40877 1176
rect 40911 1173 40923 1207
rect 40865 1167 40923 1173
rect 41414 1164 41420 1216
rect 41472 1164 41478 1216
rect 41782 1164 41788 1216
rect 41840 1164 41846 1216
rect 42058 1164 42064 1216
rect 42116 1164 42122 1216
rect 42518 1164 42524 1216
rect 42576 1164 42582 1216
rect 43272 1204 43300 1300
rect 44376 1213 44404 1300
rect 45020 1213 45048 1300
rect 43349 1207 43407 1213
rect 43349 1204 43361 1207
rect 43272 1176 43361 1204
rect 43349 1173 43361 1176
rect 43395 1173 43407 1207
rect 43349 1167 43407 1173
rect 44361 1207 44419 1213
rect 44361 1173 44373 1207
rect 44407 1173 44419 1207
rect 44361 1167 44419 1173
rect 45005 1207 45063 1213
rect 45005 1173 45017 1207
rect 45051 1173 45063 1207
rect 45005 1167 45063 1173
rect 460 1114 45540 1136
rect 460 1062 6070 1114
rect 6122 1062 6134 1114
rect 6186 1062 6198 1114
rect 6250 1062 6262 1114
rect 6314 1062 6326 1114
rect 6378 1062 11070 1114
rect 11122 1062 11134 1114
rect 11186 1062 11198 1114
rect 11250 1062 11262 1114
rect 11314 1062 11326 1114
rect 11378 1062 16070 1114
rect 16122 1062 16134 1114
rect 16186 1062 16198 1114
rect 16250 1062 16262 1114
rect 16314 1062 16326 1114
rect 16378 1062 21070 1114
rect 21122 1062 21134 1114
rect 21186 1062 21198 1114
rect 21250 1062 21262 1114
rect 21314 1062 21326 1114
rect 21378 1062 26070 1114
rect 26122 1062 26134 1114
rect 26186 1062 26198 1114
rect 26250 1062 26262 1114
rect 26314 1062 26326 1114
rect 26378 1062 31070 1114
rect 31122 1062 31134 1114
rect 31186 1062 31198 1114
rect 31250 1062 31262 1114
rect 31314 1062 31326 1114
rect 31378 1062 36070 1114
rect 36122 1062 36134 1114
rect 36186 1062 36198 1114
rect 36250 1062 36262 1114
rect 36314 1062 36326 1114
rect 36378 1062 41070 1114
rect 41122 1062 41134 1114
rect 41186 1062 41198 1114
rect 41250 1062 41262 1114
rect 41314 1062 41326 1114
rect 41378 1062 45540 1114
rect 460 1040 45540 1062
rect 14090 960 14096 1012
rect 14148 960 14154 1012
rect 14182 960 14188 1012
rect 14240 960 14246 1012
rect 20070 960 20076 1012
rect 20128 1000 20134 1012
rect 24578 1000 24584 1012
rect 20128 972 24584 1000
rect 20128 960 20134 972
rect 24578 960 24584 972
rect 24636 960 24642 1012
rect 30282 960 30288 1012
rect 30340 960 30346 1012
rect 32858 960 32864 1012
rect 32916 1000 32922 1012
rect 35618 1000 35624 1012
rect 32916 972 35624 1000
rect 32916 960 32922 972
rect 35618 960 35624 972
rect 35676 960 35682 1012
rect 38286 960 38292 1012
rect 38344 1000 38350 1012
rect 40862 1000 40868 1012
rect 38344 972 40868 1000
rect 38344 960 38350 972
rect 40862 960 40868 972
rect 40920 960 40926 1012
rect 14108 864 14136 960
rect 14200 932 14228 960
rect 25222 932 25228 944
rect 14200 904 25228 932
rect 25222 892 25228 904
rect 25280 892 25286 944
rect 30300 932 30328 960
rect 34330 932 34336 944
rect 30300 904 34336 932
rect 34330 892 34336 904
rect 34388 892 34394 944
rect 39022 892 39028 944
rect 39080 932 39086 944
rect 40126 932 40132 944
rect 39080 904 40132 932
rect 39080 892 39086 904
rect 40126 892 40132 904
rect 40184 892 40190 944
rect 21542 864 21548 876
rect 14108 836 21548 864
rect 21542 824 21548 836
rect 21600 824 21606 876
rect 27246 824 27252 876
rect 27304 864 27310 876
rect 31478 864 31484 876
rect 27304 836 31484 864
rect 27304 824 27310 836
rect 31478 824 31484 836
rect 31536 824 31542 876
rect 38470 824 38476 876
rect 38528 864 38534 876
rect 42518 864 42524 876
rect 38528 836 42524 864
rect 38528 824 38534 836
rect 42518 824 42524 836
rect 42576 824 42582 876
rect 32674 756 32680 808
rect 32732 796 32738 808
rect 36446 796 36452 808
rect 32732 768 36452 796
rect 32732 756 32738 768
rect 36446 756 36452 768
rect 36504 756 36510 808
rect 39390 756 39396 808
rect 39448 796 39454 808
rect 40954 796 40960 808
rect 39448 768 40960 796
rect 39448 756 39454 768
rect 40954 756 40960 768
rect 41012 756 41018 808
rect 34422 688 34428 740
rect 34480 728 34486 740
rect 37090 728 37096 740
rect 34480 700 37096 728
rect 34480 688 34486 700
rect 37090 688 37096 700
rect 37148 688 37154 740
rect 37826 688 37832 740
rect 37884 728 37890 740
rect 40770 728 40776 740
rect 37884 700 40776 728
rect 37884 688 37890 700
rect 40770 688 40776 700
rect 40828 688 40834 740
rect 28902 620 28908 672
rect 28960 660 28966 672
rect 30374 660 30380 672
rect 28960 632 30380 660
rect 28960 620 28966 632
rect 30374 620 30380 632
rect 30432 620 30438 672
rect 33502 620 33508 672
rect 33560 660 33566 672
rect 36814 660 36820 672
rect 33560 632 36820 660
rect 33560 620 33566 632
rect 36814 620 36820 632
rect 36872 620 36878 672
rect 40954 620 40960 672
rect 41012 660 41018 672
rect 41966 660 41972 672
rect 41012 632 41972 660
rect 41012 620 41018 632
rect 41966 620 41972 632
rect 42024 620 42030 672
<< via1 >>
rect 11704 23264 11756 23316
rect 17960 23468 18012 23520
rect 22836 23400 22888 23452
rect 14924 23332 14976 23384
rect 23480 23332 23532 23384
rect 15108 23264 15160 23316
rect 24032 23264 24084 23316
rect 6000 22992 6052 23044
rect 14556 23196 14608 23248
rect 22376 23196 22428 23248
rect 27436 23196 27488 23248
rect 23296 23128 23348 23180
rect 28172 23128 28224 23180
rect 31300 23196 31352 23248
rect 33600 23196 33652 23248
rect 34060 23196 34112 23248
rect 35072 23196 35124 23248
rect 12716 23060 12768 23112
rect 22284 23060 22336 23112
rect 28080 23060 28132 23112
rect 32864 23060 32916 23112
rect 34612 23060 34664 23112
rect 13636 22992 13688 23044
rect 24860 22992 24912 23044
rect 27896 22992 27948 23044
rect 33416 22992 33468 23044
rect 40960 22992 41012 23044
rect 8300 22924 8352 22976
rect 30656 22924 30708 22976
rect 32404 22924 32456 22976
rect 42800 22924 42852 22976
rect 6070 22822 6122 22874
rect 6134 22822 6186 22874
rect 6198 22822 6250 22874
rect 6262 22822 6314 22874
rect 6326 22822 6378 22874
rect 11070 22822 11122 22874
rect 11134 22822 11186 22874
rect 11198 22822 11250 22874
rect 11262 22822 11314 22874
rect 11326 22822 11378 22874
rect 16070 22822 16122 22874
rect 16134 22822 16186 22874
rect 16198 22822 16250 22874
rect 16262 22822 16314 22874
rect 16326 22822 16378 22874
rect 21070 22822 21122 22874
rect 21134 22822 21186 22874
rect 21198 22822 21250 22874
rect 21262 22822 21314 22874
rect 21326 22822 21378 22874
rect 26070 22822 26122 22874
rect 26134 22822 26186 22874
rect 26198 22822 26250 22874
rect 26262 22822 26314 22874
rect 26326 22822 26378 22874
rect 31070 22822 31122 22874
rect 31134 22822 31186 22874
rect 31198 22822 31250 22874
rect 31262 22822 31314 22874
rect 31326 22822 31378 22874
rect 36070 22822 36122 22874
rect 36134 22822 36186 22874
rect 36198 22822 36250 22874
rect 36262 22822 36314 22874
rect 36326 22822 36378 22874
rect 41070 22822 41122 22874
rect 41134 22822 41186 22874
rect 41198 22822 41250 22874
rect 41262 22822 41314 22874
rect 41326 22822 41378 22874
rect 848 22720 900 22772
rect 1768 22720 1820 22772
rect 2780 22720 2832 22772
rect 3608 22720 3660 22772
rect 4528 22720 4580 22772
rect 5448 22720 5500 22772
rect 6460 22720 6512 22772
rect 7288 22720 7340 22772
rect 8208 22720 8260 22772
rect 9128 22720 9180 22772
rect 10048 22720 10100 22772
rect 10968 22720 11020 22772
rect 11888 22720 11940 22772
rect 12808 22720 12860 22772
rect 13636 22763 13688 22772
rect 13636 22729 13645 22763
rect 13645 22729 13679 22763
rect 13679 22729 13688 22763
rect 13636 22720 13688 22729
rect 13820 22720 13872 22772
rect 14556 22763 14608 22772
rect 14556 22729 14565 22763
rect 14565 22729 14599 22763
rect 14599 22729 14608 22763
rect 14556 22720 14608 22729
rect 14648 22720 14700 22772
rect 15108 22720 15160 22772
rect 1952 22652 2004 22704
rect 15568 22720 15620 22772
rect 16488 22720 16540 22772
rect 17408 22720 17460 22772
rect 18328 22720 18380 22772
rect 19248 22720 19300 22772
rect 20168 22720 20220 22772
rect 20996 22720 21048 22772
rect 940 22627 992 22636
rect 940 22593 949 22627
rect 949 22593 983 22627
rect 983 22593 992 22627
rect 940 22584 992 22593
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 3976 22584 4028 22636
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6460 22627 6512 22636
rect 6460 22593 6469 22627
rect 6469 22593 6503 22627
rect 6503 22593 6512 22627
rect 6460 22584 6512 22593
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 8300 22584 8352 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 9220 22627 9272 22636
rect 9220 22593 9229 22627
rect 9229 22593 9263 22627
rect 9263 22593 9272 22627
rect 9220 22584 9272 22593
rect 10140 22627 10192 22636
rect 10140 22593 10149 22627
rect 10149 22593 10183 22627
rect 10183 22593 10192 22627
rect 10140 22584 10192 22593
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 11704 22584 11756 22636
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 12900 22627 12952 22636
rect 12900 22593 12909 22627
rect 12909 22593 12943 22627
rect 12943 22593 12952 22627
rect 12900 22584 12952 22593
rect 13452 22584 13504 22636
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 15384 22627 15436 22636
rect 15384 22593 15393 22627
rect 15393 22593 15427 22627
rect 15427 22593 15436 22627
rect 15384 22584 15436 22593
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 15660 22627 15712 22636
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 16764 22584 16816 22636
rect 17500 22627 17552 22636
rect 17500 22593 17509 22627
rect 17509 22593 17543 22627
rect 17543 22593 17552 22627
rect 17500 22584 17552 22593
rect 18236 22584 18288 22636
rect 19708 22584 19760 22636
rect 20260 22627 20312 22636
rect 20260 22593 20269 22627
rect 20269 22593 20303 22627
rect 20303 22593 20312 22627
rect 20260 22584 20312 22593
rect 22008 22720 22060 22772
rect 22928 22720 22980 22772
rect 23848 22720 23900 22772
rect 24768 22720 24820 22772
rect 25688 22720 25740 22772
rect 26608 22720 26660 22772
rect 3056 22516 3108 22568
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 17132 22516 17184 22568
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 23020 22627 23072 22636
rect 23020 22593 23029 22627
rect 23029 22593 23063 22627
rect 23063 22593 23072 22627
rect 23020 22584 23072 22593
rect 23112 22584 23164 22636
rect 24768 22627 24820 22636
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 26516 22627 26568 22636
rect 26516 22593 26525 22627
rect 26525 22593 26559 22627
rect 26559 22593 26568 22627
rect 26516 22584 26568 22593
rect 27896 22763 27948 22772
rect 27896 22729 27905 22763
rect 27905 22729 27939 22763
rect 27939 22729 27948 22763
rect 27896 22720 27948 22729
rect 28632 22720 28684 22772
rect 29736 22720 29788 22772
rect 30656 22720 30708 22772
rect 27436 22652 27488 22704
rect 27620 22652 27672 22704
rect 32404 22695 32456 22704
rect 32404 22661 32413 22695
rect 32413 22661 32447 22695
rect 32447 22661 32456 22695
rect 32404 22652 32456 22661
rect 28172 22584 28224 22636
rect 25872 22516 25924 22568
rect 28080 22559 28132 22568
rect 28080 22525 28089 22559
rect 28089 22525 28123 22559
rect 28123 22525 28132 22559
rect 28080 22516 28132 22525
rect 10600 22448 10652 22500
rect 15384 22448 15436 22500
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 9588 22380 9640 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 13360 22380 13412 22432
rect 20076 22448 20128 22500
rect 21548 22448 21600 22500
rect 21824 22448 21876 22500
rect 29000 22627 29052 22636
rect 29000 22593 29009 22627
rect 29009 22593 29043 22627
rect 29043 22593 29052 22627
rect 29000 22584 29052 22593
rect 29368 22516 29420 22568
rect 30380 22584 30432 22636
rect 30472 22627 30524 22636
rect 30472 22593 30481 22627
rect 30481 22593 30515 22627
rect 30515 22593 30524 22627
rect 30472 22584 30524 22593
rect 30932 22627 30984 22636
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 31852 22627 31904 22636
rect 31852 22593 31861 22627
rect 31861 22593 31895 22627
rect 31895 22593 31904 22627
rect 31852 22584 31904 22593
rect 32956 22584 33008 22636
rect 33416 22763 33468 22772
rect 33416 22729 33425 22763
rect 33425 22729 33459 22763
rect 33459 22729 33468 22763
rect 33416 22720 33468 22729
rect 39672 22720 39724 22772
rect 40960 22763 41012 22772
rect 40960 22729 40969 22763
rect 40969 22729 41003 22763
rect 41003 22729 41012 22763
rect 40960 22720 41012 22729
rect 42800 22763 42852 22772
rect 42800 22729 42809 22763
rect 42809 22729 42843 22763
rect 42843 22729 42852 22763
rect 42800 22720 42852 22729
rect 34888 22652 34940 22704
rect 33600 22627 33652 22636
rect 33600 22593 33609 22627
rect 33609 22593 33643 22627
rect 33643 22593 33652 22627
rect 33600 22584 33652 22593
rect 30288 22448 30340 22500
rect 32036 22516 32088 22568
rect 32128 22559 32180 22568
rect 32128 22525 32137 22559
rect 32137 22525 32171 22559
rect 32171 22525 32180 22559
rect 32128 22516 32180 22525
rect 32588 22516 32640 22568
rect 34060 22516 34112 22568
rect 34612 22559 34664 22568
rect 34612 22525 34621 22559
rect 34621 22525 34655 22559
rect 34655 22525 34664 22559
rect 34612 22516 34664 22525
rect 15844 22423 15896 22432
rect 15844 22389 15853 22423
rect 15853 22389 15887 22423
rect 15887 22389 15896 22423
rect 15844 22380 15896 22389
rect 17684 22380 17736 22432
rect 19524 22380 19576 22432
rect 21640 22380 21692 22432
rect 24308 22380 24360 22432
rect 25320 22380 25372 22432
rect 26608 22380 26660 22432
rect 27528 22423 27580 22432
rect 27528 22389 27537 22423
rect 27537 22389 27571 22423
rect 27571 22389 27580 22423
rect 27528 22380 27580 22389
rect 27620 22380 27672 22432
rect 33140 22423 33192 22432
rect 33140 22389 33149 22423
rect 33149 22389 33183 22423
rect 33183 22389 33192 22423
rect 33140 22380 33192 22389
rect 33508 22380 33560 22432
rect 33968 22380 34020 22432
rect 35072 22627 35124 22636
rect 35072 22593 35081 22627
rect 35081 22593 35115 22627
rect 35115 22593 35124 22627
rect 35072 22584 35124 22593
rect 36912 22652 36964 22704
rect 35992 22627 36044 22636
rect 35992 22593 36001 22627
rect 36001 22593 36035 22627
rect 36035 22593 36044 22627
rect 35992 22584 36044 22593
rect 37280 22584 37332 22636
rect 37648 22627 37700 22636
rect 37648 22593 37657 22627
rect 37657 22593 37691 22627
rect 37691 22593 37700 22627
rect 37648 22584 37700 22593
rect 38292 22652 38344 22704
rect 38384 22627 38436 22636
rect 38384 22593 38393 22627
rect 38393 22593 38427 22627
rect 38427 22593 38436 22627
rect 38384 22584 38436 22593
rect 38660 22652 38712 22704
rect 39488 22584 39540 22636
rect 40408 22584 40460 22636
rect 41604 22627 41656 22636
rect 41604 22593 41613 22627
rect 41613 22593 41647 22627
rect 41647 22593 41656 22627
rect 41604 22584 41656 22593
rect 42248 22584 42300 22636
rect 43168 22584 43220 22636
rect 44272 22584 44324 22636
rect 45192 22627 45244 22636
rect 45192 22593 45201 22627
rect 45201 22593 45235 22627
rect 45235 22593 45244 22627
rect 45192 22584 45244 22593
rect 37096 22559 37148 22568
rect 37096 22525 37105 22559
rect 37105 22525 37139 22559
rect 37139 22525 37148 22559
rect 37096 22516 37148 22525
rect 37556 22516 37608 22568
rect 37372 22448 37424 22500
rect 35164 22423 35216 22432
rect 35164 22389 35173 22423
rect 35173 22389 35207 22423
rect 35207 22389 35216 22423
rect 35164 22380 35216 22389
rect 35716 22423 35768 22432
rect 35716 22389 35725 22423
rect 35725 22389 35759 22423
rect 35759 22389 35768 22423
rect 35716 22380 35768 22389
rect 35808 22423 35860 22432
rect 35808 22389 35817 22423
rect 35817 22389 35851 22423
rect 35851 22389 35860 22423
rect 35808 22380 35860 22389
rect 36084 22423 36136 22432
rect 36084 22389 36093 22423
rect 36093 22389 36127 22423
rect 36127 22389 36136 22423
rect 36084 22380 36136 22389
rect 36636 22423 36688 22432
rect 36636 22389 36645 22423
rect 36645 22389 36679 22423
rect 36679 22389 36688 22423
rect 36636 22380 36688 22389
rect 37924 22448 37976 22500
rect 38016 22423 38068 22432
rect 38016 22389 38025 22423
rect 38025 22389 38059 22423
rect 38059 22389 38068 22423
rect 38016 22380 38068 22389
rect 38292 22380 38344 22432
rect 40960 22448 41012 22500
rect 38844 22423 38896 22432
rect 38844 22389 38853 22423
rect 38853 22389 38887 22423
rect 38887 22389 38896 22423
rect 38844 22380 38896 22389
rect 39212 22423 39264 22432
rect 39212 22389 39221 22423
rect 39221 22389 39255 22423
rect 39255 22389 39264 22423
rect 39212 22380 39264 22389
rect 39304 22380 39356 22432
rect 40500 22423 40552 22432
rect 40500 22389 40509 22423
rect 40509 22389 40543 22423
rect 40543 22389 40552 22423
rect 40500 22380 40552 22389
rect 41420 22423 41472 22432
rect 41420 22389 41429 22423
rect 41429 22389 41463 22423
rect 41463 22389 41472 22423
rect 41420 22380 41472 22389
rect 42156 22380 42208 22432
rect 42708 22380 42760 22432
rect 43260 22423 43312 22432
rect 43260 22389 43269 22423
rect 43269 22389 43303 22423
rect 43303 22389 43312 22423
rect 43260 22380 43312 22389
rect 43904 22380 43956 22432
rect 44180 22423 44232 22432
rect 44180 22389 44189 22423
rect 44189 22389 44223 22423
rect 44223 22389 44232 22423
rect 44180 22380 44232 22389
rect 44364 22423 44416 22432
rect 44364 22389 44373 22423
rect 44373 22389 44407 22423
rect 44407 22389 44416 22423
rect 44364 22380 44416 22389
rect 45008 22423 45060 22432
rect 45008 22389 45017 22423
rect 45017 22389 45051 22423
rect 45051 22389 45060 22423
rect 45008 22380 45060 22389
rect 3570 22278 3622 22330
rect 3634 22278 3686 22330
rect 3698 22278 3750 22330
rect 3762 22278 3814 22330
rect 3826 22278 3878 22330
rect 8570 22278 8622 22330
rect 8634 22278 8686 22330
rect 8698 22278 8750 22330
rect 8762 22278 8814 22330
rect 8826 22278 8878 22330
rect 13570 22278 13622 22330
rect 13634 22278 13686 22330
rect 13698 22278 13750 22330
rect 13762 22278 13814 22330
rect 13826 22278 13878 22330
rect 18570 22278 18622 22330
rect 18634 22278 18686 22330
rect 18698 22278 18750 22330
rect 18762 22278 18814 22330
rect 18826 22278 18878 22330
rect 23570 22278 23622 22330
rect 23634 22278 23686 22330
rect 23698 22278 23750 22330
rect 23762 22278 23814 22330
rect 23826 22278 23878 22330
rect 28570 22278 28622 22330
rect 28634 22278 28686 22330
rect 28698 22278 28750 22330
rect 28762 22278 28814 22330
rect 28826 22278 28878 22330
rect 33570 22278 33622 22330
rect 33634 22278 33686 22330
rect 33698 22278 33750 22330
rect 33762 22278 33814 22330
rect 33826 22278 33878 22330
rect 38570 22278 38622 22330
rect 38634 22278 38686 22330
rect 38698 22278 38750 22330
rect 38762 22278 38814 22330
rect 38826 22278 38878 22330
rect 43570 22278 43622 22330
rect 43634 22278 43686 22330
rect 43698 22278 43750 22330
rect 43762 22278 43814 22330
rect 43826 22278 43878 22330
rect 940 22176 992 22228
rect 1860 22176 1912 22228
rect 3240 22176 3292 22228
rect 3976 22176 4028 22228
rect 4620 22219 4672 22228
rect 4620 22185 4629 22219
rect 4629 22185 4663 22219
rect 4663 22185 4672 22219
rect 4620 22176 4672 22185
rect 5816 22176 5868 22228
rect 6000 22219 6052 22228
rect 6000 22185 6009 22219
rect 6009 22185 6043 22219
rect 6043 22185 6052 22219
rect 6000 22176 6052 22185
rect 6460 22219 6512 22228
rect 6460 22185 6469 22219
rect 6469 22185 6503 22219
rect 6503 22185 6512 22219
rect 6460 22176 6512 22185
rect 7380 22176 7432 22228
rect 8392 22176 8444 22228
rect 9220 22176 9272 22228
rect 10140 22219 10192 22228
rect 10140 22185 10149 22219
rect 10149 22185 10183 22219
rect 10183 22185 10192 22219
rect 10140 22176 10192 22185
rect 11152 22176 11204 22228
rect 11980 22176 12032 22228
rect 12900 22176 12952 22228
rect 13452 22176 13504 22228
rect 14004 22176 14056 22228
rect 14740 22176 14792 22228
rect 16764 22219 16816 22228
rect 16764 22185 16773 22219
rect 16773 22185 16807 22219
rect 16807 22185 16816 22219
rect 16764 22176 16816 22185
rect 17500 22176 17552 22228
rect 17684 22176 17736 22228
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 3056 21972 3108 22024
rect 4436 22015 4488 22024
rect 4436 21981 4445 22015
rect 4445 21981 4479 22015
rect 4479 21981 4488 22015
rect 4436 21972 4488 21981
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 16304 22108 16356 22160
rect 18236 22219 18288 22228
rect 18236 22185 18245 22219
rect 18245 22185 18279 22219
rect 18279 22185 18288 22219
rect 18236 22176 18288 22185
rect 19708 22219 19760 22228
rect 19708 22185 19717 22219
rect 19717 22185 19751 22219
rect 19751 22185 19760 22219
rect 19708 22176 19760 22185
rect 20260 22176 20312 22228
rect 5448 21904 5500 21956
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 9588 22015 9640 22024
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 12072 21972 12124 22024
rect 19524 22108 19576 22160
rect 22192 22176 22244 22228
rect 23020 22176 23072 22228
rect 23112 22219 23164 22228
rect 23112 22185 23121 22219
rect 23121 22185 23155 22219
rect 23155 22185 23164 22219
rect 23112 22176 23164 22185
rect 24768 22176 24820 22228
rect 29368 22219 29420 22228
rect 29368 22185 29377 22219
rect 29377 22185 29411 22219
rect 29411 22185 29420 22219
rect 29368 22176 29420 22185
rect 33140 22176 33192 22228
rect 33968 22176 34020 22228
rect 36452 22176 36504 22228
rect 40960 22219 41012 22228
rect 40960 22185 40969 22219
rect 40969 22185 41003 22219
rect 41003 22185 41012 22219
rect 40960 22176 41012 22185
rect 12716 21972 12768 22024
rect 13084 21972 13136 22024
rect 6460 21836 6512 21888
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 7288 21836 7340 21888
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 11612 21836 11664 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 13452 21836 13504 21888
rect 13912 21904 13964 21956
rect 14464 21972 14516 22024
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 15660 21972 15712 22024
rect 16396 21972 16448 22024
rect 15936 21904 15988 21956
rect 14096 21836 14148 21888
rect 15660 21836 15712 21888
rect 16764 21904 16816 21956
rect 17316 21972 17368 22024
rect 17500 21972 17552 22024
rect 17868 21972 17920 22024
rect 18328 21904 18380 21956
rect 18696 21972 18748 22024
rect 19064 21972 19116 22024
rect 19156 21972 19208 22024
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 18788 21947 18840 21956
rect 18788 21913 18797 21947
rect 18797 21913 18831 21947
rect 18831 21913 18840 21947
rect 18788 21904 18840 21913
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 21548 21972 21600 22024
rect 21640 21972 21692 22024
rect 22376 21972 22428 22024
rect 32036 22108 32088 22160
rect 32496 22151 32548 22160
rect 32496 22117 32505 22151
rect 32505 22117 32539 22151
rect 32539 22117 32548 22151
rect 32496 22108 32548 22117
rect 32680 22108 32732 22160
rect 35440 22108 35492 22160
rect 24768 22083 24820 22092
rect 24768 22049 24777 22083
rect 24777 22049 24811 22083
rect 24811 22049 24820 22083
rect 24768 22040 24820 22049
rect 27804 22083 27856 22092
rect 27804 22049 27813 22083
rect 27813 22049 27847 22083
rect 27847 22049 27856 22083
rect 27804 22040 27856 22049
rect 28080 22040 28132 22092
rect 28448 22040 28500 22092
rect 30012 22083 30064 22092
rect 30012 22049 30021 22083
rect 30021 22049 30055 22083
rect 30055 22049 30064 22083
rect 30012 22040 30064 22049
rect 23388 21972 23440 22024
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 17040 21836 17092 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 18236 21836 18288 21888
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 19432 21836 19484 21888
rect 19708 21836 19760 21888
rect 19800 21836 19852 21888
rect 19892 21836 19944 21888
rect 20444 21836 20496 21888
rect 22192 21836 22244 21888
rect 22284 21836 22336 21888
rect 23204 21836 23256 21888
rect 23480 21836 23532 21888
rect 23848 21879 23900 21888
rect 23848 21845 23857 21879
rect 23857 21845 23891 21879
rect 23891 21845 23900 21879
rect 23848 21836 23900 21845
rect 25136 22015 25188 22024
rect 25136 21981 25145 22015
rect 25145 21981 25179 22015
rect 25179 21981 25188 22015
rect 25136 21972 25188 21981
rect 25320 22015 25372 22024
rect 25320 21981 25329 22015
rect 25329 21981 25363 22015
rect 25363 21981 25372 22015
rect 25320 21972 25372 21981
rect 24492 21947 24544 21956
rect 24492 21913 24501 21947
rect 24501 21913 24535 21947
rect 24535 21913 24544 21947
rect 24492 21904 24544 21913
rect 25320 21836 25372 21888
rect 25596 21947 25648 21956
rect 25596 21913 25605 21947
rect 25605 21913 25639 21947
rect 25639 21913 25648 21947
rect 25596 21904 25648 21913
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 28908 22015 28960 22024
rect 28908 21981 28917 22015
rect 28917 21981 28951 22015
rect 28951 21981 28960 22015
rect 28908 21972 28960 21981
rect 30196 22015 30248 22024
rect 30196 21981 30205 22015
rect 30205 21981 30239 22015
rect 30239 21981 30248 22015
rect 30196 21972 30248 21981
rect 30288 21972 30340 22024
rect 25780 21836 25832 21888
rect 25964 21836 26016 21888
rect 27068 21879 27120 21888
rect 27068 21845 27077 21879
rect 27077 21845 27111 21879
rect 27111 21845 27120 21879
rect 27068 21836 27120 21845
rect 27896 21904 27948 21956
rect 28356 21947 28408 21956
rect 28356 21913 28365 21947
rect 28365 21913 28399 21947
rect 28399 21913 28408 21947
rect 28356 21904 28408 21913
rect 30564 21904 30616 21956
rect 27528 21836 27580 21888
rect 27988 21879 28040 21888
rect 27988 21845 27997 21879
rect 27997 21845 28031 21879
rect 28031 21845 28040 21879
rect 27988 21836 28040 21845
rect 28080 21836 28132 21888
rect 29092 21879 29144 21888
rect 29092 21845 29101 21879
rect 29101 21845 29135 21879
rect 29135 21845 29144 21879
rect 29092 21836 29144 21845
rect 30012 21836 30064 21888
rect 30932 21904 30984 21956
rect 32864 22040 32916 22092
rect 33324 22040 33376 22092
rect 37372 22108 37424 22160
rect 38200 22108 38252 22160
rect 32496 21972 32548 22024
rect 32680 21904 32732 21956
rect 32312 21836 32364 21888
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 33048 21972 33100 22024
rect 33876 22015 33928 22024
rect 33876 21981 33885 22015
rect 33885 21981 33919 22015
rect 33919 21981 33928 22015
rect 33876 21972 33928 21981
rect 35440 21972 35492 22024
rect 37372 21972 37424 22024
rect 36544 21904 36596 21956
rect 40040 22040 40092 22092
rect 43168 22040 43220 22092
rect 38936 21972 38988 22024
rect 39212 21972 39264 22024
rect 41696 21972 41748 22024
rect 43904 21972 43956 22024
rect 35624 21836 35676 21888
rect 37740 21879 37792 21888
rect 37740 21845 37749 21879
rect 37749 21845 37783 21879
rect 37783 21845 37792 21879
rect 37740 21836 37792 21845
rect 37832 21879 37884 21888
rect 37832 21845 37841 21879
rect 37841 21845 37875 21879
rect 37875 21845 37884 21879
rect 37832 21836 37884 21845
rect 38292 21879 38344 21888
rect 38292 21845 38301 21879
rect 38301 21845 38335 21879
rect 38335 21845 38344 21879
rect 38292 21836 38344 21845
rect 38384 21836 38436 21888
rect 38936 21836 38988 21888
rect 39672 21879 39724 21888
rect 39672 21845 39681 21879
rect 39681 21845 39715 21879
rect 39715 21845 39724 21879
rect 39672 21836 39724 21845
rect 39764 21836 39816 21888
rect 41972 21836 42024 21888
rect 42156 21879 42208 21888
rect 42156 21845 42165 21879
rect 42165 21845 42199 21879
rect 42199 21845 42208 21879
rect 42156 21836 42208 21845
rect 42800 21879 42852 21888
rect 42800 21845 42809 21879
rect 42809 21845 42843 21879
rect 42843 21845 42852 21879
rect 42800 21836 42852 21845
rect 6070 21734 6122 21786
rect 6134 21734 6186 21786
rect 6198 21734 6250 21786
rect 6262 21734 6314 21786
rect 6326 21734 6378 21786
rect 11070 21734 11122 21786
rect 11134 21734 11186 21786
rect 11198 21734 11250 21786
rect 11262 21734 11314 21786
rect 11326 21734 11378 21786
rect 16070 21734 16122 21786
rect 16134 21734 16186 21786
rect 16198 21734 16250 21786
rect 16262 21734 16314 21786
rect 16326 21734 16378 21786
rect 21070 21734 21122 21786
rect 21134 21734 21186 21786
rect 21198 21734 21250 21786
rect 21262 21734 21314 21786
rect 21326 21734 21378 21786
rect 26070 21734 26122 21786
rect 26134 21734 26186 21786
rect 26198 21734 26250 21786
rect 26262 21734 26314 21786
rect 26326 21734 26378 21786
rect 31070 21734 31122 21786
rect 31134 21734 31186 21786
rect 31198 21734 31250 21786
rect 31262 21734 31314 21786
rect 31326 21734 31378 21786
rect 36070 21734 36122 21786
rect 36134 21734 36186 21786
rect 36198 21734 36250 21786
rect 36262 21734 36314 21786
rect 36326 21734 36378 21786
rect 41070 21734 41122 21786
rect 41134 21734 41186 21786
rect 41198 21734 41250 21786
rect 41262 21734 41314 21786
rect 41326 21734 41378 21786
rect 10048 21632 10100 21684
rect 14280 21632 14332 21684
rect 14740 21632 14792 21684
rect 13912 21564 13964 21616
rect 13084 21496 13136 21548
rect 6736 21428 6788 21480
rect 7104 21428 7156 21480
rect 12072 21428 12124 21480
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 14464 21428 14516 21480
rect 14556 21428 14608 21480
rect 15844 21564 15896 21616
rect 16396 21607 16448 21616
rect 16396 21573 16405 21607
rect 16405 21573 16439 21607
rect 16439 21573 16448 21607
rect 16396 21564 16448 21573
rect 18696 21632 18748 21684
rect 18788 21632 18840 21684
rect 15936 21496 15988 21548
rect 5908 21292 5960 21344
rect 6828 21335 6880 21344
rect 6828 21301 6837 21335
rect 6837 21301 6871 21335
rect 6871 21301 6880 21335
rect 9312 21403 9364 21412
rect 9312 21369 9321 21403
rect 9321 21369 9355 21403
rect 9355 21369 9364 21403
rect 9312 21360 9364 21369
rect 6828 21292 6880 21301
rect 7288 21292 7340 21344
rect 10232 21292 10284 21344
rect 11060 21292 11112 21344
rect 12624 21335 12676 21344
rect 12624 21301 12633 21335
rect 12633 21301 12667 21335
rect 12667 21301 12676 21335
rect 12624 21292 12676 21301
rect 15476 21360 15528 21412
rect 15660 21360 15712 21412
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 16856 21496 16908 21548
rect 18236 21564 18288 21616
rect 16304 21428 16356 21480
rect 17684 21539 17736 21548
rect 17684 21505 17693 21539
rect 17693 21505 17727 21539
rect 17727 21505 17736 21539
rect 17684 21496 17736 21505
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 18052 21428 18104 21480
rect 18972 21428 19024 21480
rect 19432 21675 19484 21684
rect 19432 21641 19441 21675
rect 19441 21641 19475 21675
rect 19475 21641 19484 21675
rect 19432 21632 19484 21641
rect 19892 21632 19944 21684
rect 20168 21632 20220 21684
rect 20628 21632 20680 21684
rect 20812 21632 20864 21684
rect 20720 21564 20772 21616
rect 21640 21564 21692 21616
rect 19616 21428 19668 21480
rect 19892 21539 19944 21548
rect 19892 21505 19901 21539
rect 19901 21505 19935 21539
rect 19935 21505 19944 21539
rect 19892 21496 19944 21505
rect 19984 21428 20036 21480
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 20628 21539 20680 21548
rect 20628 21505 20637 21539
rect 20637 21505 20671 21539
rect 20671 21505 20680 21539
rect 20628 21496 20680 21505
rect 20444 21428 20496 21480
rect 20168 21360 20220 21412
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 17960 21292 18012 21344
rect 19984 21292 20036 21344
rect 20352 21292 20404 21344
rect 21088 21360 21140 21412
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 21548 21496 21600 21548
rect 22284 21564 22336 21616
rect 23572 21632 23624 21684
rect 25780 21675 25832 21684
rect 25780 21641 25789 21675
rect 25789 21641 25823 21675
rect 25823 21641 25832 21675
rect 25780 21632 25832 21641
rect 25872 21675 25924 21684
rect 25872 21641 25881 21675
rect 25881 21641 25915 21675
rect 25915 21641 25924 21675
rect 25872 21632 25924 21641
rect 27620 21632 27672 21684
rect 28908 21632 28960 21684
rect 30380 21675 30432 21684
rect 30380 21641 30389 21675
rect 30389 21641 30423 21675
rect 30423 21641 30432 21675
rect 30380 21632 30432 21641
rect 24124 21564 24176 21616
rect 25320 21564 25372 21616
rect 25504 21564 25556 21616
rect 26056 21564 26108 21616
rect 22008 21471 22060 21480
rect 22008 21437 22017 21471
rect 22017 21437 22051 21471
rect 22051 21437 22060 21471
rect 22008 21428 22060 21437
rect 23204 21428 23256 21480
rect 20536 21292 20588 21344
rect 23940 21428 23992 21480
rect 24492 21428 24544 21480
rect 26608 21607 26660 21616
rect 26608 21573 26617 21607
rect 26617 21573 26651 21607
rect 26651 21573 26660 21607
rect 26608 21564 26660 21573
rect 32588 21632 32640 21684
rect 33876 21632 33928 21684
rect 27160 21428 27212 21480
rect 27896 21428 27948 21480
rect 27804 21360 27856 21412
rect 21732 21292 21784 21344
rect 23848 21335 23900 21344
rect 23848 21301 23878 21335
rect 23878 21301 23900 21335
rect 23848 21292 23900 21301
rect 26976 21292 27028 21344
rect 28080 21335 28132 21344
rect 28080 21301 28089 21335
rect 28089 21301 28123 21335
rect 28123 21301 28132 21335
rect 28080 21292 28132 21301
rect 28264 21360 28316 21412
rect 29368 21496 29420 21548
rect 29920 21539 29972 21548
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 30656 21496 30708 21548
rect 30748 21539 30800 21548
rect 30748 21505 30757 21539
rect 30757 21505 30791 21539
rect 30791 21505 30800 21539
rect 30748 21496 30800 21505
rect 31024 21496 31076 21548
rect 30104 21471 30156 21480
rect 30104 21437 30113 21471
rect 30113 21437 30147 21471
rect 30147 21437 30156 21471
rect 30104 21428 30156 21437
rect 31392 21428 31444 21480
rect 30196 21360 30248 21412
rect 30748 21360 30800 21412
rect 30932 21292 30984 21344
rect 32220 21428 32272 21480
rect 32312 21428 32364 21480
rect 34060 21564 34112 21616
rect 36452 21632 36504 21684
rect 37924 21632 37976 21684
rect 40500 21632 40552 21684
rect 40960 21632 41012 21684
rect 41972 21675 42024 21684
rect 41972 21641 41981 21675
rect 41981 21641 42015 21675
rect 42015 21641 42024 21675
rect 41972 21632 42024 21641
rect 42800 21632 42852 21684
rect 44180 21675 44232 21684
rect 44180 21641 44189 21675
rect 44189 21641 44223 21675
rect 44223 21641 44232 21675
rect 44548 21675 44600 21684
rect 44180 21632 44232 21641
rect 44548 21641 44557 21675
rect 44557 21641 44591 21675
rect 44591 21641 44600 21675
rect 44548 21632 44600 21641
rect 43904 21564 43956 21616
rect 33140 21428 33192 21480
rect 33324 21471 33376 21480
rect 33324 21437 33333 21471
rect 33333 21437 33367 21471
rect 33367 21437 33376 21471
rect 33324 21428 33376 21437
rect 32864 21360 32916 21412
rect 34060 21428 34112 21480
rect 35440 21496 35492 21548
rect 35532 21539 35584 21548
rect 35532 21505 35541 21539
rect 35541 21505 35575 21539
rect 35575 21505 35584 21539
rect 35532 21496 35584 21505
rect 35900 21496 35952 21548
rect 36452 21539 36504 21548
rect 36452 21505 36461 21539
rect 36461 21505 36495 21539
rect 36495 21505 36504 21539
rect 36452 21496 36504 21505
rect 36544 21496 36596 21548
rect 37924 21496 37976 21548
rect 39764 21496 39816 21548
rect 34980 21428 35032 21480
rect 35624 21471 35676 21480
rect 35624 21437 35633 21471
rect 35633 21437 35667 21471
rect 35667 21437 35676 21471
rect 35624 21428 35676 21437
rect 35716 21471 35768 21480
rect 35716 21437 35725 21471
rect 35725 21437 35759 21471
rect 35759 21437 35768 21471
rect 35716 21428 35768 21437
rect 37464 21428 37516 21480
rect 38384 21428 38436 21480
rect 38016 21360 38068 21412
rect 40776 21471 40828 21480
rect 40776 21437 40785 21471
rect 40785 21437 40819 21471
rect 40819 21437 40828 21471
rect 40776 21428 40828 21437
rect 40868 21471 40920 21480
rect 40868 21437 40877 21471
rect 40877 21437 40911 21471
rect 40911 21437 40920 21471
rect 40868 21428 40920 21437
rect 31944 21292 31996 21344
rect 32128 21292 32180 21344
rect 33048 21292 33100 21344
rect 33232 21335 33284 21344
rect 33232 21301 33241 21335
rect 33241 21301 33275 21335
rect 33275 21301 33284 21335
rect 33232 21292 33284 21301
rect 33416 21292 33468 21344
rect 33692 21292 33744 21344
rect 36912 21292 36964 21344
rect 38476 21292 38528 21344
rect 40500 21360 40552 21412
rect 42156 21292 42208 21344
rect 44272 21292 44324 21344
rect 44916 21335 44968 21344
rect 44916 21301 44925 21335
rect 44925 21301 44959 21335
rect 44959 21301 44968 21335
rect 44916 21292 44968 21301
rect 3570 21190 3622 21242
rect 3634 21190 3686 21242
rect 3698 21190 3750 21242
rect 3762 21190 3814 21242
rect 3826 21190 3878 21242
rect 8570 21190 8622 21242
rect 8634 21190 8686 21242
rect 8698 21190 8750 21242
rect 8762 21190 8814 21242
rect 8826 21190 8878 21242
rect 13570 21190 13622 21242
rect 13634 21190 13686 21242
rect 13698 21190 13750 21242
rect 13762 21190 13814 21242
rect 13826 21190 13878 21242
rect 18570 21190 18622 21242
rect 18634 21190 18686 21242
rect 18698 21190 18750 21242
rect 18762 21190 18814 21242
rect 18826 21190 18878 21242
rect 23570 21190 23622 21242
rect 23634 21190 23686 21242
rect 23698 21190 23750 21242
rect 23762 21190 23814 21242
rect 23826 21190 23878 21242
rect 28570 21190 28622 21242
rect 28634 21190 28686 21242
rect 28698 21190 28750 21242
rect 28762 21190 28814 21242
rect 28826 21190 28878 21242
rect 33570 21190 33622 21242
rect 33634 21190 33686 21242
rect 33698 21190 33750 21242
rect 33762 21190 33814 21242
rect 33826 21190 33878 21242
rect 38570 21190 38622 21242
rect 38634 21190 38686 21242
rect 38698 21190 38750 21242
rect 38762 21190 38814 21242
rect 38826 21190 38878 21242
rect 43570 21190 43622 21242
rect 43634 21190 43686 21242
rect 43698 21190 43750 21242
rect 43762 21190 43814 21242
rect 43826 21190 43878 21242
rect 12716 21088 12768 21140
rect 14004 21088 14056 21140
rect 13360 21020 13412 21072
rect 13820 21020 13872 21072
rect 14556 21088 14608 21140
rect 15476 21088 15528 21140
rect 15568 21088 15620 21140
rect 17684 21088 17736 21140
rect 940 20927 992 20936
rect 940 20893 949 20927
rect 949 20893 983 20927
rect 983 20893 992 20927
rect 940 20884 992 20893
rect 6644 20859 6696 20868
rect 6644 20825 6653 20859
rect 6653 20825 6687 20859
rect 6687 20825 6696 20859
rect 6644 20816 6696 20825
rect 7932 20816 7984 20868
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 11888 20884 11940 20936
rect 9312 20816 9364 20868
rect 10232 20816 10284 20868
rect 14372 20884 14424 20936
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 14740 20884 14792 20893
rect 756 20791 808 20800
rect 756 20757 765 20791
rect 765 20757 799 20791
rect 799 20757 808 20791
rect 756 20748 808 20757
rect 3148 20748 3200 20800
rect 3792 20748 3844 20800
rect 5540 20791 5592 20800
rect 5540 20757 5549 20791
rect 5549 20757 5583 20791
rect 5583 20757 5592 20791
rect 5540 20748 5592 20757
rect 5632 20748 5684 20800
rect 5908 20791 5960 20800
rect 5908 20757 5917 20791
rect 5917 20757 5951 20791
rect 5951 20757 5960 20791
rect 5908 20748 5960 20757
rect 13544 20816 13596 20868
rect 14464 20816 14516 20868
rect 16120 20884 16172 20936
rect 16488 20884 16540 20936
rect 15384 20816 15436 20868
rect 22008 21088 22060 21140
rect 25872 21088 25924 21140
rect 26516 21131 26568 21140
rect 26516 21097 26525 21131
rect 26525 21097 26559 21131
rect 26559 21097 26568 21131
rect 26516 21088 26568 21097
rect 19524 21020 19576 21072
rect 19984 21020 20036 21072
rect 21732 21020 21784 21072
rect 16856 20816 16908 20868
rect 17408 20816 17460 20868
rect 18972 20884 19024 20936
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 11428 20748 11480 20800
rect 12716 20748 12768 20800
rect 15108 20748 15160 20800
rect 15936 20748 15988 20800
rect 16396 20748 16448 20800
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 17776 20748 17828 20800
rect 18328 20748 18380 20800
rect 19064 20748 19116 20800
rect 22008 20952 22060 21004
rect 23480 20952 23532 21004
rect 24768 20952 24820 21004
rect 27344 21063 27396 21072
rect 27344 21029 27353 21063
rect 27353 21029 27387 21063
rect 27387 21029 27396 21063
rect 27344 21020 27396 21029
rect 28356 21020 28408 21072
rect 28908 21020 28960 21072
rect 26976 20995 27028 21004
rect 26976 20961 26985 20995
rect 26985 20961 27019 20995
rect 27019 20961 27028 20995
rect 26976 20952 27028 20961
rect 27160 20995 27212 21004
rect 27160 20961 27169 20995
rect 27169 20961 27203 20995
rect 27203 20961 27212 20995
rect 27160 20952 27212 20961
rect 27804 20952 27856 21004
rect 30748 21131 30800 21140
rect 30748 21097 30757 21131
rect 30757 21097 30791 21131
rect 30791 21097 30800 21131
rect 30748 21088 30800 21097
rect 31944 21088 31996 21140
rect 32220 21088 32272 21140
rect 32864 21131 32916 21140
rect 32864 21097 32873 21131
rect 32873 21097 32907 21131
rect 32907 21097 32916 21131
rect 32864 21088 32916 21097
rect 33048 21088 33100 21140
rect 30564 21020 30616 21072
rect 20076 20816 20128 20868
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 21732 20884 21784 20936
rect 22468 20927 22520 20936
rect 22468 20893 22477 20927
rect 22477 20893 22511 20927
rect 22511 20893 22520 20927
rect 22468 20884 22520 20893
rect 22560 20884 22612 20936
rect 23112 20927 23164 20936
rect 23112 20893 23121 20927
rect 23121 20893 23155 20927
rect 23155 20893 23164 20927
rect 23112 20884 23164 20893
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 19984 20748 20036 20800
rect 20260 20748 20312 20800
rect 20536 20748 20588 20800
rect 20996 20816 21048 20868
rect 21180 20816 21232 20868
rect 23204 20816 23256 20868
rect 25320 20884 25372 20936
rect 27988 20884 28040 20936
rect 28172 20927 28224 20936
rect 28172 20893 28181 20927
rect 28181 20893 28215 20927
rect 28215 20893 28224 20927
rect 28172 20884 28224 20893
rect 24308 20816 24360 20868
rect 20904 20748 20956 20800
rect 21732 20748 21784 20800
rect 22468 20748 22520 20800
rect 23020 20791 23072 20800
rect 23020 20757 23029 20791
rect 23029 20757 23063 20791
rect 23063 20757 23072 20791
rect 23020 20748 23072 20757
rect 24124 20748 24176 20800
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 27068 20816 27120 20868
rect 28816 20884 28868 20936
rect 28908 20927 28960 20936
rect 28908 20893 28917 20927
rect 28917 20893 28951 20927
rect 28951 20893 28960 20927
rect 28908 20884 28960 20893
rect 30288 20884 30340 20936
rect 31484 20952 31536 21004
rect 33140 21020 33192 21072
rect 33324 20952 33376 21004
rect 33416 20952 33468 21004
rect 28356 20859 28408 20868
rect 28356 20825 28365 20859
rect 28365 20825 28399 20859
rect 28399 20825 28408 20859
rect 28356 20816 28408 20825
rect 27620 20748 27672 20800
rect 28080 20748 28132 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 29184 20859 29236 20868
rect 29184 20825 29193 20859
rect 29193 20825 29227 20859
rect 29227 20825 29236 20859
rect 29184 20816 29236 20825
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 31760 20884 31812 20936
rect 34520 21088 34572 21140
rect 35532 21088 35584 21140
rect 37280 21088 37332 21140
rect 38292 21088 38344 21140
rect 33968 20952 34020 21004
rect 36176 20995 36228 21004
rect 36176 20961 36185 20995
rect 36185 20961 36219 20995
rect 36219 20961 36228 20995
rect 36176 20952 36228 20961
rect 31852 20816 31904 20868
rect 32588 20816 32640 20868
rect 29368 20748 29420 20800
rect 30104 20748 30156 20800
rect 31760 20791 31812 20800
rect 31760 20757 31769 20791
rect 31769 20757 31803 20791
rect 31803 20757 31812 20791
rect 31760 20748 31812 20757
rect 35440 20884 35492 20936
rect 33416 20816 33468 20868
rect 33232 20748 33284 20800
rect 34060 20748 34112 20800
rect 35992 20748 36044 20800
rect 37372 20952 37424 21004
rect 40500 21088 40552 21140
rect 40776 21088 40828 21140
rect 38384 20995 38436 21004
rect 38384 20961 38393 20995
rect 38393 20961 38427 20995
rect 38427 20961 38436 20995
rect 38384 20952 38436 20961
rect 37740 20884 37792 20936
rect 37924 20884 37976 20936
rect 38108 20884 38160 20936
rect 42800 21088 42852 21140
rect 44548 21131 44600 21140
rect 44548 21097 44557 21131
rect 44557 21097 44591 21131
rect 44591 21097 44600 21131
rect 44548 21088 44600 21097
rect 41604 20995 41656 21004
rect 41604 20961 41613 20995
rect 41613 20961 41647 20995
rect 41647 20961 41656 20995
rect 41604 20952 41656 20961
rect 39212 20927 39264 20936
rect 39212 20893 39221 20927
rect 39221 20893 39255 20927
rect 39255 20893 39264 20927
rect 39212 20884 39264 20893
rect 41420 20884 41472 20936
rect 37832 20816 37884 20868
rect 38660 20816 38712 20868
rect 38568 20791 38620 20800
rect 38568 20757 38577 20791
rect 38577 20757 38611 20791
rect 38611 20757 38620 20791
rect 38568 20748 38620 20757
rect 39764 20816 39816 20868
rect 39028 20748 39080 20800
rect 40868 20816 40920 20868
rect 43168 20816 43220 20868
rect 40960 20748 41012 20800
rect 41880 20791 41932 20800
rect 41880 20757 41889 20791
rect 41889 20757 41923 20791
rect 41923 20757 41932 20791
rect 41880 20748 41932 20757
rect 42340 20791 42392 20800
rect 42340 20757 42349 20791
rect 42349 20757 42383 20791
rect 42383 20757 42392 20791
rect 42340 20748 42392 20757
rect 43444 20748 43496 20800
rect 44180 20816 44232 20868
rect 45192 20859 45244 20868
rect 45192 20825 45201 20859
rect 45201 20825 45235 20859
rect 45235 20825 45244 20859
rect 45192 20816 45244 20825
rect 44272 20748 44324 20800
rect 44732 20748 44784 20800
rect 6070 20646 6122 20698
rect 6134 20646 6186 20698
rect 6198 20646 6250 20698
rect 6262 20646 6314 20698
rect 6326 20646 6378 20698
rect 11070 20646 11122 20698
rect 11134 20646 11186 20698
rect 11198 20646 11250 20698
rect 11262 20646 11314 20698
rect 11326 20646 11378 20698
rect 16070 20646 16122 20698
rect 16134 20646 16186 20698
rect 16198 20646 16250 20698
rect 16262 20646 16314 20698
rect 16326 20646 16378 20698
rect 21070 20646 21122 20698
rect 21134 20646 21186 20698
rect 21198 20646 21250 20698
rect 21262 20646 21314 20698
rect 21326 20646 21378 20698
rect 26070 20646 26122 20698
rect 26134 20646 26186 20698
rect 26198 20646 26250 20698
rect 26262 20646 26314 20698
rect 26326 20646 26378 20698
rect 31070 20646 31122 20698
rect 31134 20646 31186 20698
rect 31198 20646 31250 20698
rect 31262 20646 31314 20698
rect 31326 20646 31378 20698
rect 36070 20646 36122 20698
rect 36134 20646 36186 20698
rect 36198 20646 36250 20698
rect 36262 20646 36314 20698
rect 36326 20646 36378 20698
rect 41070 20646 41122 20698
rect 41134 20646 41186 20698
rect 41198 20646 41250 20698
rect 41262 20646 41314 20698
rect 41326 20646 41378 20698
rect 756 20476 808 20528
rect 6644 20544 6696 20596
rect 9312 20544 9364 20596
rect 9680 20544 9732 20596
rect 12532 20587 12584 20596
rect 12532 20553 12541 20587
rect 12541 20553 12575 20587
rect 12575 20553 12584 20587
rect 13544 20587 13596 20596
rect 12532 20544 12584 20553
rect 13544 20553 13553 20587
rect 13553 20553 13587 20587
rect 13587 20553 13596 20587
rect 13544 20544 13596 20553
rect 13360 20476 13412 20528
rect 13820 20544 13872 20596
rect 14280 20544 14332 20596
rect 15108 20544 15160 20596
rect 14464 20519 14516 20528
rect 14464 20485 14473 20519
rect 14473 20485 14507 20519
rect 14507 20485 14516 20519
rect 14464 20476 14516 20485
rect 5172 20408 5224 20460
rect 3148 20340 3200 20392
rect 3332 20340 3384 20392
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 6828 20340 6880 20392
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 15936 20544 15988 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 15200 20519 15252 20528
rect 15200 20485 15209 20519
rect 15209 20485 15243 20519
rect 15243 20485 15252 20519
rect 15200 20476 15252 20485
rect 15292 20519 15344 20528
rect 15292 20485 15301 20519
rect 15301 20485 15335 20519
rect 15335 20485 15344 20519
rect 15292 20476 15344 20485
rect 16856 20544 16908 20596
rect 18788 20544 18840 20596
rect 14372 20408 14424 20417
rect 14740 20340 14792 20392
rect 15936 20408 15988 20460
rect 5632 20204 5684 20256
rect 6828 20204 6880 20256
rect 7288 20247 7340 20256
rect 7288 20213 7297 20247
rect 7297 20213 7331 20247
rect 7331 20213 7340 20247
rect 7288 20204 7340 20213
rect 7932 20204 7984 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 10232 20247 10284 20256
rect 10232 20213 10241 20247
rect 10241 20213 10275 20247
rect 10275 20213 10284 20247
rect 10232 20204 10284 20213
rect 10968 20204 11020 20256
rect 13912 20204 13964 20256
rect 14372 20272 14424 20324
rect 15476 20272 15528 20324
rect 15752 20340 15804 20392
rect 16120 20408 16172 20460
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 16488 20451 16540 20460
rect 16488 20417 16523 20451
rect 16523 20417 16540 20451
rect 16488 20408 16540 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 16948 20408 17000 20460
rect 17408 20408 17460 20460
rect 19064 20544 19116 20596
rect 19156 20544 19208 20596
rect 19892 20544 19944 20596
rect 20628 20544 20680 20596
rect 15660 20272 15712 20324
rect 16672 20272 16724 20324
rect 14188 20204 14240 20256
rect 14740 20204 14792 20256
rect 16304 20204 16356 20256
rect 17684 20340 17736 20392
rect 17776 20340 17828 20392
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 18328 20408 18380 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18972 20408 19024 20460
rect 19708 20476 19760 20528
rect 20168 20451 20220 20460
rect 20168 20417 20183 20451
rect 20183 20417 20217 20451
rect 20217 20417 20220 20451
rect 21456 20476 21508 20528
rect 20168 20408 20220 20417
rect 20444 20408 20496 20460
rect 21732 20408 21784 20460
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 23112 20544 23164 20596
rect 23388 20544 23440 20596
rect 23940 20587 23992 20596
rect 23940 20553 23949 20587
rect 23949 20553 23983 20587
rect 23983 20553 23992 20587
rect 23940 20544 23992 20553
rect 24768 20544 24820 20596
rect 25596 20587 25648 20596
rect 25596 20553 25605 20587
rect 25605 20553 25639 20587
rect 25639 20553 25648 20587
rect 25596 20544 25648 20553
rect 25688 20544 25740 20596
rect 23020 20476 23072 20528
rect 19340 20340 19392 20392
rect 19524 20340 19576 20392
rect 19156 20272 19208 20324
rect 19984 20340 20036 20392
rect 20536 20340 20588 20392
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 20812 20383 20864 20392
rect 20812 20349 20821 20383
rect 20821 20349 20855 20383
rect 20855 20349 20864 20383
rect 20812 20340 20864 20349
rect 22192 20408 22244 20460
rect 18144 20204 18196 20256
rect 18604 20204 18656 20256
rect 19064 20204 19116 20256
rect 20076 20272 20128 20324
rect 21272 20272 21324 20324
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20628 20204 20680 20256
rect 20904 20204 20956 20256
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 21916 20272 21968 20324
rect 22192 20272 22244 20324
rect 22836 20340 22888 20392
rect 24584 20408 24636 20460
rect 27344 20544 27396 20596
rect 27620 20544 27672 20596
rect 28264 20544 28316 20596
rect 28356 20544 28408 20596
rect 29092 20544 29144 20596
rect 29368 20544 29420 20596
rect 27896 20476 27948 20528
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 28172 20476 28224 20528
rect 28724 20476 28776 20528
rect 30380 20476 30432 20528
rect 30564 20476 30616 20528
rect 32036 20587 32088 20596
rect 32036 20553 32045 20587
rect 32045 20553 32079 20587
rect 32079 20553 32088 20587
rect 32036 20544 32088 20553
rect 33232 20544 33284 20596
rect 33416 20587 33468 20596
rect 33416 20553 33425 20587
rect 33425 20553 33459 20587
rect 33459 20553 33468 20587
rect 33416 20544 33468 20553
rect 32956 20519 33008 20528
rect 32956 20485 32965 20519
rect 32965 20485 32999 20519
rect 32999 20485 33008 20519
rect 32956 20476 33008 20485
rect 24216 20272 24268 20324
rect 26240 20340 26292 20392
rect 27620 20340 27672 20392
rect 27988 20340 28040 20392
rect 28172 20383 28224 20392
rect 28172 20349 28181 20383
rect 28181 20349 28215 20383
rect 28215 20349 28224 20383
rect 28172 20340 28224 20349
rect 24400 20204 24452 20256
rect 25872 20272 25924 20324
rect 29000 20340 29052 20392
rect 29184 20340 29236 20392
rect 25044 20204 25096 20256
rect 25320 20247 25372 20256
rect 25320 20213 25329 20247
rect 25329 20213 25363 20247
rect 25363 20213 25372 20247
rect 25320 20204 25372 20213
rect 28080 20247 28132 20256
rect 28080 20213 28089 20247
rect 28089 20213 28123 20247
rect 28123 20213 28132 20247
rect 28080 20204 28132 20213
rect 28264 20204 28316 20256
rect 30288 20340 30340 20392
rect 30472 20272 30524 20324
rect 30564 20272 30616 20324
rect 31116 20408 31168 20460
rect 31668 20451 31720 20460
rect 31668 20417 31677 20451
rect 31677 20417 31711 20451
rect 31711 20417 31720 20451
rect 31668 20408 31720 20417
rect 31852 20451 31904 20460
rect 31852 20417 31861 20451
rect 31861 20417 31895 20451
rect 31895 20417 31904 20451
rect 31852 20408 31904 20417
rect 31024 20340 31076 20392
rect 31392 20272 31444 20324
rect 32312 20315 32364 20324
rect 32312 20281 32321 20315
rect 32321 20281 32355 20315
rect 32355 20281 32364 20315
rect 32312 20272 32364 20281
rect 33416 20408 33468 20460
rect 34060 20587 34112 20596
rect 34060 20553 34069 20587
rect 34069 20553 34103 20587
rect 34103 20553 34112 20587
rect 34060 20544 34112 20553
rect 34520 20544 34572 20596
rect 35164 20544 35216 20596
rect 35900 20544 35952 20596
rect 36452 20544 36504 20596
rect 37280 20544 37332 20596
rect 37740 20544 37792 20596
rect 33968 20476 34020 20528
rect 34980 20519 35032 20528
rect 34980 20485 34989 20519
rect 34989 20485 35023 20519
rect 35023 20485 35032 20519
rect 34980 20476 35032 20485
rect 36820 20476 36872 20528
rect 38568 20544 38620 20596
rect 39672 20544 39724 20596
rect 39764 20544 39816 20596
rect 37924 20476 37976 20528
rect 38108 20476 38160 20528
rect 40040 20476 40092 20528
rect 40776 20544 40828 20596
rect 42340 20544 42392 20596
rect 42064 20476 42116 20528
rect 43444 20519 43496 20528
rect 43444 20485 43453 20519
rect 43453 20485 43487 20519
rect 43487 20485 43496 20519
rect 43444 20476 43496 20485
rect 36912 20408 36964 20460
rect 41420 20408 41472 20460
rect 33140 20383 33192 20392
rect 33140 20349 33149 20383
rect 33149 20349 33183 20383
rect 33183 20349 33192 20383
rect 33140 20340 33192 20349
rect 33324 20340 33376 20392
rect 34244 20383 34296 20392
rect 34244 20349 34253 20383
rect 34253 20349 34287 20383
rect 34287 20349 34296 20383
rect 34244 20340 34296 20349
rect 34612 20340 34664 20392
rect 35072 20383 35124 20392
rect 35072 20349 35081 20383
rect 35081 20349 35115 20383
rect 35115 20349 35124 20383
rect 35072 20340 35124 20349
rect 35716 20340 35768 20392
rect 34704 20272 34756 20324
rect 37188 20383 37240 20392
rect 37188 20349 37197 20383
rect 37197 20349 37231 20383
rect 37231 20349 37240 20383
rect 37188 20340 37240 20349
rect 37372 20340 37424 20392
rect 38384 20340 38436 20392
rect 39212 20340 39264 20392
rect 41788 20340 41840 20392
rect 42340 20383 42392 20392
rect 42340 20349 42349 20383
rect 42349 20349 42383 20383
rect 42383 20349 42392 20383
rect 42340 20340 42392 20349
rect 30840 20204 30892 20256
rect 35624 20247 35676 20256
rect 35624 20213 35633 20247
rect 35633 20213 35667 20247
rect 35667 20213 35676 20247
rect 39396 20272 39448 20324
rect 35624 20204 35676 20213
rect 38936 20204 38988 20256
rect 41696 20204 41748 20256
rect 42616 20247 42668 20256
rect 42616 20213 42625 20247
rect 42625 20213 42659 20247
rect 42659 20213 42668 20247
rect 42616 20204 42668 20213
rect 43812 20315 43864 20324
rect 43812 20281 43821 20315
rect 43821 20281 43855 20315
rect 43855 20281 43864 20315
rect 43812 20272 43864 20281
rect 44180 20204 44232 20256
rect 44272 20247 44324 20256
rect 44272 20213 44281 20247
rect 44281 20213 44315 20247
rect 44315 20213 44324 20247
rect 44272 20204 44324 20213
rect 3570 20102 3622 20154
rect 3634 20102 3686 20154
rect 3698 20102 3750 20154
rect 3762 20102 3814 20154
rect 3826 20102 3878 20154
rect 8570 20102 8622 20154
rect 8634 20102 8686 20154
rect 8698 20102 8750 20154
rect 8762 20102 8814 20154
rect 8826 20102 8878 20154
rect 13570 20102 13622 20154
rect 13634 20102 13686 20154
rect 13698 20102 13750 20154
rect 13762 20102 13814 20154
rect 13826 20102 13878 20154
rect 18570 20102 18622 20154
rect 18634 20102 18686 20154
rect 18698 20102 18750 20154
rect 18762 20102 18814 20154
rect 18826 20102 18878 20154
rect 23570 20102 23622 20154
rect 23634 20102 23686 20154
rect 23698 20102 23750 20154
rect 23762 20102 23814 20154
rect 23826 20102 23878 20154
rect 28570 20102 28622 20154
rect 28634 20102 28686 20154
rect 28698 20102 28750 20154
rect 28762 20102 28814 20154
rect 28826 20102 28878 20154
rect 33570 20102 33622 20154
rect 33634 20102 33686 20154
rect 33698 20102 33750 20154
rect 33762 20102 33814 20154
rect 33826 20102 33878 20154
rect 38570 20102 38622 20154
rect 38634 20102 38686 20154
rect 38698 20102 38750 20154
rect 38762 20102 38814 20154
rect 38826 20102 38878 20154
rect 43570 20102 43622 20154
rect 43634 20102 43686 20154
rect 43698 20102 43750 20154
rect 43762 20102 43814 20154
rect 43826 20102 43878 20154
rect 3332 20000 3384 20052
rect 5172 20000 5224 20052
rect 6828 20000 6880 20052
rect 8576 20000 8628 20052
rect 10140 20000 10192 20052
rect 11428 20000 11480 20052
rect 12348 20000 12400 20052
rect 12532 19975 12584 19984
rect 12532 19941 12541 19975
rect 12541 19941 12575 19975
rect 12575 19941 12584 19975
rect 12532 19932 12584 19941
rect 18052 20000 18104 20052
rect 18420 20000 18472 20052
rect 19064 20000 19116 20052
rect 21272 20000 21324 20052
rect 21456 20000 21508 20052
rect 21640 20000 21692 20052
rect 22008 20000 22060 20052
rect 22560 20000 22612 20052
rect 3976 19864 4028 19916
rect 5632 19864 5684 19916
rect 9588 19864 9640 19916
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 7288 19771 7340 19780
rect 3424 19660 3476 19712
rect 5908 19660 5960 19712
rect 7288 19737 7297 19771
rect 7297 19737 7331 19771
rect 7331 19737 7340 19771
rect 7288 19728 7340 19737
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 10968 19796 11020 19848
rect 9864 19728 9916 19780
rect 10232 19728 10284 19780
rect 11428 19864 11480 19916
rect 13360 19864 13412 19916
rect 20536 19932 20588 19984
rect 12164 19796 12216 19848
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 14464 19728 14516 19780
rect 6736 19660 6788 19712
rect 8392 19660 8444 19712
rect 9220 19660 9272 19712
rect 10876 19660 10928 19712
rect 11612 19660 11664 19712
rect 13912 19660 13964 19712
rect 14372 19703 14424 19712
rect 14372 19669 14381 19703
rect 14381 19669 14415 19703
rect 14415 19669 14424 19703
rect 14372 19660 14424 19669
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 16028 19864 16080 19916
rect 16580 19864 16632 19916
rect 17592 19864 17644 19916
rect 18328 19864 18380 19916
rect 15384 19796 15436 19848
rect 15844 19728 15896 19780
rect 15476 19660 15528 19712
rect 15936 19660 15988 19712
rect 16948 19796 17000 19848
rect 17132 19796 17184 19848
rect 16764 19660 16816 19712
rect 17776 19796 17828 19848
rect 18696 19864 18748 19916
rect 19524 19864 19576 19916
rect 20628 19907 20680 19916
rect 18052 19786 18104 19838
rect 18328 19728 18380 19780
rect 19432 19796 19484 19848
rect 19800 19796 19852 19848
rect 20628 19873 20637 19907
rect 20637 19873 20671 19907
rect 20671 19873 20680 19907
rect 20628 19864 20680 19873
rect 20996 19864 21048 19916
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 18972 19728 19024 19780
rect 19064 19728 19116 19780
rect 18144 19660 18196 19712
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 20076 19771 20128 19780
rect 20076 19737 20085 19771
rect 20085 19737 20119 19771
rect 20119 19737 20128 19771
rect 20076 19728 20128 19737
rect 20168 19728 20220 19780
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 21916 19932 21968 19984
rect 27528 20000 27580 20052
rect 24124 19932 24176 19984
rect 27620 19932 27672 19984
rect 22284 19864 22336 19916
rect 24308 19907 24360 19916
rect 24308 19873 24317 19907
rect 24317 19873 24351 19907
rect 24351 19873 24360 19907
rect 24308 19864 24360 19873
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 25964 19907 26016 19916
rect 25964 19873 25973 19907
rect 25973 19873 26007 19907
rect 26007 19873 26016 19907
rect 26240 19907 26292 19916
rect 25964 19864 26016 19873
rect 26240 19873 26249 19907
rect 26249 19873 26283 19907
rect 26283 19873 26292 19907
rect 26240 19864 26292 19873
rect 28172 19864 28224 19916
rect 30656 19975 30708 19984
rect 30656 19941 30665 19975
rect 30665 19941 30699 19975
rect 30699 19941 30708 19975
rect 30656 19932 30708 19941
rect 23296 19796 23348 19848
rect 27896 19796 27948 19848
rect 27988 19796 28040 19848
rect 20260 19660 20312 19712
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 20628 19660 20680 19712
rect 20812 19660 20864 19712
rect 22192 19728 22244 19780
rect 23480 19728 23532 19780
rect 23940 19728 23992 19780
rect 22008 19703 22060 19712
rect 22008 19669 22017 19703
rect 22017 19669 22051 19703
rect 22051 19669 22060 19703
rect 22008 19660 22060 19669
rect 22376 19703 22428 19712
rect 22376 19669 22385 19703
rect 22385 19669 22419 19703
rect 22419 19669 22428 19703
rect 22376 19660 22428 19669
rect 24032 19660 24084 19712
rect 24860 19703 24912 19712
rect 24860 19669 24869 19703
rect 24869 19669 24903 19703
rect 24903 19669 24912 19703
rect 24860 19660 24912 19669
rect 26516 19771 26568 19780
rect 26516 19737 26525 19771
rect 26525 19737 26559 19771
rect 26559 19737 26568 19771
rect 26516 19728 26568 19737
rect 28172 19728 28224 19780
rect 28264 19771 28316 19780
rect 28264 19737 28273 19771
rect 28273 19737 28307 19771
rect 28307 19737 28316 19771
rect 28264 19728 28316 19737
rect 27804 19660 27856 19712
rect 28080 19660 28132 19712
rect 30288 19796 30340 19848
rect 30748 19839 30800 19848
rect 30748 19805 30777 19839
rect 30777 19805 30800 19839
rect 31852 19864 31904 19916
rect 33140 20000 33192 20052
rect 30748 19796 30800 19805
rect 31116 19839 31168 19848
rect 31116 19805 31125 19839
rect 31125 19805 31159 19839
rect 31159 19805 31168 19839
rect 31116 19796 31168 19805
rect 35992 20000 36044 20052
rect 37648 20000 37700 20052
rect 33508 19864 33560 19916
rect 35072 19864 35124 19916
rect 37188 19907 37240 19916
rect 37188 19873 37197 19907
rect 37197 19873 37231 19907
rect 37231 19873 37240 19907
rect 37188 19864 37240 19873
rect 28540 19660 28592 19712
rect 28908 19660 28960 19712
rect 29828 19660 29880 19712
rect 30012 19660 30064 19712
rect 30748 19660 30800 19712
rect 32772 19728 32824 19780
rect 33324 19728 33376 19780
rect 34152 19771 34204 19780
rect 34152 19737 34161 19771
rect 34161 19737 34195 19771
rect 34195 19737 34204 19771
rect 34152 19728 34204 19737
rect 34888 19839 34940 19848
rect 34888 19805 34897 19839
rect 34897 19805 34931 19839
rect 34931 19805 34940 19839
rect 34888 19796 34940 19805
rect 35808 19796 35860 19848
rect 37280 19796 37332 19848
rect 38476 19932 38528 19984
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 41696 20000 41748 20052
rect 44180 20000 44232 20052
rect 44916 20043 44968 20052
rect 44916 20009 44925 20043
rect 44925 20009 44959 20043
rect 44959 20009 44968 20043
rect 44916 20000 44968 20009
rect 39396 19975 39448 19984
rect 39396 19941 39405 19975
rect 39405 19941 39439 19975
rect 39439 19941 39448 19975
rect 39396 19932 39448 19941
rect 39856 19864 39908 19916
rect 38752 19839 38804 19848
rect 38752 19805 38761 19839
rect 38761 19805 38795 19839
rect 38795 19805 38804 19839
rect 38752 19796 38804 19805
rect 41420 19864 41472 19916
rect 42616 19864 42668 19916
rect 39212 19728 39264 19780
rect 42064 19796 42116 19848
rect 31484 19703 31536 19712
rect 31484 19669 31493 19703
rect 31493 19669 31527 19703
rect 31527 19669 31536 19703
rect 31484 19660 31536 19669
rect 31944 19703 31996 19712
rect 31944 19669 31953 19703
rect 31953 19669 31987 19703
rect 31987 19669 31996 19703
rect 31944 19660 31996 19669
rect 32496 19703 32548 19712
rect 32496 19669 32505 19703
rect 32505 19669 32539 19703
rect 32539 19669 32548 19703
rect 32496 19660 32548 19669
rect 33140 19703 33192 19712
rect 33140 19669 33149 19703
rect 33149 19669 33183 19703
rect 33183 19669 33192 19703
rect 33140 19660 33192 19669
rect 34428 19660 34480 19712
rect 34704 19703 34756 19712
rect 34704 19669 34713 19703
rect 34713 19669 34747 19703
rect 34747 19669 34756 19703
rect 34704 19660 34756 19669
rect 35164 19703 35216 19712
rect 35164 19669 35173 19703
rect 35173 19669 35207 19703
rect 35207 19669 35216 19703
rect 35164 19660 35216 19669
rect 35808 19660 35860 19712
rect 37280 19660 37332 19712
rect 37924 19703 37976 19712
rect 37924 19669 37933 19703
rect 37933 19669 37967 19703
rect 37967 19669 37976 19703
rect 37924 19660 37976 19669
rect 38292 19703 38344 19712
rect 38292 19669 38301 19703
rect 38301 19669 38335 19703
rect 38335 19669 38344 19703
rect 38292 19660 38344 19669
rect 39580 19703 39632 19712
rect 39580 19669 39589 19703
rect 39589 19669 39623 19703
rect 39623 19669 39632 19703
rect 39580 19660 39632 19669
rect 39948 19703 40000 19712
rect 39948 19669 39957 19703
rect 39957 19669 39991 19703
rect 39991 19669 40000 19703
rect 39948 19660 40000 19669
rect 40776 19728 40828 19780
rect 42800 19728 42852 19780
rect 40868 19660 40920 19712
rect 42156 19703 42208 19712
rect 42156 19669 42165 19703
rect 42165 19669 42199 19703
rect 42199 19669 42208 19703
rect 42156 19660 42208 19669
rect 43996 19703 44048 19712
rect 43996 19669 44005 19703
rect 44005 19669 44039 19703
rect 44039 19669 44048 19703
rect 43996 19660 44048 19669
rect 6070 19558 6122 19610
rect 6134 19558 6186 19610
rect 6198 19558 6250 19610
rect 6262 19558 6314 19610
rect 6326 19558 6378 19610
rect 11070 19558 11122 19610
rect 11134 19558 11186 19610
rect 11198 19558 11250 19610
rect 11262 19558 11314 19610
rect 11326 19558 11378 19610
rect 16070 19558 16122 19610
rect 16134 19558 16186 19610
rect 16198 19558 16250 19610
rect 16262 19558 16314 19610
rect 16326 19558 16378 19610
rect 21070 19558 21122 19610
rect 21134 19558 21186 19610
rect 21198 19558 21250 19610
rect 21262 19558 21314 19610
rect 21326 19558 21378 19610
rect 26070 19558 26122 19610
rect 26134 19558 26186 19610
rect 26198 19558 26250 19610
rect 26262 19558 26314 19610
rect 26326 19558 26378 19610
rect 31070 19558 31122 19610
rect 31134 19558 31186 19610
rect 31198 19558 31250 19610
rect 31262 19558 31314 19610
rect 31326 19558 31378 19610
rect 36070 19558 36122 19610
rect 36134 19558 36186 19610
rect 36198 19558 36250 19610
rect 36262 19558 36314 19610
rect 36326 19558 36378 19610
rect 41070 19558 41122 19610
rect 41134 19558 41186 19610
rect 41198 19558 41250 19610
rect 41262 19558 41314 19610
rect 41326 19558 41378 19610
rect 8300 19456 8352 19508
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 9220 19456 9272 19508
rect 9588 19456 9640 19508
rect 5540 19388 5592 19440
rect 8208 19388 8260 19440
rect 5632 19320 5684 19372
rect 6000 19159 6052 19168
rect 6000 19125 6009 19159
rect 6009 19125 6043 19159
rect 6043 19125 6052 19159
rect 6828 19320 6880 19372
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 10140 19388 10192 19440
rect 10968 19456 11020 19508
rect 10876 19388 10928 19440
rect 12164 19456 12216 19508
rect 8116 19320 8168 19329
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 9864 19320 9916 19372
rect 14740 19456 14792 19508
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 13912 19388 13964 19440
rect 15016 19388 15068 19440
rect 15936 19456 15988 19508
rect 6736 19295 6788 19304
rect 6736 19261 6745 19295
rect 6745 19261 6779 19295
rect 6779 19261 6788 19295
rect 6736 19252 6788 19261
rect 6644 19184 6696 19236
rect 8392 19252 8444 19304
rect 15568 19320 15620 19372
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 16580 19456 16632 19508
rect 17408 19456 17460 19508
rect 16764 19388 16816 19440
rect 17040 19388 17092 19440
rect 17592 19388 17644 19440
rect 17684 19388 17736 19440
rect 18236 19456 18288 19508
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 19524 19456 19576 19508
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17500 19363 17552 19372
rect 17500 19329 17509 19363
rect 17509 19329 17543 19363
rect 17543 19329 17552 19363
rect 18696 19388 18748 19440
rect 17500 19320 17552 19329
rect 10692 19252 10744 19304
rect 10784 19252 10836 19304
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 6000 19116 6052 19125
rect 10416 19116 10468 19168
rect 11612 19116 11664 19168
rect 14832 19116 14884 19168
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15384 19252 15436 19304
rect 16212 19252 16264 19304
rect 17224 19252 17276 19304
rect 17684 19295 17736 19304
rect 17684 19261 17693 19295
rect 17693 19261 17727 19295
rect 17727 19261 17736 19295
rect 17684 19252 17736 19261
rect 18972 19320 19024 19372
rect 20168 19456 20220 19508
rect 20720 19456 20772 19508
rect 20812 19456 20864 19508
rect 23296 19456 23348 19508
rect 24860 19456 24912 19508
rect 26240 19456 26292 19508
rect 26516 19456 26568 19508
rect 28356 19456 28408 19508
rect 29920 19456 29972 19508
rect 15292 19184 15344 19236
rect 15752 19116 15804 19168
rect 16672 19116 16724 19168
rect 17960 19184 18012 19236
rect 19432 19252 19484 19304
rect 21732 19388 21784 19440
rect 19708 19320 19760 19372
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 17316 19116 17368 19168
rect 17776 19116 17828 19168
rect 18328 19116 18380 19168
rect 19892 19184 19944 19236
rect 21456 19363 21508 19372
rect 21456 19329 21481 19363
rect 21481 19329 21508 19363
rect 21456 19320 21508 19329
rect 22284 19320 22336 19372
rect 20536 19252 20588 19304
rect 20904 19252 20956 19304
rect 22836 19295 22888 19304
rect 20628 19159 20680 19168
rect 20628 19125 20637 19159
rect 20637 19125 20671 19159
rect 20671 19125 20680 19159
rect 20628 19116 20680 19125
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 21548 19116 21600 19168
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 21916 19116 21968 19125
rect 22836 19261 22845 19295
rect 22845 19261 22879 19295
rect 22879 19261 22888 19295
rect 22836 19252 22888 19261
rect 23112 19295 23164 19304
rect 23112 19261 23121 19295
rect 23121 19261 23155 19295
rect 23155 19261 23164 19295
rect 23112 19252 23164 19261
rect 22468 19116 22520 19168
rect 24400 19252 24452 19304
rect 25136 19184 25188 19236
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 26332 19320 26384 19372
rect 28172 19388 28224 19440
rect 27436 19320 27488 19372
rect 27620 19363 27672 19372
rect 27620 19329 27629 19363
rect 27629 19329 27663 19363
rect 27663 19329 27672 19363
rect 27620 19320 27672 19329
rect 28080 19363 28132 19372
rect 28080 19329 28089 19363
rect 28089 19329 28123 19363
rect 28123 19329 28132 19363
rect 28080 19320 28132 19329
rect 28540 19320 28592 19372
rect 28908 19320 28960 19372
rect 29644 19431 29696 19440
rect 29644 19397 29653 19431
rect 29653 19397 29687 19431
rect 29687 19397 29696 19431
rect 29644 19388 29696 19397
rect 29552 19363 29604 19372
rect 29552 19329 29561 19363
rect 29561 19329 29595 19363
rect 29595 19329 29604 19363
rect 29552 19320 29604 19329
rect 29736 19363 29788 19372
rect 29736 19329 29745 19363
rect 29745 19329 29779 19363
rect 29779 19329 29788 19363
rect 29736 19320 29788 19329
rect 30012 19363 30064 19372
rect 30012 19329 30021 19363
rect 30021 19329 30055 19363
rect 30055 19329 30064 19363
rect 30012 19320 30064 19329
rect 29460 19252 29512 19304
rect 30196 19431 30248 19440
rect 30196 19397 30205 19431
rect 30205 19397 30239 19431
rect 30239 19397 30248 19431
rect 30196 19388 30248 19397
rect 30840 19456 30892 19508
rect 31668 19499 31720 19508
rect 31668 19465 31677 19499
rect 31677 19465 31711 19499
rect 31711 19465 31720 19499
rect 31668 19456 31720 19465
rect 31852 19456 31904 19508
rect 32956 19456 33008 19508
rect 33416 19456 33468 19508
rect 32220 19388 32272 19440
rect 31300 19320 31352 19372
rect 31392 19320 31444 19372
rect 33232 19320 33284 19372
rect 34888 19456 34940 19508
rect 35716 19456 35768 19508
rect 34612 19388 34664 19440
rect 30840 19252 30892 19304
rect 31116 19295 31168 19304
rect 31116 19261 31125 19295
rect 31125 19261 31159 19295
rect 31159 19261 31168 19295
rect 31116 19252 31168 19261
rect 31576 19184 31628 19236
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 26424 19116 26476 19168
rect 26608 19159 26660 19168
rect 26608 19125 26617 19159
rect 26617 19125 26651 19159
rect 26651 19125 26660 19159
rect 26608 19116 26660 19125
rect 27160 19116 27212 19168
rect 28264 19116 28316 19168
rect 29644 19116 29696 19168
rect 30564 19159 30616 19168
rect 30564 19125 30573 19159
rect 30573 19125 30607 19159
rect 30607 19125 30616 19159
rect 30564 19116 30616 19125
rect 31300 19116 31352 19168
rect 31852 19295 31904 19304
rect 31852 19261 31861 19295
rect 31861 19261 31895 19295
rect 31895 19261 31904 19295
rect 31852 19252 31904 19261
rect 33140 19184 33192 19236
rect 34060 19295 34112 19304
rect 34060 19261 34069 19295
rect 34069 19261 34103 19295
rect 34103 19261 34112 19295
rect 34060 19252 34112 19261
rect 34520 19252 34572 19304
rect 34244 19184 34296 19236
rect 35532 19252 35584 19304
rect 35808 19295 35860 19304
rect 35808 19261 35817 19295
rect 35817 19261 35851 19295
rect 35851 19261 35860 19295
rect 35808 19252 35860 19261
rect 37280 19456 37332 19508
rect 38292 19456 38344 19508
rect 39580 19456 39632 19508
rect 38108 19388 38160 19440
rect 35992 19320 36044 19372
rect 37280 19295 37332 19304
rect 36084 19184 36136 19236
rect 37280 19261 37289 19295
rect 37289 19261 37323 19295
rect 37323 19261 37332 19295
rect 37280 19252 37332 19261
rect 38016 19252 38068 19304
rect 38108 19252 38160 19304
rect 39764 19388 39816 19440
rect 40868 19456 40920 19508
rect 41696 19456 41748 19508
rect 41788 19499 41840 19508
rect 41788 19465 41797 19499
rect 41797 19465 41831 19499
rect 41831 19465 41840 19499
rect 41788 19456 41840 19465
rect 42156 19499 42208 19508
rect 42156 19465 42165 19499
rect 42165 19465 42199 19499
rect 42199 19465 42208 19499
rect 42156 19456 42208 19465
rect 43996 19456 44048 19508
rect 41512 19363 41564 19372
rect 41512 19329 41521 19363
rect 41521 19329 41555 19363
rect 41555 19329 41564 19363
rect 41512 19320 41564 19329
rect 39212 19295 39264 19304
rect 39212 19261 39228 19295
rect 39228 19261 39262 19295
rect 39262 19261 39264 19295
rect 39212 19252 39264 19261
rect 41604 19252 41656 19304
rect 42340 19295 42392 19304
rect 42340 19261 42349 19295
rect 42349 19261 42383 19295
rect 42383 19261 42392 19295
rect 42340 19252 42392 19261
rect 41420 19184 41472 19236
rect 42708 19388 42760 19440
rect 43444 19388 43496 19440
rect 43168 19295 43220 19304
rect 43168 19261 43177 19295
rect 43177 19261 43211 19295
rect 43211 19261 43220 19295
rect 43168 19252 43220 19261
rect 44732 19295 44784 19304
rect 44732 19261 44741 19295
rect 44741 19261 44775 19295
rect 44775 19261 44784 19295
rect 44732 19252 44784 19261
rect 42800 19184 42852 19236
rect 32772 19116 32824 19168
rect 35348 19159 35400 19168
rect 35348 19125 35357 19159
rect 35357 19125 35391 19159
rect 35391 19125 35400 19159
rect 35348 19116 35400 19125
rect 35900 19116 35952 19168
rect 36176 19159 36228 19168
rect 36176 19125 36185 19159
rect 36185 19125 36219 19159
rect 36219 19125 36228 19159
rect 36176 19116 36228 19125
rect 36268 19116 36320 19168
rect 36912 19159 36964 19168
rect 36912 19125 36921 19159
rect 36921 19125 36955 19159
rect 36955 19125 36964 19159
rect 36912 19116 36964 19125
rect 37096 19116 37148 19168
rect 39028 19159 39080 19168
rect 39028 19125 39037 19159
rect 39037 19125 39071 19159
rect 39071 19125 39080 19159
rect 39028 19116 39080 19125
rect 3570 19014 3622 19066
rect 3634 19014 3686 19066
rect 3698 19014 3750 19066
rect 3762 19014 3814 19066
rect 3826 19014 3878 19066
rect 8570 19014 8622 19066
rect 8634 19014 8686 19066
rect 8698 19014 8750 19066
rect 8762 19014 8814 19066
rect 8826 19014 8878 19066
rect 13570 19014 13622 19066
rect 13634 19014 13686 19066
rect 13698 19014 13750 19066
rect 13762 19014 13814 19066
rect 13826 19014 13878 19066
rect 18570 19014 18622 19066
rect 18634 19014 18686 19066
rect 18698 19014 18750 19066
rect 18762 19014 18814 19066
rect 18826 19014 18878 19066
rect 23570 19014 23622 19066
rect 23634 19014 23686 19066
rect 23698 19014 23750 19066
rect 23762 19014 23814 19066
rect 23826 19014 23878 19066
rect 28570 19014 28622 19066
rect 28634 19014 28686 19066
rect 28698 19014 28750 19066
rect 28762 19014 28814 19066
rect 28826 19014 28878 19066
rect 33570 19014 33622 19066
rect 33634 19014 33686 19066
rect 33698 19014 33750 19066
rect 33762 19014 33814 19066
rect 33826 19014 33878 19066
rect 38570 19014 38622 19066
rect 38634 19014 38686 19066
rect 38698 19014 38750 19066
rect 38762 19014 38814 19066
rect 38826 19014 38878 19066
rect 43570 19014 43622 19066
rect 43634 19014 43686 19066
rect 43698 19014 43750 19066
rect 43762 19014 43814 19066
rect 43826 19014 43878 19066
rect 6644 18912 6696 18964
rect 6000 18887 6052 18896
rect 6000 18853 6009 18887
rect 6009 18853 6043 18887
rect 6043 18853 6052 18887
rect 6000 18844 6052 18853
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 5448 18708 5500 18760
rect 5632 18708 5684 18760
rect 7104 18912 7156 18964
rect 10232 18912 10284 18964
rect 7012 18844 7064 18896
rect 7748 18844 7800 18896
rect 9128 18776 9180 18828
rect 11428 18912 11480 18964
rect 11888 18912 11940 18964
rect 14556 18912 14608 18964
rect 14740 18912 14792 18964
rect 18236 18887 18288 18896
rect 18236 18853 18245 18887
rect 18245 18853 18279 18887
rect 18279 18853 18288 18887
rect 18236 18844 18288 18853
rect 18420 18912 18472 18964
rect 19340 18912 19392 18964
rect 19432 18912 19484 18964
rect 8392 18708 8444 18760
rect 7840 18640 7892 18692
rect 4896 18615 4948 18624
rect 4896 18581 4905 18615
rect 4905 18581 4939 18615
rect 4939 18581 4948 18615
rect 4896 18572 4948 18581
rect 5540 18572 5592 18624
rect 6552 18572 6604 18624
rect 6920 18572 6972 18624
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 10140 18708 10192 18760
rect 10416 18708 10468 18760
rect 14372 18776 14424 18828
rect 14556 18776 14608 18828
rect 14832 18776 14884 18828
rect 15200 18776 15252 18828
rect 15568 18776 15620 18828
rect 10692 18708 10744 18760
rect 10876 18708 10928 18760
rect 12992 18708 13044 18760
rect 11612 18640 11664 18692
rect 13176 18640 13228 18692
rect 8576 18572 8628 18624
rect 10784 18572 10836 18624
rect 12072 18572 12124 18624
rect 15292 18708 15344 18760
rect 15752 18819 15804 18828
rect 15752 18785 15761 18819
rect 15761 18785 15795 18819
rect 15795 18785 15804 18819
rect 15752 18776 15804 18785
rect 16948 18776 17000 18828
rect 18328 18776 18380 18828
rect 14740 18640 14792 18692
rect 16212 18708 16264 18760
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 17224 18708 17276 18760
rect 17500 18708 17552 18760
rect 17868 18708 17920 18760
rect 18052 18708 18104 18760
rect 18972 18708 19024 18760
rect 20444 18912 20496 18964
rect 20168 18844 20220 18896
rect 23480 18912 23532 18964
rect 24032 18912 24084 18964
rect 25596 18912 25648 18964
rect 26240 18912 26292 18964
rect 27804 18912 27856 18964
rect 28172 18955 28224 18964
rect 28172 18921 28181 18955
rect 28181 18921 28215 18955
rect 28215 18921 28224 18955
rect 28172 18912 28224 18921
rect 28908 18912 28960 18964
rect 21916 18776 21968 18828
rect 24032 18776 24084 18828
rect 24308 18819 24360 18828
rect 24308 18785 24317 18819
rect 24317 18785 24351 18819
rect 24351 18785 24360 18819
rect 24308 18776 24360 18785
rect 27988 18844 28040 18896
rect 29184 18887 29236 18896
rect 29184 18853 29193 18887
rect 29193 18853 29227 18887
rect 29227 18853 29236 18887
rect 31944 18912 31996 18964
rect 29184 18844 29236 18853
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 19892 18640 19944 18692
rect 20168 18683 20220 18692
rect 20168 18649 20177 18683
rect 20177 18649 20211 18683
rect 20211 18649 20220 18683
rect 20168 18640 20220 18649
rect 15016 18572 15068 18624
rect 15660 18615 15712 18624
rect 15660 18581 15669 18615
rect 15669 18581 15703 18615
rect 15703 18581 15712 18615
rect 15660 18572 15712 18581
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 16764 18572 16816 18624
rect 17408 18572 17460 18624
rect 17960 18572 18012 18624
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 24124 18751 24176 18760
rect 24124 18717 24133 18751
rect 24133 18717 24167 18751
rect 24167 18717 24176 18751
rect 24124 18708 24176 18717
rect 24492 18708 24544 18760
rect 25964 18708 26016 18760
rect 30380 18776 30432 18828
rect 31852 18844 31904 18896
rect 32036 18844 32088 18896
rect 30840 18776 30892 18828
rect 31760 18776 31812 18828
rect 33140 18912 33192 18964
rect 36176 18912 36228 18964
rect 38476 18912 38528 18964
rect 39948 18912 40000 18964
rect 40960 18955 41012 18964
rect 40960 18921 40969 18955
rect 40969 18921 41003 18955
rect 41003 18921 41012 18955
rect 40960 18912 41012 18921
rect 41512 18912 41564 18964
rect 41604 18912 41656 18964
rect 33416 18819 33468 18828
rect 33416 18785 33425 18819
rect 33425 18785 33459 18819
rect 33459 18785 33468 18819
rect 33416 18776 33468 18785
rect 33508 18819 33560 18828
rect 33508 18785 33517 18819
rect 33517 18785 33551 18819
rect 33551 18785 33560 18819
rect 33508 18776 33560 18785
rect 26424 18751 26476 18760
rect 26424 18717 26433 18751
rect 26433 18717 26467 18751
rect 26467 18717 26476 18751
rect 26424 18708 26476 18717
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28448 18751 28500 18760
rect 28448 18717 28457 18751
rect 28457 18717 28491 18751
rect 28491 18717 28500 18751
rect 28448 18708 28500 18717
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 29920 18751 29972 18760
rect 29920 18717 29929 18751
rect 29929 18717 29963 18751
rect 29963 18717 29972 18751
rect 29920 18708 29972 18717
rect 32404 18708 32456 18760
rect 22468 18640 22520 18692
rect 21548 18572 21600 18624
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 23204 18615 23256 18624
rect 23204 18581 23213 18615
rect 23213 18581 23247 18615
rect 23247 18581 23256 18615
rect 23204 18572 23256 18581
rect 24308 18572 24360 18624
rect 24860 18683 24912 18692
rect 24860 18649 24869 18683
rect 24869 18649 24903 18683
rect 24903 18649 24912 18683
rect 24860 18640 24912 18649
rect 26792 18640 26844 18692
rect 27160 18640 27212 18692
rect 30748 18683 30800 18692
rect 30748 18649 30757 18683
rect 30757 18649 30791 18683
rect 30791 18649 30800 18683
rect 30748 18640 30800 18649
rect 32496 18640 32548 18692
rect 32864 18708 32916 18760
rect 34704 18819 34756 18828
rect 34704 18785 34713 18819
rect 34713 18785 34747 18819
rect 34747 18785 34756 18819
rect 34704 18776 34756 18785
rect 37004 18776 37056 18828
rect 37280 18776 37332 18828
rect 37556 18776 37608 18828
rect 38384 18776 38436 18828
rect 39028 18776 39080 18828
rect 39212 18819 39264 18828
rect 39212 18785 39221 18819
rect 39221 18785 39255 18819
rect 39255 18785 39264 18819
rect 39212 18776 39264 18785
rect 40960 18776 41012 18828
rect 25136 18572 25188 18624
rect 26332 18615 26384 18624
rect 26332 18581 26341 18615
rect 26341 18581 26375 18615
rect 26375 18581 26384 18615
rect 26332 18572 26384 18581
rect 28356 18572 28408 18624
rect 31116 18572 31168 18624
rect 32128 18572 32180 18624
rect 32312 18615 32364 18624
rect 32312 18581 32321 18615
rect 32321 18581 32355 18615
rect 32355 18581 32364 18615
rect 32312 18572 32364 18581
rect 34152 18640 34204 18692
rect 36268 18751 36320 18760
rect 36268 18717 36277 18751
rect 36277 18717 36311 18751
rect 36311 18717 36320 18751
rect 36268 18708 36320 18717
rect 37924 18708 37976 18760
rect 38476 18751 38528 18760
rect 38476 18717 38485 18751
rect 38485 18717 38519 18751
rect 38519 18717 38528 18751
rect 38476 18708 38528 18717
rect 34060 18572 34112 18624
rect 34244 18615 34296 18624
rect 34244 18581 34253 18615
rect 34253 18581 34287 18615
rect 34287 18581 34296 18615
rect 34244 18572 34296 18581
rect 34612 18572 34664 18624
rect 34888 18572 34940 18624
rect 37004 18640 37056 18692
rect 38108 18640 38160 18692
rect 41420 18751 41472 18760
rect 41420 18717 41429 18751
rect 41429 18717 41463 18751
rect 41463 18717 41472 18751
rect 41420 18708 41472 18717
rect 41512 18751 41564 18760
rect 41512 18717 41521 18751
rect 41521 18717 41555 18751
rect 41555 18717 41564 18751
rect 42156 18776 42208 18828
rect 41512 18708 41564 18717
rect 36084 18572 36136 18624
rect 36452 18572 36504 18624
rect 36820 18572 36872 18624
rect 39488 18683 39540 18692
rect 39488 18649 39497 18683
rect 39497 18649 39531 18683
rect 39531 18649 39540 18683
rect 39488 18640 39540 18649
rect 39764 18640 39816 18692
rect 41696 18572 41748 18624
rect 42984 18640 43036 18692
rect 42248 18615 42300 18624
rect 42248 18581 42257 18615
rect 42257 18581 42291 18615
rect 42291 18581 42300 18615
rect 42248 18572 42300 18581
rect 42708 18615 42760 18624
rect 42708 18581 42717 18615
rect 42717 18581 42751 18615
rect 42751 18581 42760 18615
rect 42708 18572 42760 18581
rect 43720 18572 43772 18624
rect 43812 18572 43864 18624
rect 44824 18572 44876 18624
rect 6070 18470 6122 18522
rect 6134 18470 6186 18522
rect 6198 18470 6250 18522
rect 6262 18470 6314 18522
rect 6326 18470 6378 18522
rect 11070 18470 11122 18522
rect 11134 18470 11186 18522
rect 11198 18470 11250 18522
rect 11262 18470 11314 18522
rect 11326 18470 11378 18522
rect 16070 18470 16122 18522
rect 16134 18470 16186 18522
rect 16198 18470 16250 18522
rect 16262 18470 16314 18522
rect 16326 18470 16378 18522
rect 21070 18470 21122 18522
rect 21134 18470 21186 18522
rect 21198 18470 21250 18522
rect 21262 18470 21314 18522
rect 21326 18470 21378 18522
rect 26070 18470 26122 18522
rect 26134 18470 26186 18522
rect 26198 18470 26250 18522
rect 26262 18470 26314 18522
rect 26326 18470 26378 18522
rect 31070 18470 31122 18522
rect 31134 18470 31186 18522
rect 31198 18470 31250 18522
rect 31262 18470 31314 18522
rect 31326 18470 31378 18522
rect 36070 18470 36122 18522
rect 36134 18470 36186 18522
rect 36198 18470 36250 18522
rect 36262 18470 36314 18522
rect 36326 18470 36378 18522
rect 41070 18470 41122 18522
rect 41134 18470 41186 18522
rect 41198 18470 41250 18522
rect 41262 18470 41314 18522
rect 41326 18470 41378 18522
rect 4896 18368 4948 18420
rect 5448 18368 5500 18420
rect 4620 18300 4672 18352
rect 3792 18275 3844 18284
rect 3792 18241 3801 18275
rect 3801 18241 3835 18275
rect 3835 18241 3844 18275
rect 3792 18232 3844 18241
rect 5632 18368 5684 18420
rect 7380 18368 7432 18420
rect 7840 18368 7892 18420
rect 8392 18368 8444 18420
rect 11612 18368 11664 18420
rect 12992 18411 13044 18420
rect 12992 18377 13001 18411
rect 13001 18377 13035 18411
rect 13035 18377 13044 18411
rect 12992 18368 13044 18377
rect 8300 18300 8352 18352
rect 10140 18300 10192 18352
rect 5632 18232 5684 18284
rect 5816 18164 5868 18216
rect 6552 18232 6604 18284
rect 8116 18232 8168 18284
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 7104 18164 7156 18216
rect 10784 18164 10836 18216
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 11980 18232 12032 18284
rect 12164 18232 12216 18284
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 13360 18232 13412 18284
rect 15844 18368 15896 18420
rect 11612 18164 11664 18216
rect 5724 18028 5776 18080
rect 6000 18071 6052 18080
rect 6000 18037 6009 18071
rect 6009 18037 6043 18071
rect 6043 18037 6052 18071
rect 6000 18028 6052 18037
rect 7012 18028 7064 18080
rect 8116 18028 8168 18080
rect 9956 18028 10008 18080
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 11520 18028 11572 18080
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 13176 18028 13228 18080
rect 14740 18028 14792 18080
rect 15936 18300 15988 18352
rect 16488 18368 16540 18420
rect 17960 18368 18012 18420
rect 19616 18368 19668 18420
rect 19892 18368 19944 18420
rect 20168 18368 20220 18420
rect 16580 18300 16632 18352
rect 16672 18300 16724 18352
rect 16764 18343 16816 18352
rect 16764 18309 16773 18343
rect 16773 18309 16807 18343
rect 16807 18309 16816 18343
rect 16764 18300 16816 18309
rect 17132 18343 17184 18352
rect 15016 18232 15068 18284
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 15844 18164 15896 18216
rect 16488 18232 16540 18284
rect 17132 18309 17141 18343
rect 17141 18309 17175 18343
rect 17175 18309 17184 18343
rect 17132 18300 17184 18309
rect 17316 18343 17368 18352
rect 17316 18309 17341 18343
rect 17341 18309 17368 18343
rect 17316 18300 17368 18309
rect 17500 18232 17552 18284
rect 17684 18232 17736 18284
rect 19340 18300 19392 18352
rect 20628 18368 20680 18420
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 22560 18368 22612 18420
rect 22744 18368 22796 18420
rect 24768 18368 24820 18420
rect 24860 18368 24912 18420
rect 25688 18368 25740 18420
rect 29184 18368 29236 18420
rect 20996 18300 21048 18352
rect 21548 18300 21600 18352
rect 17960 18275 18012 18284
rect 17960 18241 17969 18275
rect 17969 18241 18003 18275
rect 18003 18241 18012 18275
rect 17960 18232 18012 18241
rect 20260 18232 20312 18284
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 20444 18275 20496 18284
rect 20444 18241 20453 18275
rect 20453 18241 20487 18275
rect 20487 18241 20496 18275
rect 20444 18232 20496 18241
rect 15108 18096 15160 18148
rect 16028 18028 16080 18080
rect 21180 18275 21232 18284
rect 21180 18241 21189 18275
rect 21189 18241 21223 18275
rect 21223 18241 21232 18275
rect 21180 18232 21232 18241
rect 21364 18275 21416 18284
rect 21364 18241 21373 18275
rect 21373 18241 21407 18275
rect 21407 18241 21416 18275
rect 21364 18232 21416 18241
rect 17040 18139 17092 18148
rect 17040 18105 17049 18139
rect 17049 18105 17083 18139
rect 17083 18105 17092 18139
rect 17040 18096 17092 18105
rect 17868 18096 17920 18148
rect 20444 18096 20496 18148
rect 21548 18164 21600 18216
rect 22744 18275 22796 18284
rect 22744 18241 22753 18275
rect 22753 18241 22787 18275
rect 22787 18241 22796 18275
rect 22744 18232 22796 18241
rect 22836 18275 22888 18284
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 24216 18232 24268 18284
rect 24400 18232 24452 18284
rect 24860 18232 24912 18284
rect 24952 18232 25004 18284
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 25596 18232 25648 18284
rect 26976 18232 27028 18284
rect 27528 18300 27580 18352
rect 27620 18300 27672 18352
rect 23112 18164 23164 18216
rect 25964 18096 26016 18148
rect 26976 18139 27028 18148
rect 26976 18105 26985 18139
rect 26985 18105 27019 18139
rect 27019 18105 27028 18139
rect 26976 18096 27028 18105
rect 27896 18232 27948 18284
rect 29276 18300 29328 18352
rect 29644 18300 29696 18352
rect 30196 18368 30248 18420
rect 30748 18368 30800 18420
rect 32312 18368 32364 18420
rect 30840 18300 30892 18352
rect 28908 18164 28960 18216
rect 30012 18164 30064 18216
rect 31484 18232 31536 18284
rect 31668 18275 31720 18284
rect 31668 18241 31677 18275
rect 31677 18241 31711 18275
rect 31711 18241 31720 18275
rect 31668 18232 31720 18241
rect 31760 18275 31812 18284
rect 31760 18241 31769 18275
rect 31769 18241 31803 18275
rect 31803 18241 31812 18275
rect 31760 18232 31812 18241
rect 32128 18300 32180 18352
rect 32496 18300 32548 18352
rect 33416 18368 33468 18420
rect 34520 18411 34572 18420
rect 34520 18377 34529 18411
rect 34529 18377 34563 18411
rect 34563 18377 34572 18411
rect 34520 18368 34572 18377
rect 35808 18368 35860 18420
rect 33232 18300 33284 18352
rect 30932 18164 30984 18216
rect 32036 18164 32088 18216
rect 32312 18207 32364 18216
rect 32312 18173 32321 18207
rect 32321 18173 32355 18207
rect 32355 18173 32364 18207
rect 32312 18164 32364 18173
rect 32680 18164 32732 18216
rect 34244 18300 34296 18352
rect 34888 18300 34940 18352
rect 34520 18164 34572 18216
rect 34980 18207 35032 18216
rect 34980 18173 34989 18207
rect 34989 18173 35023 18207
rect 35023 18173 35032 18207
rect 34980 18164 35032 18173
rect 34152 18096 34204 18148
rect 17132 18028 17184 18080
rect 17316 18071 17368 18080
rect 17316 18037 17325 18071
rect 17325 18037 17359 18071
rect 17359 18037 17368 18071
rect 17316 18028 17368 18037
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 18144 18028 18196 18080
rect 19984 18028 20036 18080
rect 20812 18028 20864 18080
rect 20904 18028 20956 18080
rect 24860 18028 24912 18080
rect 24952 18028 25004 18080
rect 25136 18028 25188 18080
rect 26424 18071 26476 18080
rect 26424 18037 26433 18071
rect 26433 18037 26467 18071
rect 26467 18037 26476 18071
rect 26424 18028 26476 18037
rect 26608 18028 26660 18080
rect 27160 18028 27212 18080
rect 29000 18071 29052 18080
rect 29000 18037 29009 18071
rect 29009 18037 29043 18071
rect 29043 18037 29052 18071
rect 29000 18028 29052 18037
rect 31116 18071 31168 18080
rect 31116 18037 31125 18071
rect 31125 18037 31159 18071
rect 31159 18037 31168 18071
rect 31116 18028 31168 18037
rect 33232 18028 33284 18080
rect 39028 18368 39080 18420
rect 39304 18368 39356 18420
rect 40040 18411 40092 18420
rect 40040 18377 40049 18411
rect 40049 18377 40083 18411
rect 40083 18377 40092 18411
rect 40040 18368 40092 18377
rect 41512 18368 41564 18420
rect 37096 18300 37148 18352
rect 37280 18300 37332 18352
rect 36912 18207 36964 18216
rect 36912 18173 36921 18207
rect 36921 18173 36955 18207
rect 36955 18173 36964 18207
rect 36912 18164 36964 18173
rect 38476 18096 38528 18148
rect 40960 18300 41012 18352
rect 42708 18368 42760 18420
rect 42984 18368 43036 18420
rect 43720 18368 43772 18420
rect 44824 18368 44876 18420
rect 38936 18164 38988 18216
rect 39856 18164 39908 18216
rect 40316 18164 40368 18216
rect 42800 18300 42852 18352
rect 41696 18232 41748 18284
rect 42064 18164 42116 18216
rect 42800 18164 42852 18216
rect 43812 18207 43864 18216
rect 43812 18173 43821 18207
rect 43821 18173 43855 18207
rect 43855 18173 43864 18207
rect 43812 18164 43864 18173
rect 37280 18028 37332 18080
rect 38936 18028 38988 18080
rect 39028 18028 39080 18080
rect 40592 18071 40644 18080
rect 40592 18037 40601 18071
rect 40601 18037 40635 18071
rect 40635 18037 40644 18071
rect 40592 18028 40644 18037
rect 41512 18028 41564 18080
rect 42248 18028 42300 18080
rect 3570 17926 3622 17978
rect 3634 17926 3686 17978
rect 3698 17926 3750 17978
rect 3762 17926 3814 17978
rect 3826 17926 3878 17978
rect 8570 17926 8622 17978
rect 8634 17926 8686 17978
rect 8698 17926 8750 17978
rect 8762 17926 8814 17978
rect 8826 17926 8878 17978
rect 13570 17926 13622 17978
rect 13634 17926 13686 17978
rect 13698 17926 13750 17978
rect 13762 17926 13814 17978
rect 13826 17926 13878 17978
rect 18570 17926 18622 17978
rect 18634 17926 18686 17978
rect 18698 17926 18750 17978
rect 18762 17926 18814 17978
rect 18826 17926 18878 17978
rect 23570 17926 23622 17978
rect 23634 17926 23686 17978
rect 23698 17926 23750 17978
rect 23762 17926 23814 17978
rect 23826 17926 23878 17978
rect 28570 17926 28622 17978
rect 28634 17926 28686 17978
rect 28698 17926 28750 17978
rect 28762 17926 28814 17978
rect 28826 17926 28878 17978
rect 33570 17926 33622 17978
rect 33634 17926 33686 17978
rect 33698 17926 33750 17978
rect 33762 17926 33814 17978
rect 33826 17926 33878 17978
rect 38570 17926 38622 17978
rect 38634 17926 38686 17978
rect 38698 17926 38750 17978
rect 38762 17926 38814 17978
rect 38826 17926 38878 17978
rect 43570 17926 43622 17978
rect 43634 17926 43686 17978
rect 43698 17926 43750 17978
rect 43762 17926 43814 17978
rect 43826 17926 43878 17978
rect 4436 17867 4488 17876
rect 4436 17833 4445 17867
rect 4445 17833 4479 17867
rect 4479 17833 4488 17867
rect 4436 17824 4488 17833
rect 6368 17824 6420 17876
rect 6828 17824 6880 17876
rect 7748 17824 7800 17876
rect 8392 17867 8444 17876
rect 8392 17833 8401 17867
rect 8401 17833 8435 17867
rect 8435 17833 8444 17867
rect 8392 17824 8444 17833
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 9588 17867 9640 17876
rect 9588 17833 9597 17867
rect 9597 17833 9631 17867
rect 9631 17833 9640 17867
rect 9588 17824 9640 17833
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 12716 17824 12768 17876
rect 12992 17824 13044 17876
rect 13360 17824 13412 17876
rect 16304 17824 16356 17876
rect 5540 17688 5592 17740
rect 4160 17552 4212 17604
rect 4436 17620 4488 17672
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 8024 17620 8076 17672
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 3976 17484 4028 17536
rect 6644 17595 6696 17604
rect 6644 17561 6653 17595
rect 6653 17561 6687 17595
rect 6687 17561 6696 17595
rect 6644 17552 6696 17561
rect 5632 17484 5684 17536
rect 5816 17484 5868 17536
rect 6552 17484 6604 17536
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 11336 17756 11388 17808
rect 10140 17688 10192 17740
rect 12256 17688 12308 17740
rect 12532 17731 12584 17740
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 15200 17756 15252 17808
rect 12348 17620 12400 17672
rect 13360 17620 13412 17672
rect 15108 17688 15160 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 16028 17731 16080 17740
rect 16028 17697 16037 17731
rect 16037 17697 16071 17731
rect 16071 17697 16080 17731
rect 16028 17688 16080 17697
rect 16764 17756 16816 17808
rect 16948 17756 17000 17808
rect 17960 17824 18012 17876
rect 19616 17824 19668 17876
rect 19984 17824 20036 17876
rect 20352 17824 20404 17876
rect 20812 17867 20864 17876
rect 20812 17833 20821 17867
rect 20821 17833 20855 17867
rect 20855 17833 20864 17867
rect 20812 17824 20864 17833
rect 21916 17824 21968 17876
rect 22376 17824 22428 17876
rect 22744 17824 22796 17876
rect 27528 17824 27580 17876
rect 9772 17552 9824 17604
rect 8852 17484 8904 17536
rect 9956 17484 10008 17536
rect 10784 17484 10836 17536
rect 12992 17552 13044 17604
rect 13912 17620 13964 17672
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 16856 17688 16908 17740
rect 17316 17688 17368 17740
rect 17684 17688 17736 17740
rect 16580 17620 16632 17672
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 17500 17620 17552 17672
rect 17592 17620 17644 17672
rect 18144 17620 18196 17672
rect 19708 17688 19760 17740
rect 20996 17756 21048 17808
rect 21180 17688 21232 17740
rect 22008 17688 22060 17740
rect 12440 17484 12492 17536
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 14280 17484 14332 17536
rect 14740 17484 14792 17536
rect 16488 17484 16540 17536
rect 16856 17595 16908 17604
rect 16856 17561 16865 17595
rect 16865 17561 16899 17595
rect 16899 17561 16908 17595
rect 16856 17552 16908 17561
rect 17040 17552 17092 17604
rect 19340 17552 19392 17604
rect 17316 17527 17368 17536
rect 17316 17493 17325 17527
rect 17325 17493 17359 17527
rect 17359 17493 17368 17527
rect 17316 17484 17368 17493
rect 18880 17484 18932 17536
rect 19432 17484 19484 17536
rect 19524 17527 19576 17536
rect 19524 17493 19533 17527
rect 19533 17493 19567 17527
rect 19567 17493 19576 17527
rect 19524 17484 19576 17493
rect 20444 17620 20496 17672
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 23296 17731 23348 17740
rect 23296 17697 23305 17731
rect 23305 17697 23339 17731
rect 23339 17697 23348 17731
rect 23296 17688 23348 17697
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 24860 17688 24912 17740
rect 19984 17595 20036 17604
rect 19984 17561 19993 17595
rect 19993 17561 20027 17595
rect 20027 17561 20036 17595
rect 19984 17552 20036 17561
rect 20628 17552 20680 17604
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 26792 17620 26844 17672
rect 27160 17663 27212 17672
rect 27160 17629 27183 17663
rect 27183 17629 27212 17663
rect 27160 17620 27212 17629
rect 29920 17824 29972 17876
rect 31116 17824 31168 17876
rect 31208 17867 31260 17876
rect 31208 17833 31217 17867
rect 31217 17833 31251 17867
rect 31251 17833 31260 17867
rect 31208 17824 31260 17833
rect 31576 17824 31628 17876
rect 32864 17824 32916 17876
rect 32956 17824 33008 17876
rect 34980 17824 35032 17876
rect 35992 17824 36044 17876
rect 36912 17824 36964 17876
rect 38200 17824 38252 17876
rect 39488 17824 39540 17876
rect 40040 17824 40092 17876
rect 40316 17867 40368 17876
rect 40316 17833 40325 17867
rect 40325 17833 40359 17867
rect 40359 17833 40368 17867
rect 40316 17824 40368 17833
rect 28448 17756 28500 17808
rect 30564 17756 30616 17808
rect 28540 17688 28592 17740
rect 31668 17756 31720 17808
rect 31852 17756 31904 17808
rect 42248 17824 42300 17876
rect 44916 17824 44968 17876
rect 32220 17731 32272 17740
rect 32220 17697 32229 17731
rect 32229 17697 32263 17731
rect 32263 17697 32272 17731
rect 32220 17688 32272 17697
rect 32588 17688 32640 17740
rect 33784 17688 33836 17740
rect 35624 17688 35676 17740
rect 24308 17552 24360 17604
rect 20352 17484 20404 17536
rect 20996 17484 21048 17536
rect 21640 17527 21692 17536
rect 21640 17493 21649 17527
rect 21649 17493 21683 17527
rect 21683 17493 21692 17527
rect 21640 17484 21692 17493
rect 21916 17484 21968 17536
rect 22560 17527 22612 17536
rect 22560 17493 22569 17527
rect 22569 17493 22603 17527
rect 22603 17493 22612 17527
rect 22560 17484 22612 17493
rect 23204 17527 23256 17536
rect 23204 17493 23213 17527
rect 23213 17493 23247 17527
rect 23247 17493 23256 17527
rect 23204 17484 23256 17493
rect 23480 17484 23532 17536
rect 26608 17552 26660 17604
rect 25412 17484 25464 17536
rect 27344 17484 27396 17536
rect 27620 17484 27672 17536
rect 28724 17484 28776 17536
rect 30472 17620 30524 17672
rect 30196 17552 30248 17604
rect 30840 17595 30892 17604
rect 30840 17561 30849 17595
rect 30849 17561 30883 17595
rect 30883 17561 30892 17595
rect 30840 17552 30892 17561
rect 30564 17484 30616 17536
rect 31484 17484 31536 17536
rect 31760 17663 31812 17672
rect 31760 17629 31769 17663
rect 31769 17629 31803 17663
rect 31803 17629 31812 17663
rect 31760 17620 31812 17629
rect 32312 17552 32364 17604
rect 34520 17552 34572 17604
rect 35348 17620 35400 17672
rect 35532 17620 35584 17672
rect 37188 17688 37240 17740
rect 36176 17663 36228 17672
rect 36176 17629 36185 17663
rect 36185 17629 36219 17663
rect 36219 17629 36228 17663
rect 36176 17620 36228 17629
rect 37740 17620 37792 17672
rect 39028 17688 39080 17740
rect 39488 17688 39540 17740
rect 41328 17688 41380 17740
rect 42984 17731 43036 17740
rect 42984 17697 42993 17731
rect 42993 17697 43027 17731
rect 43027 17697 43036 17731
rect 42984 17688 43036 17697
rect 43076 17731 43128 17740
rect 43076 17697 43085 17731
rect 43085 17697 43119 17731
rect 43119 17697 43128 17731
rect 43076 17688 43128 17697
rect 32128 17484 32180 17536
rect 32404 17484 32456 17536
rect 33048 17484 33100 17536
rect 34796 17527 34848 17536
rect 34796 17493 34805 17527
rect 34805 17493 34839 17527
rect 34839 17493 34848 17527
rect 34796 17484 34848 17493
rect 35900 17552 35952 17604
rect 35992 17552 36044 17604
rect 37280 17552 37332 17604
rect 36452 17484 36504 17536
rect 36912 17484 36964 17536
rect 37464 17484 37516 17536
rect 39120 17484 39172 17536
rect 40132 17552 40184 17604
rect 39396 17484 39448 17536
rect 40040 17484 40092 17536
rect 40592 17620 40644 17672
rect 43260 17620 43312 17672
rect 41420 17552 41472 17604
rect 42432 17552 42484 17604
rect 43536 17527 43588 17536
rect 43536 17493 43545 17527
rect 43545 17493 43579 17527
rect 43579 17493 43588 17527
rect 43904 17527 43956 17536
rect 43536 17484 43588 17493
rect 43904 17493 43913 17527
rect 43913 17493 43947 17527
rect 43947 17493 43956 17527
rect 43904 17484 43956 17493
rect 44916 17527 44968 17536
rect 44916 17493 44925 17527
rect 44925 17493 44959 17527
rect 44959 17493 44968 17527
rect 44916 17484 44968 17493
rect 6070 17382 6122 17434
rect 6134 17382 6186 17434
rect 6198 17382 6250 17434
rect 6262 17382 6314 17434
rect 6326 17382 6378 17434
rect 11070 17382 11122 17434
rect 11134 17382 11186 17434
rect 11198 17382 11250 17434
rect 11262 17382 11314 17434
rect 11326 17382 11378 17434
rect 16070 17382 16122 17434
rect 16134 17382 16186 17434
rect 16198 17382 16250 17434
rect 16262 17382 16314 17434
rect 16326 17382 16378 17434
rect 21070 17382 21122 17434
rect 21134 17382 21186 17434
rect 21198 17382 21250 17434
rect 21262 17382 21314 17434
rect 21326 17382 21378 17434
rect 26070 17382 26122 17434
rect 26134 17382 26186 17434
rect 26198 17382 26250 17434
rect 26262 17382 26314 17434
rect 26326 17382 26378 17434
rect 31070 17382 31122 17434
rect 31134 17382 31186 17434
rect 31198 17382 31250 17434
rect 31262 17382 31314 17434
rect 31326 17382 31378 17434
rect 36070 17382 36122 17434
rect 36134 17382 36186 17434
rect 36198 17382 36250 17434
rect 36262 17382 36314 17434
rect 36326 17382 36378 17434
rect 41070 17382 41122 17434
rect 41134 17382 41186 17434
rect 41198 17382 41250 17434
rect 41262 17382 41314 17434
rect 41326 17382 41378 17434
rect 5632 17280 5684 17332
rect 6552 17280 6604 17332
rect 6644 17280 6696 17332
rect 7564 17280 7616 17332
rect 7840 17280 7892 17332
rect 8024 17280 8076 17332
rect 8852 17280 8904 17332
rect 9772 17323 9824 17332
rect 9772 17289 9781 17323
rect 9781 17289 9815 17323
rect 9815 17289 9824 17323
rect 9772 17280 9824 17289
rect 4528 17212 4580 17264
rect 4620 17212 4672 17264
rect 5448 17144 5500 17196
rect 5908 17144 5960 17196
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 3332 17076 3384 17128
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 4160 17076 4212 17128
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 5816 17076 5868 17085
rect 7012 17076 7064 17128
rect 12808 17280 12860 17332
rect 13360 17280 13412 17332
rect 14832 17255 14884 17264
rect 14832 17221 14841 17255
rect 14841 17221 14875 17255
rect 14875 17221 14884 17255
rect 14832 17212 14884 17221
rect 15200 17280 15252 17332
rect 16672 17280 16724 17332
rect 17040 17280 17092 17332
rect 18880 17280 18932 17332
rect 9680 17144 9732 17196
rect 9956 17076 10008 17128
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10784 17144 10836 17196
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 12256 17144 12308 17196
rect 14280 17144 14332 17196
rect 15568 17187 15620 17196
rect 15568 17153 15583 17187
rect 15583 17153 15617 17187
rect 15617 17153 15620 17187
rect 15568 17144 15620 17153
rect 15844 17144 15896 17196
rect 16580 17144 16632 17196
rect 16948 17144 17000 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 16304 17119 16356 17128
rect 16304 17085 16313 17119
rect 16313 17085 16347 17119
rect 16347 17085 16356 17119
rect 16304 17076 16356 17085
rect 15292 17008 15344 17060
rect 15568 17008 15620 17060
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 8116 16940 8168 16992
rect 8576 16940 8628 16992
rect 9036 16940 9088 16992
rect 10048 16940 10100 16992
rect 10784 16940 10836 16992
rect 12440 16940 12492 16992
rect 15016 16983 15068 16992
rect 15016 16949 15025 16983
rect 15025 16949 15059 16983
rect 15059 16949 15068 16983
rect 15016 16940 15068 16949
rect 15476 16940 15528 16992
rect 15936 16940 15988 16992
rect 16396 17008 16448 17060
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 17868 17144 17920 17196
rect 18236 17144 18288 17196
rect 19524 17280 19576 17332
rect 19432 17212 19484 17264
rect 19984 17280 20036 17332
rect 20260 17280 20312 17332
rect 20444 17323 20496 17332
rect 20444 17289 20453 17323
rect 20453 17289 20487 17323
rect 20487 17289 20496 17323
rect 20444 17280 20496 17289
rect 20628 17323 20680 17332
rect 20628 17289 20637 17323
rect 20637 17289 20671 17323
rect 20671 17289 20680 17323
rect 20628 17280 20680 17289
rect 22376 17323 22428 17332
rect 22376 17289 22385 17323
rect 22385 17289 22419 17323
rect 22419 17289 22428 17323
rect 22376 17280 22428 17289
rect 22560 17280 22612 17332
rect 17132 17008 17184 17060
rect 19708 17187 19760 17196
rect 19708 17153 19717 17187
rect 19717 17153 19751 17187
rect 19751 17153 19760 17187
rect 19708 17144 19760 17153
rect 19892 17187 19944 17230
rect 19892 17178 19902 17187
rect 19902 17178 19936 17187
rect 19936 17178 19944 17187
rect 18420 17008 18472 17060
rect 19340 17008 19392 17060
rect 20168 17119 20220 17128
rect 20168 17085 20177 17119
rect 20177 17085 20211 17119
rect 20211 17085 20220 17119
rect 20168 17076 20220 17085
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 20996 17144 21048 17196
rect 24308 17323 24360 17332
rect 24308 17289 24317 17323
rect 24317 17289 24351 17323
rect 24351 17289 24360 17323
rect 24308 17280 24360 17289
rect 24952 17280 25004 17332
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 27896 17323 27948 17332
rect 27896 17289 27905 17323
rect 27905 17289 27939 17323
rect 27939 17289 27948 17323
rect 27896 17280 27948 17289
rect 24216 17212 24268 17264
rect 26424 17212 26476 17264
rect 24400 17187 24452 17196
rect 24400 17153 24409 17187
rect 24409 17153 24443 17187
rect 24443 17153 24452 17187
rect 24400 17144 24452 17153
rect 24952 17187 25004 17196
rect 24952 17153 24961 17187
rect 24961 17153 24995 17187
rect 24995 17153 25004 17187
rect 24952 17144 25004 17153
rect 29000 17280 29052 17332
rect 29552 17280 29604 17332
rect 30380 17280 30432 17332
rect 30472 17280 30524 17332
rect 30840 17280 30892 17332
rect 28356 17212 28408 17264
rect 20536 17076 20588 17128
rect 25228 17076 25280 17128
rect 20352 17008 20404 17060
rect 20904 17051 20956 17060
rect 20904 17017 20913 17051
rect 20913 17017 20947 17051
rect 20947 17017 20956 17051
rect 20904 17008 20956 17017
rect 22284 17008 22336 17060
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 17684 16940 17736 16992
rect 18328 16940 18380 16992
rect 19524 16983 19576 16992
rect 19524 16949 19533 16983
rect 19533 16949 19567 16983
rect 19567 16949 19576 16983
rect 19524 16940 19576 16949
rect 21640 16940 21692 16992
rect 22376 16940 22428 16992
rect 23940 16940 23992 16992
rect 24768 16983 24820 16992
rect 24768 16949 24777 16983
rect 24777 16949 24811 16983
rect 24811 16949 24820 16983
rect 24768 16940 24820 16949
rect 26792 16940 26844 16992
rect 28264 17187 28316 17196
rect 28264 17153 28298 17187
rect 28298 17153 28316 17187
rect 28264 17144 28316 17153
rect 28540 17212 28592 17264
rect 31760 17280 31812 17332
rect 29276 17144 29328 17196
rect 28724 16940 28776 16992
rect 29000 16940 29052 16992
rect 29276 16940 29328 16992
rect 29368 16983 29420 16992
rect 29368 16949 29377 16983
rect 29377 16949 29411 16983
rect 29411 16949 29420 16983
rect 29368 16940 29420 16949
rect 29920 17008 29972 17060
rect 30564 17187 30616 17196
rect 30564 17153 30573 17187
rect 30573 17153 30607 17187
rect 30607 17153 30616 17187
rect 30564 17144 30616 17153
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 32036 17280 32088 17332
rect 32312 17280 32364 17332
rect 31024 17144 31076 17196
rect 32588 17212 32640 17264
rect 32680 17255 32732 17264
rect 32680 17221 32689 17255
rect 32689 17221 32723 17255
rect 32723 17221 32732 17255
rect 32680 17212 32732 17221
rect 32864 17323 32916 17332
rect 32864 17289 32889 17323
rect 32889 17289 32916 17323
rect 32864 17280 32916 17289
rect 33140 17280 33192 17332
rect 33784 17323 33836 17332
rect 33784 17289 33793 17323
rect 33793 17289 33827 17323
rect 33827 17289 33836 17323
rect 33784 17280 33836 17289
rect 34520 17280 34572 17332
rect 34796 17280 34848 17332
rect 34888 17280 34940 17332
rect 39028 17280 39080 17332
rect 31760 17187 31812 17196
rect 31760 17153 31769 17187
rect 31769 17153 31803 17187
rect 31803 17153 31812 17187
rect 31760 17144 31812 17153
rect 31852 17144 31904 17196
rect 32312 17119 32364 17128
rect 30564 17008 30616 17060
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 32496 17119 32548 17128
rect 32496 17085 32505 17119
rect 32505 17085 32539 17119
rect 32539 17085 32548 17119
rect 32496 17076 32548 17085
rect 32772 17144 32824 17196
rect 34060 17144 34112 17196
rect 38200 17255 38252 17264
rect 38200 17221 38209 17255
rect 38209 17221 38243 17255
rect 38243 17221 38252 17255
rect 38200 17212 38252 17221
rect 38936 17212 38988 17264
rect 40040 17255 40092 17264
rect 40040 17221 40049 17255
rect 40049 17221 40083 17255
rect 40083 17221 40092 17255
rect 41512 17280 41564 17332
rect 42800 17323 42852 17332
rect 42800 17289 42809 17323
rect 42809 17289 42843 17323
rect 42843 17289 42852 17323
rect 42800 17280 42852 17289
rect 43168 17280 43220 17332
rect 43904 17323 43956 17332
rect 43904 17289 43913 17323
rect 43913 17289 43947 17323
rect 43947 17289 43956 17323
rect 43904 17280 43956 17289
rect 40040 17212 40092 17221
rect 42432 17212 42484 17264
rect 36820 17187 36872 17196
rect 36820 17153 36829 17187
rect 36829 17153 36863 17187
rect 36863 17153 36872 17187
rect 36820 17144 36872 17153
rect 37464 17144 37516 17196
rect 39580 17144 39632 17196
rect 40132 17187 40184 17196
rect 40132 17153 40141 17187
rect 40141 17153 40175 17187
rect 40175 17153 40184 17187
rect 40132 17144 40184 17153
rect 37280 17008 37332 17060
rect 39764 17051 39816 17060
rect 39764 17017 39773 17051
rect 39773 17017 39807 17051
rect 39807 17017 39816 17051
rect 39764 17008 39816 17017
rect 40960 17144 41012 17196
rect 41604 17144 41656 17196
rect 43352 17144 43404 17196
rect 44916 17144 44968 17196
rect 41052 17076 41104 17128
rect 41512 17076 41564 17128
rect 41880 17076 41932 17128
rect 31116 16983 31168 16992
rect 31116 16949 31125 16983
rect 31125 16949 31159 16983
rect 31159 16949 31168 16983
rect 31116 16940 31168 16949
rect 33232 16940 33284 16992
rect 34520 16940 34572 16992
rect 36176 16983 36228 16992
rect 36176 16949 36185 16983
rect 36185 16949 36219 16983
rect 36219 16949 36228 16983
rect 36176 16940 36228 16949
rect 36636 16983 36688 16992
rect 36636 16949 36645 16983
rect 36645 16949 36679 16983
rect 36679 16949 36688 16983
rect 36636 16940 36688 16949
rect 37188 16983 37240 16992
rect 37188 16949 37197 16983
rect 37197 16949 37231 16983
rect 37231 16949 37240 16983
rect 37188 16940 37240 16949
rect 37464 16983 37516 16992
rect 37464 16949 37473 16983
rect 37473 16949 37507 16983
rect 37507 16949 37516 16983
rect 37464 16940 37516 16949
rect 38936 16940 38988 16992
rect 39580 16940 39632 16992
rect 39856 16940 39908 16992
rect 40592 16983 40644 16992
rect 40592 16949 40601 16983
rect 40601 16949 40635 16983
rect 40635 16949 40644 16983
rect 40592 16940 40644 16949
rect 41788 16983 41840 16992
rect 41788 16949 41797 16983
rect 41797 16949 41831 16983
rect 41831 16949 41840 16983
rect 41788 16940 41840 16949
rect 42800 16940 42852 16992
rect 43536 16983 43588 16992
rect 43536 16949 43545 16983
rect 43545 16949 43579 16983
rect 43579 16949 43588 16983
rect 44640 16983 44692 16992
rect 43536 16940 43588 16949
rect 44640 16949 44649 16983
rect 44649 16949 44683 16983
rect 44683 16949 44692 16983
rect 44640 16940 44692 16949
rect 3570 16838 3622 16890
rect 3634 16838 3686 16890
rect 3698 16838 3750 16890
rect 3762 16838 3814 16890
rect 3826 16838 3878 16890
rect 8570 16838 8622 16890
rect 8634 16838 8686 16890
rect 8698 16838 8750 16890
rect 8762 16838 8814 16890
rect 8826 16838 8878 16890
rect 13570 16838 13622 16890
rect 13634 16838 13686 16890
rect 13698 16838 13750 16890
rect 13762 16838 13814 16890
rect 13826 16838 13878 16890
rect 18570 16838 18622 16890
rect 18634 16838 18686 16890
rect 18698 16838 18750 16890
rect 18762 16838 18814 16890
rect 18826 16838 18878 16890
rect 23570 16838 23622 16890
rect 23634 16838 23686 16890
rect 23698 16838 23750 16890
rect 23762 16838 23814 16890
rect 23826 16838 23878 16890
rect 28570 16838 28622 16890
rect 28634 16838 28686 16890
rect 28698 16838 28750 16890
rect 28762 16838 28814 16890
rect 28826 16838 28878 16890
rect 33570 16838 33622 16890
rect 33634 16838 33686 16890
rect 33698 16838 33750 16890
rect 33762 16838 33814 16890
rect 33826 16838 33878 16890
rect 38570 16838 38622 16890
rect 38634 16838 38686 16890
rect 38698 16838 38750 16890
rect 38762 16838 38814 16890
rect 38826 16838 38878 16890
rect 43570 16838 43622 16890
rect 43634 16838 43686 16890
rect 43698 16838 43750 16890
rect 43762 16838 43814 16890
rect 43826 16838 43878 16890
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 8024 16736 8076 16788
rect 4620 16600 4672 16652
rect 3332 16396 3384 16448
rect 4436 16532 4488 16584
rect 6644 16532 6696 16584
rect 9680 16668 9732 16720
rect 9956 16736 10008 16788
rect 10140 16736 10192 16788
rect 10416 16736 10468 16788
rect 10692 16736 10744 16788
rect 12992 16736 13044 16788
rect 10048 16600 10100 16652
rect 10416 16600 10468 16652
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 5080 16507 5132 16516
rect 5080 16473 5089 16507
rect 5089 16473 5123 16507
rect 5123 16473 5132 16507
rect 5080 16464 5132 16473
rect 6552 16439 6604 16448
rect 6552 16405 6561 16439
rect 6561 16405 6595 16439
rect 6595 16405 6604 16439
rect 6552 16396 6604 16405
rect 6828 16396 6880 16448
rect 8116 16439 8168 16448
rect 8116 16405 8125 16439
rect 8125 16405 8159 16439
rect 8159 16405 8168 16439
rect 8116 16396 8168 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 8576 16396 8628 16405
rect 9588 16532 9640 16584
rect 11888 16600 11940 16652
rect 11428 16532 11480 16584
rect 14556 16600 14608 16652
rect 15292 16600 15344 16652
rect 16304 16736 16356 16788
rect 16488 16736 16540 16788
rect 17040 16736 17092 16788
rect 19616 16736 19668 16788
rect 20168 16736 20220 16788
rect 20996 16736 21048 16788
rect 17408 16600 17460 16652
rect 17684 16600 17736 16652
rect 19524 16600 19576 16652
rect 12164 16532 12216 16584
rect 18144 16532 18196 16584
rect 9220 16439 9272 16448
rect 9220 16405 9229 16439
rect 9229 16405 9263 16439
rect 9263 16405 9272 16439
rect 9220 16396 9272 16405
rect 11612 16464 11664 16516
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 11796 16396 11848 16448
rect 12440 16396 12492 16448
rect 13360 16396 13412 16448
rect 14280 16396 14332 16448
rect 19340 16464 19392 16516
rect 20352 16464 20404 16516
rect 18328 16396 18380 16448
rect 18512 16396 18564 16448
rect 20168 16396 20220 16448
rect 20812 16532 20864 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 23204 16736 23256 16788
rect 24952 16736 25004 16788
rect 28264 16736 28316 16788
rect 30656 16736 30708 16788
rect 21272 16532 21324 16584
rect 21456 16532 21508 16584
rect 24400 16643 24452 16652
rect 22284 16532 22336 16584
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 25136 16600 25188 16652
rect 25228 16643 25280 16652
rect 25228 16609 25237 16643
rect 25237 16609 25271 16643
rect 25271 16609 25280 16643
rect 25228 16600 25280 16609
rect 26424 16600 26476 16652
rect 26608 16600 26660 16652
rect 27344 16600 27396 16652
rect 24032 16532 24084 16584
rect 26976 16532 27028 16584
rect 21732 16464 21784 16516
rect 27896 16532 27948 16584
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 28172 16532 28224 16541
rect 28356 16532 28408 16584
rect 28632 16532 28684 16584
rect 29000 16668 29052 16720
rect 30656 16600 30708 16652
rect 31116 16736 31168 16788
rect 31668 16736 31720 16788
rect 32220 16736 32272 16788
rect 32312 16736 32364 16788
rect 35900 16779 35952 16788
rect 35900 16745 35909 16779
rect 35909 16745 35943 16779
rect 35943 16745 35952 16779
rect 35900 16736 35952 16745
rect 36820 16736 36872 16788
rect 37188 16736 37240 16788
rect 32128 16668 32180 16720
rect 33324 16668 33376 16720
rect 31484 16600 31536 16652
rect 32312 16600 32364 16652
rect 32496 16600 32548 16652
rect 33416 16600 33468 16652
rect 29368 16532 29420 16584
rect 29920 16575 29972 16584
rect 29920 16541 29929 16575
rect 29929 16541 29963 16575
rect 29963 16541 29972 16575
rect 29920 16532 29972 16541
rect 21272 16396 21324 16448
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 22376 16439 22428 16448
rect 22376 16405 22385 16439
rect 22385 16405 22419 16439
rect 22419 16405 22428 16439
rect 22376 16396 22428 16405
rect 23020 16396 23072 16448
rect 23296 16396 23348 16448
rect 23756 16439 23808 16448
rect 23756 16405 23765 16439
rect 23765 16405 23799 16439
rect 23799 16405 23808 16439
rect 23756 16396 23808 16405
rect 24124 16439 24176 16448
rect 24124 16405 24133 16439
rect 24133 16405 24167 16439
rect 24167 16405 24176 16439
rect 24124 16396 24176 16405
rect 24952 16439 25004 16448
rect 24952 16405 24961 16439
rect 24961 16405 24995 16439
rect 24995 16405 25004 16439
rect 24952 16396 25004 16405
rect 25412 16439 25464 16448
rect 25412 16405 25421 16439
rect 25421 16405 25455 16439
rect 25455 16405 25464 16439
rect 25412 16396 25464 16405
rect 25504 16396 25556 16448
rect 26884 16439 26936 16448
rect 26884 16405 26893 16439
rect 26893 16405 26927 16439
rect 26927 16405 26936 16439
rect 26884 16396 26936 16405
rect 28908 16464 28960 16516
rect 27620 16396 27672 16448
rect 27712 16439 27764 16448
rect 27712 16405 27721 16439
rect 27721 16405 27755 16439
rect 27755 16405 27764 16439
rect 27712 16396 27764 16405
rect 29184 16396 29236 16448
rect 29552 16464 29604 16516
rect 30564 16532 30616 16584
rect 30288 16396 30340 16448
rect 30840 16396 30892 16448
rect 30932 16396 30984 16448
rect 35992 16600 36044 16652
rect 34060 16575 34112 16584
rect 34060 16541 34069 16575
rect 34069 16541 34103 16575
rect 34103 16541 34112 16575
rect 34060 16532 34112 16541
rect 35808 16532 35860 16584
rect 37188 16600 37240 16652
rect 38200 16736 38252 16788
rect 39120 16736 39172 16788
rect 33692 16464 33744 16516
rect 34796 16464 34848 16516
rect 36452 16464 36504 16516
rect 38292 16532 38344 16584
rect 32956 16396 33008 16448
rect 33048 16439 33100 16448
rect 33048 16405 33057 16439
rect 33057 16405 33091 16439
rect 33091 16405 33100 16439
rect 33048 16396 33100 16405
rect 35716 16396 35768 16448
rect 35900 16396 35952 16448
rect 36176 16396 36228 16448
rect 36912 16396 36964 16448
rect 37924 16396 37976 16448
rect 38016 16439 38068 16448
rect 38016 16405 38025 16439
rect 38025 16405 38059 16439
rect 38059 16405 38068 16439
rect 38016 16396 38068 16405
rect 38844 16643 38896 16652
rect 38844 16609 38853 16643
rect 38853 16609 38887 16643
rect 38887 16609 38896 16643
rect 38844 16600 38896 16609
rect 39028 16600 39080 16652
rect 39948 16736 40000 16788
rect 40592 16736 40644 16788
rect 40960 16779 41012 16788
rect 40960 16745 40969 16779
rect 40969 16745 41003 16779
rect 41003 16745 41012 16779
rect 40960 16736 41012 16745
rect 43076 16736 43128 16788
rect 43904 16779 43956 16788
rect 43904 16745 43913 16779
rect 43913 16745 43947 16779
rect 43947 16745 43956 16779
rect 43904 16736 43956 16745
rect 44640 16736 44692 16788
rect 39212 16668 39264 16720
rect 38936 16532 38988 16584
rect 39120 16532 39172 16584
rect 40960 16532 41012 16584
rect 38844 16464 38896 16516
rect 39488 16464 39540 16516
rect 39948 16464 40000 16516
rect 41328 16464 41380 16516
rect 42708 16464 42760 16516
rect 43352 16643 43404 16652
rect 43352 16609 43361 16643
rect 43361 16609 43395 16643
rect 43395 16609 43404 16643
rect 43352 16600 43404 16609
rect 44180 16600 44232 16652
rect 44364 16532 44416 16584
rect 40776 16396 40828 16448
rect 41604 16396 41656 16448
rect 42892 16439 42944 16448
rect 42892 16405 42901 16439
rect 42901 16405 42935 16439
rect 42935 16405 42944 16439
rect 42892 16396 42944 16405
rect 6070 16294 6122 16346
rect 6134 16294 6186 16346
rect 6198 16294 6250 16346
rect 6262 16294 6314 16346
rect 6326 16294 6378 16346
rect 11070 16294 11122 16346
rect 11134 16294 11186 16346
rect 11198 16294 11250 16346
rect 11262 16294 11314 16346
rect 11326 16294 11378 16346
rect 16070 16294 16122 16346
rect 16134 16294 16186 16346
rect 16198 16294 16250 16346
rect 16262 16294 16314 16346
rect 16326 16294 16378 16346
rect 21070 16294 21122 16346
rect 21134 16294 21186 16346
rect 21198 16294 21250 16346
rect 21262 16294 21314 16346
rect 21326 16294 21378 16346
rect 26070 16294 26122 16346
rect 26134 16294 26186 16346
rect 26198 16294 26250 16346
rect 26262 16294 26314 16346
rect 26326 16294 26378 16346
rect 31070 16294 31122 16346
rect 31134 16294 31186 16346
rect 31198 16294 31250 16346
rect 31262 16294 31314 16346
rect 31326 16294 31378 16346
rect 36070 16294 36122 16346
rect 36134 16294 36186 16346
rect 36198 16294 36250 16346
rect 36262 16294 36314 16346
rect 36326 16294 36378 16346
rect 41070 16294 41122 16346
rect 41134 16294 41186 16346
rect 41198 16294 41250 16346
rect 41262 16294 41314 16346
rect 41326 16294 41378 16346
rect 4344 16192 4396 16244
rect 4620 16192 4672 16244
rect 5080 16192 5132 16244
rect 5448 16192 5500 16244
rect 7380 16235 7432 16244
rect 7380 16201 7389 16235
rect 7389 16201 7423 16235
rect 7423 16201 7432 16235
rect 7380 16192 7432 16201
rect 5448 16099 5500 16108
rect 5448 16065 5457 16099
rect 5457 16065 5491 16099
rect 5491 16065 5500 16099
rect 5448 16056 5500 16065
rect 3332 15988 3384 16040
rect 5448 15920 5500 15972
rect 5816 16031 5868 16040
rect 5816 15997 5825 16031
rect 5825 15997 5859 16031
rect 5859 15997 5868 16031
rect 5816 15988 5868 15997
rect 6552 16031 6604 16040
rect 6552 15997 6561 16031
rect 6561 15997 6595 16031
rect 6595 15997 6604 16031
rect 6552 15988 6604 15997
rect 8576 16192 8628 16244
rect 9220 16192 9272 16244
rect 8116 16124 8168 16176
rect 10324 16192 10376 16244
rect 11428 16124 11480 16176
rect 12256 16056 12308 16108
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 16396 16192 16448 16244
rect 16856 16192 16908 16244
rect 17224 16192 17276 16244
rect 17592 16192 17644 16244
rect 19708 16192 19760 16244
rect 21548 16235 21600 16244
rect 21548 16201 21557 16235
rect 21557 16201 21591 16235
rect 21591 16201 21600 16235
rect 21548 16192 21600 16201
rect 24032 16192 24084 16244
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 14280 16056 14332 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 15568 16099 15620 16108
rect 15568 16065 15577 16099
rect 15577 16065 15611 16099
rect 15611 16065 15620 16099
rect 15568 16056 15620 16065
rect 15936 16056 15988 16108
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 16580 16056 16632 16108
rect 16948 16124 17000 16176
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 18420 16167 18472 16176
rect 18420 16133 18429 16167
rect 18429 16133 18463 16167
rect 18463 16133 18472 16167
rect 18420 16124 18472 16133
rect 18512 16124 18564 16176
rect 20260 16167 20312 16176
rect 20260 16133 20269 16167
rect 20269 16133 20303 16167
rect 20303 16133 20312 16167
rect 20260 16124 20312 16133
rect 21732 16124 21784 16176
rect 24216 16124 24268 16176
rect 24768 16124 24820 16176
rect 27620 16192 27672 16244
rect 28724 16192 28776 16244
rect 29552 16192 29604 16244
rect 30104 16192 30156 16244
rect 32036 16192 32088 16244
rect 33048 16192 33100 16244
rect 3424 15852 3476 15904
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 9680 15895 9732 15904
rect 9680 15861 9689 15895
rect 9689 15861 9723 15895
rect 9723 15861 9732 15895
rect 9680 15852 9732 15861
rect 10140 15852 10192 15904
rect 10416 15852 10468 15904
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 14188 15988 14240 16040
rect 14740 15988 14792 16040
rect 16488 15988 16540 16040
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 17684 16056 17736 16108
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 20168 16056 20220 16108
rect 12716 15920 12768 15972
rect 16672 15920 16724 15972
rect 16764 15920 16816 15972
rect 17592 15920 17644 15972
rect 12164 15852 12216 15904
rect 12624 15895 12676 15904
rect 12624 15861 12633 15895
rect 12633 15861 12667 15895
rect 12667 15861 12676 15895
rect 12624 15852 12676 15861
rect 14280 15852 14332 15904
rect 16948 15852 17000 15904
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 20812 16056 20864 16108
rect 19892 15963 19944 15972
rect 19892 15929 19901 15963
rect 19901 15929 19935 15963
rect 19935 15929 19944 15963
rect 19892 15920 19944 15929
rect 18236 15852 18288 15904
rect 21088 15920 21140 15972
rect 21916 16099 21968 16108
rect 21916 16065 21925 16099
rect 21925 16065 21959 16099
rect 21959 16065 21968 16099
rect 21916 16056 21968 16065
rect 26332 16056 26384 16108
rect 27068 16099 27120 16108
rect 27068 16065 27077 16099
rect 27077 16065 27111 16099
rect 27111 16065 27120 16099
rect 27068 16056 27120 16065
rect 27712 16056 27764 16108
rect 28264 16056 28316 16108
rect 28724 16056 28776 16108
rect 30196 16124 30248 16176
rect 22100 15988 22152 16040
rect 22284 15988 22336 16040
rect 20812 15852 20864 15904
rect 21916 15852 21968 15904
rect 22652 16031 22704 16040
rect 22652 15997 22661 16031
rect 22661 15997 22695 16031
rect 22695 15997 22704 16031
rect 22652 15988 22704 15997
rect 22468 15852 22520 15904
rect 24860 15988 24912 16040
rect 24952 15988 25004 16040
rect 26884 15988 26936 16040
rect 26516 15963 26568 15972
rect 26516 15929 26525 15963
rect 26525 15929 26559 15963
rect 26559 15929 26568 15963
rect 26516 15920 26568 15929
rect 29276 16056 29328 16108
rect 32312 16124 32364 16176
rect 34060 16124 34112 16176
rect 29092 15988 29144 16040
rect 29092 15852 29144 15904
rect 29736 16031 29788 16040
rect 29736 15997 29745 16031
rect 29745 15997 29779 16031
rect 29779 15997 29788 16031
rect 29736 15988 29788 15997
rect 30932 15988 30984 16040
rect 34796 16056 34848 16108
rect 35992 16192 36044 16244
rect 36636 16124 36688 16176
rect 39212 16124 39264 16176
rect 40132 16192 40184 16244
rect 40684 16235 40736 16244
rect 40684 16201 40693 16235
rect 40693 16201 40727 16235
rect 40727 16201 40736 16235
rect 40684 16192 40736 16201
rect 42892 16192 42944 16244
rect 43352 16192 43404 16244
rect 35716 16099 35768 16108
rect 35716 16065 35725 16099
rect 35725 16065 35759 16099
rect 35759 16065 35768 16099
rect 35716 16056 35768 16065
rect 32772 15988 32824 16040
rect 33416 15988 33468 16040
rect 35256 15988 35308 16040
rect 35440 15988 35492 16040
rect 35808 15988 35860 16040
rect 37924 16056 37976 16108
rect 40776 16099 40828 16108
rect 40776 16065 40785 16099
rect 40785 16065 40819 16099
rect 40819 16065 40828 16099
rect 40776 16056 40828 16065
rect 36636 16031 36688 16040
rect 36636 15997 36645 16031
rect 36645 15997 36679 16031
rect 36679 15997 36688 16031
rect 36636 15988 36688 15997
rect 37464 15988 37516 16040
rect 38476 16031 38528 16040
rect 38476 15997 38485 16031
rect 38485 15997 38519 16031
rect 38519 15997 38528 16031
rect 38476 15988 38528 15997
rect 38016 15920 38068 15972
rect 39488 15988 39540 16040
rect 41604 16099 41656 16108
rect 41604 16065 41613 16099
rect 41613 16065 41647 16099
rect 41647 16065 41656 16099
rect 41604 16056 41656 16065
rect 43168 16056 43220 16108
rect 41788 16031 41840 16040
rect 41788 15997 41797 16031
rect 41797 15997 41831 16031
rect 41831 15997 41840 16031
rect 41788 15988 41840 15997
rect 32956 15852 33008 15904
rect 35072 15852 35124 15904
rect 38200 15852 38252 15904
rect 39764 15852 39816 15904
rect 40500 15852 40552 15904
rect 43904 15895 43956 15904
rect 43904 15861 43913 15895
rect 43913 15861 43947 15895
rect 43947 15861 43956 15895
rect 43904 15852 43956 15861
rect 44364 15852 44416 15904
rect 3570 15750 3622 15802
rect 3634 15750 3686 15802
rect 3698 15750 3750 15802
rect 3762 15750 3814 15802
rect 3826 15750 3878 15802
rect 8570 15750 8622 15802
rect 8634 15750 8686 15802
rect 8698 15750 8750 15802
rect 8762 15750 8814 15802
rect 8826 15750 8878 15802
rect 13570 15750 13622 15802
rect 13634 15750 13686 15802
rect 13698 15750 13750 15802
rect 13762 15750 13814 15802
rect 13826 15750 13878 15802
rect 18570 15750 18622 15802
rect 18634 15750 18686 15802
rect 18698 15750 18750 15802
rect 18762 15750 18814 15802
rect 18826 15750 18878 15802
rect 23570 15750 23622 15802
rect 23634 15750 23686 15802
rect 23698 15750 23750 15802
rect 23762 15750 23814 15802
rect 23826 15750 23878 15802
rect 28570 15750 28622 15802
rect 28634 15750 28686 15802
rect 28698 15750 28750 15802
rect 28762 15750 28814 15802
rect 28826 15750 28878 15802
rect 33570 15750 33622 15802
rect 33634 15750 33686 15802
rect 33698 15750 33750 15802
rect 33762 15750 33814 15802
rect 33826 15750 33878 15802
rect 38570 15750 38622 15802
rect 38634 15750 38686 15802
rect 38698 15750 38750 15802
rect 38762 15750 38814 15802
rect 38826 15750 38878 15802
rect 43570 15750 43622 15802
rect 43634 15750 43686 15802
rect 43698 15750 43750 15802
rect 43762 15750 43814 15802
rect 43826 15750 43878 15802
rect 4344 15648 4396 15700
rect 5816 15648 5868 15700
rect 4528 15512 4580 15564
rect 5448 15512 5500 15564
rect 6644 15444 6696 15496
rect 10140 15648 10192 15700
rect 9588 15580 9640 15632
rect 10416 15580 10468 15632
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8116 15444 8168 15496
rect 8208 15444 8260 15496
rect 9772 15512 9824 15564
rect 3424 15308 3476 15360
rect 11520 15648 11572 15700
rect 12624 15648 12676 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 14556 15648 14608 15700
rect 16764 15648 16816 15700
rect 17040 15648 17092 15700
rect 12256 15444 12308 15496
rect 10784 15376 10836 15428
rect 11152 15376 11204 15428
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 13360 15444 13412 15496
rect 14740 15512 14792 15564
rect 16856 15623 16908 15632
rect 16856 15589 16865 15623
rect 16865 15589 16899 15623
rect 16899 15589 16908 15623
rect 16856 15580 16908 15589
rect 9956 15308 10008 15360
rect 11796 15308 11848 15360
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 13084 15351 13136 15360
rect 13084 15317 13093 15351
rect 13093 15317 13127 15351
rect 13127 15317 13136 15351
rect 13084 15308 13136 15317
rect 13268 15376 13320 15428
rect 13912 15376 13964 15428
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 14924 15376 14976 15428
rect 15660 15376 15712 15428
rect 19432 15648 19484 15700
rect 20904 15648 20956 15700
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21456 15648 21508 15700
rect 21916 15648 21968 15700
rect 22560 15648 22612 15700
rect 23020 15648 23072 15700
rect 25504 15648 25556 15700
rect 20812 15580 20864 15632
rect 23664 15580 23716 15632
rect 26976 15580 27028 15632
rect 27160 15648 27212 15700
rect 28172 15580 28224 15632
rect 17776 15444 17828 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 19892 15444 19944 15496
rect 15384 15308 15436 15360
rect 16488 15308 16540 15360
rect 17224 15351 17276 15360
rect 17224 15317 17233 15351
rect 17233 15317 17267 15351
rect 17267 15317 17276 15351
rect 17224 15308 17276 15317
rect 18420 15308 18472 15360
rect 18788 15308 18840 15360
rect 20168 15376 20220 15428
rect 20720 15444 20772 15496
rect 22284 15512 22336 15564
rect 22468 15512 22520 15564
rect 23296 15555 23348 15564
rect 23296 15521 23305 15555
rect 23305 15521 23339 15555
rect 23339 15521 23348 15555
rect 23296 15512 23348 15521
rect 23388 15555 23440 15564
rect 23388 15521 23397 15555
rect 23397 15521 23431 15555
rect 23431 15521 23440 15555
rect 23388 15512 23440 15521
rect 22100 15444 22152 15496
rect 26608 15512 26660 15564
rect 20996 15376 21048 15428
rect 22008 15376 22060 15428
rect 22376 15376 22428 15428
rect 20444 15308 20496 15360
rect 23480 15308 23532 15360
rect 25320 15444 25372 15496
rect 24032 15419 24084 15428
rect 24032 15385 24041 15419
rect 24041 15385 24075 15419
rect 24075 15385 24084 15419
rect 24032 15376 24084 15385
rect 26332 15376 26384 15428
rect 26424 15376 26476 15428
rect 27620 15512 27672 15564
rect 27804 15512 27856 15564
rect 28908 15648 28960 15700
rect 29000 15580 29052 15632
rect 28172 15487 28224 15496
rect 28172 15453 28181 15487
rect 28181 15453 28215 15487
rect 28215 15453 28224 15487
rect 28172 15444 28224 15453
rect 28448 15444 28500 15496
rect 29092 15444 29144 15496
rect 29736 15648 29788 15700
rect 30656 15691 30708 15700
rect 30656 15657 30665 15691
rect 30665 15657 30699 15691
rect 30699 15657 30708 15691
rect 30656 15648 30708 15657
rect 33140 15648 33192 15700
rect 33416 15648 33468 15700
rect 37924 15691 37976 15700
rect 37924 15657 37933 15691
rect 37933 15657 37967 15691
rect 37967 15657 37976 15691
rect 37924 15648 37976 15657
rect 38292 15691 38344 15700
rect 38292 15657 38301 15691
rect 38301 15657 38335 15691
rect 38335 15657 38344 15691
rect 38292 15648 38344 15657
rect 40500 15648 40552 15700
rect 40684 15648 40736 15700
rect 32220 15580 32272 15632
rect 32864 15580 32916 15632
rect 30656 15512 30708 15564
rect 30932 15555 30984 15564
rect 30932 15521 30941 15555
rect 30941 15521 30975 15555
rect 30975 15521 30984 15555
rect 30932 15512 30984 15521
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 29644 15487 29696 15496
rect 29644 15453 29653 15487
rect 29653 15453 29687 15487
rect 29687 15453 29696 15487
rect 29644 15444 29696 15453
rect 29736 15444 29788 15496
rect 30104 15444 30156 15496
rect 32312 15444 32364 15496
rect 24860 15308 24912 15360
rect 25320 15308 25372 15360
rect 25504 15308 25556 15360
rect 25780 15308 25832 15360
rect 26516 15308 26568 15360
rect 27160 15308 27212 15360
rect 28816 15308 28868 15360
rect 29736 15308 29788 15360
rect 30196 15376 30248 15428
rect 30472 15419 30524 15428
rect 30472 15385 30481 15419
rect 30481 15385 30515 15419
rect 30515 15385 30524 15419
rect 30472 15376 30524 15385
rect 30380 15308 30432 15360
rect 31852 15308 31904 15360
rect 32588 15308 32640 15360
rect 32772 15308 32824 15360
rect 33324 15444 33376 15496
rect 35348 15512 35400 15564
rect 36636 15512 36688 15564
rect 37188 15512 37240 15564
rect 38936 15580 38988 15632
rect 40776 15580 40828 15632
rect 42248 15580 42300 15632
rect 41420 15512 41472 15564
rect 42064 15512 42116 15564
rect 42708 15555 42760 15564
rect 42708 15521 42717 15555
rect 42717 15521 42751 15555
rect 42751 15521 42760 15555
rect 42708 15512 42760 15521
rect 33876 15487 33928 15496
rect 33876 15453 33885 15487
rect 33885 15453 33919 15487
rect 33919 15453 33928 15487
rect 33876 15444 33928 15453
rect 34060 15487 34112 15496
rect 34060 15453 34069 15487
rect 34069 15453 34103 15487
rect 34103 15453 34112 15487
rect 34060 15444 34112 15453
rect 38200 15444 38252 15496
rect 38752 15444 38804 15496
rect 39120 15444 39172 15496
rect 36452 15376 36504 15428
rect 37556 15376 37608 15428
rect 40040 15376 40092 15428
rect 34704 15308 34756 15360
rect 35808 15351 35860 15360
rect 35808 15317 35817 15351
rect 35817 15317 35851 15351
rect 35851 15317 35860 15351
rect 35808 15308 35860 15317
rect 37648 15351 37700 15360
rect 37648 15317 37657 15351
rect 37657 15317 37691 15351
rect 37691 15317 37700 15351
rect 37648 15308 37700 15317
rect 38108 15351 38160 15360
rect 38108 15317 38117 15351
rect 38117 15317 38151 15351
rect 38151 15317 38160 15351
rect 38108 15308 38160 15317
rect 39120 15308 39172 15360
rect 39856 15308 39908 15360
rect 41052 15351 41104 15360
rect 41052 15317 41061 15351
rect 41061 15317 41095 15351
rect 41095 15317 41104 15351
rect 41052 15308 41104 15317
rect 41696 15487 41748 15496
rect 41696 15453 41705 15487
rect 41705 15453 41739 15487
rect 41739 15453 41748 15487
rect 41696 15444 41748 15453
rect 42800 15444 42852 15496
rect 43444 15444 43496 15496
rect 45008 15444 45060 15496
rect 41512 15308 41564 15360
rect 41604 15308 41656 15360
rect 42616 15351 42668 15360
rect 42616 15317 42625 15351
rect 42625 15317 42659 15351
rect 42659 15317 42668 15351
rect 42616 15308 42668 15317
rect 42984 15351 43036 15360
rect 42984 15317 42993 15351
rect 42993 15317 43027 15351
rect 43027 15317 43036 15351
rect 42984 15308 43036 15317
rect 43076 15308 43128 15360
rect 43904 15351 43956 15360
rect 43904 15317 43913 15351
rect 43913 15317 43947 15351
rect 43947 15317 43956 15351
rect 43904 15308 43956 15317
rect 44364 15308 44416 15360
rect 6070 15206 6122 15258
rect 6134 15206 6186 15258
rect 6198 15206 6250 15258
rect 6262 15206 6314 15258
rect 6326 15206 6378 15258
rect 11070 15206 11122 15258
rect 11134 15206 11186 15258
rect 11198 15206 11250 15258
rect 11262 15206 11314 15258
rect 11326 15206 11378 15258
rect 16070 15206 16122 15258
rect 16134 15206 16186 15258
rect 16198 15206 16250 15258
rect 16262 15206 16314 15258
rect 16326 15206 16378 15258
rect 21070 15206 21122 15258
rect 21134 15206 21186 15258
rect 21198 15206 21250 15258
rect 21262 15206 21314 15258
rect 21326 15206 21378 15258
rect 26070 15206 26122 15258
rect 26134 15206 26186 15258
rect 26198 15206 26250 15258
rect 26262 15206 26314 15258
rect 26326 15206 26378 15258
rect 31070 15206 31122 15258
rect 31134 15206 31186 15258
rect 31198 15206 31250 15258
rect 31262 15206 31314 15258
rect 31326 15206 31378 15258
rect 36070 15206 36122 15258
rect 36134 15206 36186 15258
rect 36198 15206 36250 15258
rect 36262 15206 36314 15258
rect 36326 15206 36378 15258
rect 41070 15206 41122 15258
rect 41134 15206 41186 15258
rect 41198 15206 41250 15258
rect 41262 15206 41314 15258
rect 41326 15206 41378 15258
rect 4344 15147 4396 15156
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 9772 15104 9824 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10324 15104 10376 15156
rect 6644 15036 6696 15088
rect 8300 15036 8352 15088
rect 940 15011 992 15020
rect 940 14977 949 15011
rect 949 14977 983 15011
rect 983 14977 992 15011
rect 940 14968 992 14977
rect 4528 14968 4580 15020
rect 4896 14968 4948 15020
rect 11612 15104 11664 15156
rect 13268 15104 13320 15156
rect 14556 15104 14608 15156
rect 14832 15104 14884 15156
rect 18236 15104 18288 15156
rect 12808 15036 12860 15088
rect 4804 14900 4856 14952
rect 5632 14900 5684 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 8116 14900 8168 14952
rect 9036 14900 9088 14952
rect 756 14807 808 14816
rect 756 14773 765 14807
rect 765 14773 799 14807
rect 799 14773 808 14807
rect 756 14764 808 14773
rect 4620 14764 4672 14816
rect 5448 14807 5500 14816
rect 5448 14773 5457 14807
rect 5457 14773 5491 14807
rect 5491 14773 5500 14807
rect 5448 14764 5500 14773
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 11428 15011 11480 15020
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 14096 14968 14148 15020
rect 14188 14968 14240 15020
rect 12348 14900 12400 14952
rect 15752 14943 15804 14952
rect 15752 14909 15761 14943
rect 15761 14909 15795 14943
rect 15795 14909 15804 14943
rect 15752 14900 15804 14909
rect 16212 14968 16264 15020
rect 16488 14968 16540 15020
rect 16856 15036 16908 15088
rect 17132 15079 17184 15088
rect 17132 15045 17157 15079
rect 17157 15045 17184 15079
rect 17500 15079 17552 15088
rect 17132 15036 17184 15045
rect 17500 15045 17509 15079
rect 17509 15045 17543 15079
rect 17543 15045 17552 15079
rect 17500 15036 17552 15045
rect 22652 15104 22704 15156
rect 19984 14968 20036 15020
rect 20076 14968 20128 15020
rect 23388 15104 23440 15156
rect 23664 15104 23716 15156
rect 23940 15104 23992 15156
rect 24032 15104 24084 15156
rect 24400 15104 24452 15156
rect 25228 15104 25280 15156
rect 25412 15104 25464 15156
rect 26516 15104 26568 15156
rect 26608 15147 26660 15156
rect 26608 15113 26617 15147
rect 26617 15113 26651 15147
rect 26651 15113 26660 15147
rect 26608 15104 26660 15113
rect 20720 14968 20772 15020
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 17960 14900 18012 14952
rect 18420 14832 18472 14884
rect 20904 14968 20956 15020
rect 21456 14968 21508 15020
rect 21548 15011 21600 15020
rect 21548 14977 21557 15011
rect 21557 14977 21591 15011
rect 21591 14977 21600 15011
rect 21548 14968 21600 14977
rect 22192 14968 22244 15020
rect 21180 14900 21232 14952
rect 21916 14832 21968 14884
rect 22560 14900 22612 14952
rect 23388 15011 23440 15020
rect 23388 14977 23397 15011
rect 23397 14977 23431 15011
rect 23431 14977 23440 15011
rect 23388 14968 23440 14977
rect 22468 14832 22520 14884
rect 24400 14968 24452 15020
rect 25780 15036 25832 15088
rect 26792 15104 26844 15156
rect 27160 15104 27212 15156
rect 29368 15104 29420 15156
rect 30012 15104 30064 15156
rect 30472 15104 30524 15156
rect 30656 15147 30708 15156
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 24216 14900 24268 14952
rect 24768 14900 24820 14952
rect 24124 14832 24176 14884
rect 25412 14900 25464 14952
rect 25688 14943 25740 14952
rect 25688 14909 25697 14943
rect 25697 14909 25731 14943
rect 25731 14909 25740 14943
rect 25688 14900 25740 14909
rect 8208 14764 8260 14816
rect 10048 14764 10100 14816
rect 11888 14764 11940 14816
rect 13268 14764 13320 14816
rect 14372 14764 14424 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15844 14764 15896 14816
rect 16672 14764 16724 14816
rect 17040 14764 17092 14816
rect 17592 14764 17644 14816
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 18788 14764 18840 14816
rect 19432 14764 19484 14816
rect 19892 14764 19944 14816
rect 20168 14807 20220 14816
rect 20168 14773 20177 14807
rect 20177 14773 20211 14807
rect 20211 14773 20220 14807
rect 20168 14764 20220 14773
rect 20444 14764 20496 14816
rect 20996 14764 21048 14816
rect 22836 14764 22888 14816
rect 23940 14764 23992 14816
rect 24492 14764 24544 14816
rect 24860 14807 24912 14816
rect 24860 14773 24869 14807
rect 24869 14773 24903 14807
rect 24903 14773 24912 14807
rect 24860 14764 24912 14773
rect 26240 14968 26292 15020
rect 26608 14900 26660 14952
rect 27068 15011 27120 15020
rect 27068 14977 27077 15011
rect 27077 14977 27111 15011
rect 27111 14977 27120 15011
rect 27068 14968 27120 14977
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 30288 15079 30340 15088
rect 30288 15045 30297 15079
rect 30297 15045 30331 15079
rect 30331 15045 30340 15079
rect 30288 15036 30340 15045
rect 31024 15036 31076 15088
rect 28264 15011 28316 15020
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 29644 14968 29696 15020
rect 26884 14900 26936 14952
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 25412 14764 25464 14816
rect 25964 14807 26016 14816
rect 25964 14773 25973 14807
rect 25973 14773 26007 14807
rect 26007 14773 26016 14807
rect 25964 14764 26016 14773
rect 26424 14764 26476 14816
rect 26884 14807 26936 14816
rect 26884 14773 26893 14807
rect 26893 14773 26927 14807
rect 26927 14773 26936 14807
rect 26884 14764 26936 14773
rect 27528 14807 27580 14816
rect 27528 14773 27537 14807
rect 27537 14773 27571 14807
rect 27571 14773 27580 14807
rect 27528 14764 27580 14773
rect 28172 14764 28224 14816
rect 29920 14968 29972 15020
rect 32680 15147 32732 15156
rect 32680 15113 32689 15147
rect 32689 15113 32723 15147
rect 32723 15113 32732 15147
rect 32680 15104 32732 15113
rect 33876 15104 33928 15156
rect 35072 15104 35124 15156
rect 35348 15104 35400 15156
rect 35808 15104 35860 15156
rect 36452 15104 36504 15156
rect 37648 15104 37700 15156
rect 38660 15104 38712 15156
rect 32220 15079 32272 15088
rect 32220 15045 32229 15079
rect 32229 15045 32263 15079
rect 32263 15045 32272 15079
rect 32220 15036 32272 15045
rect 32588 15036 32640 15088
rect 34060 15036 34112 15088
rect 35440 15036 35492 15088
rect 30196 14900 30248 14952
rect 32036 14968 32088 15020
rect 32864 15011 32916 15020
rect 30656 14900 30708 14952
rect 32864 14977 32873 15011
rect 32873 14977 32907 15011
rect 32907 14977 32916 15011
rect 32864 14968 32916 14977
rect 32956 15011 33008 15020
rect 32956 14977 32965 15011
rect 32965 14977 32999 15011
rect 32999 14977 33008 15011
rect 32956 14968 33008 14977
rect 33140 15011 33192 15020
rect 33140 14977 33149 15011
rect 33149 14977 33183 15011
rect 33183 14977 33192 15011
rect 33140 14968 33192 14977
rect 33232 14968 33284 15020
rect 32496 14943 32548 14952
rect 32496 14909 32505 14943
rect 32505 14909 32539 14943
rect 32539 14909 32548 14943
rect 32496 14900 32548 14909
rect 32680 14900 32732 14952
rect 33324 14900 33376 14952
rect 34152 14900 34204 14952
rect 31760 14875 31812 14884
rect 31760 14841 31769 14875
rect 31769 14841 31803 14875
rect 31803 14841 31812 14875
rect 31760 14832 31812 14841
rect 32588 14832 32640 14884
rect 37556 15036 37608 15088
rect 38200 15036 38252 15088
rect 39396 15079 39448 15088
rect 39396 15045 39405 15079
rect 39405 15045 39439 15079
rect 39439 15045 39448 15079
rect 39396 15036 39448 15045
rect 30564 14764 30616 14816
rect 31208 14764 31260 14816
rect 32772 14764 32824 14816
rect 33048 14764 33100 14816
rect 35072 14900 35124 14952
rect 37740 14968 37792 15020
rect 39212 14968 39264 15020
rect 39672 14968 39724 15020
rect 40960 15104 41012 15156
rect 40224 15036 40276 15088
rect 41604 15036 41656 15088
rect 42984 15104 43036 15156
rect 37188 14943 37240 14952
rect 37188 14909 37197 14943
rect 37197 14909 37231 14943
rect 37231 14909 37240 14943
rect 37188 14900 37240 14909
rect 39028 14900 39080 14952
rect 36820 14832 36872 14884
rect 41788 14943 41840 14952
rect 41788 14909 41797 14943
rect 41797 14909 41831 14943
rect 41831 14909 41840 14943
rect 41788 14900 41840 14909
rect 41236 14832 41288 14884
rect 45192 15011 45244 15020
rect 45192 14977 45201 15011
rect 45201 14977 45235 15011
rect 45235 14977 45244 15011
rect 45192 14968 45244 14977
rect 36912 14764 36964 14816
rect 37280 14764 37332 14816
rect 38660 14764 38712 14816
rect 38936 14807 38988 14816
rect 38936 14773 38945 14807
rect 38945 14773 38979 14807
rect 38979 14773 38988 14807
rect 38936 14764 38988 14773
rect 39212 14764 39264 14816
rect 40776 14764 40828 14816
rect 41144 14764 41196 14816
rect 41420 14764 41472 14816
rect 41512 14764 41564 14816
rect 42616 14764 42668 14816
rect 43904 14807 43956 14816
rect 43904 14773 43913 14807
rect 43913 14773 43947 14807
rect 43947 14773 43956 14807
rect 43904 14764 43956 14773
rect 44364 14764 44416 14816
rect 45008 14807 45060 14816
rect 45008 14773 45017 14807
rect 45017 14773 45051 14807
rect 45051 14773 45060 14807
rect 45008 14764 45060 14773
rect 3570 14662 3622 14714
rect 3634 14662 3686 14714
rect 3698 14662 3750 14714
rect 3762 14662 3814 14714
rect 3826 14662 3878 14714
rect 8570 14662 8622 14714
rect 8634 14662 8686 14714
rect 8698 14662 8750 14714
rect 8762 14662 8814 14714
rect 8826 14662 8878 14714
rect 13570 14662 13622 14714
rect 13634 14662 13686 14714
rect 13698 14662 13750 14714
rect 13762 14662 13814 14714
rect 13826 14662 13878 14714
rect 18570 14662 18622 14714
rect 18634 14662 18686 14714
rect 18698 14662 18750 14714
rect 18762 14662 18814 14714
rect 18826 14662 18878 14714
rect 23570 14662 23622 14714
rect 23634 14662 23686 14714
rect 23698 14662 23750 14714
rect 23762 14662 23814 14714
rect 23826 14662 23878 14714
rect 28570 14662 28622 14714
rect 28634 14662 28686 14714
rect 28698 14662 28750 14714
rect 28762 14662 28814 14714
rect 28826 14662 28878 14714
rect 33570 14662 33622 14714
rect 33634 14662 33686 14714
rect 33698 14662 33750 14714
rect 33762 14662 33814 14714
rect 33826 14662 33878 14714
rect 38570 14662 38622 14714
rect 38634 14662 38686 14714
rect 38698 14662 38750 14714
rect 38762 14662 38814 14714
rect 38826 14662 38878 14714
rect 43570 14662 43622 14714
rect 43634 14662 43686 14714
rect 43698 14662 43750 14714
rect 43762 14662 43814 14714
rect 43826 14662 43878 14714
rect 4344 14560 4396 14612
rect 4804 14560 4856 14612
rect 5632 14560 5684 14612
rect 9680 14560 9732 14612
rect 6644 14492 6696 14544
rect 7748 14492 7800 14544
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 4896 14424 4948 14476
rect 5724 14424 5776 14476
rect 8208 14424 8260 14476
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 9588 14356 9640 14408
rect 9772 14424 9824 14476
rect 10048 14424 10100 14476
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 9864 14288 9916 14340
rect 10324 14356 10376 14408
rect 13084 14560 13136 14612
rect 13544 14560 13596 14612
rect 15752 14560 15804 14612
rect 16948 14560 17000 14612
rect 17776 14560 17828 14612
rect 18420 14560 18472 14612
rect 18696 14560 18748 14612
rect 19248 14560 19300 14612
rect 12348 14424 12400 14476
rect 14832 14424 14884 14476
rect 11888 14331 11940 14340
rect 11888 14297 11897 14331
rect 11897 14297 11931 14331
rect 11931 14297 11940 14331
rect 11888 14288 11940 14297
rect 14004 14288 14056 14340
rect 15108 14492 15160 14544
rect 16396 14492 16448 14544
rect 19616 14492 19668 14544
rect 20076 14560 20128 14612
rect 20444 14560 20496 14612
rect 21272 14560 21324 14612
rect 21548 14560 21600 14612
rect 23204 14560 23256 14612
rect 19892 14492 19944 14544
rect 21456 14492 21508 14544
rect 22744 14492 22796 14544
rect 23756 14535 23808 14544
rect 23756 14501 23765 14535
rect 23765 14501 23799 14535
rect 23799 14501 23808 14535
rect 23756 14492 23808 14501
rect 23940 14492 23992 14544
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 24860 14560 24912 14612
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 16856 14424 16908 14476
rect 22192 14424 22244 14476
rect 25228 14492 25280 14544
rect 27068 14560 27120 14612
rect 28264 14560 28316 14612
rect 28356 14560 28408 14612
rect 14740 14288 14792 14340
rect 17684 14356 17736 14408
rect 18236 14356 18288 14408
rect 18696 14356 18748 14408
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 18972 14399 19024 14408
rect 18972 14365 18981 14399
rect 18981 14365 19015 14399
rect 19015 14365 19024 14399
rect 18972 14356 19024 14365
rect 19064 14356 19116 14408
rect 19248 14356 19300 14408
rect 19708 14356 19760 14408
rect 8392 14220 8444 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 10140 14220 10192 14272
rect 10692 14263 10744 14272
rect 10692 14229 10701 14263
rect 10701 14229 10735 14263
rect 10735 14229 10744 14263
rect 10692 14220 10744 14229
rect 11428 14220 11480 14272
rect 11520 14220 11572 14272
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 13544 14220 13596 14272
rect 13912 14263 13964 14272
rect 13912 14229 13921 14263
rect 13921 14229 13955 14263
rect 13955 14229 13964 14263
rect 13912 14220 13964 14229
rect 14188 14220 14240 14272
rect 14556 14220 14608 14272
rect 15660 14288 15712 14340
rect 16856 14288 16908 14340
rect 17868 14288 17920 14340
rect 17776 14263 17828 14272
rect 17776 14229 17785 14263
rect 17785 14229 17819 14263
rect 17819 14229 17828 14263
rect 17776 14220 17828 14229
rect 18328 14220 18380 14272
rect 18696 14220 18748 14272
rect 19340 14331 19392 14340
rect 19340 14297 19349 14331
rect 19349 14297 19383 14331
rect 19383 14297 19392 14331
rect 19340 14288 19392 14297
rect 19432 14288 19484 14340
rect 20168 14356 20220 14408
rect 21180 14356 21232 14408
rect 19892 14220 19944 14272
rect 21272 14288 21324 14340
rect 21456 14356 21508 14408
rect 21916 14356 21968 14408
rect 22652 14356 22704 14408
rect 22928 14356 22980 14408
rect 23940 14399 23992 14408
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 26700 14424 26752 14476
rect 27160 14424 27212 14476
rect 27804 14467 27856 14476
rect 27804 14433 27813 14467
rect 27813 14433 27847 14467
rect 27847 14433 27856 14467
rect 27804 14424 27856 14433
rect 29092 14560 29144 14612
rect 29276 14560 29328 14612
rect 24216 14399 24268 14408
rect 24216 14365 24225 14399
rect 24225 14365 24259 14399
rect 24259 14365 24268 14399
rect 24216 14356 24268 14365
rect 20352 14220 20404 14272
rect 21916 14220 21968 14272
rect 22008 14263 22060 14272
rect 22008 14229 22017 14263
rect 22017 14229 22051 14263
rect 22051 14229 22060 14263
rect 22008 14220 22060 14229
rect 22284 14220 22336 14272
rect 23296 14220 23348 14272
rect 24032 14220 24084 14272
rect 25412 14399 25464 14408
rect 25412 14365 25421 14399
rect 25421 14365 25455 14399
rect 25455 14365 25464 14399
rect 25412 14356 25464 14365
rect 26792 14356 26844 14408
rect 26976 14356 27028 14408
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 29000 14356 29052 14408
rect 30748 14560 30800 14612
rect 30656 14424 30708 14476
rect 31116 14492 31168 14544
rect 31300 14560 31352 14612
rect 31668 14560 31720 14612
rect 32128 14560 32180 14612
rect 32496 14560 32548 14612
rect 35624 14560 35676 14612
rect 36636 14603 36688 14612
rect 36636 14569 36645 14603
rect 36645 14569 36679 14603
rect 36679 14569 36688 14603
rect 36636 14560 36688 14569
rect 37096 14560 37148 14612
rect 40132 14560 40184 14612
rect 42800 14560 42852 14612
rect 31484 14492 31536 14544
rect 32956 14535 33008 14544
rect 32956 14501 32965 14535
rect 32965 14501 32999 14535
rect 32999 14501 33008 14535
rect 32956 14492 33008 14501
rect 33324 14535 33376 14544
rect 33324 14501 33333 14535
rect 33333 14501 33367 14535
rect 33367 14501 33376 14535
rect 33324 14492 33376 14501
rect 33508 14492 33560 14544
rect 34336 14492 34388 14544
rect 32956 14356 33008 14408
rect 35532 14492 35584 14544
rect 25228 14220 25280 14272
rect 25688 14220 25740 14272
rect 26608 14220 26660 14272
rect 27436 14288 27488 14340
rect 30840 14288 30892 14340
rect 31024 14288 31076 14340
rect 32128 14288 32180 14340
rect 33692 14356 33744 14408
rect 33784 14399 33836 14408
rect 33784 14365 33793 14399
rect 33793 14365 33827 14399
rect 33827 14365 33836 14399
rect 33784 14356 33836 14365
rect 34888 14399 34940 14408
rect 34888 14365 34897 14399
rect 34897 14365 34931 14399
rect 34931 14365 34940 14399
rect 34888 14356 34940 14365
rect 35164 14356 35216 14408
rect 35716 14467 35768 14476
rect 35716 14433 35725 14467
rect 35725 14433 35759 14467
rect 35759 14433 35768 14467
rect 35716 14424 35768 14433
rect 35808 14424 35860 14476
rect 36544 14424 36596 14476
rect 35992 14356 36044 14408
rect 39028 14424 39080 14476
rect 41420 14492 41472 14544
rect 44272 14560 44324 14612
rect 39856 14424 39908 14476
rect 40040 14424 40092 14476
rect 40960 14467 41012 14476
rect 40960 14433 40969 14467
rect 40969 14433 41003 14467
rect 41003 14433 41012 14467
rect 40960 14424 41012 14433
rect 41880 14424 41932 14476
rect 38016 14399 38068 14408
rect 38016 14365 38025 14399
rect 38025 14365 38059 14399
rect 38059 14365 38068 14399
rect 38016 14356 38068 14365
rect 38108 14356 38160 14408
rect 38476 14356 38528 14408
rect 38844 14356 38896 14408
rect 42616 14356 42668 14408
rect 34980 14288 35032 14340
rect 35808 14331 35860 14340
rect 35808 14297 35842 14331
rect 35842 14297 35860 14331
rect 35808 14288 35860 14297
rect 28080 14263 28132 14272
rect 28080 14229 28089 14263
rect 28089 14229 28123 14263
rect 28123 14229 28132 14263
rect 28080 14220 28132 14229
rect 28908 14220 28960 14272
rect 29000 14220 29052 14272
rect 30288 14263 30340 14272
rect 30288 14229 30297 14263
rect 30297 14229 30331 14263
rect 30331 14229 30340 14263
rect 30288 14220 30340 14229
rect 30564 14263 30616 14272
rect 30564 14229 30573 14263
rect 30573 14229 30607 14263
rect 30607 14229 30616 14263
rect 30564 14220 30616 14229
rect 30932 14220 30984 14272
rect 32404 14220 32456 14272
rect 33968 14220 34020 14272
rect 35072 14263 35124 14272
rect 35072 14229 35081 14263
rect 35081 14229 35115 14263
rect 35115 14229 35124 14263
rect 35072 14220 35124 14229
rect 35716 14220 35768 14272
rect 36452 14220 36504 14272
rect 37372 14263 37424 14272
rect 37372 14229 37381 14263
rect 37381 14229 37415 14263
rect 37415 14229 37424 14263
rect 37372 14220 37424 14229
rect 37556 14263 37608 14272
rect 37556 14229 37565 14263
rect 37565 14229 37599 14263
rect 37599 14229 37608 14263
rect 37556 14220 37608 14229
rect 37832 14263 37884 14272
rect 37832 14229 37841 14263
rect 37841 14229 37875 14263
rect 37875 14229 37884 14263
rect 37832 14220 37884 14229
rect 39120 14220 39172 14272
rect 39488 14331 39540 14340
rect 39488 14297 39497 14331
rect 39497 14297 39531 14331
rect 39531 14297 39540 14331
rect 39488 14288 39540 14297
rect 40224 14288 40276 14340
rect 44180 14288 44232 14340
rect 39764 14220 39816 14272
rect 40868 14220 40920 14272
rect 41236 14263 41288 14272
rect 41236 14229 41245 14263
rect 41245 14229 41279 14263
rect 41279 14229 41288 14263
rect 41236 14220 41288 14229
rect 41512 14220 41564 14272
rect 42800 14263 42852 14272
rect 42800 14229 42809 14263
rect 42809 14229 42843 14263
rect 42843 14229 42852 14263
rect 42800 14220 42852 14229
rect 43076 14263 43128 14272
rect 43076 14229 43085 14263
rect 43085 14229 43119 14263
rect 43119 14229 43128 14263
rect 43076 14220 43128 14229
rect 43444 14263 43496 14272
rect 43444 14229 43453 14263
rect 43453 14229 43487 14263
rect 43487 14229 43496 14263
rect 43444 14220 43496 14229
rect 44364 14220 44416 14272
rect 44732 14220 44784 14272
rect 6070 14118 6122 14170
rect 6134 14118 6186 14170
rect 6198 14118 6250 14170
rect 6262 14118 6314 14170
rect 6326 14118 6378 14170
rect 11070 14118 11122 14170
rect 11134 14118 11186 14170
rect 11198 14118 11250 14170
rect 11262 14118 11314 14170
rect 11326 14118 11378 14170
rect 16070 14118 16122 14170
rect 16134 14118 16186 14170
rect 16198 14118 16250 14170
rect 16262 14118 16314 14170
rect 16326 14118 16378 14170
rect 21070 14118 21122 14170
rect 21134 14118 21186 14170
rect 21198 14118 21250 14170
rect 21262 14118 21314 14170
rect 21326 14118 21378 14170
rect 26070 14118 26122 14170
rect 26134 14118 26186 14170
rect 26198 14118 26250 14170
rect 26262 14118 26314 14170
rect 26326 14118 26378 14170
rect 31070 14118 31122 14170
rect 31134 14118 31186 14170
rect 31198 14118 31250 14170
rect 31262 14118 31314 14170
rect 31326 14118 31378 14170
rect 36070 14118 36122 14170
rect 36134 14118 36186 14170
rect 36198 14118 36250 14170
rect 36262 14118 36314 14170
rect 36326 14118 36378 14170
rect 41070 14118 41122 14170
rect 41134 14118 41186 14170
rect 41198 14118 41250 14170
rect 41262 14118 41314 14170
rect 41326 14118 41378 14170
rect 756 13744 808 13796
rect 6644 14016 6696 14068
rect 8116 14016 8168 14068
rect 4344 13948 4396 14000
rect 10048 14016 10100 14068
rect 10692 14016 10744 14068
rect 8392 13948 8444 14000
rect 3424 13812 3476 13864
rect 3792 13855 3844 13864
rect 3792 13821 3801 13855
rect 3801 13821 3835 13855
rect 3835 13821 3844 13855
rect 3792 13812 3844 13821
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 9588 13880 9640 13932
rect 10140 13880 10192 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 13360 14016 13412 14068
rect 13544 14016 13596 14068
rect 14004 14016 14056 14068
rect 9772 13812 9824 13864
rect 13636 13948 13688 14000
rect 14740 13948 14792 14000
rect 15108 13991 15160 14000
rect 15108 13957 15117 13991
rect 15117 13957 15151 13991
rect 15151 13957 15160 13991
rect 15108 13948 15160 13957
rect 18420 14016 18472 14068
rect 18788 14016 18840 14068
rect 19984 14016 20036 14068
rect 18236 13948 18288 14000
rect 18696 13948 18748 14000
rect 19156 13948 19208 14000
rect 11336 13812 11388 13864
rect 13912 13812 13964 13864
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 17316 13880 17368 13932
rect 14832 13812 14884 13864
rect 16580 13855 16632 13864
rect 16580 13821 16589 13855
rect 16589 13821 16623 13855
rect 16623 13821 16632 13855
rect 16580 13812 16632 13821
rect 16672 13812 16724 13864
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 18144 13880 18196 13932
rect 17960 13812 18012 13864
rect 20996 13948 21048 14000
rect 24124 14016 24176 14068
rect 24676 14016 24728 14068
rect 23756 13948 23808 14000
rect 26700 14016 26752 14068
rect 26884 14016 26936 14068
rect 27160 14016 27212 14068
rect 20536 13812 20588 13864
rect 19708 13744 19760 13796
rect 22100 13880 22152 13932
rect 21548 13812 21600 13864
rect 22468 13880 22520 13932
rect 22652 13923 22704 13932
rect 22652 13889 22661 13923
rect 22661 13889 22695 13923
rect 22695 13889 22704 13923
rect 22652 13880 22704 13889
rect 23112 13923 23164 13932
rect 23112 13889 23121 13923
rect 23121 13889 23155 13923
rect 23155 13889 23164 13923
rect 23112 13880 23164 13889
rect 23204 13880 23256 13932
rect 22192 13787 22244 13796
rect 22192 13753 22201 13787
rect 22201 13753 22235 13787
rect 22235 13753 22244 13787
rect 22192 13744 22244 13753
rect 4252 13676 4304 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 12440 13676 12492 13728
rect 14188 13676 14240 13728
rect 15568 13719 15620 13728
rect 15568 13685 15577 13719
rect 15577 13685 15611 13719
rect 15611 13685 15620 13719
rect 15568 13676 15620 13685
rect 16488 13719 16540 13728
rect 16488 13685 16497 13719
rect 16497 13685 16531 13719
rect 16531 13685 16540 13719
rect 16488 13676 16540 13685
rect 17592 13676 17644 13728
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 20444 13676 20496 13728
rect 22928 13812 22980 13864
rect 23480 13880 23532 13932
rect 23940 13880 23992 13932
rect 28172 14059 28224 14068
rect 28172 14025 28181 14059
rect 28181 14025 28215 14059
rect 28215 14025 28224 14059
rect 28172 14016 28224 14025
rect 28356 14016 28408 14068
rect 28448 14016 28500 14068
rect 29000 14059 29052 14068
rect 29000 14025 29009 14059
rect 29009 14025 29043 14059
rect 29043 14025 29052 14059
rect 29000 14016 29052 14025
rect 30472 14016 30524 14068
rect 29736 13948 29788 14000
rect 29920 13948 29972 14000
rect 31392 13948 31444 14000
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 24124 13744 24176 13796
rect 24952 13744 25004 13796
rect 27068 13880 27120 13932
rect 28448 13880 28500 13932
rect 29000 13880 29052 13932
rect 29092 13880 29144 13932
rect 30840 13880 30892 13932
rect 31484 13880 31536 13932
rect 24768 13676 24820 13728
rect 25136 13719 25188 13728
rect 25136 13685 25145 13719
rect 25145 13685 25179 13719
rect 25179 13685 25188 13719
rect 25136 13676 25188 13685
rect 25320 13719 25372 13728
rect 25320 13685 25329 13719
rect 25329 13685 25363 13719
rect 25363 13685 25372 13719
rect 25320 13676 25372 13685
rect 25412 13676 25464 13728
rect 27804 13812 27856 13864
rect 27344 13744 27396 13796
rect 28172 13744 28224 13796
rect 28816 13744 28868 13796
rect 32588 14016 32640 14068
rect 32864 14016 32916 14068
rect 32496 13948 32548 14000
rect 33324 14016 33376 14068
rect 33784 14016 33836 14068
rect 35992 14016 36044 14068
rect 36544 14016 36596 14068
rect 36912 14016 36964 14068
rect 38476 14016 38528 14068
rect 39488 14016 39540 14068
rect 32588 13880 32640 13932
rect 33416 13948 33468 14000
rect 37832 13948 37884 14000
rect 38200 13948 38252 14000
rect 40224 13948 40276 14000
rect 35072 13923 35124 13932
rect 35072 13889 35081 13923
rect 35081 13889 35115 13923
rect 35115 13889 35124 13923
rect 35072 13880 35124 13889
rect 31944 13744 31996 13796
rect 34428 13812 34480 13864
rect 34796 13812 34848 13864
rect 35716 13812 35768 13864
rect 36360 13855 36412 13864
rect 36360 13821 36369 13855
rect 36369 13821 36403 13855
rect 36403 13821 36412 13855
rect 36360 13812 36412 13821
rect 30564 13676 30616 13728
rect 36544 13880 36596 13932
rect 37188 13923 37240 13932
rect 37188 13889 37197 13923
rect 37197 13889 37231 13923
rect 37231 13889 37240 13923
rect 37188 13880 37240 13889
rect 37280 13880 37332 13932
rect 40960 13880 41012 13932
rect 37096 13855 37148 13864
rect 37096 13821 37105 13855
rect 37105 13821 37139 13855
rect 37139 13821 37148 13855
rect 37096 13812 37148 13821
rect 39212 13812 39264 13864
rect 33232 13676 33284 13728
rect 33508 13676 33560 13728
rect 34428 13676 34480 13728
rect 38844 13744 38896 13796
rect 39580 13855 39632 13864
rect 39580 13821 39589 13855
rect 39589 13821 39623 13855
rect 39623 13821 39632 13855
rect 39580 13812 39632 13821
rect 39672 13812 39724 13864
rect 42248 14059 42300 14068
rect 42248 14025 42257 14059
rect 42257 14025 42291 14059
rect 42291 14025 42300 14059
rect 42248 14016 42300 14025
rect 34612 13719 34664 13728
rect 34612 13685 34621 13719
rect 34621 13685 34655 13719
rect 34655 13685 34664 13719
rect 34612 13676 34664 13685
rect 37280 13676 37332 13728
rect 37556 13676 37608 13728
rect 39212 13719 39264 13728
rect 39212 13685 39221 13719
rect 39221 13685 39255 13719
rect 39255 13685 39264 13719
rect 39212 13676 39264 13685
rect 39304 13676 39356 13728
rect 42800 13855 42852 13864
rect 42800 13821 42809 13855
rect 42809 13821 42843 13855
rect 42843 13821 42852 13855
rect 42800 13812 42852 13821
rect 43352 13744 43404 13796
rect 43904 13787 43956 13796
rect 43904 13753 43913 13787
rect 43913 13753 43947 13787
rect 43947 13753 43956 13787
rect 44732 13787 44784 13796
rect 43904 13744 43956 13753
rect 44732 13753 44741 13787
rect 44741 13753 44775 13787
rect 44775 13753 44784 13787
rect 44732 13744 44784 13753
rect 43076 13676 43128 13728
rect 44364 13676 44416 13728
rect 44548 13676 44600 13728
rect 3570 13574 3622 13626
rect 3634 13574 3686 13626
rect 3698 13574 3750 13626
rect 3762 13574 3814 13626
rect 3826 13574 3878 13626
rect 8570 13574 8622 13626
rect 8634 13574 8686 13626
rect 8698 13574 8750 13626
rect 8762 13574 8814 13626
rect 8826 13574 8878 13626
rect 13570 13574 13622 13626
rect 13634 13574 13686 13626
rect 13698 13574 13750 13626
rect 13762 13574 13814 13626
rect 13826 13574 13878 13626
rect 18570 13574 18622 13626
rect 18634 13574 18686 13626
rect 18698 13574 18750 13626
rect 18762 13574 18814 13626
rect 18826 13574 18878 13626
rect 23570 13574 23622 13626
rect 23634 13574 23686 13626
rect 23698 13574 23750 13626
rect 23762 13574 23814 13626
rect 23826 13574 23878 13626
rect 28570 13574 28622 13626
rect 28634 13574 28686 13626
rect 28698 13574 28750 13626
rect 28762 13574 28814 13626
rect 28826 13574 28878 13626
rect 33570 13574 33622 13626
rect 33634 13574 33686 13626
rect 33698 13574 33750 13626
rect 33762 13574 33814 13626
rect 33826 13574 33878 13626
rect 38570 13574 38622 13626
rect 38634 13574 38686 13626
rect 38698 13574 38750 13626
rect 38762 13574 38814 13626
rect 38826 13574 38878 13626
rect 43570 13574 43622 13626
rect 43634 13574 43686 13626
rect 43698 13574 43750 13626
rect 43762 13574 43814 13626
rect 43826 13574 43878 13626
rect 4252 13472 4304 13524
rect 5632 13472 5684 13524
rect 7012 13472 7064 13524
rect 10232 13472 10284 13524
rect 11428 13472 11480 13524
rect 12256 13472 12308 13524
rect 5264 13404 5316 13456
rect 9588 13404 9640 13456
rect 12900 13472 12952 13524
rect 17040 13472 17092 13524
rect 17960 13472 18012 13524
rect 18696 13472 18748 13524
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 5540 13268 5592 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 6920 13336 6972 13388
rect 10508 13336 10560 13388
rect 15660 13404 15712 13456
rect 14280 13336 14332 13388
rect 6184 13268 6236 13320
rect 9496 13268 9548 13320
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 11336 13268 11388 13320
rect 6644 13200 6696 13252
rect 3424 13132 3476 13141
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 9956 13200 10008 13252
rect 10140 13200 10192 13252
rect 11704 13243 11756 13252
rect 11704 13209 11713 13243
rect 11713 13209 11747 13243
rect 11747 13209 11756 13243
rect 11704 13200 11756 13209
rect 12164 13200 12216 13252
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 11520 13132 11572 13184
rect 11612 13132 11664 13184
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 19432 13472 19484 13524
rect 19984 13472 20036 13524
rect 20904 13472 20956 13524
rect 21916 13472 21968 13524
rect 18512 13336 18564 13388
rect 21916 13379 21968 13388
rect 16488 13268 16540 13320
rect 18696 13268 18748 13320
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 18972 13311 19024 13320
rect 18972 13277 18981 13311
rect 18981 13277 19015 13311
rect 19015 13277 19024 13311
rect 18972 13268 19024 13277
rect 14004 13200 14056 13252
rect 14372 13200 14424 13252
rect 19156 13200 19208 13252
rect 19248 13243 19300 13252
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 19340 13200 19392 13252
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22284 13404 22336 13456
rect 22560 13404 22612 13456
rect 23112 13472 23164 13524
rect 24032 13472 24084 13524
rect 24400 13472 24452 13524
rect 25504 13472 25556 13524
rect 26608 13515 26660 13524
rect 26608 13481 26617 13515
rect 26617 13481 26651 13515
rect 26651 13481 26660 13515
rect 26608 13472 26660 13481
rect 26884 13515 26936 13524
rect 26884 13481 26893 13515
rect 26893 13481 26927 13515
rect 26927 13481 26936 13515
rect 26884 13472 26936 13481
rect 27068 13515 27120 13524
rect 27068 13481 27077 13515
rect 27077 13481 27111 13515
rect 27111 13481 27120 13515
rect 27068 13472 27120 13481
rect 27160 13472 27212 13524
rect 28448 13472 28500 13524
rect 28724 13472 28776 13524
rect 29644 13515 29696 13524
rect 29644 13481 29653 13515
rect 29653 13481 29687 13515
rect 29687 13481 29696 13515
rect 29644 13472 29696 13481
rect 29828 13472 29880 13524
rect 31484 13472 31536 13524
rect 32220 13472 32272 13524
rect 32588 13515 32640 13524
rect 32588 13481 32597 13515
rect 32597 13481 32631 13515
rect 32631 13481 32640 13515
rect 32588 13472 32640 13481
rect 34520 13472 34572 13524
rect 24676 13404 24728 13456
rect 28356 13404 28408 13456
rect 22192 13311 22244 13320
rect 22192 13277 22195 13311
rect 22195 13277 22229 13311
rect 22229 13277 22244 13311
rect 18420 13132 18472 13184
rect 18696 13132 18748 13184
rect 19800 13132 19852 13184
rect 22192 13268 22244 13277
rect 22836 13268 22888 13320
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 23848 13311 23900 13320
rect 23848 13277 23857 13311
rect 23857 13277 23891 13311
rect 23891 13277 23900 13311
rect 23848 13268 23900 13277
rect 24584 13336 24636 13388
rect 24768 13336 24820 13388
rect 26424 13336 26476 13388
rect 26516 13336 26568 13388
rect 27068 13336 27120 13388
rect 27344 13379 27396 13388
rect 27344 13345 27353 13379
rect 27353 13345 27387 13379
rect 27387 13345 27396 13379
rect 27344 13336 27396 13345
rect 28540 13336 28592 13388
rect 28908 13336 28960 13388
rect 30472 13404 30524 13456
rect 33416 13404 33468 13456
rect 33876 13404 33928 13456
rect 24492 13268 24544 13320
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 26884 13268 26936 13320
rect 26976 13268 27028 13320
rect 28080 13268 28132 13320
rect 28632 13268 28684 13320
rect 21548 13200 21600 13252
rect 23204 13200 23256 13252
rect 20352 13132 20404 13184
rect 20812 13132 20864 13184
rect 22468 13175 22520 13184
rect 22468 13141 22477 13175
rect 22477 13141 22511 13175
rect 22511 13141 22520 13175
rect 22468 13132 22520 13141
rect 23480 13132 23532 13184
rect 24032 13132 24084 13184
rect 24676 13132 24728 13184
rect 24860 13132 24912 13184
rect 25136 13132 25188 13184
rect 25412 13132 25464 13184
rect 26424 13200 26476 13252
rect 26792 13132 26844 13184
rect 27620 13132 27672 13184
rect 27896 13132 27948 13184
rect 28080 13132 28132 13184
rect 28632 13132 28684 13184
rect 28724 13175 28776 13184
rect 28724 13141 28733 13175
rect 28733 13141 28767 13175
rect 28767 13141 28776 13175
rect 28724 13132 28776 13141
rect 29092 13200 29144 13252
rect 29368 13311 29420 13320
rect 29368 13277 29377 13311
rect 29377 13277 29411 13311
rect 29411 13277 29420 13311
rect 29368 13268 29420 13277
rect 33048 13336 33100 13388
rect 33232 13379 33284 13388
rect 33232 13345 33241 13379
rect 33241 13345 33275 13379
rect 33275 13345 33284 13379
rect 33232 13336 33284 13345
rect 33324 13336 33376 13388
rect 29736 13268 29788 13320
rect 30472 13268 30524 13320
rect 30564 13268 30616 13320
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 33968 13268 34020 13320
rect 35900 13472 35952 13524
rect 35992 13472 36044 13524
rect 36360 13472 36412 13524
rect 37372 13472 37424 13524
rect 38016 13472 38068 13524
rect 39304 13472 39356 13524
rect 40224 13472 40276 13524
rect 35624 13336 35676 13388
rect 36544 13336 36596 13388
rect 31392 13200 31444 13252
rect 30932 13132 30984 13184
rect 31484 13132 31536 13184
rect 33876 13200 33928 13252
rect 34336 13243 34388 13252
rect 34336 13209 34345 13243
rect 34345 13209 34379 13243
rect 34379 13209 34388 13243
rect 34336 13200 34388 13209
rect 37556 13268 37608 13320
rect 33048 13175 33100 13184
rect 33048 13141 33057 13175
rect 33057 13141 33091 13175
rect 33091 13141 33100 13175
rect 33048 13132 33100 13141
rect 33508 13175 33560 13184
rect 33508 13141 33517 13175
rect 33517 13141 33551 13175
rect 33551 13141 33560 13175
rect 33508 13132 33560 13141
rect 34704 13132 34756 13184
rect 35072 13132 35124 13184
rect 37648 13200 37700 13252
rect 38200 13336 38252 13388
rect 39028 13404 39080 13456
rect 40776 13336 40828 13388
rect 39028 13268 39080 13320
rect 38844 13132 38896 13184
rect 39488 13243 39540 13252
rect 39488 13209 39497 13243
rect 39497 13209 39531 13243
rect 39531 13209 39540 13243
rect 39488 13200 39540 13209
rect 39764 13200 39816 13252
rect 40224 13200 40276 13252
rect 41328 13515 41380 13524
rect 41328 13481 41337 13515
rect 41337 13481 41371 13515
rect 41371 13481 41380 13515
rect 41328 13472 41380 13481
rect 40960 13404 41012 13456
rect 43076 13447 43128 13456
rect 43076 13413 43085 13447
rect 43085 13413 43119 13447
rect 43119 13413 43128 13447
rect 43076 13404 43128 13413
rect 39212 13132 39264 13184
rect 41972 13175 42024 13184
rect 41972 13141 41981 13175
rect 41981 13141 42015 13175
rect 42015 13141 42024 13175
rect 41972 13132 42024 13141
rect 43352 13132 43404 13184
rect 44548 13175 44600 13184
rect 44548 13141 44557 13175
rect 44557 13141 44591 13175
rect 44591 13141 44600 13175
rect 44548 13132 44600 13141
rect 6070 13030 6122 13082
rect 6134 13030 6186 13082
rect 6198 13030 6250 13082
rect 6262 13030 6314 13082
rect 6326 13030 6378 13082
rect 11070 13030 11122 13082
rect 11134 13030 11186 13082
rect 11198 13030 11250 13082
rect 11262 13030 11314 13082
rect 11326 13030 11378 13082
rect 16070 13030 16122 13082
rect 16134 13030 16186 13082
rect 16198 13030 16250 13082
rect 16262 13030 16314 13082
rect 16326 13030 16378 13082
rect 21070 13030 21122 13082
rect 21134 13030 21186 13082
rect 21198 13030 21250 13082
rect 21262 13030 21314 13082
rect 21326 13030 21378 13082
rect 26070 13030 26122 13082
rect 26134 13030 26186 13082
rect 26198 13030 26250 13082
rect 26262 13030 26314 13082
rect 26326 13030 26378 13082
rect 31070 13030 31122 13082
rect 31134 13030 31186 13082
rect 31198 13030 31250 13082
rect 31262 13030 31314 13082
rect 31326 13030 31378 13082
rect 36070 13030 36122 13082
rect 36134 13030 36186 13082
rect 36198 13030 36250 13082
rect 36262 13030 36314 13082
rect 36326 13030 36378 13082
rect 41070 13030 41122 13082
rect 41134 13030 41186 13082
rect 41198 13030 41250 13082
rect 41262 13030 41314 13082
rect 41326 13030 41378 13082
rect 5908 12928 5960 12980
rect 6920 12928 6972 12980
rect 7288 12928 7340 12980
rect 8484 12928 8536 12980
rect 9956 12928 10008 12980
rect 6644 12860 6696 12912
rect 11428 12971 11480 12980
rect 11428 12937 11437 12971
rect 11437 12937 11471 12971
rect 11471 12937 11480 12971
rect 11428 12928 11480 12937
rect 12900 12928 12952 12980
rect 13912 12928 13964 12980
rect 14004 12928 14056 12980
rect 16948 12928 17000 12980
rect 17868 12928 17920 12980
rect 17960 12928 18012 12980
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 5632 12792 5684 12844
rect 8208 12792 8260 12844
rect 10140 12792 10192 12844
rect 11336 12792 11388 12844
rect 5080 12724 5132 12776
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5632 12656 5684 12708
rect 6000 12724 6052 12776
rect 6644 12724 6696 12776
rect 8024 12724 8076 12776
rect 9128 12724 9180 12776
rect 9772 12724 9824 12776
rect 5172 12588 5224 12640
rect 7840 12631 7892 12640
rect 7840 12597 7849 12631
rect 7849 12597 7883 12631
rect 7883 12597 7892 12631
rect 7840 12588 7892 12597
rect 8208 12588 8260 12640
rect 13176 12860 13228 12912
rect 13360 12903 13412 12912
rect 13360 12869 13369 12903
rect 13369 12869 13403 12903
rect 13403 12869 13412 12903
rect 13360 12860 13412 12869
rect 14372 12860 14424 12912
rect 19156 12928 19208 12980
rect 18236 12903 18288 12912
rect 18236 12869 18245 12903
rect 18245 12869 18279 12903
rect 18279 12869 18288 12903
rect 18236 12860 18288 12869
rect 19616 12928 19668 12980
rect 20444 12860 20496 12912
rect 12624 12792 12676 12844
rect 12716 12792 12768 12844
rect 13268 12792 13320 12844
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 15476 12724 15528 12776
rect 16488 12792 16540 12844
rect 17592 12792 17644 12844
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 19984 12792 20036 12844
rect 20168 12792 20220 12844
rect 17776 12724 17828 12776
rect 18236 12724 18288 12776
rect 18880 12724 18932 12776
rect 18972 12724 19024 12776
rect 19248 12724 19300 12776
rect 9404 12588 9456 12640
rect 9680 12588 9732 12640
rect 19616 12656 19668 12708
rect 20904 12928 20956 12980
rect 22744 12928 22796 12980
rect 24584 12928 24636 12980
rect 22468 12792 22520 12844
rect 23296 12792 23348 12844
rect 23756 12835 23808 12844
rect 23756 12801 23765 12835
rect 23765 12801 23799 12835
rect 23799 12801 23808 12835
rect 23756 12792 23808 12801
rect 20812 12724 20864 12776
rect 20904 12656 20956 12708
rect 21548 12724 21600 12776
rect 23204 12656 23256 12708
rect 23296 12656 23348 12708
rect 24032 12724 24084 12776
rect 24400 12792 24452 12844
rect 24952 12860 25004 12912
rect 25320 12860 25372 12912
rect 25412 12860 25464 12912
rect 26424 12860 26476 12912
rect 26792 12860 26844 12912
rect 27620 12928 27672 12980
rect 28356 12928 28408 12980
rect 29368 12928 29420 12980
rect 29552 12928 29604 12980
rect 29828 12928 29880 12980
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 14096 12588 14148 12640
rect 15292 12588 15344 12640
rect 19708 12631 19760 12640
rect 19708 12597 19717 12631
rect 19717 12597 19751 12631
rect 19751 12597 19760 12631
rect 19708 12588 19760 12597
rect 19892 12588 19944 12640
rect 20628 12588 20680 12640
rect 24124 12631 24176 12640
rect 24124 12597 24133 12631
rect 24133 12597 24167 12631
rect 24167 12597 24176 12631
rect 24124 12588 24176 12597
rect 24584 12631 24636 12640
rect 24584 12597 24593 12631
rect 24593 12597 24627 12631
rect 24627 12597 24636 12631
rect 24584 12588 24636 12597
rect 24860 12656 24912 12708
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 27160 12792 27212 12844
rect 28080 12860 28132 12912
rect 28908 12860 28960 12912
rect 25228 12724 25280 12733
rect 25688 12724 25740 12776
rect 26516 12724 26568 12776
rect 26608 12724 26660 12776
rect 27528 12792 27580 12844
rect 28540 12792 28592 12844
rect 28632 12835 28684 12844
rect 28632 12801 28641 12835
rect 28641 12801 28675 12835
rect 28675 12801 28684 12835
rect 28632 12792 28684 12801
rect 30012 12860 30064 12912
rect 30472 12928 30524 12980
rect 30748 12928 30800 12980
rect 26424 12656 26476 12708
rect 25780 12588 25832 12640
rect 26976 12699 27028 12708
rect 26976 12665 26985 12699
rect 26985 12665 27019 12699
rect 27019 12665 27028 12699
rect 26976 12656 27028 12665
rect 27804 12724 27856 12776
rect 29736 12835 29788 12844
rect 29736 12801 29745 12835
rect 29745 12801 29779 12835
rect 29779 12801 29788 12835
rect 29736 12792 29788 12801
rect 30288 12835 30340 12844
rect 30288 12801 30297 12835
rect 30297 12801 30331 12835
rect 30331 12801 30340 12835
rect 30288 12792 30340 12801
rect 31484 12860 31536 12912
rect 32220 12860 32272 12912
rect 33232 12860 33284 12912
rect 33508 12860 33560 12912
rect 33876 12860 33928 12912
rect 34980 12928 35032 12980
rect 35808 12928 35860 12980
rect 36544 12928 36596 12980
rect 37280 12928 37332 12980
rect 37648 12928 37700 12980
rect 38936 12928 38988 12980
rect 39488 12928 39540 12980
rect 40132 12928 40184 12980
rect 42432 12971 42484 12980
rect 42432 12937 42441 12971
rect 42441 12937 42475 12971
rect 42475 12937 42484 12971
rect 42432 12928 42484 12937
rect 35348 12860 35400 12912
rect 38200 12860 38252 12912
rect 26700 12631 26752 12640
rect 26700 12597 26709 12631
rect 26709 12597 26743 12631
rect 26743 12597 26752 12631
rect 26700 12588 26752 12597
rect 26792 12588 26844 12640
rect 27436 12588 27488 12640
rect 27896 12588 27948 12640
rect 29276 12724 29328 12776
rect 30104 12724 30156 12776
rect 33324 12835 33376 12844
rect 33324 12801 33333 12835
rect 33333 12801 33367 12835
rect 33367 12801 33376 12835
rect 33324 12792 33376 12801
rect 28816 12656 28868 12708
rect 30840 12724 30892 12776
rect 31484 12767 31536 12776
rect 31484 12733 31493 12767
rect 31493 12733 31527 12767
rect 31527 12733 31536 12767
rect 31484 12724 31536 12733
rect 35624 12792 35676 12844
rect 39672 12903 39724 12912
rect 39672 12869 39681 12903
rect 39681 12869 39715 12903
rect 39715 12869 39724 12903
rect 39672 12860 39724 12869
rect 39764 12903 39816 12912
rect 39764 12869 39773 12903
rect 39773 12869 39807 12903
rect 39807 12869 39816 12903
rect 39764 12860 39816 12869
rect 39856 12860 39908 12912
rect 40040 12792 40092 12844
rect 35992 12724 36044 12776
rect 36912 12767 36964 12776
rect 36912 12733 36921 12767
rect 36921 12733 36955 12767
rect 36955 12733 36964 12767
rect 36912 12724 36964 12733
rect 39580 12724 39632 12776
rect 39212 12699 39264 12708
rect 39212 12665 39221 12699
rect 39221 12665 39255 12699
rect 39255 12665 39264 12699
rect 39212 12656 39264 12665
rect 40960 12724 41012 12776
rect 42892 12724 42944 12776
rect 29092 12588 29144 12640
rect 29828 12588 29880 12640
rect 29920 12631 29972 12640
rect 29920 12597 29929 12631
rect 29929 12597 29963 12631
rect 29963 12597 29972 12631
rect 29920 12588 29972 12597
rect 30380 12588 30432 12640
rect 30748 12588 30800 12640
rect 32312 12588 32364 12640
rect 32772 12588 32824 12640
rect 32864 12588 32916 12640
rect 33048 12588 33100 12640
rect 33416 12588 33468 12640
rect 34152 12588 34204 12640
rect 39028 12588 39080 12640
rect 40500 12588 40552 12640
rect 41972 12588 42024 12640
rect 42616 12588 42668 12640
rect 44364 12588 44416 12640
rect 3570 12486 3622 12538
rect 3634 12486 3686 12538
rect 3698 12486 3750 12538
rect 3762 12486 3814 12538
rect 3826 12486 3878 12538
rect 8570 12486 8622 12538
rect 8634 12486 8686 12538
rect 8698 12486 8750 12538
rect 8762 12486 8814 12538
rect 8826 12486 8878 12538
rect 13570 12486 13622 12538
rect 13634 12486 13686 12538
rect 13698 12486 13750 12538
rect 13762 12486 13814 12538
rect 13826 12486 13878 12538
rect 18570 12486 18622 12538
rect 18634 12486 18686 12538
rect 18698 12486 18750 12538
rect 18762 12486 18814 12538
rect 18826 12486 18878 12538
rect 23570 12486 23622 12538
rect 23634 12486 23686 12538
rect 23698 12486 23750 12538
rect 23762 12486 23814 12538
rect 23826 12486 23878 12538
rect 28570 12486 28622 12538
rect 28634 12486 28686 12538
rect 28698 12486 28750 12538
rect 28762 12486 28814 12538
rect 28826 12486 28878 12538
rect 33570 12486 33622 12538
rect 33634 12486 33686 12538
rect 33698 12486 33750 12538
rect 33762 12486 33814 12538
rect 33826 12486 33878 12538
rect 38570 12486 38622 12538
rect 38634 12486 38686 12538
rect 38698 12486 38750 12538
rect 38762 12486 38814 12538
rect 38826 12486 38878 12538
rect 43570 12486 43622 12538
rect 43634 12486 43686 12538
rect 43698 12486 43750 12538
rect 43762 12486 43814 12538
rect 43826 12486 43878 12538
rect 5264 12384 5316 12436
rect 5080 12316 5132 12368
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 8024 12427 8076 12436
rect 8024 12393 8033 12427
rect 8033 12393 8067 12427
rect 8067 12393 8076 12427
rect 8024 12384 8076 12393
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 11704 12384 11756 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 17132 12384 17184 12436
rect 17776 12384 17828 12436
rect 17868 12384 17920 12436
rect 18880 12384 18932 12436
rect 19064 12384 19116 12436
rect 19892 12384 19944 12436
rect 20352 12384 20404 12436
rect 22928 12384 22980 12436
rect 23388 12427 23440 12436
rect 23388 12393 23397 12427
rect 23397 12393 23431 12427
rect 23431 12393 23440 12427
rect 23388 12384 23440 12393
rect 23940 12384 23992 12436
rect 24216 12384 24268 12436
rect 24492 12384 24544 12436
rect 5540 12248 5592 12300
rect 6000 12248 6052 12300
rect 7104 12248 7156 12300
rect 7288 12291 7340 12300
rect 7288 12257 7297 12291
rect 7297 12257 7331 12291
rect 7331 12257 7340 12291
rect 7288 12248 7340 12257
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 16856 12359 16908 12368
rect 16856 12325 16865 12359
rect 16865 12325 16899 12359
rect 16899 12325 16908 12359
rect 16856 12316 16908 12325
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 17408 12359 17460 12368
rect 17408 12325 17417 12359
rect 17417 12325 17451 12359
rect 17451 12325 17460 12359
rect 17408 12316 17460 12325
rect 17684 12248 17736 12300
rect 7380 12223 7432 12232
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 9588 12223 9640 12232
rect 4988 12155 5040 12164
rect 4988 12121 4997 12155
rect 4997 12121 5031 12155
rect 5031 12121 5040 12155
rect 4988 12112 5040 12121
rect 5080 12112 5132 12164
rect 5264 12044 5316 12096
rect 6828 12112 6880 12164
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12992 12180 13044 12232
rect 14280 12180 14332 12232
rect 15292 12180 15344 12232
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15568 12180 15620 12232
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 18420 12248 18472 12300
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18328 12180 18380 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19064 12223 19116 12232
rect 19064 12189 19078 12223
rect 19078 12189 19112 12223
rect 19112 12189 19116 12223
rect 19064 12180 19116 12189
rect 19248 12180 19300 12232
rect 19524 12316 19576 12368
rect 10140 12112 10192 12164
rect 15016 12112 15068 12164
rect 18052 12155 18104 12164
rect 18052 12121 18061 12155
rect 18061 12121 18095 12155
rect 18095 12121 18104 12155
rect 18052 12112 18104 12121
rect 9036 12044 9088 12053
rect 12164 12044 12216 12096
rect 12624 12044 12676 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 16580 12044 16632 12096
rect 17960 12044 18012 12096
rect 18236 12044 18288 12096
rect 18420 12087 18472 12096
rect 18420 12053 18429 12087
rect 18429 12053 18463 12087
rect 18463 12053 18472 12087
rect 18420 12044 18472 12053
rect 18696 12044 18748 12096
rect 19156 12112 19208 12164
rect 19616 12155 19668 12164
rect 19616 12121 19625 12155
rect 19625 12121 19659 12155
rect 19659 12121 19668 12155
rect 19616 12112 19668 12121
rect 19708 12112 19760 12164
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 20352 12248 20404 12300
rect 22836 12359 22888 12368
rect 22836 12325 22845 12359
rect 22845 12325 22879 12359
rect 22879 12325 22888 12359
rect 22836 12316 22888 12325
rect 24676 12384 24728 12436
rect 25596 12384 25648 12436
rect 27160 12384 27212 12436
rect 28908 12384 28960 12436
rect 30656 12384 30708 12436
rect 30840 12384 30892 12436
rect 33324 12384 33376 12436
rect 33876 12427 33928 12436
rect 33876 12393 33885 12427
rect 33885 12393 33919 12427
rect 33919 12393 33928 12427
rect 33876 12384 33928 12393
rect 34060 12427 34112 12436
rect 34060 12393 34069 12427
rect 34069 12393 34103 12427
rect 34103 12393 34112 12427
rect 34060 12384 34112 12393
rect 34428 12316 34480 12368
rect 34612 12384 34664 12436
rect 34796 12316 34848 12368
rect 20628 12180 20680 12232
rect 20812 12180 20864 12232
rect 22468 12180 22520 12232
rect 21456 12112 21508 12164
rect 19432 12044 19484 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 22744 12180 22796 12232
rect 22836 12180 22888 12232
rect 23112 12223 23164 12232
rect 23112 12189 23121 12223
rect 23121 12189 23155 12223
rect 23155 12189 23164 12223
rect 23112 12180 23164 12189
rect 23388 12180 23440 12232
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 24768 12291 24820 12300
rect 24768 12257 24777 12291
rect 24777 12257 24811 12291
rect 24811 12257 24820 12291
rect 24768 12248 24820 12257
rect 25044 12248 25096 12300
rect 25964 12248 26016 12300
rect 26884 12248 26936 12300
rect 27712 12248 27764 12300
rect 27896 12291 27948 12300
rect 27896 12257 27905 12291
rect 27905 12257 27939 12291
rect 27939 12257 27948 12291
rect 27896 12248 27948 12257
rect 28448 12248 28500 12300
rect 29644 12248 29696 12300
rect 29828 12248 29880 12300
rect 24308 12180 24360 12232
rect 24400 12223 24452 12232
rect 24400 12189 24409 12223
rect 24409 12189 24443 12223
rect 24443 12189 24452 12223
rect 24400 12180 24452 12189
rect 25136 12223 25188 12232
rect 25136 12189 25145 12223
rect 25145 12189 25179 12223
rect 25179 12189 25188 12223
rect 25136 12180 25188 12189
rect 26516 12180 26568 12232
rect 26700 12180 26752 12232
rect 25688 12112 25740 12164
rect 27896 12112 27948 12164
rect 30656 12180 30708 12232
rect 32864 12248 32916 12300
rect 33324 12291 33376 12300
rect 33324 12257 33333 12291
rect 33333 12257 33367 12291
rect 33367 12257 33376 12291
rect 33324 12248 33376 12257
rect 31576 12223 31628 12232
rect 31576 12189 31585 12223
rect 31585 12189 31619 12223
rect 31619 12189 31628 12223
rect 31576 12180 31628 12189
rect 31668 12180 31720 12232
rect 32496 12223 32548 12232
rect 32496 12189 32505 12223
rect 32505 12189 32539 12223
rect 32539 12189 32548 12223
rect 32496 12180 32548 12189
rect 33876 12180 33928 12232
rect 34980 12291 35032 12300
rect 34980 12257 34989 12291
rect 34989 12257 35023 12291
rect 35023 12257 35032 12291
rect 34980 12248 35032 12257
rect 35716 12384 35768 12436
rect 37096 12384 37148 12436
rect 37188 12427 37240 12436
rect 37188 12393 37197 12427
rect 37197 12393 37231 12427
rect 37231 12393 37240 12427
rect 37188 12384 37240 12393
rect 43444 12384 43496 12436
rect 36452 12248 36504 12300
rect 37740 12291 37792 12300
rect 37740 12257 37749 12291
rect 37749 12257 37783 12291
rect 37783 12257 37792 12291
rect 37740 12248 37792 12257
rect 35164 12223 35216 12232
rect 35164 12189 35173 12223
rect 35173 12189 35207 12223
rect 35207 12189 35216 12223
rect 35164 12180 35216 12189
rect 37556 12180 37608 12232
rect 37648 12223 37700 12232
rect 37648 12189 37657 12223
rect 37657 12189 37691 12223
rect 37691 12189 37700 12223
rect 37648 12180 37700 12189
rect 38568 12291 38620 12300
rect 38568 12257 38577 12291
rect 38577 12257 38611 12291
rect 38611 12257 38620 12291
rect 38568 12248 38620 12257
rect 38752 12316 38804 12368
rect 42248 12316 42300 12368
rect 44548 12316 44600 12368
rect 39304 12248 39356 12300
rect 41604 12248 41656 12300
rect 38292 12180 38344 12232
rect 39120 12180 39172 12232
rect 41420 12180 41472 12232
rect 26976 12087 27028 12096
rect 26976 12053 26985 12087
rect 26985 12053 27019 12087
rect 27019 12053 27028 12087
rect 26976 12044 27028 12053
rect 27620 12044 27672 12096
rect 28080 12044 28132 12096
rect 30012 12044 30064 12096
rect 30196 12044 30248 12096
rect 32312 12044 32364 12096
rect 33140 12044 33192 12096
rect 33324 12044 33376 12096
rect 33508 12087 33560 12096
rect 33508 12053 33517 12087
rect 33517 12053 33551 12087
rect 33551 12053 33560 12087
rect 33508 12044 33560 12053
rect 34244 12044 34296 12096
rect 37096 12112 37148 12164
rect 36452 12044 36504 12096
rect 37280 12087 37332 12096
rect 37280 12053 37289 12087
rect 37289 12053 37323 12087
rect 37323 12053 37332 12087
rect 37280 12044 37332 12053
rect 38200 12112 38252 12164
rect 39120 12044 39172 12096
rect 43076 12112 43128 12164
rect 39948 12044 40000 12096
rect 40500 12044 40552 12096
rect 40960 12044 41012 12096
rect 41788 12087 41840 12096
rect 41788 12053 41797 12087
rect 41797 12053 41831 12087
rect 41831 12053 41840 12087
rect 41788 12044 41840 12053
rect 42616 12044 42668 12096
rect 44364 12044 44416 12096
rect 44640 12044 44692 12096
rect 6070 11942 6122 11994
rect 6134 11942 6186 11994
rect 6198 11942 6250 11994
rect 6262 11942 6314 11994
rect 6326 11942 6378 11994
rect 11070 11942 11122 11994
rect 11134 11942 11186 11994
rect 11198 11942 11250 11994
rect 11262 11942 11314 11994
rect 11326 11942 11378 11994
rect 16070 11942 16122 11994
rect 16134 11942 16186 11994
rect 16198 11942 16250 11994
rect 16262 11942 16314 11994
rect 16326 11942 16378 11994
rect 21070 11942 21122 11994
rect 21134 11942 21186 11994
rect 21198 11942 21250 11994
rect 21262 11942 21314 11994
rect 21326 11942 21378 11994
rect 26070 11942 26122 11994
rect 26134 11942 26186 11994
rect 26198 11942 26250 11994
rect 26262 11942 26314 11994
rect 26326 11942 26378 11994
rect 31070 11942 31122 11994
rect 31134 11942 31186 11994
rect 31198 11942 31250 11994
rect 31262 11942 31314 11994
rect 31326 11942 31378 11994
rect 36070 11942 36122 11994
rect 36134 11942 36186 11994
rect 36198 11942 36250 11994
rect 36262 11942 36314 11994
rect 36326 11942 36378 11994
rect 41070 11942 41122 11994
rect 41134 11942 41186 11994
rect 41198 11942 41250 11994
rect 41262 11942 41314 11994
rect 41326 11942 41378 11994
rect 4068 11840 4120 11892
rect 5080 11840 5132 11892
rect 5172 11815 5224 11824
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 5908 11840 5960 11892
rect 6828 11840 6880 11892
rect 8024 11840 8076 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 9680 11840 9732 11892
rect 9772 11840 9824 11892
rect 10140 11840 10192 11892
rect 12164 11840 12216 11892
rect 13820 11840 13872 11892
rect 5272 11747 5324 11756
rect 5272 11713 5281 11747
rect 5281 11713 5315 11747
rect 5315 11713 5324 11747
rect 5272 11704 5324 11713
rect 5724 11772 5776 11824
rect 12992 11772 13044 11824
rect 15752 11840 15804 11892
rect 16856 11840 16908 11892
rect 14464 11772 14516 11824
rect 18420 11840 18472 11892
rect 19156 11840 19208 11892
rect 20352 11840 20404 11892
rect 20904 11840 20956 11892
rect 21456 11840 21508 11892
rect 22192 11840 22244 11892
rect 22836 11840 22888 11892
rect 18236 11772 18288 11824
rect 5540 11745 5592 11754
rect 5540 11711 5549 11745
rect 5549 11711 5583 11745
rect 5583 11711 5592 11745
rect 5540 11702 5592 11711
rect 7104 11704 7156 11756
rect 11888 11704 11940 11756
rect 15752 11704 15804 11756
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 5540 11568 5592 11620
rect 7380 11636 7432 11688
rect 10232 11636 10284 11688
rect 11612 11636 11664 11688
rect 7656 11500 7708 11552
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 9036 11500 9088 11552
rect 11520 11568 11572 11620
rect 12532 11679 12584 11688
rect 12532 11645 12541 11679
rect 12541 11645 12575 11679
rect 12575 11645 12584 11679
rect 12532 11636 12584 11645
rect 14004 11636 14056 11688
rect 15016 11636 15068 11688
rect 15844 11636 15896 11688
rect 16580 11679 16632 11688
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 19708 11772 19760 11824
rect 19800 11704 19852 11756
rect 19984 11704 20036 11756
rect 20168 11704 20220 11756
rect 20536 11704 20588 11756
rect 20628 11747 20680 11756
rect 20628 11713 20637 11747
rect 20637 11713 20671 11747
rect 20671 11713 20680 11747
rect 20628 11704 20680 11713
rect 22468 11772 22520 11824
rect 28080 11883 28132 11892
rect 28080 11849 28089 11883
rect 28089 11849 28123 11883
rect 28123 11849 28132 11883
rect 28080 11840 28132 11849
rect 24492 11772 24544 11824
rect 26516 11772 26568 11824
rect 26608 11815 26660 11824
rect 26608 11781 26617 11815
rect 26617 11781 26651 11815
rect 26651 11781 26660 11815
rect 26608 11772 26660 11781
rect 19524 11636 19576 11688
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 21640 11704 21692 11756
rect 25688 11704 25740 11756
rect 27712 11704 27764 11756
rect 28448 11815 28500 11824
rect 28448 11781 28457 11815
rect 28457 11781 28491 11815
rect 28491 11781 28500 11815
rect 28448 11772 28500 11781
rect 30012 11840 30064 11892
rect 30104 11840 30156 11892
rect 29828 11772 29880 11824
rect 30380 11840 30432 11892
rect 30564 11840 30616 11892
rect 30748 11840 30800 11892
rect 11704 11543 11756 11552
rect 11704 11509 11713 11543
rect 11713 11509 11747 11543
rect 11747 11509 11756 11543
rect 11704 11500 11756 11509
rect 12624 11500 12676 11552
rect 13912 11500 13964 11552
rect 15660 11500 15712 11552
rect 15936 11500 15988 11552
rect 17224 11500 17276 11552
rect 18972 11500 19024 11552
rect 19892 11568 19944 11620
rect 19984 11611 20036 11620
rect 19984 11577 19993 11611
rect 19993 11577 20027 11611
rect 20027 11577 20036 11611
rect 19984 11568 20036 11577
rect 20260 11568 20312 11620
rect 20720 11568 20772 11620
rect 22008 11679 22060 11688
rect 22008 11645 22017 11679
rect 22017 11645 22051 11679
rect 22051 11645 22060 11679
rect 22008 11636 22060 11645
rect 25136 11636 25188 11688
rect 25412 11636 25464 11688
rect 25780 11636 25832 11688
rect 26240 11636 26292 11688
rect 28080 11636 28132 11688
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 21548 11500 21600 11552
rect 23112 11500 23164 11552
rect 24124 11500 24176 11552
rect 29552 11568 29604 11620
rect 29736 11636 29788 11688
rect 30196 11568 30248 11620
rect 24400 11500 24452 11552
rect 25688 11500 25740 11552
rect 29828 11500 29880 11552
rect 30012 11500 30064 11552
rect 30656 11704 30708 11756
rect 30840 11772 30892 11824
rect 32128 11840 32180 11892
rect 32312 11840 32364 11892
rect 33232 11840 33284 11892
rect 33324 11840 33376 11892
rect 34612 11840 34664 11892
rect 35440 11840 35492 11892
rect 35716 11840 35768 11892
rect 32220 11772 32272 11824
rect 32588 11772 32640 11824
rect 33324 11747 33376 11756
rect 33324 11713 33333 11747
rect 33333 11713 33367 11747
rect 33367 11713 33376 11747
rect 33324 11704 33376 11713
rect 32864 11636 32916 11688
rect 32680 11568 32732 11620
rect 34520 11772 34572 11824
rect 34704 11747 34756 11756
rect 34704 11713 34713 11747
rect 34713 11713 34747 11747
rect 34747 11713 34756 11747
rect 34704 11704 34756 11713
rect 35900 11704 35952 11756
rect 33968 11636 34020 11688
rect 34428 11679 34480 11688
rect 34428 11645 34437 11679
rect 34437 11645 34471 11679
rect 34471 11645 34480 11679
rect 34428 11636 34480 11645
rect 34520 11636 34572 11688
rect 37096 11840 37148 11892
rect 37280 11840 37332 11892
rect 37648 11840 37700 11892
rect 37464 11772 37516 11824
rect 38292 11840 38344 11892
rect 40776 11883 40828 11892
rect 40776 11849 40785 11883
rect 40785 11849 40819 11883
rect 40819 11849 40828 11883
rect 40776 11840 40828 11849
rect 41604 11840 41656 11892
rect 42340 11883 42392 11892
rect 42340 11849 42349 11883
rect 42349 11849 42383 11883
rect 42383 11849 42392 11883
rect 42340 11840 42392 11849
rect 39212 11772 39264 11824
rect 44732 11772 44784 11824
rect 36544 11636 36596 11688
rect 35716 11568 35768 11620
rect 37004 11636 37056 11688
rect 38200 11636 38252 11688
rect 38476 11679 38528 11688
rect 38476 11645 38485 11679
rect 38485 11645 38519 11679
rect 38519 11645 38528 11679
rect 38476 11636 38528 11645
rect 37924 11568 37976 11620
rect 39764 11636 39816 11688
rect 41420 11704 41472 11756
rect 43076 11747 43128 11756
rect 43076 11713 43085 11747
rect 43085 11713 43119 11747
rect 43119 11713 43128 11747
rect 43076 11704 43128 11713
rect 40408 11679 40460 11688
rect 40408 11645 40417 11679
rect 40417 11645 40451 11679
rect 40451 11645 40460 11679
rect 40408 11636 40460 11645
rect 41604 11636 41656 11688
rect 42432 11636 42484 11688
rect 42708 11636 42760 11688
rect 45008 11704 45060 11756
rect 44824 11679 44876 11688
rect 44824 11645 44833 11679
rect 44833 11645 44867 11679
rect 44867 11645 44876 11679
rect 44824 11636 44876 11645
rect 33048 11500 33100 11552
rect 33140 11543 33192 11552
rect 33140 11509 33149 11543
rect 33149 11509 33183 11543
rect 33183 11509 33192 11543
rect 33140 11500 33192 11509
rect 33232 11500 33284 11552
rect 34060 11500 34112 11552
rect 35072 11543 35124 11552
rect 35072 11509 35081 11543
rect 35081 11509 35115 11543
rect 35115 11509 35124 11543
rect 35072 11500 35124 11509
rect 36912 11500 36964 11552
rect 37096 11500 37148 11552
rect 38752 11500 38804 11552
rect 38936 11500 38988 11552
rect 40960 11500 41012 11552
rect 3570 11398 3622 11450
rect 3634 11398 3686 11450
rect 3698 11398 3750 11450
rect 3762 11398 3814 11450
rect 3826 11398 3878 11450
rect 8570 11398 8622 11450
rect 8634 11398 8686 11450
rect 8698 11398 8750 11450
rect 8762 11398 8814 11450
rect 8826 11398 8878 11450
rect 13570 11398 13622 11450
rect 13634 11398 13686 11450
rect 13698 11398 13750 11450
rect 13762 11398 13814 11450
rect 13826 11398 13878 11450
rect 18570 11398 18622 11450
rect 18634 11398 18686 11450
rect 18698 11398 18750 11450
rect 18762 11398 18814 11450
rect 18826 11398 18878 11450
rect 23570 11398 23622 11450
rect 23634 11398 23686 11450
rect 23698 11398 23750 11450
rect 23762 11398 23814 11450
rect 23826 11398 23878 11450
rect 28570 11398 28622 11450
rect 28634 11398 28686 11450
rect 28698 11398 28750 11450
rect 28762 11398 28814 11450
rect 28826 11398 28878 11450
rect 33570 11398 33622 11450
rect 33634 11398 33686 11450
rect 33698 11398 33750 11450
rect 33762 11398 33814 11450
rect 33826 11398 33878 11450
rect 38570 11398 38622 11450
rect 38634 11398 38686 11450
rect 38698 11398 38750 11450
rect 38762 11398 38814 11450
rect 38826 11398 38878 11450
rect 43570 11398 43622 11450
rect 43634 11398 43686 11450
rect 43698 11398 43750 11450
rect 43762 11398 43814 11450
rect 43826 11398 43878 11450
rect 7104 11296 7156 11348
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 11704 11296 11756 11348
rect 12532 11296 12584 11348
rect 4160 11024 4212 11076
rect 4988 11092 5040 11144
rect 5356 11092 5408 11144
rect 8392 11024 8444 11076
rect 9036 11024 9088 11076
rect 9680 11092 9732 11144
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 9496 11067 9548 11076
rect 9496 11033 9505 11067
rect 9505 11033 9539 11067
rect 9539 11033 9548 11067
rect 9496 11024 9548 11033
rect 11428 11092 11480 11144
rect 12624 11228 12676 11280
rect 12992 11228 13044 11280
rect 13084 11228 13136 11280
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 13820 11160 13872 11212
rect 16948 11296 17000 11348
rect 19064 11296 19116 11348
rect 20720 11339 20772 11348
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 20904 11296 20956 11348
rect 21364 11296 21416 11348
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 24124 11296 24176 11348
rect 25964 11296 26016 11348
rect 26240 11296 26292 11348
rect 27620 11296 27672 11348
rect 27896 11339 27948 11348
rect 27896 11305 27905 11339
rect 27905 11305 27939 11339
rect 27939 11305 27948 11339
rect 27896 11296 27948 11305
rect 28448 11296 28500 11348
rect 29644 11296 29696 11348
rect 14372 11228 14424 11280
rect 17684 11228 17736 11280
rect 17776 11228 17828 11280
rect 21640 11228 21692 11280
rect 23388 11228 23440 11280
rect 13728 11092 13780 11144
rect 4344 10956 4396 11008
rect 5172 10956 5224 11008
rect 5540 10956 5592 11008
rect 5724 10999 5776 11008
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 5724 10956 5776 10965
rect 6000 10956 6052 11008
rect 9312 10999 9364 11008
rect 9312 10965 9321 10999
rect 9321 10965 9355 10999
rect 9355 10965 9364 10999
rect 9312 10956 9364 10965
rect 10232 10999 10284 11008
rect 10232 10965 10241 10999
rect 10241 10965 10275 10999
rect 10275 10965 10284 10999
rect 10232 10956 10284 10965
rect 11428 10956 11480 11008
rect 11704 10999 11756 11008
rect 11704 10965 11713 10999
rect 11713 10965 11747 10999
rect 11747 10965 11756 10999
rect 11704 10956 11756 10965
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15016 11092 15068 11144
rect 19340 11160 19392 11212
rect 19524 11160 19576 11212
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 15660 11024 15712 11076
rect 15844 11024 15896 11076
rect 19248 11092 19300 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20260 11160 20312 11212
rect 20352 11092 20404 11144
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 22468 11203 22520 11212
rect 22468 11169 22477 11203
rect 22477 11169 22511 11203
rect 22511 11169 22520 11203
rect 22468 11160 22520 11169
rect 22652 11160 22704 11212
rect 22836 11160 22888 11212
rect 25688 11228 25740 11280
rect 24584 11160 24636 11212
rect 25964 11160 26016 11212
rect 26976 11160 27028 11212
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 13636 10956 13688 11008
rect 13912 10956 13964 11008
rect 14004 10956 14056 11008
rect 14280 10956 14332 11008
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 18972 10956 19024 11008
rect 20260 10956 20312 11008
rect 21548 10999 21600 11008
rect 21548 10965 21557 10999
rect 21557 10965 21591 10999
rect 21591 10965 21600 10999
rect 21548 10956 21600 10965
rect 21640 10999 21692 11008
rect 21640 10965 21649 10999
rect 21649 10965 21683 10999
rect 21683 10965 21692 10999
rect 21640 10956 21692 10965
rect 21916 10956 21968 11008
rect 22744 11092 22796 11144
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24032 11092 24084 11101
rect 24400 11092 24452 11144
rect 29460 11228 29512 11280
rect 29184 11160 29236 11212
rect 29644 11160 29696 11212
rect 31760 11296 31812 11348
rect 32680 11296 32732 11348
rect 31852 11228 31904 11280
rect 30748 11160 30800 11212
rect 31668 11160 31720 11212
rect 29736 11092 29788 11144
rect 32036 11092 32088 11144
rect 32312 11092 32364 11144
rect 33324 11296 33376 11348
rect 32680 11160 32732 11212
rect 32864 11160 32916 11212
rect 32956 11160 33008 11212
rect 37004 11296 37056 11348
rect 37924 11296 37976 11348
rect 33968 11160 34020 11212
rect 34060 11160 34112 11212
rect 34428 11203 34480 11212
rect 34428 11169 34437 11203
rect 34437 11169 34471 11203
rect 34471 11169 34480 11203
rect 34428 11160 34480 11169
rect 35440 11160 35492 11212
rect 35716 11160 35768 11212
rect 38844 11296 38896 11348
rect 39304 11296 39356 11348
rect 39948 11296 40000 11348
rect 27712 11024 27764 11076
rect 29368 11024 29420 11076
rect 29552 11067 29604 11076
rect 29552 11033 29561 11067
rect 29561 11033 29595 11067
rect 29595 11033 29604 11067
rect 29552 11024 29604 11033
rect 30656 11024 30708 11076
rect 22928 10956 22980 11008
rect 25596 10956 25648 11008
rect 28448 10956 28500 11008
rect 32312 10956 32364 11008
rect 32404 10999 32456 11008
rect 32404 10965 32434 10999
rect 32434 10965 32456 10999
rect 34336 11024 34388 11076
rect 34980 11024 35032 11076
rect 32404 10956 32456 10965
rect 33324 10956 33376 11008
rect 33876 10956 33928 11008
rect 34888 10956 34940 11008
rect 36084 10956 36136 11008
rect 36636 11092 36688 11144
rect 38844 11203 38896 11212
rect 38844 11169 38853 11203
rect 38853 11169 38887 11203
rect 38887 11169 38896 11203
rect 38844 11160 38896 11169
rect 41972 11228 42024 11280
rect 39028 11160 39080 11212
rect 41604 11160 41656 11212
rect 42064 11160 42116 11212
rect 38660 11135 38712 11144
rect 38660 11101 38669 11135
rect 38669 11101 38703 11135
rect 38703 11101 38712 11135
rect 38660 11092 38712 11101
rect 37096 11024 37148 11076
rect 37464 10999 37516 11008
rect 37464 10965 37473 10999
rect 37473 10965 37507 10999
rect 37507 10965 37516 10999
rect 37464 10956 37516 10965
rect 38568 11024 38620 11076
rect 38476 10956 38528 11008
rect 41512 11135 41564 11144
rect 41512 11101 41521 11135
rect 41521 11101 41555 11135
rect 41555 11101 41564 11135
rect 41512 11092 41564 11101
rect 42800 11296 42852 11348
rect 44548 11296 44600 11348
rect 42708 11228 42760 11280
rect 43444 11092 43496 11144
rect 39028 11024 39080 11076
rect 39948 11024 40000 11076
rect 40776 11024 40828 11076
rect 42800 11024 42852 11076
rect 39672 10956 39724 11008
rect 40316 10956 40368 11008
rect 41880 10956 41932 11008
rect 42984 10999 43036 11008
rect 42984 10965 42993 10999
rect 42993 10965 43027 10999
rect 43027 10965 43036 10999
rect 42984 10956 43036 10965
rect 44548 10999 44600 11008
rect 44548 10965 44557 10999
rect 44557 10965 44591 10999
rect 44591 10965 44600 10999
rect 44548 10956 44600 10965
rect 44732 10956 44784 11008
rect 6070 10854 6122 10906
rect 6134 10854 6186 10906
rect 6198 10854 6250 10906
rect 6262 10854 6314 10906
rect 6326 10854 6378 10906
rect 11070 10854 11122 10906
rect 11134 10854 11186 10906
rect 11198 10854 11250 10906
rect 11262 10854 11314 10906
rect 11326 10854 11378 10906
rect 16070 10854 16122 10906
rect 16134 10854 16186 10906
rect 16198 10854 16250 10906
rect 16262 10854 16314 10906
rect 16326 10854 16378 10906
rect 21070 10854 21122 10906
rect 21134 10854 21186 10906
rect 21198 10854 21250 10906
rect 21262 10854 21314 10906
rect 21326 10854 21378 10906
rect 26070 10854 26122 10906
rect 26134 10854 26186 10906
rect 26198 10854 26250 10906
rect 26262 10854 26314 10906
rect 26326 10854 26378 10906
rect 31070 10854 31122 10906
rect 31134 10854 31186 10906
rect 31198 10854 31250 10906
rect 31262 10854 31314 10906
rect 31326 10854 31378 10906
rect 36070 10854 36122 10906
rect 36134 10854 36186 10906
rect 36198 10854 36250 10906
rect 36262 10854 36314 10906
rect 36326 10854 36378 10906
rect 41070 10854 41122 10906
rect 41134 10854 41186 10906
rect 41198 10854 41250 10906
rect 41262 10854 41314 10906
rect 41326 10854 41378 10906
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 9312 10752 9364 10804
rect 11520 10752 11572 10804
rect 11796 10752 11848 10804
rect 13084 10752 13136 10804
rect 14280 10752 14332 10804
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 5356 10548 5408 10600
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 9036 10684 9088 10736
rect 10232 10684 10284 10736
rect 11428 10684 11480 10736
rect 12164 10684 12216 10736
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17776 10752 17828 10804
rect 18972 10795 19024 10804
rect 18972 10761 18981 10795
rect 18981 10761 19015 10795
rect 19015 10761 19024 10795
rect 18972 10752 19024 10761
rect 19248 10752 19300 10804
rect 15108 10684 15160 10736
rect 15936 10684 15988 10736
rect 16856 10684 16908 10736
rect 18236 10684 18288 10736
rect 20260 10684 20312 10736
rect 21640 10727 21692 10736
rect 21640 10693 21649 10727
rect 21649 10693 21683 10727
rect 21683 10693 21692 10727
rect 21640 10684 21692 10693
rect 22192 10752 22244 10804
rect 22468 10752 22520 10804
rect 24860 10752 24912 10804
rect 25320 10795 25372 10804
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 25688 10795 25740 10804
rect 25688 10761 25697 10795
rect 25697 10761 25731 10795
rect 25731 10761 25740 10795
rect 25688 10752 25740 10761
rect 27620 10752 27672 10804
rect 28080 10752 28132 10804
rect 28172 10752 28224 10804
rect 28356 10752 28408 10804
rect 29368 10795 29420 10804
rect 29368 10761 29393 10795
rect 29393 10761 29420 10795
rect 29368 10752 29420 10761
rect 29552 10752 29604 10804
rect 30196 10752 30248 10804
rect 25596 10684 25648 10736
rect 29184 10727 29236 10736
rect 29184 10693 29193 10727
rect 29193 10693 29227 10727
rect 29227 10693 29236 10727
rect 29184 10684 29236 10693
rect 29644 10684 29696 10736
rect 29920 10684 29972 10736
rect 3424 10412 3476 10464
rect 3976 10412 4028 10464
rect 6000 10480 6052 10532
rect 7840 10523 7892 10532
rect 7840 10489 7849 10523
rect 7849 10489 7883 10523
rect 7883 10489 7892 10523
rect 7840 10480 7892 10489
rect 8484 10616 8536 10668
rect 10048 10616 10100 10668
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 8392 10412 8444 10464
rect 8484 10412 8536 10464
rect 8944 10412 8996 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 10784 10548 10836 10600
rect 11612 10548 11664 10600
rect 11796 10548 11848 10600
rect 11888 10412 11940 10464
rect 12716 10412 12768 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13360 10548 13412 10600
rect 13636 10548 13688 10600
rect 15752 10616 15804 10668
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 25044 10659 25096 10668
rect 25044 10625 25053 10659
rect 25053 10625 25087 10659
rect 25087 10625 25096 10659
rect 25044 10616 25096 10625
rect 25964 10616 26016 10668
rect 26148 10616 26200 10668
rect 27712 10616 27764 10668
rect 28264 10659 28316 10668
rect 28264 10625 28273 10659
rect 28273 10625 28307 10659
rect 28307 10625 28316 10659
rect 28264 10616 28316 10625
rect 17132 10548 17184 10600
rect 15660 10480 15712 10532
rect 14004 10412 14056 10464
rect 14556 10412 14608 10464
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 16580 10455 16632 10464
rect 16580 10421 16589 10455
rect 16589 10421 16623 10455
rect 16623 10421 16632 10455
rect 16580 10412 16632 10421
rect 17500 10591 17552 10600
rect 17500 10557 17509 10591
rect 17509 10557 17543 10591
rect 17543 10557 17552 10591
rect 17500 10548 17552 10557
rect 19984 10412 20036 10464
rect 20812 10412 20864 10464
rect 21180 10412 21232 10464
rect 21548 10412 21600 10464
rect 22008 10412 22060 10464
rect 23204 10591 23256 10600
rect 23204 10557 23213 10591
rect 23213 10557 23247 10591
rect 23247 10557 23256 10591
rect 23204 10548 23256 10557
rect 23940 10548 23992 10600
rect 25596 10548 25648 10600
rect 29276 10616 29328 10668
rect 29736 10659 29788 10668
rect 29736 10625 29745 10659
rect 29745 10625 29779 10659
rect 29779 10625 29788 10659
rect 29736 10616 29788 10625
rect 30932 10684 30984 10736
rect 30472 10616 30524 10668
rect 30840 10616 30892 10668
rect 30288 10548 30340 10600
rect 31668 10684 31720 10736
rect 32588 10752 32640 10804
rect 31484 10659 31536 10668
rect 31484 10625 31493 10659
rect 31493 10625 31527 10659
rect 31527 10625 31536 10659
rect 31484 10616 31536 10625
rect 28264 10480 28316 10532
rect 29276 10480 29328 10532
rect 23940 10412 23992 10464
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 25780 10412 25832 10464
rect 28080 10455 28132 10464
rect 28080 10421 28089 10455
rect 28089 10421 28123 10455
rect 28123 10421 28132 10455
rect 28080 10412 28132 10421
rect 29828 10480 29880 10532
rect 32496 10548 32548 10600
rect 34428 10752 34480 10804
rect 34520 10752 34572 10804
rect 33876 10684 33928 10736
rect 35992 10752 36044 10804
rect 36452 10795 36504 10804
rect 36452 10761 36461 10795
rect 36461 10761 36495 10795
rect 36495 10761 36504 10795
rect 36452 10752 36504 10761
rect 34980 10684 35032 10736
rect 37464 10752 37516 10804
rect 36268 10659 36320 10668
rect 36268 10625 36277 10659
rect 36277 10625 36311 10659
rect 36311 10625 36320 10659
rect 36268 10616 36320 10625
rect 36544 10616 36596 10668
rect 34888 10548 34940 10600
rect 35624 10591 35676 10600
rect 35624 10557 35633 10591
rect 35633 10557 35667 10591
rect 35667 10557 35676 10591
rect 35624 10548 35676 10557
rect 35716 10591 35768 10600
rect 35716 10557 35725 10591
rect 35725 10557 35759 10591
rect 35759 10557 35768 10591
rect 35716 10548 35768 10557
rect 35808 10548 35860 10600
rect 29644 10412 29696 10464
rect 38752 10752 38804 10804
rect 39764 10752 39816 10804
rect 39212 10616 39264 10668
rect 39948 10684 40000 10736
rect 37096 10548 37148 10600
rect 39672 10591 39724 10600
rect 39672 10557 39681 10591
rect 39681 10557 39715 10591
rect 39715 10557 39724 10591
rect 39672 10548 39724 10557
rect 39948 10591 40000 10600
rect 39948 10557 39957 10591
rect 39957 10557 39991 10591
rect 39991 10557 40000 10591
rect 39948 10548 40000 10557
rect 41420 10795 41472 10804
rect 41420 10761 41429 10795
rect 41429 10761 41463 10795
rect 41463 10761 41472 10795
rect 41420 10752 41472 10761
rect 42340 10795 42392 10804
rect 42340 10761 42349 10795
rect 42349 10761 42383 10795
rect 42383 10761 42392 10795
rect 42340 10752 42392 10761
rect 43260 10752 43312 10804
rect 44272 10752 44324 10804
rect 44548 10752 44600 10804
rect 42984 10684 43036 10736
rect 41972 10659 42024 10668
rect 41972 10625 41981 10659
rect 41981 10625 42015 10659
rect 42015 10625 42024 10659
rect 41972 10616 42024 10625
rect 41788 10548 41840 10600
rect 42524 10548 42576 10600
rect 30564 10412 30616 10464
rect 30748 10412 30800 10464
rect 31484 10412 31536 10464
rect 32128 10412 32180 10464
rect 35992 10412 36044 10464
rect 36084 10455 36136 10464
rect 36084 10421 36093 10455
rect 36093 10421 36127 10455
rect 36127 10421 36136 10455
rect 36084 10412 36136 10421
rect 41788 10455 41840 10464
rect 41788 10421 41797 10455
rect 41797 10421 41831 10455
rect 41831 10421 41840 10455
rect 41788 10412 41840 10421
rect 44732 10412 44784 10464
rect 44824 10455 44876 10464
rect 44824 10421 44833 10455
rect 44833 10421 44867 10455
rect 44867 10421 44876 10455
rect 44824 10412 44876 10421
rect 3570 10310 3622 10362
rect 3634 10310 3686 10362
rect 3698 10310 3750 10362
rect 3762 10310 3814 10362
rect 3826 10310 3878 10362
rect 8570 10310 8622 10362
rect 8634 10310 8686 10362
rect 8698 10310 8750 10362
rect 8762 10310 8814 10362
rect 8826 10310 8878 10362
rect 13570 10310 13622 10362
rect 13634 10310 13686 10362
rect 13698 10310 13750 10362
rect 13762 10310 13814 10362
rect 13826 10310 13878 10362
rect 18570 10310 18622 10362
rect 18634 10310 18686 10362
rect 18698 10310 18750 10362
rect 18762 10310 18814 10362
rect 18826 10310 18878 10362
rect 23570 10310 23622 10362
rect 23634 10310 23686 10362
rect 23698 10310 23750 10362
rect 23762 10310 23814 10362
rect 23826 10310 23878 10362
rect 28570 10310 28622 10362
rect 28634 10310 28686 10362
rect 28698 10310 28750 10362
rect 28762 10310 28814 10362
rect 28826 10310 28878 10362
rect 33570 10310 33622 10362
rect 33634 10310 33686 10362
rect 33698 10310 33750 10362
rect 33762 10310 33814 10362
rect 33826 10310 33878 10362
rect 38570 10310 38622 10362
rect 38634 10310 38686 10362
rect 38698 10310 38750 10362
rect 38762 10310 38814 10362
rect 38826 10310 38878 10362
rect 43570 10310 43622 10362
rect 43634 10310 43686 10362
rect 43698 10310 43750 10362
rect 43762 10310 43814 10362
rect 43826 10310 43878 10362
rect 3332 10208 3384 10260
rect 4344 10208 4396 10260
rect 3884 10004 3936 10056
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4344 10004 4396 10056
rect 5540 10208 5592 10260
rect 5816 10208 5868 10260
rect 9680 10208 9732 10260
rect 10508 10208 10560 10260
rect 11704 10208 11756 10260
rect 11796 10208 11848 10260
rect 12348 10208 12400 10260
rect 12808 10208 12860 10260
rect 13360 10208 13412 10260
rect 6000 10072 6052 10124
rect 7012 10072 7064 10124
rect 7748 10004 7800 10056
rect 8024 10004 8076 10056
rect 9036 10072 9088 10124
rect 10048 10004 10100 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 12164 10140 12216 10192
rect 13084 10140 13136 10192
rect 13176 10140 13228 10192
rect 14096 10208 14148 10260
rect 14464 10208 14516 10260
rect 15108 10208 15160 10260
rect 16580 10208 16632 10260
rect 17408 10208 17460 10260
rect 17500 10208 17552 10260
rect 18052 10208 18104 10260
rect 5080 9936 5132 9988
rect 6920 9936 6972 9988
rect 8484 9936 8536 9988
rect 11980 10004 12032 10056
rect 10784 9936 10836 9988
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 13176 10004 13228 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 14372 10072 14424 10124
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 14280 10004 14332 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 16672 10004 16724 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 4160 9868 4212 9920
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 5724 9868 5776 9920
rect 6184 9868 6236 9920
rect 6552 9868 6604 9920
rect 8392 9868 8444 9920
rect 9588 9868 9640 9920
rect 11520 9868 11572 9920
rect 14096 9936 14148 9988
rect 14188 9936 14240 9988
rect 12716 9868 12768 9920
rect 13544 9868 13596 9920
rect 13912 9868 13964 9920
rect 15016 9868 15068 9920
rect 15844 9936 15896 9988
rect 17776 10004 17828 10056
rect 19248 10208 19300 10260
rect 19616 10183 19668 10192
rect 19616 10149 19625 10183
rect 19625 10149 19659 10183
rect 19659 10149 19668 10183
rect 19616 10140 19668 10149
rect 20628 10208 20680 10260
rect 18972 10072 19024 10124
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18880 10004 18932 10056
rect 20168 10072 20220 10124
rect 20904 10208 20956 10260
rect 22468 10208 22520 10260
rect 23204 10208 23256 10260
rect 23296 10208 23348 10260
rect 24860 10208 24912 10260
rect 22008 10140 22060 10192
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 19432 9868 19484 9920
rect 20628 10004 20680 10056
rect 20168 9979 20220 9988
rect 20168 9945 20177 9979
rect 20177 9945 20211 9979
rect 20211 9945 20220 9979
rect 21088 10072 21140 10124
rect 21640 10072 21692 10124
rect 21180 10004 21232 10056
rect 21456 10004 21508 10056
rect 20168 9936 20220 9945
rect 21548 9936 21600 9988
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 22836 10115 22888 10124
rect 22836 10081 22845 10115
rect 22845 10081 22879 10115
rect 22879 10081 22888 10115
rect 22836 10072 22888 10081
rect 22928 10047 22980 10056
rect 22928 10013 22937 10047
rect 22937 10013 22971 10047
rect 22971 10013 22980 10047
rect 22928 10004 22980 10013
rect 23204 10047 23256 10056
rect 23204 10013 23214 10047
rect 23214 10013 23248 10047
rect 23248 10013 23256 10047
rect 23204 10004 23256 10013
rect 23388 10072 23440 10124
rect 25412 10140 25464 10192
rect 24308 10072 24360 10124
rect 28448 10208 28500 10260
rect 29092 10208 29144 10260
rect 23756 10047 23808 10056
rect 23756 10013 23765 10047
rect 23765 10013 23799 10047
rect 23799 10013 23808 10047
rect 23756 10004 23808 10013
rect 24032 10047 24084 10056
rect 24032 10013 24041 10047
rect 24041 10013 24075 10047
rect 24075 10013 24084 10047
rect 24032 10004 24084 10013
rect 28264 10072 28316 10124
rect 28540 10072 28592 10124
rect 26148 10047 26200 10056
rect 26148 10013 26157 10047
rect 26157 10013 26191 10047
rect 26191 10013 26200 10047
rect 26148 10004 26200 10013
rect 27712 10004 27764 10056
rect 28356 10004 28408 10056
rect 29368 10004 29420 10056
rect 29920 10072 29972 10124
rect 30656 10208 30708 10260
rect 33048 10208 33100 10260
rect 33140 10208 33192 10260
rect 33232 10208 33284 10260
rect 34060 10208 34112 10260
rect 34336 10208 34388 10260
rect 35808 10251 35860 10260
rect 35808 10217 35817 10251
rect 35817 10217 35851 10251
rect 35851 10217 35860 10251
rect 35808 10208 35860 10217
rect 35900 10251 35952 10260
rect 35900 10217 35909 10251
rect 35909 10217 35943 10251
rect 35943 10217 35952 10251
rect 35900 10208 35952 10217
rect 35992 10208 36044 10260
rect 36544 10208 36596 10260
rect 38384 10208 38436 10260
rect 39948 10208 40000 10260
rect 41788 10208 41840 10260
rect 41880 10208 41932 10260
rect 42984 10251 43036 10260
rect 29552 10004 29604 10056
rect 21732 9911 21784 9920
rect 21732 9877 21741 9911
rect 21741 9877 21775 9911
rect 21775 9877 21784 9911
rect 21732 9868 21784 9877
rect 21824 9868 21876 9920
rect 22284 9868 22336 9920
rect 23296 9868 23348 9920
rect 25688 9936 25740 9988
rect 23848 9868 23900 9920
rect 24400 9868 24452 9920
rect 25136 9868 25188 9920
rect 29000 9936 29052 9988
rect 29276 9936 29328 9988
rect 30288 10115 30340 10124
rect 30288 10081 30297 10115
rect 30297 10081 30331 10115
rect 30331 10081 30340 10115
rect 30288 10072 30340 10081
rect 31760 10072 31812 10124
rect 32864 10140 32916 10192
rect 30288 9936 30340 9988
rect 27988 9868 28040 9920
rect 30656 10004 30708 10056
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 32036 10004 32088 10056
rect 30932 9936 30984 9988
rect 32772 10004 32824 10056
rect 32864 9936 32916 9988
rect 33600 10072 33652 10124
rect 35716 10072 35768 10124
rect 32588 9911 32640 9920
rect 32588 9877 32597 9911
rect 32597 9877 32631 9911
rect 32631 9877 32640 9911
rect 32588 9868 32640 9877
rect 32956 9911 33008 9920
rect 32956 9877 32965 9911
rect 32965 9877 32999 9911
rect 32999 9877 33008 9911
rect 32956 9868 33008 9877
rect 33508 9936 33560 9988
rect 36268 10047 36320 10056
rect 36268 10013 36277 10047
rect 36277 10013 36311 10047
rect 36311 10013 36320 10047
rect 36268 10004 36320 10013
rect 36912 10047 36964 10056
rect 36912 10013 36921 10047
rect 36921 10013 36955 10047
rect 36955 10013 36964 10047
rect 36912 10004 36964 10013
rect 39028 10140 39080 10192
rect 38660 10004 38712 10056
rect 39304 10072 39356 10124
rect 39396 10072 39448 10124
rect 39120 10004 39172 10056
rect 40316 10004 40368 10056
rect 40408 10004 40460 10056
rect 34428 9936 34480 9988
rect 34888 9936 34940 9988
rect 35624 9936 35676 9988
rect 40776 9936 40828 9988
rect 42524 9936 42576 9988
rect 35348 9868 35400 9920
rect 36728 9911 36780 9920
rect 36728 9877 36737 9911
rect 36737 9877 36771 9911
rect 36771 9877 36780 9911
rect 36728 9868 36780 9877
rect 37004 9911 37056 9920
rect 37004 9877 37013 9911
rect 37013 9877 37047 9911
rect 37047 9877 37056 9911
rect 37004 9868 37056 9877
rect 37280 9911 37332 9920
rect 37280 9877 37289 9911
rect 37289 9877 37323 9911
rect 37323 9877 37332 9911
rect 37280 9868 37332 9877
rect 37924 9911 37976 9920
rect 37924 9877 37933 9911
rect 37933 9877 37967 9911
rect 37967 9877 37976 9911
rect 37924 9868 37976 9877
rect 38016 9911 38068 9920
rect 38016 9877 38025 9911
rect 38025 9877 38059 9911
rect 38059 9877 38068 9911
rect 38016 9868 38068 9877
rect 39672 9868 39724 9920
rect 40408 9868 40460 9920
rect 40960 9868 41012 9920
rect 42984 10217 42993 10251
rect 42993 10217 43027 10251
rect 43027 10217 43036 10251
rect 42984 10208 43036 10217
rect 44548 10251 44600 10260
rect 44548 10217 44557 10251
rect 44557 10217 44591 10251
rect 44591 10217 44600 10251
rect 44548 10208 44600 10217
rect 43260 10183 43312 10192
rect 43260 10149 43269 10183
rect 43269 10149 43303 10183
rect 43303 10149 43312 10183
rect 43260 10140 43312 10149
rect 44824 10140 44876 10192
rect 6070 9766 6122 9818
rect 6134 9766 6186 9818
rect 6198 9766 6250 9818
rect 6262 9766 6314 9818
rect 6326 9766 6378 9818
rect 11070 9766 11122 9818
rect 11134 9766 11186 9818
rect 11198 9766 11250 9818
rect 11262 9766 11314 9818
rect 11326 9766 11378 9818
rect 16070 9766 16122 9818
rect 16134 9766 16186 9818
rect 16198 9766 16250 9818
rect 16262 9766 16314 9818
rect 16326 9766 16378 9818
rect 21070 9766 21122 9818
rect 21134 9766 21186 9818
rect 21198 9766 21250 9818
rect 21262 9766 21314 9818
rect 21326 9766 21378 9818
rect 26070 9766 26122 9818
rect 26134 9766 26186 9818
rect 26198 9766 26250 9818
rect 26262 9766 26314 9818
rect 26326 9766 26378 9818
rect 31070 9766 31122 9818
rect 31134 9766 31186 9818
rect 31198 9766 31250 9818
rect 31262 9766 31314 9818
rect 31326 9766 31378 9818
rect 36070 9766 36122 9818
rect 36134 9766 36186 9818
rect 36198 9766 36250 9818
rect 36262 9766 36314 9818
rect 36326 9766 36378 9818
rect 41070 9766 41122 9818
rect 41134 9766 41186 9818
rect 41198 9766 41250 9818
rect 41262 9766 41314 9818
rect 41326 9766 41378 9818
rect 3424 9664 3476 9716
rect 4344 9664 4396 9716
rect 4436 9664 4488 9716
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 5908 9664 5960 9716
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 7748 9596 7800 9648
rect 5264 9460 5316 9512
rect 5356 9460 5408 9512
rect 8024 9664 8076 9716
rect 8300 9664 8352 9716
rect 9128 9664 9180 9716
rect 10140 9707 10192 9716
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 13268 9664 13320 9716
rect 13452 9664 13504 9716
rect 13544 9664 13596 9716
rect 14188 9664 14240 9716
rect 15108 9664 15160 9716
rect 5080 9324 5132 9376
rect 6092 9324 6144 9376
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 8208 9460 8260 9512
rect 9588 9528 9640 9580
rect 10600 9596 10652 9648
rect 12072 9596 12124 9648
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12532 9596 12584 9648
rect 10048 9460 10100 9512
rect 12716 9528 12768 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 12900 9528 12952 9580
rect 13360 9639 13412 9648
rect 13360 9605 13369 9639
rect 13369 9605 13403 9639
rect 13403 9605 13412 9639
rect 13360 9596 13412 9605
rect 16580 9664 16632 9716
rect 17132 9664 17184 9716
rect 16948 9596 17000 9648
rect 12348 9460 12400 9512
rect 13360 9460 13412 9512
rect 7012 9324 7064 9333
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 11520 9324 11572 9376
rect 11980 9324 12032 9376
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 12900 9324 12952 9376
rect 14004 9324 14056 9376
rect 15384 9460 15436 9512
rect 16856 9528 16908 9580
rect 18420 9664 18472 9716
rect 20812 9664 20864 9716
rect 17684 9596 17736 9648
rect 18052 9596 18104 9648
rect 19156 9596 19208 9648
rect 20352 9639 20404 9648
rect 20352 9605 20361 9639
rect 20361 9605 20395 9639
rect 20395 9605 20404 9639
rect 20352 9596 20404 9605
rect 21272 9596 21324 9648
rect 15016 9392 15068 9444
rect 19248 9503 19300 9512
rect 19248 9469 19257 9503
rect 19257 9469 19291 9503
rect 19291 9469 19300 9503
rect 19248 9460 19300 9469
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 20904 9528 20956 9580
rect 21824 9664 21876 9716
rect 19340 9435 19392 9444
rect 19340 9401 19349 9435
rect 19349 9401 19383 9435
rect 19383 9401 19392 9435
rect 19340 9392 19392 9401
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 18972 9324 19024 9376
rect 19984 9392 20036 9444
rect 21732 9460 21784 9512
rect 21180 9435 21232 9444
rect 21180 9401 21189 9435
rect 21189 9401 21223 9435
rect 21223 9401 21232 9435
rect 21180 9392 21232 9401
rect 21548 9392 21600 9444
rect 20444 9324 20496 9376
rect 21824 9324 21876 9376
rect 22284 9664 22336 9716
rect 23756 9664 23808 9716
rect 24400 9707 24452 9716
rect 24400 9673 24409 9707
rect 24409 9673 24443 9707
rect 24443 9673 24452 9707
rect 24400 9664 24452 9673
rect 24584 9664 24636 9716
rect 24952 9664 25004 9716
rect 25412 9664 25464 9716
rect 23112 9596 23164 9648
rect 22008 9528 22060 9580
rect 23848 9596 23900 9648
rect 22376 9460 22428 9512
rect 23020 9460 23072 9512
rect 23204 9392 23256 9444
rect 22192 9324 22244 9376
rect 22836 9324 22888 9376
rect 23940 9460 23992 9512
rect 23480 9392 23532 9444
rect 24768 9460 24820 9512
rect 25596 9639 25648 9648
rect 25596 9605 25605 9639
rect 25605 9605 25639 9639
rect 25639 9605 25648 9639
rect 25596 9596 25648 9605
rect 25688 9596 25740 9648
rect 27712 9664 27764 9716
rect 29736 9664 29788 9716
rect 25044 9460 25096 9512
rect 25228 9460 25280 9512
rect 26700 9503 26752 9512
rect 26700 9469 26709 9503
rect 26709 9469 26743 9503
rect 26743 9469 26752 9503
rect 26700 9460 26752 9469
rect 27620 9503 27672 9512
rect 27620 9469 27629 9503
rect 27629 9469 27663 9503
rect 27663 9469 27672 9503
rect 27620 9460 27672 9469
rect 27988 9571 28040 9580
rect 27988 9537 27997 9571
rect 27997 9537 28031 9571
rect 28031 9537 28040 9571
rect 27988 9528 28040 9537
rect 28172 9460 28224 9512
rect 29368 9460 29420 9512
rect 30196 9596 30248 9648
rect 30380 9639 30432 9648
rect 30380 9605 30389 9639
rect 30389 9605 30423 9639
rect 30423 9605 30432 9639
rect 30380 9596 30432 9605
rect 30472 9596 30524 9648
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 29920 9528 29972 9580
rect 30012 9460 30064 9512
rect 23940 9324 23992 9376
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 29920 9392 29972 9444
rect 30380 9392 30432 9444
rect 31944 9664 31996 9716
rect 32496 9707 32548 9716
rect 32496 9673 32505 9707
rect 32505 9673 32539 9707
rect 32539 9673 32548 9707
rect 32496 9664 32548 9673
rect 32956 9707 33008 9716
rect 32956 9673 32965 9707
rect 32965 9673 32999 9707
rect 32999 9673 33008 9707
rect 32956 9664 33008 9673
rect 33048 9664 33100 9716
rect 34520 9664 34572 9716
rect 34888 9664 34940 9716
rect 31576 9596 31628 9648
rect 33968 9639 34020 9648
rect 33968 9605 33993 9639
rect 33993 9605 34020 9639
rect 33968 9596 34020 9605
rect 35072 9596 35124 9648
rect 36452 9664 36504 9716
rect 38660 9664 38712 9716
rect 40408 9664 40460 9716
rect 32036 9528 32088 9580
rect 33232 9528 33284 9580
rect 33324 9571 33376 9580
rect 33324 9537 33333 9571
rect 33333 9537 33367 9571
rect 33367 9537 33376 9571
rect 33324 9528 33376 9537
rect 32772 9460 32824 9512
rect 34336 9460 34388 9512
rect 30748 9435 30800 9444
rect 30748 9401 30757 9435
rect 30757 9401 30791 9435
rect 30791 9401 30800 9435
rect 30748 9392 30800 9401
rect 31208 9435 31260 9444
rect 31208 9401 31217 9435
rect 31217 9401 31251 9435
rect 31251 9401 31260 9435
rect 31208 9392 31260 9401
rect 29736 9324 29788 9376
rect 29828 9324 29880 9376
rect 31852 9367 31904 9376
rect 31852 9333 31861 9367
rect 31861 9333 31895 9367
rect 31895 9333 31904 9367
rect 31852 9324 31904 9333
rect 32036 9367 32088 9376
rect 32036 9333 32045 9367
rect 32045 9333 32079 9367
rect 32079 9333 32088 9367
rect 32036 9324 32088 9333
rect 32128 9324 32180 9376
rect 32864 9324 32916 9376
rect 33968 9367 34020 9376
rect 33968 9333 33977 9367
rect 33977 9333 34011 9367
rect 34011 9333 34020 9367
rect 33968 9324 34020 9333
rect 34796 9460 34848 9512
rect 34888 9460 34940 9512
rect 35808 9460 35860 9512
rect 36820 9639 36872 9648
rect 36820 9605 36845 9639
rect 36845 9605 36872 9639
rect 36820 9596 36872 9605
rect 37280 9596 37332 9648
rect 37464 9596 37516 9648
rect 41788 9664 41840 9716
rect 42984 9707 43036 9716
rect 42984 9673 42993 9707
rect 42993 9673 43027 9707
rect 43027 9673 43036 9707
rect 42984 9664 43036 9673
rect 43260 9664 43312 9716
rect 41512 9596 41564 9648
rect 37096 9571 37148 9580
rect 37096 9537 37105 9571
rect 37105 9537 37139 9571
rect 37139 9537 37148 9571
rect 37096 9528 37148 9537
rect 36636 9460 36688 9512
rect 40132 9460 40184 9512
rect 40868 9528 40920 9580
rect 42708 9528 42760 9580
rect 44640 9528 44692 9580
rect 38476 9392 38528 9444
rect 41696 9460 41748 9512
rect 41972 9503 42024 9512
rect 41972 9469 41981 9503
rect 41981 9469 42015 9503
rect 42015 9469 42024 9503
rect 41972 9460 42024 9469
rect 42616 9460 42668 9512
rect 42064 9392 42116 9444
rect 35900 9324 35952 9376
rect 37188 9324 37240 9376
rect 39764 9367 39816 9376
rect 39764 9333 39773 9367
rect 39773 9333 39807 9367
rect 39807 9333 39816 9367
rect 39764 9324 39816 9333
rect 44732 9435 44784 9444
rect 44732 9401 44741 9435
rect 44741 9401 44775 9435
rect 44775 9401 44784 9435
rect 44732 9392 44784 9401
rect 44548 9324 44600 9376
rect 3570 9222 3622 9274
rect 3634 9222 3686 9274
rect 3698 9222 3750 9274
rect 3762 9222 3814 9274
rect 3826 9222 3878 9274
rect 8570 9222 8622 9274
rect 8634 9222 8686 9274
rect 8698 9222 8750 9274
rect 8762 9222 8814 9274
rect 8826 9222 8878 9274
rect 13570 9222 13622 9274
rect 13634 9222 13686 9274
rect 13698 9222 13750 9274
rect 13762 9222 13814 9274
rect 13826 9222 13878 9274
rect 18570 9222 18622 9274
rect 18634 9222 18686 9274
rect 18698 9222 18750 9274
rect 18762 9222 18814 9274
rect 18826 9222 18878 9274
rect 23570 9222 23622 9274
rect 23634 9222 23686 9274
rect 23698 9222 23750 9274
rect 23762 9222 23814 9274
rect 23826 9222 23878 9274
rect 28570 9222 28622 9274
rect 28634 9222 28686 9274
rect 28698 9222 28750 9274
rect 28762 9222 28814 9274
rect 28826 9222 28878 9274
rect 33570 9222 33622 9274
rect 33634 9222 33686 9274
rect 33698 9222 33750 9274
rect 33762 9222 33814 9274
rect 33826 9222 33878 9274
rect 38570 9222 38622 9274
rect 38634 9222 38686 9274
rect 38698 9222 38750 9274
rect 38762 9222 38814 9274
rect 38826 9222 38878 9274
rect 43570 9222 43622 9274
rect 43634 9222 43686 9274
rect 43698 9222 43750 9274
rect 43762 9222 43814 9274
rect 43826 9222 43878 9274
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 6644 9163 6696 9172
rect 6644 9129 6653 9163
rect 6653 9129 6687 9163
rect 6687 9129 6696 9163
rect 6644 9120 6696 9129
rect 6920 9120 6972 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8208 9120 8260 9172
rect 8484 9120 8536 9172
rect 9036 9120 9088 9172
rect 10508 9120 10560 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11980 9120 12032 9172
rect 12716 9120 12768 9172
rect 13360 9120 13412 9172
rect 9956 9095 10008 9104
rect 9956 9061 9965 9095
rect 9965 9061 9999 9095
rect 9999 9061 10008 9095
rect 9956 9052 10008 9061
rect 10048 9052 10100 9104
rect 10324 9052 10376 9104
rect 12992 9095 13044 9104
rect 12992 9061 13001 9095
rect 13001 9061 13035 9095
rect 13035 9061 13044 9095
rect 12992 9052 13044 9061
rect 15016 9120 15068 9172
rect 19248 9120 19300 9172
rect 21548 9163 21600 9172
rect 14188 9095 14240 9104
rect 14188 9061 14197 9095
rect 14197 9061 14231 9095
rect 14231 9061 14240 9095
rect 14188 9052 14240 9061
rect 13452 8984 13504 9036
rect 13820 8984 13872 9036
rect 15200 8984 15252 9036
rect 18236 8984 18288 9036
rect 18972 8984 19024 9036
rect 4160 8916 4212 8968
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 6000 8848 6052 8900
rect 8392 8848 8444 8900
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 8944 8916 8996 8968
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 9496 8916 9548 8968
rect 9680 8916 9732 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 940 8823 992 8832
rect 940 8789 949 8823
rect 949 8789 983 8823
rect 983 8789 992 8823
rect 940 8780 992 8789
rect 7012 8780 7064 8832
rect 8484 8780 8536 8832
rect 9312 8848 9364 8900
rect 9588 8780 9640 8832
rect 10140 8823 10192 8832
rect 10140 8789 10149 8823
rect 10149 8789 10183 8823
rect 10183 8789 10192 8823
rect 10140 8780 10192 8789
rect 12900 8916 12952 8968
rect 13360 8916 13412 8968
rect 14004 8959 14056 8968
rect 14004 8925 14013 8959
rect 14013 8925 14047 8959
rect 14047 8925 14056 8959
rect 14004 8916 14056 8925
rect 11704 8848 11756 8900
rect 11888 8848 11940 8900
rect 12716 8848 12768 8900
rect 13084 8848 13136 8900
rect 13176 8891 13228 8900
rect 13176 8857 13185 8891
rect 13185 8857 13219 8891
rect 13219 8857 13228 8891
rect 13176 8848 13228 8857
rect 13544 8848 13596 8900
rect 12440 8780 12492 8832
rect 12808 8780 12860 8832
rect 14464 8780 14516 8832
rect 15016 8780 15068 8832
rect 15108 8780 15160 8832
rect 15384 8780 15436 8832
rect 16580 8916 16632 8968
rect 19432 8916 19484 8968
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 22928 9120 22980 9172
rect 23020 9120 23072 9172
rect 19616 9052 19668 9104
rect 23296 9095 23348 9104
rect 23296 9061 23305 9095
rect 23305 9061 23339 9095
rect 23339 9061 23348 9095
rect 23296 9052 23348 9061
rect 23664 9120 23716 9172
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 25320 9120 25372 9172
rect 25964 9120 26016 9172
rect 26700 9120 26752 9172
rect 27528 9120 27580 9172
rect 27896 9120 27948 9172
rect 29184 9163 29236 9172
rect 29184 9129 29193 9163
rect 29193 9129 29227 9163
rect 29227 9129 29236 9163
rect 29184 9120 29236 9129
rect 29552 9120 29604 9172
rect 29920 9120 29972 9172
rect 30472 9120 30524 9172
rect 31576 9120 31628 9172
rect 25136 9052 25188 9104
rect 31668 9052 31720 9104
rect 32036 9052 32088 9104
rect 19800 8959 19852 8968
rect 19800 8925 19809 8959
rect 19809 8925 19843 8959
rect 19843 8925 19852 8959
rect 19800 8916 19852 8925
rect 21548 8916 21600 8968
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 22376 8916 22428 8968
rect 22560 8916 22612 8968
rect 22652 8916 22704 8968
rect 23940 8984 23992 9036
rect 24860 8984 24912 9036
rect 25780 8984 25832 9036
rect 27436 8984 27488 9036
rect 28080 8984 28132 9036
rect 22836 8916 22888 8968
rect 16856 8848 16908 8900
rect 17500 8848 17552 8900
rect 15844 8823 15896 8832
rect 15844 8789 15853 8823
rect 15853 8789 15887 8823
rect 15887 8789 15896 8823
rect 15844 8780 15896 8789
rect 15936 8780 15988 8832
rect 20168 8848 20220 8900
rect 18512 8780 18564 8832
rect 21732 8848 21784 8900
rect 23204 8916 23256 8968
rect 25228 8959 25280 8968
rect 25228 8925 25237 8959
rect 25237 8925 25271 8959
rect 25271 8925 25280 8959
rect 25228 8916 25280 8925
rect 23388 8780 23440 8832
rect 24492 8848 24544 8900
rect 25504 8848 25556 8900
rect 24400 8780 24452 8832
rect 24952 8823 25004 8832
rect 24952 8789 24961 8823
rect 24961 8789 24995 8823
rect 24995 8789 25004 8823
rect 24952 8780 25004 8789
rect 25320 8780 25372 8832
rect 25964 8823 26016 8832
rect 25964 8789 25973 8823
rect 25973 8789 26007 8823
rect 26007 8789 26016 8823
rect 25964 8780 26016 8789
rect 29828 8984 29880 9036
rect 30288 8984 30340 9036
rect 31300 8984 31352 9036
rect 31484 8984 31536 9036
rect 31852 8984 31904 9036
rect 32772 9120 32824 9172
rect 33140 9120 33192 9172
rect 33416 9120 33468 9172
rect 33968 9120 34020 9172
rect 35900 9163 35952 9172
rect 35900 9129 35909 9163
rect 35909 9129 35943 9163
rect 35943 9129 35952 9163
rect 35900 9120 35952 9129
rect 35992 9120 36044 9172
rect 36176 9120 36228 9172
rect 32220 9052 32272 9104
rect 32404 8984 32456 9036
rect 34336 9052 34388 9104
rect 34888 9095 34940 9104
rect 34888 9061 34897 9095
rect 34897 9061 34931 9095
rect 34931 9061 34940 9095
rect 34888 9052 34940 9061
rect 34980 9052 35032 9104
rect 26516 8891 26568 8900
rect 26516 8857 26525 8891
rect 26525 8857 26559 8891
rect 26559 8857 26568 8891
rect 26516 8848 26568 8857
rect 26884 8848 26936 8900
rect 26976 8891 27028 8900
rect 26976 8857 26985 8891
rect 26985 8857 27019 8891
rect 27019 8857 27028 8891
rect 26976 8848 27028 8857
rect 27988 8848 28040 8900
rect 27620 8780 27672 8832
rect 30012 8848 30064 8900
rect 28448 8823 28500 8832
rect 28448 8789 28457 8823
rect 28457 8789 28491 8823
rect 28491 8789 28500 8823
rect 28448 8780 28500 8789
rect 28724 8780 28776 8832
rect 29184 8780 29236 8832
rect 30104 8780 30156 8832
rect 30380 8780 30432 8832
rect 32588 8916 32640 8968
rect 33232 8984 33284 9036
rect 33600 8984 33652 9036
rect 34428 8984 34480 9036
rect 35532 9027 35584 9036
rect 35532 8993 35541 9027
rect 35541 8993 35575 9027
rect 35575 8993 35584 9027
rect 35532 8984 35584 8993
rect 38016 9120 38068 9172
rect 39764 9120 39816 9172
rect 43260 9120 43312 9172
rect 35440 8916 35492 8968
rect 31484 8780 31536 8832
rect 32128 8780 32180 8832
rect 32496 8823 32548 8832
rect 32496 8789 32505 8823
rect 32505 8789 32539 8823
rect 32539 8789 32548 8823
rect 32496 8780 32548 8789
rect 33048 8848 33100 8900
rect 33600 8848 33652 8900
rect 34336 8848 34388 8900
rect 34980 8848 35032 8900
rect 37004 9027 37056 9036
rect 37004 8993 37013 9027
rect 37013 8993 37047 9027
rect 37047 8993 37056 9027
rect 37004 8984 37056 8993
rect 37096 8984 37148 9036
rect 33232 8780 33284 8832
rect 34428 8823 34480 8832
rect 34428 8789 34437 8823
rect 34437 8789 34471 8823
rect 34471 8789 34480 8823
rect 34428 8780 34480 8789
rect 35808 8848 35860 8900
rect 36544 8916 36596 8968
rect 36636 8916 36688 8968
rect 38292 8916 38344 8968
rect 40592 8984 40644 9036
rect 39672 8916 39724 8968
rect 39764 8959 39816 8968
rect 39764 8925 39773 8959
rect 39773 8925 39807 8959
rect 39807 8925 39816 8959
rect 39764 8916 39816 8925
rect 36176 8891 36228 8900
rect 36176 8857 36185 8891
rect 36185 8857 36219 8891
rect 36219 8857 36228 8891
rect 36176 8848 36228 8857
rect 37464 8848 37516 8900
rect 41512 8916 41564 8968
rect 35624 8780 35676 8832
rect 36544 8780 36596 8832
rect 38844 8823 38896 8832
rect 38844 8789 38853 8823
rect 38853 8789 38887 8823
rect 38887 8789 38896 8823
rect 38844 8780 38896 8789
rect 42524 8848 42576 8900
rect 40960 8780 41012 8832
rect 41880 8780 41932 8832
rect 44548 8823 44600 8832
rect 44548 8789 44557 8823
rect 44557 8789 44591 8823
rect 44591 8789 44600 8823
rect 44548 8780 44600 8789
rect 44916 8823 44968 8832
rect 44916 8789 44925 8823
rect 44925 8789 44959 8823
rect 44959 8789 44968 8823
rect 44916 8780 44968 8789
rect 6070 8678 6122 8730
rect 6134 8678 6186 8730
rect 6198 8678 6250 8730
rect 6262 8678 6314 8730
rect 6326 8678 6378 8730
rect 11070 8678 11122 8730
rect 11134 8678 11186 8730
rect 11198 8678 11250 8730
rect 11262 8678 11314 8730
rect 11326 8678 11378 8730
rect 16070 8678 16122 8730
rect 16134 8678 16186 8730
rect 16198 8678 16250 8730
rect 16262 8678 16314 8730
rect 16326 8678 16378 8730
rect 21070 8678 21122 8730
rect 21134 8678 21186 8730
rect 21198 8678 21250 8730
rect 21262 8678 21314 8730
rect 21326 8678 21378 8730
rect 26070 8678 26122 8730
rect 26134 8678 26186 8730
rect 26198 8678 26250 8730
rect 26262 8678 26314 8730
rect 26326 8678 26378 8730
rect 31070 8678 31122 8730
rect 31134 8678 31186 8730
rect 31198 8678 31250 8730
rect 31262 8678 31314 8730
rect 31326 8678 31378 8730
rect 36070 8678 36122 8730
rect 36134 8678 36186 8730
rect 36198 8678 36250 8730
rect 36262 8678 36314 8730
rect 36326 8678 36378 8730
rect 41070 8678 41122 8730
rect 41134 8678 41186 8730
rect 41198 8678 41250 8730
rect 41262 8678 41314 8730
rect 41326 8678 41378 8730
rect 6000 8619 6052 8628
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 6644 8576 6696 8628
rect 7656 8619 7708 8628
rect 7656 8585 7665 8619
rect 7665 8585 7699 8619
rect 7699 8585 7708 8619
rect 7656 8576 7708 8585
rect 8208 8576 8260 8628
rect 10140 8576 10192 8628
rect 8944 8508 8996 8560
rect 10324 8440 10376 8492
rect 11244 8576 11296 8628
rect 12072 8576 12124 8628
rect 13268 8576 13320 8628
rect 11796 8508 11848 8560
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 9312 8372 9364 8424
rect 9588 8372 9640 8424
rect 10416 8304 10468 8356
rect 12440 8483 12492 8492
rect 11704 8372 11756 8424
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 12716 8440 12768 8492
rect 13084 8508 13136 8560
rect 13452 8508 13504 8560
rect 13636 8508 13688 8560
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 17224 8576 17276 8628
rect 18052 8576 18104 8628
rect 16580 8508 16632 8560
rect 12532 8372 12584 8424
rect 13636 8372 13688 8424
rect 14188 8372 14240 8424
rect 12808 8304 12860 8356
rect 15292 8440 15344 8492
rect 16672 8440 16724 8492
rect 17224 8440 17276 8492
rect 17316 8440 17368 8492
rect 17960 8508 18012 8560
rect 19156 8619 19208 8628
rect 19156 8585 19165 8619
rect 19165 8585 19199 8619
rect 19199 8585 19208 8619
rect 19156 8576 19208 8585
rect 20260 8576 20312 8628
rect 21548 8576 21600 8628
rect 25228 8576 25280 8628
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 19524 8551 19576 8560
rect 19524 8517 19533 8551
rect 19533 8517 19567 8551
rect 19567 8517 19576 8551
rect 19524 8508 19576 8517
rect 19984 8508 20036 8560
rect 15016 8372 15068 8424
rect 15936 8372 15988 8424
rect 19616 8440 19668 8492
rect 20812 8508 20864 8560
rect 22100 8508 22152 8560
rect 22468 8508 22520 8560
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 23112 8508 23164 8560
rect 9220 8236 9272 8288
rect 10784 8236 10836 8288
rect 10876 8279 10928 8288
rect 10876 8245 10885 8279
rect 10885 8245 10919 8279
rect 10919 8245 10928 8279
rect 10876 8236 10928 8245
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 13176 8236 13228 8288
rect 14280 8236 14332 8288
rect 14740 8304 14792 8356
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 20168 8372 20220 8424
rect 19616 8304 19668 8356
rect 22008 8372 22060 8424
rect 22376 8372 22428 8424
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 15384 8279 15436 8288
rect 15384 8245 15393 8279
rect 15393 8245 15427 8279
rect 15427 8245 15436 8279
rect 15384 8236 15436 8245
rect 16028 8236 16080 8288
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 19524 8236 19576 8288
rect 20168 8279 20220 8288
rect 20168 8245 20177 8279
rect 20177 8245 20211 8279
rect 20211 8245 20220 8279
rect 20168 8236 20220 8245
rect 20720 8304 20772 8356
rect 20996 8304 21048 8356
rect 21916 8347 21968 8356
rect 21916 8313 21925 8347
rect 21925 8313 21959 8347
rect 21959 8313 21968 8347
rect 21916 8304 21968 8313
rect 23480 8415 23532 8424
rect 23480 8381 23489 8415
rect 23489 8381 23523 8415
rect 23523 8381 23532 8415
rect 23480 8372 23532 8381
rect 24400 8508 24452 8560
rect 26792 8508 26844 8560
rect 22744 8347 22796 8356
rect 22744 8313 22753 8347
rect 22753 8313 22787 8347
rect 22787 8313 22796 8347
rect 22744 8304 22796 8313
rect 25688 8440 25740 8492
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 24768 8372 24820 8424
rect 25964 8372 26016 8424
rect 26976 8372 27028 8424
rect 28264 8508 28316 8560
rect 29920 8576 29972 8628
rect 30472 8508 30524 8560
rect 30748 8551 30800 8560
rect 30748 8517 30757 8551
rect 30757 8517 30791 8551
rect 30791 8517 30800 8551
rect 30748 8508 30800 8517
rect 30840 8508 30892 8560
rect 32496 8576 32548 8628
rect 31668 8508 31720 8560
rect 31852 8508 31904 8560
rect 33048 8576 33100 8628
rect 34152 8576 34204 8628
rect 34336 8619 34388 8628
rect 34336 8585 34345 8619
rect 34345 8585 34379 8619
rect 34379 8585 34388 8619
rect 34336 8576 34388 8585
rect 34520 8576 34572 8628
rect 27620 8440 27672 8492
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 27436 8415 27488 8424
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 28356 8372 28408 8424
rect 28540 8372 28592 8424
rect 29828 8440 29880 8492
rect 30012 8440 30064 8492
rect 30380 8483 30432 8492
rect 30380 8449 30389 8483
rect 30389 8449 30423 8483
rect 30423 8449 30432 8483
rect 30380 8440 30432 8449
rect 30656 8440 30708 8492
rect 31392 8440 31444 8492
rect 32404 8440 32456 8492
rect 34060 8508 34112 8560
rect 34520 8483 34572 8492
rect 34520 8449 34529 8483
rect 34529 8449 34563 8483
rect 34563 8449 34572 8483
rect 34520 8440 34572 8449
rect 34796 8508 34848 8560
rect 34888 8551 34940 8560
rect 34888 8517 34897 8551
rect 34897 8517 34931 8551
rect 34931 8517 34940 8551
rect 34888 8508 34940 8517
rect 35808 8576 35860 8628
rect 35348 8508 35400 8560
rect 36176 8508 36228 8560
rect 38752 8576 38804 8628
rect 40960 8576 41012 8628
rect 37372 8508 37424 8560
rect 40040 8508 40092 8560
rect 36636 8483 36688 8492
rect 36636 8449 36645 8483
rect 36645 8449 36679 8483
rect 36679 8449 36688 8483
rect 36636 8440 36688 8449
rect 30288 8415 30340 8424
rect 30288 8381 30297 8415
rect 30297 8381 30331 8415
rect 30331 8381 30340 8415
rect 30288 8372 30340 8381
rect 30840 8372 30892 8424
rect 24032 8236 24084 8288
rect 24124 8236 24176 8288
rect 25044 8236 25096 8288
rect 26884 8279 26936 8288
rect 26884 8245 26893 8279
rect 26893 8245 26927 8279
rect 26927 8245 26936 8279
rect 26884 8236 26936 8245
rect 27252 8236 27304 8288
rect 28448 8236 28500 8288
rect 31668 8304 31720 8356
rect 32220 8415 32272 8424
rect 32220 8381 32229 8415
rect 32229 8381 32263 8415
rect 32263 8381 32272 8415
rect 32220 8372 32272 8381
rect 32312 8415 32364 8424
rect 32312 8381 32321 8415
rect 32321 8381 32355 8415
rect 32355 8381 32364 8415
rect 32312 8372 32364 8381
rect 32864 8372 32916 8424
rect 36084 8372 36136 8424
rect 40224 8508 40276 8560
rect 40592 8440 40644 8492
rect 42524 8508 42576 8560
rect 40776 8483 40828 8492
rect 40776 8449 40785 8483
rect 40785 8449 40819 8483
rect 40819 8449 40828 8483
rect 40776 8440 40828 8449
rect 41420 8483 41472 8492
rect 41420 8449 41429 8483
rect 41429 8449 41463 8483
rect 41463 8449 41472 8483
rect 41420 8440 41472 8449
rect 38200 8372 38252 8424
rect 29368 8236 29420 8288
rect 31208 8236 31260 8288
rect 31760 8236 31812 8288
rect 31852 8279 31904 8288
rect 31852 8245 31861 8279
rect 31861 8245 31895 8279
rect 31895 8245 31904 8279
rect 31852 8236 31904 8245
rect 31944 8236 31996 8288
rect 37096 8236 37148 8288
rect 37556 8236 37608 8288
rect 37924 8236 37976 8288
rect 40132 8372 40184 8424
rect 40684 8372 40736 8424
rect 43444 8372 43496 8424
rect 44916 8415 44968 8424
rect 44916 8381 44925 8415
rect 44925 8381 44959 8415
rect 44959 8381 44968 8415
rect 44916 8372 44968 8381
rect 39764 8304 39816 8356
rect 38384 8279 38436 8288
rect 38384 8245 38393 8279
rect 38393 8245 38427 8279
rect 38427 8245 38436 8279
rect 38384 8236 38436 8245
rect 38844 8236 38896 8288
rect 42800 8236 42852 8288
rect 44548 8236 44600 8288
rect 3570 8134 3622 8186
rect 3634 8134 3686 8186
rect 3698 8134 3750 8186
rect 3762 8134 3814 8186
rect 3826 8134 3878 8186
rect 8570 8134 8622 8186
rect 8634 8134 8686 8186
rect 8698 8134 8750 8186
rect 8762 8134 8814 8186
rect 8826 8134 8878 8186
rect 13570 8134 13622 8186
rect 13634 8134 13686 8186
rect 13698 8134 13750 8186
rect 13762 8134 13814 8186
rect 13826 8134 13878 8186
rect 18570 8134 18622 8186
rect 18634 8134 18686 8186
rect 18698 8134 18750 8186
rect 18762 8134 18814 8186
rect 18826 8134 18878 8186
rect 23570 8134 23622 8186
rect 23634 8134 23686 8186
rect 23698 8134 23750 8186
rect 23762 8134 23814 8186
rect 23826 8134 23878 8186
rect 28570 8134 28622 8186
rect 28634 8134 28686 8186
rect 28698 8134 28750 8186
rect 28762 8134 28814 8186
rect 28826 8134 28878 8186
rect 33570 8134 33622 8186
rect 33634 8134 33686 8186
rect 33698 8134 33750 8186
rect 33762 8134 33814 8186
rect 33826 8134 33878 8186
rect 38570 8134 38622 8186
rect 38634 8134 38686 8186
rect 38698 8134 38750 8186
rect 38762 8134 38814 8186
rect 38826 8134 38878 8186
rect 43570 8134 43622 8186
rect 43634 8134 43686 8186
rect 43698 8134 43750 8186
rect 43762 8134 43814 8186
rect 43826 8134 43878 8186
rect 8484 8032 8536 8084
rect 8944 8032 8996 8084
rect 8392 7828 8444 7880
rect 9312 7964 9364 8016
rect 10140 8032 10192 8084
rect 10508 8032 10560 8084
rect 10048 7964 10100 8016
rect 9588 7896 9640 7948
rect 10876 7896 10928 7948
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 11888 8032 11940 8084
rect 12900 8032 12952 8084
rect 13360 8032 13412 8084
rect 12716 7964 12768 8016
rect 14924 8032 14976 8084
rect 18236 8075 18288 8084
rect 18236 8041 18245 8075
rect 18245 8041 18279 8075
rect 18279 8041 18288 8075
rect 18236 8032 18288 8041
rect 20628 8032 20680 8084
rect 22192 8032 22244 8084
rect 23296 8032 23348 8084
rect 24860 8032 24912 8084
rect 25504 8032 25556 8084
rect 27620 8032 27672 8084
rect 12440 7828 12492 7880
rect 12624 7828 12676 7880
rect 22560 8007 22612 8016
rect 22560 7973 22569 8007
rect 22569 7973 22603 8007
rect 22603 7973 22612 8007
rect 22560 7964 22612 7973
rect 10600 7760 10652 7812
rect 13176 7896 13228 7948
rect 14280 7896 14332 7948
rect 16764 7896 16816 7948
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 20628 7896 20680 7948
rect 21456 7896 21508 7948
rect 15384 7828 15436 7880
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 17408 7828 17460 7880
rect 17500 7828 17552 7880
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 20536 7828 20588 7880
rect 13176 7760 13228 7812
rect 10416 7692 10468 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 12532 7735 12584 7744
rect 12532 7701 12541 7735
rect 12541 7701 12575 7735
rect 12575 7701 12584 7735
rect 12532 7692 12584 7701
rect 12992 7692 13044 7744
rect 14464 7760 14516 7812
rect 15200 7760 15252 7812
rect 16488 7760 16540 7812
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 15844 7735 15896 7744
rect 15844 7701 15859 7735
rect 15859 7701 15893 7735
rect 15893 7701 15896 7735
rect 15844 7692 15896 7701
rect 16764 7692 16816 7744
rect 17408 7692 17460 7744
rect 18880 7803 18932 7812
rect 18880 7769 18889 7803
rect 18889 7769 18923 7803
rect 18923 7769 18932 7803
rect 18880 7760 18932 7769
rect 19892 7760 19944 7812
rect 20444 7760 20496 7812
rect 20904 7760 20956 7812
rect 22284 7760 22336 7812
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 22836 7828 22888 7880
rect 24124 7939 24176 7948
rect 24124 7905 24133 7939
rect 24133 7905 24167 7939
rect 24167 7905 24176 7939
rect 24124 7896 24176 7905
rect 24492 7896 24544 7948
rect 28448 8032 28500 8084
rect 22652 7760 22704 7812
rect 18052 7692 18104 7744
rect 21824 7692 21876 7744
rect 23020 7692 23072 7744
rect 23480 7692 23532 7744
rect 24216 7692 24268 7744
rect 25688 7828 25740 7880
rect 27988 7828 28040 7880
rect 28448 7871 28500 7880
rect 28448 7837 28457 7871
rect 28457 7837 28491 7871
rect 28491 7837 28500 7871
rect 29184 7964 29236 8016
rect 28816 7896 28868 7948
rect 29092 7939 29144 7948
rect 29092 7905 29101 7939
rect 29101 7905 29135 7939
rect 29135 7905 29144 7939
rect 29092 7896 29144 7905
rect 31208 8032 31260 8084
rect 31668 8032 31720 8084
rect 31852 8032 31904 8084
rect 32864 8032 32916 8084
rect 34244 8032 34296 8084
rect 36728 8032 36780 8084
rect 36912 8032 36964 8084
rect 37464 8032 37516 8084
rect 38476 8032 38528 8084
rect 41420 8032 41472 8084
rect 43260 8032 43312 8084
rect 29644 7896 29696 7948
rect 30380 7964 30432 8016
rect 30840 7964 30892 8016
rect 28448 7828 28500 7837
rect 29276 7871 29328 7880
rect 29276 7837 29285 7871
rect 29285 7837 29319 7871
rect 29319 7837 29328 7871
rect 29276 7828 29328 7837
rect 29736 7871 29788 7880
rect 29736 7837 29745 7871
rect 29745 7837 29779 7871
rect 29779 7837 29788 7871
rect 29736 7828 29788 7837
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 30288 7896 30340 7948
rect 31760 7964 31812 8016
rect 31300 7896 31352 7948
rect 31392 7896 31444 7948
rect 32036 7896 32088 7948
rect 34060 7964 34112 8016
rect 32956 7896 33008 7948
rect 30748 7871 30800 7880
rect 30748 7837 30757 7871
rect 30757 7837 30791 7871
rect 30791 7837 30800 7871
rect 30748 7828 30800 7837
rect 30840 7871 30892 7880
rect 30840 7837 30849 7871
rect 30849 7837 30883 7871
rect 30883 7837 30892 7871
rect 30840 7828 30892 7837
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 37004 7896 37056 7948
rect 37556 7896 37608 7948
rect 37648 7939 37700 7948
rect 37648 7905 37657 7939
rect 37657 7905 37691 7939
rect 37691 7905 37700 7939
rect 37648 7896 37700 7905
rect 29092 7760 29144 7812
rect 31484 7760 31536 7812
rect 32036 7760 32088 7812
rect 26424 7692 26476 7744
rect 26608 7692 26660 7744
rect 28172 7692 28224 7744
rect 29552 7735 29604 7744
rect 29552 7701 29561 7735
rect 29561 7701 29595 7735
rect 29595 7701 29604 7735
rect 29552 7692 29604 7701
rect 30380 7735 30432 7744
rect 30380 7701 30389 7735
rect 30389 7701 30423 7735
rect 30423 7701 30432 7735
rect 30380 7692 30432 7701
rect 30564 7735 30616 7744
rect 30564 7701 30573 7735
rect 30573 7701 30607 7735
rect 30607 7701 30616 7735
rect 30564 7692 30616 7701
rect 34060 7871 34112 7880
rect 34060 7837 34069 7871
rect 34069 7837 34103 7871
rect 34103 7837 34112 7871
rect 34060 7828 34112 7837
rect 34428 7828 34480 7880
rect 35072 7828 35124 7880
rect 37464 7828 37516 7880
rect 38384 7828 38436 7880
rect 37096 7760 37148 7812
rect 39580 7871 39632 7880
rect 39580 7837 39589 7871
rect 39589 7837 39623 7871
rect 39623 7837 39632 7871
rect 39580 7828 39632 7837
rect 39672 7871 39724 7880
rect 39672 7837 39681 7871
rect 39681 7837 39715 7871
rect 39715 7837 39724 7871
rect 39672 7828 39724 7837
rect 34428 7692 34480 7744
rect 35716 7692 35768 7744
rect 35808 7692 35860 7744
rect 36176 7692 36228 7744
rect 36728 7692 36780 7744
rect 38200 7692 38252 7744
rect 39212 7760 39264 7812
rect 40592 7760 40644 7812
rect 40776 7692 40828 7744
rect 42064 7939 42116 7948
rect 42064 7905 42073 7939
rect 42073 7905 42107 7939
rect 42107 7905 42116 7939
rect 42064 7896 42116 7905
rect 42708 7896 42760 7948
rect 42800 7939 42852 7948
rect 42800 7905 42809 7939
rect 42809 7905 42843 7939
rect 42843 7905 42852 7939
rect 42800 7896 42852 7905
rect 41880 7871 41932 7880
rect 41880 7837 41889 7871
rect 41889 7837 41923 7871
rect 41923 7837 41932 7871
rect 41880 7828 41932 7837
rect 41328 7692 41380 7744
rect 45008 7760 45060 7812
rect 43444 7692 43496 7744
rect 44180 7735 44232 7744
rect 44180 7701 44189 7735
rect 44189 7701 44223 7735
rect 44223 7701 44232 7735
rect 44180 7692 44232 7701
rect 44548 7735 44600 7744
rect 44548 7701 44557 7735
rect 44557 7701 44591 7735
rect 44591 7701 44600 7735
rect 44916 7735 44968 7744
rect 44548 7692 44600 7701
rect 44916 7701 44925 7735
rect 44925 7701 44959 7735
rect 44959 7701 44968 7735
rect 44916 7692 44968 7701
rect 6070 7590 6122 7642
rect 6134 7590 6186 7642
rect 6198 7590 6250 7642
rect 6262 7590 6314 7642
rect 6326 7590 6378 7642
rect 11070 7590 11122 7642
rect 11134 7590 11186 7642
rect 11198 7590 11250 7642
rect 11262 7590 11314 7642
rect 11326 7590 11378 7642
rect 16070 7590 16122 7642
rect 16134 7590 16186 7642
rect 16198 7590 16250 7642
rect 16262 7590 16314 7642
rect 16326 7590 16378 7642
rect 21070 7590 21122 7642
rect 21134 7590 21186 7642
rect 21198 7590 21250 7642
rect 21262 7590 21314 7642
rect 21326 7590 21378 7642
rect 26070 7590 26122 7642
rect 26134 7590 26186 7642
rect 26198 7590 26250 7642
rect 26262 7590 26314 7642
rect 26326 7590 26378 7642
rect 31070 7590 31122 7642
rect 31134 7590 31186 7642
rect 31198 7590 31250 7642
rect 31262 7590 31314 7642
rect 31326 7590 31378 7642
rect 36070 7590 36122 7642
rect 36134 7590 36186 7642
rect 36198 7590 36250 7642
rect 36262 7590 36314 7642
rect 36326 7590 36378 7642
rect 41070 7590 41122 7642
rect 41134 7590 41186 7642
rect 41198 7590 41250 7642
rect 41262 7590 41314 7642
rect 41326 7590 41378 7642
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 7748 7488 7800 7540
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 9220 7488 9272 7540
rect 10048 7488 10100 7540
rect 10600 7488 10652 7540
rect 11428 7488 11480 7540
rect 11888 7488 11940 7540
rect 14464 7488 14516 7540
rect 16672 7488 16724 7540
rect 17592 7488 17644 7540
rect 18880 7488 18932 7540
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 10508 7352 10560 7404
rect 11796 7352 11848 7404
rect 15844 7420 15896 7472
rect 16580 7420 16632 7472
rect 9956 7284 10008 7336
rect 10416 7284 10468 7336
rect 13084 7216 13136 7268
rect 14648 7216 14700 7268
rect 15200 7352 15252 7404
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 17408 7352 17460 7404
rect 17684 7352 17736 7404
rect 17960 7352 18012 7404
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 18604 7420 18656 7472
rect 20168 7488 20220 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 22468 7488 22520 7540
rect 22560 7488 22612 7540
rect 24308 7531 24360 7540
rect 24308 7497 24317 7531
rect 24317 7497 24351 7531
rect 24351 7497 24360 7531
rect 24308 7488 24360 7497
rect 24400 7531 24452 7540
rect 24400 7497 24409 7531
rect 24409 7497 24443 7531
rect 24443 7497 24452 7531
rect 24400 7488 24452 7497
rect 20904 7420 20956 7472
rect 21824 7420 21876 7472
rect 22008 7420 22060 7472
rect 15568 7284 15620 7336
rect 15660 7284 15712 7336
rect 15936 7216 15988 7268
rect 10600 7148 10652 7200
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 13176 7148 13228 7200
rect 15108 7191 15160 7200
rect 15108 7157 15117 7191
rect 15117 7157 15151 7191
rect 15151 7157 15160 7191
rect 15108 7148 15160 7157
rect 15292 7148 15344 7200
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 17040 7148 17092 7200
rect 19800 7284 19852 7336
rect 19892 7284 19944 7336
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 24216 7420 24268 7472
rect 22468 7352 22520 7404
rect 24952 7488 25004 7540
rect 25412 7488 25464 7540
rect 26516 7531 26568 7540
rect 26516 7497 26525 7531
rect 26525 7497 26559 7531
rect 26559 7497 26568 7531
rect 26516 7488 26568 7497
rect 26884 7488 26936 7540
rect 28172 7488 28224 7540
rect 28356 7531 28408 7540
rect 28356 7497 28365 7531
rect 28365 7497 28399 7531
rect 28399 7497 28408 7531
rect 28356 7488 28408 7497
rect 28632 7488 28684 7540
rect 24768 7352 24820 7404
rect 25228 7420 25280 7472
rect 27988 7352 28040 7404
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 23204 7284 23256 7336
rect 24032 7284 24084 7336
rect 25044 7284 25096 7336
rect 25228 7284 25280 7336
rect 26608 7327 26660 7336
rect 26608 7293 26617 7327
rect 26617 7293 26651 7327
rect 26651 7293 26660 7327
rect 26608 7284 26660 7293
rect 29552 7488 29604 7540
rect 30380 7488 30432 7540
rect 31668 7488 31720 7540
rect 31944 7488 31996 7540
rect 32864 7488 32916 7540
rect 34060 7488 34112 7540
rect 34152 7531 34204 7540
rect 34152 7497 34161 7531
rect 34161 7497 34195 7531
rect 34195 7497 34204 7531
rect 34152 7488 34204 7497
rect 34244 7488 34296 7540
rect 34520 7488 34572 7540
rect 35992 7531 36044 7540
rect 35992 7497 36001 7531
rect 36001 7497 36035 7531
rect 36035 7497 36044 7531
rect 35992 7488 36044 7497
rect 38292 7488 38344 7540
rect 30104 7420 30156 7472
rect 31484 7352 31536 7404
rect 32956 7352 33008 7404
rect 18328 7148 18380 7200
rect 22100 7148 22152 7200
rect 22192 7148 22244 7200
rect 23388 7148 23440 7200
rect 27988 7216 28040 7268
rect 25688 7148 25740 7200
rect 28908 7148 28960 7200
rect 29828 7148 29880 7200
rect 30840 7216 30892 7268
rect 31116 7216 31168 7268
rect 34152 7284 34204 7336
rect 34888 7395 34940 7404
rect 34888 7361 34897 7395
rect 34897 7361 34931 7395
rect 34931 7361 34940 7395
rect 34888 7352 34940 7361
rect 37096 7352 37148 7404
rect 35164 7327 35216 7336
rect 35164 7293 35173 7327
rect 35173 7293 35207 7327
rect 35207 7293 35216 7327
rect 35164 7284 35216 7293
rect 37004 7284 37056 7336
rect 37372 7420 37424 7472
rect 39580 7488 39632 7540
rect 40776 7488 40828 7540
rect 43260 7488 43312 7540
rect 44548 7488 44600 7540
rect 37372 7284 37424 7336
rect 37648 7284 37700 7336
rect 37740 7284 37792 7336
rect 33416 7148 33468 7200
rect 34060 7148 34112 7200
rect 36176 7216 36228 7268
rect 34980 7148 35032 7200
rect 37188 7148 37240 7200
rect 38200 7148 38252 7200
rect 40500 7463 40552 7472
rect 40500 7429 40509 7463
rect 40509 7429 40543 7463
rect 40543 7429 40552 7463
rect 40500 7420 40552 7429
rect 44180 7420 44232 7472
rect 44732 7420 44784 7472
rect 39120 7352 39172 7404
rect 39580 7327 39632 7336
rect 39580 7293 39589 7327
rect 39589 7293 39623 7327
rect 39623 7293 39632 7327
rect 39580 7284 39632 7293
rect 41420 7352 41472 7404
rect 41512 7395 41564 7404
rect 41512 7361 41521 7395
rect 41521 7361 41555 7395
rect 41555 7361 41564 7395
rect 41512 7352 41564 7361
rect 43076 7352 43128 7404
rect 40684 7327 40736 7336
rect 40684 7293 40693 7327
rect 40693 7293 40727 7327
rect 40727 7293 40736 7327
rect 40684 7284 40736 7293
rect 42064 7284 42116 7336
rect 44548 7216 44600 7268
rect 39856 7191 39908 7200
rect 39856 7157 39865 7191
rect 39865 7157 39899 7191
rect 39899 7157 39908 7191
rect 39856 7148 39908 7157
rect 40960 7148 41012 7200
rect 41328 7191 41380 7200
rect 41328 7157 41337 7191
rect 41337 7157 41371 7191
rect 41371 7157 41380 7191
rect 41328 7148 41380 7157
rect 41420 7148 41472 7200
rect 41880 7148 41932 7200
rect 43444 7148 43496 7200
rect 3570 7046 3622 7098
rect 3634 7046 3686 7098
rect 3698 7046 3750 7098
rect 3762 7046 3814 7098
rect 3826 7046 3878 7098
rect 8570 7046 8622 7098
rect 8634 7046 8686 7098
rect 8698 7046 8750 7098
rect 8762 7046 8814 7098
rect 8826 7046 8878 7098
rect 13570 7046 13622 7098
rect 13634 7046 13686 7098
rect 13698 7046 13750 7098
rect 13762 7046 13814 7098
rect 13826 7046 13878 7098
rect 18570 7046 18622 7098
rect 18634 7046 18686 7098
rect 18698 7046 18750 7098
rect 18762 7046 18814 7098
rect 18826 7046 18878 7098
rect 23570 7046 23622 7098
rect 23634 7046 23686 7098
rect 23698 7046 23750 7098
rect 23762 7046 23814 7098
rect 23826 7046 23878 7098
rect 28570 7046 28622 7098
rect 28634 7046 28686 7098
rect 28698 7046 28750 7098
rect 28762 7046 28814 7098
rect 28826 7046 28878 7098
rect 33570 7046 33622 7098
rect 33634 7046 33686 7098
rect 33698 7046 33750 7098
rect 33762 7046 33814 7098
rect 33826 7046 33878 7098
rect 38570 7046 38622 7098
rect 38634 7046 38686 7098
rect 38698 7046 38750 7098
rect 38762 7046 38814 7098
rect 38826 7046 38878 7098
rect 43570 7046 43622 7098
rect 43634 7046 43686 7098
rect 43698 7046 43750 7098
rect 43762 7046 43814 7098
rect 43826 7046 43878 7098
rect 7656 6944 7708 6996
rect 10048 6944 10100 6996
rect 10600 6944 10652 6996
rect 11888 6944 11940 6996
rect 15108 6987 15160 6996
rect 15108 6953 15138 6987
rect 15138 6953 15160 6987
rect 15108 6944 15160 6953
rect 16580 6987 16632 6996
rect 16580 6953 16589 6987
rect 16589 6953 16623 6987
rect 16623 6953 16632 6987
rect 16580 6944 16632 6953
rect 17040 6987 17092 6996
rect 17040 6953 17049 6987
rect 17049 6953 17083 6987
rect 17083 6953 17092 6987
rect 17040 6944 17092 6953
rect 17316 6944 17368 6996
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 18420 6944 18472 6996
rect 20628 6987 20680 6996
rect 20628 6953 20637 6987
rect 20637 6953 20671 6987
rect 20671 6953 20680 6987
rect 20628 6944 20680 6953
rect 20904 6944 20956 6996
rect 8944 6876 8996 6928
rect 9588 6876 9640 6928
rect 9404 6808 9456 6860
rect 8484 6740 8536 6792
rect 15752 6808 15804 6860
rect 17868 6876 17920 6928
rect 20536 6876 20588 6928
rect 16764 6808 16816 6860
rect 17684 6851 17736 6860
rect 17684 6817 17693 6851
rect 17693 6817 17727 6851
rect 17727 6817 17736 6851
rect 17684 6808 17736 6817
rect 10416 6672 10468 6724
rect 7656 6604 7708 6656
rect 10232 6604 10284 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 12532 6672 12584 6724
rect 14648 6715 14700 6724
rect 14648 6681 14657 6715
rect 14657 6681 14691 6715
rect 14691 6681 14700 6715
rect 16488 6740 16540 6792
rect 14648 6672 14700 6681
rect 15384 6672 15436 6724
rect 15660 6672 15712 6724
rect 16764 6672 16816 6724
rect 10600 6604 10652 6613
rect 12624 6604 12676 6656
rect 13084 6604 13136 6656
rect 15844 6604 15896 6656
rect 17592 6740 17644 6792
rect 18328 6740 18380 6792
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19524 6808 19576 6860
rect 20444 6808 20496 6860
rect 20720 6808 20772 6860
rect 22376 6876 22428 6928
rect 22836 6987 22888 6996
rect 22836 6953 22845 6987
rect 22845 6953 22879 6987
rect 22879 6953 22888 6987
rect 22836 6944 22888 6953
rect 24216 6944 24268 6996
rect 24308 6944 24360 6996
rect 26424 6944 26476 6996
rect 27712 6944 27764 6996
rect 27988 6987 28040 6996
rect 27988 6953 27997 6987
rect 27997 6953 28031 6987
rect 28031 6953 28040 6987
rect 27988 6944 28040 6953
rect 28724 6944 28776 6996
rect 23204 6876 23256 6928
rect 22008 6808 22060 6860
rect 18420 6672 18472 6724
rect 22376 6740 22428 6792
rect 22652 6740 22704 6792
rect 23296 6851 23348 6860
rect 23296 6817 23305 6851
rect 23305 6817 23339 6851
rect 23339 6817 23348 6851
rect 23296 6808 23348 6817
rect 20996 6672 21048 6724
rect 21548 6672 21600 6724
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 17408 6604 17460 6656
rect 18512 6604 18564 6656
rect 19156 6604 19208 6656
rect 19248 6604 19300 6656
rect 19432 6604 19484 6656
rect 19892 6604 19944 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 20352 6604 20404 6656
rect 22192 6604 22244 6656
rect 25320 6876 25372 6928
rect 25596 6808 25648 6860
rect 26608 6876 26660 6928
rect 25964 6783 26016 6792
rect 25964 6749 25973 6783
rect 25973 6749 26007 6783
rect 26007 6749 26016 6783
rect 25964 6740 26016 6749
rect 27436 6783 27488 6792
rect 27436 6749 27445 6783
rect 27445 6749 27479 6783
rect 27479 6749 27488 6783
rect 27436 6740 27488 6749
rect 30288 6876 30340 6928
rect 31484 6876 31536 6928
rect 27804 6672 27856 6724
rect 24216 6604 24268 6656
rect 25044 6604 25096 6656
rect 25596 6604 25648 6656
rect 26148 6647 26200 6656
rect 26148 6613 26157 6647
rect 26157 6613 26191 6647
rect 26191 6613 26200 6647
rect 26148 6604 26200 6613
rect 27436 6604 27488 6656
rect 28540 6783 28592 6792
rect 28540 6749 28549 6783
rect 28549 6749 28583 6783
rect 28583 6749 28592 6783
rect 28540 6740 28592 6749
rect 28724 6740 28776 6792
rect 30288 6740 30340 6792
rect 30472 6740 30524 6792
rect 30748 6740 30800 6792
rect 30840 6740 30892 6792
rect 29460 6672 29512 6724
rect 31024 6672 31076 6724
rect 31392 6672 31444 6724
rect 33968 6944 34020 6996
rect 34428 6987 34480 6996
rect 34428 6953 34437 6987
rect 34437 6953 34471 6987
rect 34471 6953 34480 6987
rect 34428 6944 34480 6953
rect 34888 6944 34940 6996
rect 32864 6808 32916 6860
rect 33692 6808 33744 6860
rect 34980 6876 35032 6928
rect 31944 6740 31996 6792
rect 29552 6604 29604 6656
rect 30748 6647 30800 6656
rect 30748 6613 30757 6647
rect 30757 6613 30791 6647
rect 30791 6613 30800 6647
rect 30748 6604 30800 6613
rect 31576 6604 31628 6656
rect 32496 6604 32548 6656
rect 33416 6672 33468 6724
rect 35992 6740 36044 6792
rect 36912 6851 36964 6860
rect 36912 6817 36921 6851
rect 36921 6817 36955 6851
rect 36955 6817 36964 6851
rect 36912 6808 36964 6817
rect 37740 6876 37792 6928
rect 37924 6851 37976 6860
rect 37924 6817 37933 6851
rect 37933 6817 37967 6851
rect 37967 6817 37976 6851
rect 37924 6808 37976 6817
rect 39212 6851 39264 6860
rect 39212 6817 39221 6851
rect 39221 6817 39255 6851
rect 39255 6817 39264 6851
rect 39212 6808 39264 6817
rect 39856 6944 39908 6996
rect 40500 6944 40552 6996
rect 41328 6987 41380 6996
rect 41328 6953 41358 6987
rect 41358 6953 41380 6987
rect 41328 6944 41380 6953
rect 43444 6944 43496 6996
rect 44916 6987 44968 6996
rect 44916 6953 44925 6987
rect 44925 6953 44959 6987
rect 44959 6953 44968 6987
rect 44916 6944 44968 6953
rect 40684 6808 40736 6860
rect 41880 6808 41932 6860
rect 36728 6783 36780 6792
rect 36728 6749 36737 6783
rect 36737 6749 36771 6783
rect 36771 6749 36780 6783
rect 36728 6740 36780 6749
rect 34060 6715 34112 6724
rect 34060 6681 34069 6715
rect 34069 6681 34103 6715
rect 34103 6681 34112 6715
rect 34060 6672 34112 6681
rect 34612 6672 34664 6724
rect 35256 6672 35308 6724
rect 33784 6604 33836 6656
rect 33968 6604 34020 6656
rect 34704 6647 34756 6656
rect 34704 6613 34713 6647
rect 34713 6613 34747 6647
rect 34747 6613 34756 6647
rect 34704 6604 34756 6613
rect 34888 6604 34940 6656
rect 35532 6647 35584 6656
rect 35532 6613 35541 6647
rect 35541 6613 35575 6647
rect 35575 6613 35584 6647
rect 35532 6604 35584 6613
rect 36176 6672 36228 6724
rect 38016 6672 38068 6724
rect 36452 6604 36504 6656
rect 36820 6647 36872 6656
rect 36820 6613 36829 6647
rect 36829 6613 36863 6647
rect 36863 6613 36872 6647
rect 36820 6604 36872 6613
rect 37280 6647 37332 6656
rect 37280 6613 37289 6647
rect 37289 6613 37323 6647
rect 37323 6613 37332 6647
rect 37280 6604 37332 6613
rect 39120 6740 39172 6792
rect 40868 6740 40920 6792
rect 38844 6604 38896 6656
rect 40316 6604 40368 6656
rect 42524 6808 42576 6860
rect 42800 6851 42852 6860
rect 42800 6817 42809 6851
rect 42809 6817 42843 6851
rect 42843 6817 42852 6851
rect 42800 6808 42852 6817
rect 44180 6808 44232 6860
rect 42892 6740 42944 6792
rect 43260 6647 43312 6656
rect 43260 6613 43269 6647
rect 43269 6613 43303 6647
rect 43303 6613 43312 6647
rect 43260 6604 43312 6613
rect 6070 6502 6122 6554
rect 6134 6502 6186 6554
rect 6198 6502 6250 6554
rect 6262 6502 6314 6554
rect 6326 6502 6378 6554
rect 11070 6502 11122 6554
rect 11134 6502 11186 6554
rect 11198 6502 11250 6554
rect 11262 6502 11314 6554
rect 11326 6502 11378 6554
rect 16070 6502 16122 6554
rect 16134 6502 16186 6554
rect 16198 6502 16250 6554
rect 16262 6502 16314 6554
rect 16326 6502 16378 6554
rect 21070 6502 21122 6554
rect 21134 6502 21186 6554
rect 21198 6502 21250 6554
rect 21262 6502 21314 6554
rect 21326 6502 21378 6554
rect 26070 6502 26122 6554
rect 26134 6502 26186 6554
rect 26198 6502 26250 6554
rect 26262 6502 26314 6554
rect 26326 6502 26378 6554
rect 31070 6502 31122 6554
rect 31134 6502 31186 6554
rect 31198 6502 31250 6554
rect 31262 6502 31314 6554
rect 31326 6502 31378 6554
rect 36070 6502 36122 6554
rect 36134 6502 36186 6554
rect 36198 6502 36250 6554
rect 36262 6502 36314 6554
rect 36326 6502 36378 6554
rect 41070 6502 41122 6554
rect 41134 6502 41186 6554
rect 41198 6502 41250 6554
rect 41262 6502 41314 6554
rect 41326 6502 41378 6554
rect 1308 6264 1360 6316
rect 15016 6400 15068 6452
rect 15936 6400 15988 6452
rect 16580 6400 16632 6452
rect 16948 6400 17000 6452
rect 7656 6375 7708 6384
rect 7656 6341 7665 6375
rect 7665 6341 7699 6375
rect 7699 6341 7708 6375
rect 7656 6332 7708 6341
rect 9404 6332 9456 6384
rect 10508 6332 10560 6384
rect 8484 6264 8536 6316
rect 9128 6264 9180 6316
rect 4988 6196 5040 6248
rect 7656 6128 7708 6180
rect 15660 6264 15712 6316
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 16580 6264 16632 6316
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17684 6264 17736 6316
rect 17960 6400 18012 6452
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 19156 6400 19208 6452
rect 20996 6400 21048 6452
rect 21548 6443 21600 6452
rect 21548 6409 21557 6443
rect 21557 6409 21591 6443
rect 21591 6409 21600 6443
rect 21548 6400 21600 6409
rect 17868 6332 17920 6384
rect 19892 6332 19944 6384
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 10600 6060 10652 6112
rect 13176 6128 13228 6180
rect 13636 6171 13688 6180
rect 13636 6137 13645 6171
rect 13645 6137 13679 6171
rect 13679 6137 13688 6171
rect 13636 6128 13688 6137
rect 15568 6196 15620 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16304 6196 16356 6248
rect 18052 6196 18104 6248
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 20904 6264 20956 6316
rect 18972 6196 19024 6248
rect 19340 6196 19392 6248
rect 21456 6264 21508 6316
rect 21916 6400 21968 6452
rect 23388 6400 23440 6452
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 25504 6400 25556 6452
rect 25780 6400 25832 6452
rect 25964 6400 26016 6452
rect 27804 6400 27856 6452
rect 28356 6400 28408 6452
rect 22008 6332 22060 6384
rect 22560 6332 22612 6384
rect 22744 6332 22796 6384
rect 25320 6375 25372 6384
rect 25320 6341 25329 6375
rect 25329 6341 25363 6375
rect 25363 6341 25372 6375
rect 25320 6332 25372 6341
rect 25412 6332 25464 6384
rect 24124 6264 24176 6316
rect 24676 6264 24728 6316
rect 24768 6264 24820 6316
rect 23112 6196 23164 6248
rect 25872 6196 25924 6248
rect 16764 6128 16816 6180
rect 20352 6171 20404 6180
rect 20352 6137 20361 6171
rect 20361 6137 20395 6171
rect 20395 6137 20404 6171
rect 20352 6128 20404 6137
rect 21640 6128 21692 6180
rect 21916 6128 21968 6180
rect 11796 6060 11848 6112
rect 12624 6060 12676 6112
rect 14096 6060 14148 6112
rect 16212 6103 16264 6112
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 16672 6060 16724 6112
rect 17500 6060 17552 6112
rect 19248 6060 19300 6112
rect 21088 6060 21140 6112
rect 21180 6060 21232 6112
rect 22192 6103 22244 6112
rect 22192 6069 22201 6103
rect 22201 6069 22235 6103
rect 22235 6069 22244 6103
rect 22192 6060 22244 6069
rect 22836 6060 22888 6112
rect 24032 6128 24084 6180
rect 27620 6332 27672 6384
rect 28908 6400 28960 6452
rect 30748 6400 30800 6452
rect 30840 6400 30892 6452
rect 26700 6264 26752 6316
rect 27896 6264 27948 6316
rect 26424 6196 26476 6248
rect 27068 6239 27120 6248
rect 27068 6205 27077 6239
rect 27077 6205 27111 6239
rect 27111 6205 27120 6239
rect 27068 6196 27120 6205
rect 23756 6060 23808 6112
rect 24400 6060 24452 6112
rect 25228 6060 25280 6112
rect 25872 6103 25924 6112
rect 25872 6069 25881 6103
rect 25881 6069 25915 6103
rect 25915 6069 25924 6103
rect 25872 6060 25924 6069
rect 26516 6128 26568 6180
rect 26608 6128 26660 6180
rect 27712 6196 27764 6248
rect 30104 6332 30156 6384
rect 30288 6332 30340 6384
rect 34704 6400 34756 6452
rect 35256 6400 35308 6452
rect 36452 6400 36504 6452
rect 36912 6400 36964 6452
rect 29276 6264 29328 6316
rect 29460 6196 29512 6248
rect 32956 6332 33008 6384
rect 34152 6332 34204 6384
rect 31576 6264 31628 6316
rect 35992 6264 36044 6316
rect 37280 6332 37332 6384
rect 38844 6443 38896 6452
rect 38844 6409 38853 6443
rect 38853 6409 38887 6443
rect 38887 6409 38896 6443
rect 38844 6400 38896 6409
rect 39120 6400 39172 6452
rect 41512 6400 41564 6452
rect 42800 6400 42852 6452
rect 43076 6443 43128 6452
rect 43076 6409 43085 6443
rect 43085 6409 43119 6443
rect 43119 6409 43128 6443
rect 43076 6400 43128 6409
rect 43352 6400 43404 6452
rect 44732 6443 44784 6452
rect 44732 6409 44741 6443
rect 44741 6409 44775 6443
rect 44775 6409 44784 6443
rect 44732 6400 44784 6409
rect 37004 6307 37056 6316
rect 37004 6273 37013 6307
rect 37013 6273 37047 6307
rect 37047 6273 37056 6307
rect 37004 6264 37056 6273
rect 38476 6264 38528 6316
rect 38660 6264 38712 6316
rect 39212 6332 39264 6384
rect 40500 6332 40552 6384
rect 33232 6196 33284 6248
rect 34244 6196 34296 6248
rect 34612 6239 34664 6248
rect 34612 6205 34621 6239
rect 34621 6205 34655 6239
rect 34655 6205 34664 6239
rect 34612 6196 34664 6205
rect 35256 6196 35308 6248
rect 37096 6239 37148 6248
rect 37096 6205 37105 6239
rect 37105 6205 37139 6239
rect 37139 6205 37148 6239
rect 37096 6196 37148 6205
rect 40316 6264 40368 6316
rect 40592 6264 40644 6316
rect 27436 6060 27488 6112
rect 28356 6060 28408 6112
rect 33416 6103 33468 6112
rect 33416 6069 33425 6103
rect 33425 6069 33459 6103
rect 33459 6069 33468 6103
rect 33416 6060 33468 6069
rect 33692 6103 33744 6112
rect 33692 6069 33701 6103
rect 33701 6069 33735 6103
rect 33735 6069 33744 6103
rect 33692 6060 33744 6069
rect 34152 6060 34204 6112
rect 35808 6128 35860 6180
rect 35992 6128 36044 6180
rect 36176 6103 36228 6112
rect 36176 6069 36185 6103
rect 36185 6069 36219 6103
rect 36219 6069 36228 6103
rect 36176 6060 36228 6069
rect 38660 6128 38712 6180
rect 40684 6196 40736 6248
rect 40776 6171 40828 6180
rect 40776 6137 40785 6171
rect 40785 6137 40819 6171
rect 40819 6137 40828 6171
rect 40776 6128 40828 6137
rect 39304 6060 39356 6112
rect 39580 6060 39632 6112
rect 42064 6196 42116 6248
rect 44364 6264 44416 6316
rect 42708 6196 42760 6248
rect 44180 6196 44232 6248
rect 42984 6060 43036 6112
rect 43996 6103 44048 6112
rect 43996 6069 44005 6103
rect 44005 6069 44039 6103
rect 44039 6069 44048 6103
rect 43996 6060 44048 6069
rect 3570 5958 3622 6010
rect 3634 5958 3686 6010
rect 3698 5958 3750 6010
rect 3762 5958 3814 6010
rect 3826 5958 3878 6010
rect 8570 5958 8622 6010
rect 8634 5958 8686 6010
rect 8698 5958 8750 6010
rect 8762 5958 8814 6010
rect 8826 5958 8878 6010
rect 13570 5958 13622 6010
rect 13634 5958 13686 6010
rect 13698 5958 13750 6010
rect 13762 5958 13814 6010
rect 13826 5958 13878 6010
rect 18570 5958 18622 6010
rect 18634 5958 18686 6010
rect 18698 5958 18750 6010
rect 18762 5958 18814 6010
rect 18826 5958 18878 6010
rect 23570 5958 23622 6010
rect 23634 5958 23686 6010
rect 23698 5958 23750 6010
rect 23762 5958 23814 6010
rect 23826 5958 23878 6010
rect 28570 5958 28622 6010
rect 28634 5958 28686 6010
rect 28698 5958 28750 6010
rect 28762 5958 28814 6010
rect 28826 5958 28878 6010
rect 33570 5958 33622 6010
rect 33634 5958 33686 6010
rect 33698 5958 33750 6010
rect 33762 5958 33814 6010
rect 33826 5958 33878 6010
rect 38570 5958 38622 6010
rect 38634 5958 38686 6010
rect 38698 5958 38750 6010
rect 38762 5958 38814 6010
rect 38826 5958 38878 6010
rect 43570 5958 43622 6010
rect 43634 5958 43686 6010
rect 43698 5958 43750 6010
rect 43762 5958 43814 6010
rect 43826 5958 43878 6010
rect 2504 5856 2556 5908
rect 3056 5856 3108 5908
rect 4252 5856 4304 5908
rect 5448 5856 5500 5908
rect 7196 5856 7248 5908
rect 7656 5856 7708 5908
rect 8300 5856 8352 5908
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 10508 5856 10560 5908
rect 13176 5899 13228 5908
rect 13176 5865 13185 5899
rect 13185 5865 13219 5899
rect 13219 5865 13228 5899
rect 13176 5856 13228 5865
rect 14372 5856 14424 5908
rect 5724 5788 5776 5840
rect 12808 5788 12860 5840
rect 13360 5788 13412 5840
rect 14464 5788 14516 5840
rect 15200 5856 15252 5908
rect 16028 5899 16080 5908
rect 16028 5865 16037 5899
rect 16037 5865 16071 5899
rect 16071 5865 16080 5899
rect 16028 5856 16080 5865
rect 16948 5856 17000 5908
rect 17132 5856 17184 5908
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 17776 5856 17828 5908
rect 19800 5856 19852 5908
rect 20260 5856 20312 5908
rect 20444 5856 20496 5908
rect 21456 5856 21508 5908
rect 7288 5720 7340 5772
rect 4988 5652 5040 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 2596 5516 2648 5568
rect 2872 5516 2924 5568
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 7748 5516 7800 5568
rect 9128 5516 9180 5568
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 10416 5516 10468 5568
rect 11520 5516 11572 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 14188 5516 14240 5568
rect 15568 5720 15620 5772
rect 14464 5627 14516 5636
rect 14464 5593 14473 5627
rect 14473 5593 14507 5627
rect 14507 5593 14516 5627
rect 14464 5584 14516 5593
rect 14648 5584 14700 5636
rect 15108 5584 15160 5636
rect 15200 5627 15252 5636
rect 15200 5593 15227 5627
rect 15227 5593 15252 5627
rect 15200 5584 15252 5593
rect 14924 5516 14976 5568
rect 15844 5627 15896 5636
rect 15844 5593 15853 5627
rect 15853 5593 15887 5627
rect 15887 5593 15896 5627
rect 15844 5584 15896 5593
rect 16764 5720 16816 5772
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 17960 5831 18012 5840
rect 17960 5797 17969 5831
rect 17969 5797 18003 5831
rect 18003 5797 18012 5831
rect 17960 5788 18012 5797
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 18420 5720 18472 5772
rect 17500 5652 17552 5661
rect 18052 5652 18104 5704
rect 19248 5720 19300 5772
rect 19524 5763 19576 5772
rect 19524 5729 19533 5763
rect 19533 5729 19567 5763
rect 19567 5729 19576 5763
rect 19524 5720 19576 5729
rect 20168 5720 20220 5772
rect 20260 5720 20312 5772
rect 20996 5720 21048 5772
rect 21640 5720 21692 5772
rect 23020 5720 23072 5772
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 24584 5856 24636 5908
rect 25136 5899 25188 5908
rect 25136 5865 25145 5899
rect 25145 5865 25179 5899
rect 25179 5865 25188 5899
rect 25136 5856 25188 5865
rect 17868 5584 17920 5636
rect 16396 5516 16448 5568
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 16580 5516 16632 5568
rect 16856 5516 16908 5568
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 18328 5584 18380 5636
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18512 5584 18564 5636
rect 18696 5584 18748 5636
rect 18972 5695 19024 5704
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 19156 5695 19208 5704
rect 19156 5661 19165 5695
rect 19165 5661 19199 5695
rect 19199 5661 19208 5695
rect 19156 5652 19208 5661
rect 19340 5652 19392 5704
rect 21088 5652 21140 5704
rect 21824 5652 21876 5704
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 22836 5652 22888 5704
rect 21548 5584 21600 5636
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 19524 5516 19576 5568
rect 19708 5516 19760 5568
rect 19800 5516 19852 5568
rect 22376 5516 22428 5568
rect 24308 5695 24360 5704
rect 24308 5661 24317 5695
rect 24317 5661 24351 5695
rect 24351 5661 24360 5695
rect 24308 5652 24360 5661
rect 24400 5652 24452 5704
rect 25228 5720 25280 5772
rect 26056 5720 26108 5772
rect 27068 5856 27120 5908
rect 28080 5899 28132 5908
rect 28080 5865 28089 5899
rect 28089 5865 28123 5899
rect 28123 5865 28132 5899
rect 28080 5856 28132 5865
rect 28908 5856 28960 5908
rect 27988 5788 28040 5840
rect 25044 5652 25096 5704
rect 26792 5652 26844 5704
rect 27068 5652 27120 5704
rect 27436 5652 27488 5704
rect 25596 5584 25648 5636
rect 22928 5516 22980 5568
rect 24400 5516 24452 5568
rect 24860 5516 24912 5568
rect 25412 5516 25464 5568
rect 27252 5584 27304 5636
rect 27988 5584 28040 5636
rect 28908 5763 28960 5772
rect 28908 5729 28917 5763
rect 28917 5729 28951 5763
rect 28951 5729 28960 5763
rect 28908 5720 28960 5729
rect 29276 5720 29328 5772
rect 30564 5856 30616 5908
rect 30380 5788 30432 5840
rect 31024 5856 31076 5908
rect 31760 5856 31812 5908
rect 33232 5899 33284 5908
rect 33232 5865 33241 5899
rect 33241 5865 33275 5899
rect 33275 5865 33284 5899
rect 33232 5856 33284 5865
rect 34612 5856 34664 5908
rect 32404 5720 32456 5772
rect 32680 5720 32732 5772
rect 33140 5720 33192 5772
rect 33968 5720 34020 5772
rect 34060 5763 34112 5772
rect 34060 5729 34069 5763
rect 34069 5729 34103 5763
rect 34103 5729 34112 5763
rect 34060 5720 34112 5729
rect 30288 5652 30340 5704
rect 29092 5584 29144 5636
rect 29184 5627 29236 5636
rect 29184 5593 29193 5627
rect 29193 5593 29227 5627
rect 29227 5593 29236 5627
rect 29184 5584 29236 5593
rect 28264 5559 28316 5568
rect 28264 5525 28273 5559
rect 28273 5525 28307 5559
rect 28307 5525 28316 5559
rect 28264 5516 28316 5525
rect 28448 5516 28500 5568
rect 32680 5584 32732 5636
rect 33324 5652 33376 5704
rect 34520 5763 34572 5772
rect 34520 5729 34529 5763
rect 34529 5729 34563 5763
rect 34563 5729 34572 5763
rect 34520 5720 34572 5729
rect 34336 5695 34388 5704
rect 34336 5661 34345 5695
rect 34345 5661 34379 5695
rect 34379 5661 34388 5695
rect 34336 5652 34388 5661
rect 34704 5652 34756 5704
rect 35532 5856 35584 5908
rect 36820 5856 36872 5908
rect 37096 5856 37148 5908
rect 37280 5856 37332 5908
rect 38108 5899 38160 5908
rect 38108 5865 38117 5899
rect 38117 5865 38151 5899
rect 38151 5865 38160 5899
rect 38108 5856 38160 5865
rect 38476 5856 38528 5908
rect 39028 5856 39080 5908
rect 43076 5856 43128 5908
rect 43352 5856 43404 5908
rect 44916 5899 44968 5908
rect 44916 5865 44925 5899
rect 44925 5865 44959 5899
rect 44959 5865 44968 5899
rect 44916 5856 44968 5865
rect 40960 5788 41012 5840
rect 36176 5720 36228 5772
rect 36820 5720 36872 5772
rect 35256 5695 35308 5704
rect 35256 5661 35265 5695
rect 35265 5661 35299 5695
rect 35299 5661 35308 5695
rect 35256 5652 35308 5661
rect 36636 5652 36688 5704
rect 36912 5652 36964 5704
rect 37188 5652 37240 5704
rect 37924 5720 37976 5772
rect 38200 5652 38252 5704
rect 39856 5720 39908 5772
rect 36820 5584 36872 5636
rect 32588 5559 32640 5568
rect 32588 5525 32597 5559
rect 32597 5525 32631 5559
rect 32631 5525 32640 5559
rect 32588 5516 32640 5525
rect 32772 5516 32824 5568
rect 32864 5516 32916 5568
rect 36452 5516 36504 5568
rect 37096 5559 37148 5568
rect 37096 5525 37105 5559
rect 37105 5525 37139 5559
rect 37139 5525 37148 5559
rect 37096 5516 37148 5525
rect 37280 5516 37332 5568
rect 39120 5584 39172 5636
rect 38476 5559 38528 5568
rect 38476 5525 38485 5559
rect 38485 5525 38519 5559
rect 38519 5525 38528 5559
rect 38476 5516 38528 5525
rect 38936 5516 38988 5568
rect 39488 5627 39540 5636
rect 39488 5593 39497 5627
rect 39497 5593 39531 5627
rect 39531 5593 39540 5627
rect 39488 5584 39540 5593
rect 40224 5584 40276 5636
rect 40868 5652 40920 5704
rect 42524 5720 42576 5772
rect 40868 5516 40920 5568
rect 43076 5559 43128 5568
rect 43076 5525 43085 5559
rect 43085 5525 43119 5559
rect 43119 5525 43128 5559
rect 43076 5516 43128 5525
rect 6070 5414 6122 5466
rect 6134 5414 6186 5466
rect 6198 5414 6250 5466
rect 6262 5414 6314 5466
rect 6326 5414 6378 5466
rect 11070 5414 11122 5466
rect 11134 5414 11186 5466
rect 11198 5414 11250 5466
rect 11262 5414 11314 5466
rect 11326 5414 11378 5466
rect 16070 5414 16122 5466
rect 16134 5414 16186 5466
rect 16198 5414 16250 5466
rect 16262 5414 16314 5466
rect 16326 5414 16378 5466
rect 21070 5414 21122 5466
rect 21134 5414 21186 5466
rect 21198 5414 21250 5466
rect 21262 5414 21314 5466
rect 21326 5414 21378 5466
rect 26070 5414 26122 5466
rect 26134 5414 26186 5466
rect 26198 5414 26250 5466
rect 26262 5414 26314 5466
rect 26326 5414 26378 5466
rect 31070 5414 31122 5466
rect 31134 5414 31186 5466
rect 31198 5414 31250 5466
rect 31262 5414 31314 5466
rect 31326 5414 31378 5466
rect 36070 5414 36122 5466
rect 36134 5414 36186 5466
rect 36198 5414 36250 5466
rect 36262 5414 36314 5466
rect 36326 5414 36378 5466
rect 41070 5414 41122 5466
rect 41134 5414 41186 5466
rect 41198 5414 41250 5466
rect 41262 5414 41314 5466
rect 41326 5414 41378 5466
rect 3424 5355 3476 5364
rect 3424 5321 3433 5355
rect 3433 5321 3467 5355
rect 3467 5321 3476 5355
rect 3424 5312 3476 5321
rect 4620 5312 4672 5364
rect 5448 5312 5500 5364
rect 6460 5312 6512 5364
rect 7748 5312 7800 5364
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 11796 5312 11848 5364
rect 13176 5312 13228 5364
rect 8392 5244 8444 5296
rect 9128 5287 9180 5296
rect 9128 5253 9137 5287
rect 9137 5253 9171 5287
rect 9171 5253 9180 5287
rect 9128 5244 9180 5253
rect 11520 5287 11572 5296
rect 11520 5253 11529 5287
rect 11529 5253 11563 5287
rect 11563 5253 11572 5287
rect 11520 5244 11572 5253
rect 5356 5176 5408 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13268 5176 13320 5228
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 1584 4972 1636 5024
rect 2320 4972 2372 5024
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 6736 5108 6788 5160
rect 10692 5108 10744 5160
rect 12532 5108 12584 5160
rect 12624 5108 12676 5160
rect 13728 5176 13780 5228
rect 15108 5312 15160 5364
rect 14372 5287 14424 5296
rect 14372 5253 14381 5287
rect 14381 5253 14415 5287
rect 14415 5253 14424 5287
rect 14372 5244 14424 5253
rect 15752 5244 15804 5296
rect 16028 5287 16080 5296
rect 16028 5253 16037 5287
rect 16037 5253 16071 5287
rect 16071 5253 16080 5287
rect 16028 5244 16080 5253
rect 15660 5176 15712 5228
rect 16488 5312 16540 5364
rect 16580 5287 16632 5296
rect 16580 5253 16587 5287
rect 16587 5253 16621 5287
rect 16621 5253 16632 5287
rect 16580 5244 16632 5253
rect 16764 5244 16816 5296
rect 17040 5244 17092 5296
rect 17132 5287 17184 5296
rect 17132 5253 17141 5287
rect 17141 5253 17175 5287
rect 17175 5253 17184 5287
rect 17132 5244 17184 5253
rect 18144 5312 18196 5364
rect 19800 5312 19852 5364
rect 20076 5312 20128 5364
rect 14740 5108 14792 5160
rect 15568 5108 15620 5160
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 19340 5244 19392 5296
rect 21824 5244 21876 5296
rect 22560 5244 22612 5296
rect 18696 5176 18748 5185
rect 21916 5176 21968 5228
rect 22744 5176 22796 5228
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 23112 5176 23164 5228
rect 23296 5219 23348 5228
rect 23296 5185 23305 5219
rect 23305 5185 23339 5219
rect 23339 5185 23348 5219
rect 23296 5176 23348 5185
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 20812 5108 20864 5160
rect 7288 5040 7340 5092
rect 4068 4972 4120 5024
rect 4344 5015 4396 5024
rect 4344 4981 4353 5015
rect 4353 4981 4387 5015
rect 4387 4981 4396 5015
rect 4344 4972 4396 4981
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 8300 4972 8352 5024
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 11612 4972 11664 5024
rect 12072 5015 12124 5024
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 14004 5083 14056 5092
rect 14004 5049 14013 5083
rect 14013 5049 14047 5083
rect 14047 5049 14056 5083
rect 14004 5040 14056 5049
rect 16672 4972 16724 5024
rect 17224 4972 17276 5024
rect 19064 5015 19116 5024
rect 19064 4981 19073 5015
rect 19073 4981 19107 5015
rect 19107 4981 19116 5015
rect 19064 4972 19116 4981
rect 19432 4972 19484 5024
rect 21548 5040 21600 5092
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 20904 4972 20956 4981
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 25780 5312 25832 5364
rect 26148 5312 26200 5364
rect 26792 5312 26844 5364
rect 27620 5312 27672 5364
rect 25044 5108 25096 5160
rect 25688 5176 25740 5228
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 25964 5176 26016 5228
rect 26332 5219 26384 5228
rect 26332 5185 26341 5219
rect 26341 5185 26375 5219
rect 26375 5185 26384 5219
rect 26332 5176 26384 5185
rect 27896 5244 27948 5296
rect 29092 5355 29144 5364
rect 29092 5321 29101 5355
rect 29101 5321 29135 5355
rect 29135 5321 29144 5355
rect 29092 5312 29144 5321
rect 29552 5355 29604 5364
rect 29552 5321 29561 5355
rect 29561 5321 29595 5355
rect 29595 5321 29604 5355
rect 29552 5312 29604 5321
rect 30380 5355 30432 5364
rect 30380 5321 30389 5355
rect 30389 5321 30423 5355
rect 30423 5321 30432 5355
rect 30380 5312 30432 5321
rect 30748 5312 30800 5364
rect 31576 5312 31628 5364
rect 28356 5219 28408 5228
rect 28356 5185 28365 5219
rect 28365 5185 28399 5219
rect 28399 5185 28408 5219
rect 28356 5176 28408 5185
rect 22008 4972 22060 5024
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 24308 5015 24360 5024
rect 24308 4981 24317 5015
rect 24317 4981 24351 5015
rect 24351 4981 24360 5015
rect 24308 4972 24360 4981
rect 24492 4972 24544 5024
rect 25228 5015 25280 5024
rect 25228 4981 25237 5015
rect 25237 4981 25271 5015
rect 25271 4981 25280 5015
rect 25228 4972 25280 4981
rect 25780 4972 25832 5024
rect 26056 5015 26108 5024
rect 26056 4981 26065 5015
rect 26065 4981 26099 5015
rect 26099 4981 26108 5015
rect 26056 4972 26108 4981
rect 26148 4972 26200 5024
rect 30288 5219 30340 5228
rect 30288 5185 30297 5219
rect 30297 5185 30331 5219
rect 30331 5185 30340 5219
rect 30288 5176 30340 5185
rect 32588 5312 32640 5364
rect 32680 5312 32732 5364
rect 34336 5312 34388 5364
rect 36360 5312 36412 5364
rect 36820 5312 36872 5364
rect 40040 5355 40092 5364
rect 40040 5321 40049 5355
rect 40049 5321 40083 5355
rect 40083 5321 40092 5355
rect 40040 5312 40092 5321
rect 40592 5312 40644 5364
rect 40960 5312 41012 5364
rect 41788 5312 41840 5364
rect 43076 5355 43128 5364
rect 43076 5321 43085 5355
rect 43085 5321 43119 5355
rect 43119 5321 43128 5355
rect 43076 5312 43128 5321
rect 43996 5312 44048 5364
rect 44548 5355 44600 5364
rect 44548 5321 44557 5355
rect 44557 5321 44591 5355
rect 44591 5321 44600 5355
rect 44548 5312 44600 5321
rect 40132 5244 40184 5296
rect 42892 5244 42944 5296
rect 43352 5244 43404 5296
rect 32864 5176 32916 5228
rect 34520 5176 34572 5228
rect 36084 5176 36136 5228
rect 36636 5176 36688 5228
rect 37096 5176 37148 5228
rect 37280 5176 37332 5228
rect 39028 5176 39080 5228
rect 39396 5176 39448 5228
rect 39948 5219 40000 5228
rect 39948 5185 39957 5219
rect 39957 5185 39991 5219
rect 39991 5185 40000 5219
rect 39948 5176 40000 5185
rect 42064 5176 42116 5228
rect 29552 5108 29604 5160
rect 30196 5108 30248 5160
rect 30564 5108 30616 5160
rect 31392 5108 31444 5160
rect 34152 5108 34204 5160
rect 34244 5108 34296 5160
rect 34704 5151 34756 5160
rect 34704 5117 34713 5151
rect 34713 5117 34747 5151
rect 34747 5117 34756 5151
rect 34704 5108 34756 5117
rect 36728 5108 36780 5160
rect 38016 5151 38068 5160
rect 38016 5117 38025 5151
rect 38025 5117 38059 5151
rect 38059 5117 38068 5151
rect 38016 5108 38068 5117
rect 39304 5108 39356 5160
rect 39580 5108 39632 5160
rect 40868 5151 40920 5160
rect 40868 5117 40877 5151
rect 40877 5117 40911 5151
rect 40911 5117 40920 5151
rect 40868 5108 40920 5117
rect 40960 5151 41012 5160
rect 40960 5117 40969 5151
rect 40969 5117 41003 5151
rect 41003 5117 41012 5151
rect 40960 5108 41012 5117
rect 28264 5015 28316 5024
rect 28264 4981 28273 5015
rect 28273 4981 28307 5015
rect 28307 4981 28316 5015
rect 28264 4972 28316 4981
rect 29184 4972 29236 5024
rect 31392 4972 31444 5024
rect 32864 4972 32916 5024
rect 33324 5015 33376 5024
rect 33324 4981 33333 5015
rect 33333 4981 33367 5015
rect 33367 4981 33376 5015
rect 33324 4972 33376 4981
rect 34152 4972 34204 5024
rect 34428 5015 34480 5024
rect 34428 4981 34437 5015
rect 34437 4981 34471 5015
rect 34471 4981 34480 5015
rect 34428 4972 34480 4981
rect 35348 4972 35400 5024
rect 36452 4972 36504 5024
rect 39212 4972 39264 5024
rect 41972 5015 42024 5024
rect 41972 4981 41981 5015
rect 41981 4981 42015 5015
rect 42015 4981 42024 5015
rect 41972 4972 42024 4981
rect 44088 4972 44140 5024
rect 44180 5015 44232 5024
rect 44180 4981 44189 5015
rect 44189 4981 44223 5015
rect 44223 4981 44232 5015
rect 44180 4972 44232 4981
rect 3570 4870 3622 4922
rect 3634 4870 3686 4922
rect 3698 4870 3750 4922
rect 3762 4870 3814 4922
rect 3826 4870 3878 4922
rect 8570 4870 8622 4922
rect 8634 4870 8686 4922
rect 8698 4870 8750 4922
rect 8762 4870 8814 4922
rect 8826 4870 8878 4922
rect 13570 4870 13622 4922
rect 13634 4870 13686 4922
rect 13698 4870 13750 4922
rect 13762 4870 13814 4922
rect 13826 4870 13878 4922
rect 18570 4870 18622 4922
rect 18634 4870 18686 4922
rect 18698 4870 18750 4922
rect 18762 4870 18814 4922
rect 18826 4870 18878 4922
rect 23570 4870 23622 4922
rect 23634 4870 23686 4922
rect 23698 4870 23750 4922
rect 23762 4870 23814 4922
rect 23826 4870 23878 4922
rect 28570 4870 28622 4922
rect 28634 4870 28686 4922
rect 28698 4870 28750 4922
rect 28762 4870 28814 4922
rect 28826 4870 28878 4922
rect 33570 4870 33622 4922
rect 33634 4870 33686 4922
rect 33698 4870 33750 4922
rect 33762 4870 33814 4922
rect 33826 4870 33878 4922
rect 38570 4870 38622 4922
rect 38634 4870 38686 4922
rect 38698 4870 38750 4922
rect 38762 4870 38814 4922
rect 38826 4870 38878 4922
rect 43570 4870 43622 4922
rect 43634 4870 43686 4922
rect 43698 4870 43750 4922
rect 43762 4870 43814 4922
rect 43826 4870 43878 4922
rect 11796 4768 11848 4820
rect 12256 4768 12308 4820
rect 14096 4768 14148 4820
rect 1584 4632 1636 4684
rect 4068 4632 4120 4684
rect 5264 4632 5316 4684
rect 8300 4632 8352 4684
rect 8484 4632 8536 4684
rect 9312 4632 9364 4684
rect 2596 4564 2648 4616
rect 3516 4607 3568 4616
rect 3516 4573 3525 4607
rect 3525 4573 3559 4607
rect 3559 4573 3568 4607
rect 3516 4564 3568 4573
rect 3976 4564 4028 4616
rect 4620 4564 4672 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 1492 4496 1544 4548
rect 2780 4496 2832 4548
rect 4712 4496 4764 4548
rect 5540 4496 5592 4548
rect 940 4471 992 4480
rect 940 4437 949 4471
rect 949 4437 983 4471
rect 983 4437 992 4471
rect 940 4428 992 4437
rect 2320 4428 2372 4480
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 6920 4428 6972 4480
rect 7932 4428 7984 4480
rect 8392 4564 8444 4616
rect 13912 4700 13964 4752
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 14004 4632 14056 4684
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16396 4768 16448 4820
rect 17132 4768 17184 4820
rect 19432 4811 19484 4820
rect 19432 4777 19441 4811
rect 19441 4777 19475 4811
rect 19475 4777 19484 4811
rect 19432 4768 19484 4777
rect 19708 4811 19760 4820
rect 19708 4777 19717 4811
rect 19717 4777 19751 4811
rect 19751 4777 19760 4811
rect 19708 4768 19760 4777
rect 20996 4768 21048 4820
rect 21824 4768 21876 4820
rect 13176 4564 13228 4616
rect 15752 4564 15804 4616
rect 15936 4743 15988 4752
rect 15936 4709 15945 4743
rect 15945 4709 15979 4743
rect 15979 4709 15988 4743
rect 15936 4700 15988 4709
rect 17960 4700 18012 4752
rect 18052 4700 18104 4752
rect 19524 4700 19576 4752
rect 11612 4496 11664 4548
rect 8392 4428 8444 4480
rect 9588 4471 9640 4480
rect 9588 4437 9597 4471
rect 9597 4437 9631 4471
rect 9631 4437 9640 4471
rect 9588 4428 9640 4437
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 10692 4428 10744 4480
rect 11520 4428 11572 4480
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 12808 4428 12860 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 14372 4539 14424 4548
rect 14372 4505 14381 4539
rect 14381 4505 14415 4539
rect 14415 4505 14424 4539
rect 14372 4496 14424 4505
rect 15660 4496 15712 4548
rect 15844 4496 15896 4548
rect 16028 4496 16080 4548
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 19064 4564 19116 4616
rect 16580 4496 16632 4548
rect 16948 4496 17000 4548
rect 17132 4496 17184 4548
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 20444 4632 20496 4684
rect 20996 4632 21048 4684
rect 22560 4768 22612 4820
rect 22652 4768 22704 4820
rect 23848 4768 23900 4820
rect 24584 4768 24636 4820
rect 20904 4564 20956 4616
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 22100 4632 22152 4641
rect 19984 4496 20036 4548
rect 21640 4496 21692 4548
rect 23112 4564 23164 4616
rect 24676 4700 24728 4752
rect 25136 4700 25188 4752
rect 23296 4632 23348 4684
rect 23940 4632 23992 4684
rect 24952 4632 25004 4684
rect 27436 4700 27488 4752
rect 30012 4743 30064 4752
rect 30012 4709 30021 4743
rect 30021 4709 30055 4743
rect 30055 4709 30064 4743
rect 30012 4700 30064 4709
rect 30288 4768 30340 4820
rect 32956 4768 33008 4820
rect 34336 4768 34388 4820
rect 34520 4768 34572 4820
rect 38016 4768 38068 4820
rect 38384 4768 38436 4820
rect 39488 4768 39540 4820
rect 31852 4700 31904 4752
rect 34060 4700 34112 4752
rect 35348 4700 35400 4752
rect 35992 4700 36044 4752
rect 36452 4700 36504 4752
rect 26792 4632 26844 4684
rect 22376 4496 22428 4548
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 22468 4428 22520 4480
rect 24124 4471 24176 4480
rect 24124 4437 24133 4471
rect 24133 4437 24167 4471
rect 24167 4437 24176 4471
rect 24768 4496 24820 4548
rect 25596 4496 25648 4548
rect 27712 4607 27764 4616
rect 27712 4573 27721 4607
rect 27721 4573 27755 4607
rect 27755 4573 27764 4607
rect 27712 4564 27764 4573
rect 27988 4632 28040 4684
rect 28448 4632 28500 4684
rect 28724 4632 28776 4684
rect 28356 4564 28408 4616
rect 24124 4428 24176 4437
rect 25688 4471 25740 4480
rect 25688 4437 25697 4471
rect 25697 4437 25731 4471
rect 25731 4437 25740 4471
rect 25688 4428 25740 4437
rect 25964 4496 26016 4548
rect 26332 4496 26384 4548
rect 27620 4496 27672 4548
rect 29276 4607 29328 4616
rect 29276 4573 29285 4607
rect 29285 4573 29319 4607
rect 29319 4573 29328 4607
rect 29276 4564 29328 4573
rect 30196 4632 30248 4684
rect 31392 4632 31444 4684
rect 31576 4632 31628 4684
rect 37924 4700 37976 4752
rect 40592 4768 40644 4820
rect 41788 4811 41840 4820
rect 41788 4777 41797 4811
rect 41797 4777 41831 4811
rect 41831 4777 41840 4811
rect 41788 4768 41840 4777
rect 42248 4811 42300 4820
rect 42248 4777 42257 4811
rect 42257 4777 42291 4811
rect 42291 4777 42300 4811
rect 42892 4811 42944 4820
rect 42248 4768 42300 4777
rect 42892 4777 42901 4811
rect 42901 4777 42935 4811
rect 42935 4777 42944 4811
rect 42892 4768 42944 4777
rect 42984 4768 43036 4820
rect 44088 4768 44140 4820
rect 34428 4632 34480 4684
rect 36360 4675 36412 4684
rect 36360 4641 36369 4675
rect 36369 4641 36403 4675
rect 36403 4641 36412 4675
rect 36360 4632 36412 4641
rect 36544 4675 36596 4684
rect 36544 4641 36553 4675
rect 36553 4641 36587 4675
rect 36587 4641 36596 4675
rect 36544 4632 36596 4641
rect 37004 4632 37056 4684
rect 26792 4428 26844 4480
rect 29092 4428 29144 4480
rect 30840 4496 30892 4548
rect 34060 4607 34112 4616
rect 34060 4573 34069 4607
rect 34069 4573 34103 4607
rect 34103 4573 34112 4607
rect 34060 4564 34112 4573
rect 36084 4564 36136 4616
rect 36912 4564 36964 4616
rect 37188 4564 37240 4616
rect 39212 4632 39264 4684
rect 39856 4700 39908 4752
rect 40408 4700 40460 4752
rect 30656 4428 30708 4480
rect 30932 4471 30984 4480
rect 30932 4437 30941 4471
rect 30941 4437 30975 4471
rect 30975 4437 30984 4471
rect 30932 4428 30984 4437
rect 31392 4471 31444 4480
rect 31392 4437 31401 4471
rect 31401 4437 31435 4471
rect 31435 4437 31444 4471
rect 31392 4428 31444 4437
rect 32588 4428 32640 4480
rect 33048 4496 33100 4548
rect 35716 4496 35768 4548
rect 37740 4539 37792 4548
rect 37740 4505 37749 4539
rect 37749 4505 37783 4539
rect 37783 4505 37792 4539
rect 37740 4496 37792 4505
rect 35348 4428 35400 4480
rect 35808 4471 35860 4480
rect 35808 4437 35817 4471
rect 35817 4437 35851 4471
rect 35851 4437 35860 4471
rect 40040 4632 40092 4684
rect 43996 4743 44048 4752
rect 43996 4709 44005 4743
rect 44005 4709 44039 4743
rect 44039 4709 44048 4743
rect 43996 4700 44048 4709
rect 42524 4632 42576 4684
rect 43444 4632 43496 4684
rect 39948 4564 40000 4616
rect 40868 4496 40920 4548
rect 41512 4539 41564 4548
rect 41512 4505 41521 4539
rect 41521 4505 41555 4539
rect 41555 4505 41564 4539
rect 41512 4496 41564 4505
rect 35808 4428 35860 4437
rect 40040 4471 40092 4480
rect 40040 4437 40049 4471
rect 40049 4437 40083 4471
rect 40083 4437 40092 4471
rect 40040 4428 40092 4437
rect 40500 4471 40552 4480
rect 40500 4437 40509 4471
rect 40509 4437 40543 4471
rect 40543 4437 40552 4471
rect 40500 4428 40552 4437
rect 6070 4326 6122 4378
rect 6134 4326 6186 4378
rect 6198 4326 6250 4378
rect 6262 4326 6314 4378
rect 6326 4326 6378 4378
rect 11070 4326 11122 4378
rect 11134 4326 11186 4378
rect 11198 4326 11250 4378
rect 11262 4326 11314 4378
rect 11326 4326 11378 4378
rect 16070 4326 16122 4378
rect 16134 4326 16186 4378
rect 16198 4326 16250 4378
rect 16262 4326 16314 4378
rect 16326 4326 16378 4378
rect 21070 4326 21122 4378
rect 21134 4326 21186 4378
rect 21198 4326 21250 4378
rect 21262 4326 21314 4378
rect 21326 4326 21378 4378
rect 26070 4326 26122 4378
rect 26134 4326 26186 4378
rect 26198 4326 26250 4378
rect 26262 4326 26314 4378
rect 26326 4326 26378 4378
rect 31070 4326 31122 4378
rect 31134 4326 31186 4378
rect 31198 4326 31250 4378
rect 31262 4326 31314 4378
rect 31326 4326 31378 4378
rect 36070 4326 36122 4378
rect 36134 4326 36186 4378
rect 36198 4326 36250 4378
rect 36262 4326 36314 4378
rect 36326 4326 36378 4378
rect 41070 4326 41122 4378
rect 41134 4326 41186 4378
rect 41198 4326 41250 4378
rect 41262 4326 41314 4378
rect 41326 4326 41378 4378
rect 1492 4156 1544 4208
rect 2596 4088 2648 4140
rect 4344 4156 4396 4208
rect 4712 4224 4764 4276
rect 5540 4224 5592 4276
rect 5908 4224 5960 4276
rect 940 3952 992 4004
rect 5080 4088 5132 4140
rect 9128 4224 9180 4276
rect 9588 4224 9640 4276
rect 11704 4224 11756 4276
rect 12532 4224 12584 4276
rect 14280 4224 14332 4276
rect 14372 4224 14424 4276
rect 15752 4224 15804 4276
rect 22284 4224 22336 4276
rect 22376 4224 22428 4276
rect 23480 4224 23532 4276
rect 24124 4224 24176 4276
rect 25596 4224 25648 4276
rect 26424 4224 26476 4276
rect 26700 4224 26752 4276
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 8300 4156 8352 4208
rect 6460 4088 6512 4097
rect 7932 4088 7984 4140
rect 3332 3995 3384 4004
rect 3332 3961 3341 3995
rect 3341 3961 3375 3995
rect 3375 3961 3384 3995
rect 5356 4020 5408 4072
rect 6920 4020 6972 4072
rect 3332 3952 3384 3961
rect 2780 3884 2832 3936
rect 6644 3884 6696 3936
rect 10232 4088 10284 4140
rect 12072 4156 12124 4208
rect 12900 4088 12952 4140
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 13268 4020 13320 4072
rect 8392 3884 8444 3936
rect 8944 3884 8996 3936
rect 9036 3884 9088 3936
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 12532 3884 12584 3936
rect 12992 3884 13044 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 14464 4088 14516 4140
rect 15936 4156 15988 4208
rect 15200 4088 15252 4140
rect 16212 4088 16264 4140
rect 16580 4156 16632 4208
rect 16764 4156 16816 4208
rect 17132 4156 17184 4208
rect 19064 4156 19116 4208
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 20352 4156 20404 4208
rect 20076 4088 20128 4140
rect 20444 4088 20496 4140
rect 20536 4088 20588 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 23112 4088 23164 4140
rect 23848 4088 23900 4140
rect 24308 4088 24360 4140
rect 24400 4088 24452 4140
rect 25136 4156 25188 4208
rect 25872 4156 25924 4208
rect 14004 4020 14056 4072
rect 16304 4063 16356 4072
rect 16304 4029 16313 4063
rect 16313 4029 16347 4063
rect 16347 4029 16356 4063
rect 16304 4020 16356 4029
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 17684 4020 17736 4072
rect 19156 4020 19208 4072
rect 20720 4020 20772 4072
rect 21548 4063 21600 4072
rect 21548 4029 21557 4063
rect 21557 4029 21591 4063
rect 21591 4029 21600 4063
rect 21548 4020 21600 4029
rect 13912 3952 13964 4004
rect 14096 3884 14148 3936
rect 15844 3884 15896 3936
rect 19708 3884 19760 3936
rect 22192 3884 22244 3936
rect 22284 3884 22336 3936
rect 23940 4020 23992 4072
rect 23112 3952 23164 4004
rect 25688 4131 25740 4140
rect 25688 4097 25697 4131
rect 25697 4097 25731 4131
rect 25731 4097 25740 4131
rect 25688 4088 25740 4097
rect 25780 4131 25832 4140
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 25964 4020 26016 4072
rect 25872 3952 25924 4004
rect 27620 4224 27672 4276
rect 28264 4224 28316 4276
rect 27712 4199 27764 4208
rect 27712 4165 27721 4199
rect 27721 4165 27755 4199
rect 27755 4165 27764 4199
rect 27712 4156 27764 4165
rect 28080 4156 28132 4208
rect 26700 4131 26752 4140
rect 26700 4097 26709 4131
rect 26709 4097 26743 4131
rect 26743 4097 26752 4131
rect 26700 4088 26752 4097
rect 26608 3952 26660 4004
rect 27252 4131 27304 4140
rect 27252 4097 27261 4131
rect 27261 4097 27295 4131
rect 27295 4097 27304 4131
rect 27252 4088 27304 4097
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 28172 4088 28224 4140
rect 28724 4156 28776 4208
rect 29184 4224 29236 4276
rect 29644 4224 29696 4276
rect 30932 4224 30984 4276
rect 31024 4267 31076 4276
rect 31024 4233 31033 4267
rect 31033 4233 31067 4267
rect 31067 4233 31076 4267
rect 31024 4224 31076 4233
rect 33324 4224 33376 4276
rect 28632 4088 28684 4140
rect 27528 4020 27580 4072
rect 27988 4020 28040 4072
rect 29276 4131 29328 4140
rect 29276 4097 29285 4131
rect 29285 4097 29319 4131
rect 29319 4097 29328 4131
rect 29276 4088 29328 4097
rect 29736 4131 29788 4140
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 29368 4020 29420 4072
rect 32404 4156 32456 4208
rect 30196 4131 30248 4140
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 30840 4088 30892 4140
rect 30932 4088 30984 4140
rect 32220 4131 32272 4140
rect 32220 4097 32229 4131
rect 32229 4097 32263 4131
rect 32263 4097 32272 4131
rect 32220 4088 32272 4097
rect 33416 4088 33468 4140
rect 34152 4156 34204 4208
rect 35992 4156 36044 4208
rect 30656 4020 30708 4072
rect 31208 3952 31260 4004
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 26424 3884 26476 3936
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 28448 3884 28500 3936
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 29460 3884 29512 3936
rect 29552 3927 29604 3936
rect 29552 3893 29561 3927
rect 29561 3893 29595 3927
rect 29595 3893 29604 3927
rect 29552 3884 29604 3893
rect 30012 3927 30064 3936
rect 30012 3893 30021 3927
rect 30021 3893 30055 3927
rect 30055 3893 30064 3927
rect 30012 3884 30064 3893
rect 30472 3884 30524 3936
rect 30564 3927 30616 3936
rect 30564 3893 30573 3927
rect 30573 3893 30607 3927
rect 30607 3893 30616 3927
rect 30564 3884 30616 3893
rect 31852 3995 31904 4004
rect 31852 3961 31861 3995
rect 31861 3961 31895 3995
rect 31895 3961 31904 3995
rect 31852 3952 31904 3961
rect 33140 4020 33192 4072
rect 35900 4088 35952 4140
rect 37280 4156 37332 4208
rect 37464 4088 37516 4140
rect 38292 4156 38344 4208
rect 39948 4224 40000 4276
rect 40500 4224 40552 4276
rect 40960 4224 41012 4276
rect 41880 4224 41932 4276
rect 41972 4267 42024 4276
rect 41972 4233 41981 4267
rect 41981 4233 42015 4267
rect 42015 4233 42024 4267
rect 41972 4224 42024 4233
rect 42984 4224 43036 4276
rect 43444 4267 43496 4276
rect 43444 4233 43453 4267
rect 43453 4233 43487 4267
rect 43487 4233 43496 4267
rect 43444 4224 43496 4233
rect 43996 4224 44048 4276
rect 44732 4224 44784 4276
rect 39396 4088 39448 4140
rect 40224 4088 40276 4140
rect 40316 4131 40368 4140
rect 40316 4097 40325 4131
rect 40325 4097 40359 4131
rect 40359 4097 40368 4131
rect 40316 4088 40368 4097
rect 41788 4156 41840 4208
rect 34152 4063 34204 4072
rect 34152 4029 34161 4063
rect 34161 4029 34195 4063
rect 34195 4029 34204 4063
rect 34152 4020 34204 4029
rect 34428 4063 34480 4072
rect 34428 4029 34437 4063
rect 34437 4029 34471 4063
rect 34471 4029 34480 4063
rect 34428 4020 34480 4029
rect 36452 4020 36504 4072
rect 38384 4063 38436 4072
rect 38384 4029 38393 4063
rect 38393 4029 38427 4063
rect 38427 4029 38436 4063
rect 38384 4020 38436 4029
rect 39764 4020 39816 4072
rect 33968 3995 34020 4004
rect 33968 3961 33977 3995
rect 33977 3961 34011 3995
rect 34011 3961 34020 3995
rect 33968 3952 34020 3961
rect 35900 3927 35952 3936
rect 35900 3893 35909 3927
rect 35909 3893 35943 3927
rect 35943 3893 35952 3927
rect 35900 3884 35952 3893
rect 36820 3995 36872 4004
rect 36820 3961 36829 3995
rect 36829 3961 36863 3995
rect 36863 3961 36872 3995
rect 36820 3952 36872 3961
rect 37924 3927 37976 3936
rect 37924 3893 37933 3927
rect 37933 3893 37967 3927
rect 37967 3893 37976 3927
rect 37924 3884 37976 3893
rect 38200 3884 38252 3936
rect 39948 3927 40000 3936
rect 39948 3893 39957 3927
rect 39957 3893 39991 3927
rect 39991 3893 40000 3927
rect 39948 3884 40000 3893
rect 40868 3884 40920 3936
rect 3570 3782 3622 3834
rect 3634 3782 3686 3834
rect 3698 3782 3750 3834
rect 3762 3782 3814 3834
rect 3826 3782 3878 3834
rect 8570 3782 8622 3834
rect 8634 3782 8686 3834
rect 8698 3782 8750 3834
rect 8762 3782 8814 3834
rect 8826 3782 8878 3834
rect 13570 3782 13622 3834
rect 13634 3782 13686 3834
rect 13698 3782 13750 3834
rect 13762 3782 13814 3834
rect 13826 3782 13878 3834
rect 18570 3782 18622 3834
rect 18634 3782 18686 3834
rect 18698 3782 18750 3834
rect 18762 3782 18814 3834
rect 18826 3782 18878 3834
rect 23570 3782 23622 3834
rect 23634 3782 23686 3834
rect 23698 3782 23750 3834
rect 23762 3782 23814 3834
rect 23826 3782 23878 3834
rect 28570 3782 28622 3834
rect 28634 3782 28686 3834
rect 28698 3782 28750 3834
rect 28762 3782 28814 3834
rect 28826 3782 28878 3834
rect 33570 3782 33622 3834
rect 33634 3782 33686 3834
rect 33698 3782 33750 3834
rect 33762 3782 33814 3834
rect 33826 3782 33878 3834
rect 38570 3782 38622 3834
rect 38634 3782 38686 3834
rect 38698 3782 38750 3834
rect 38762 3782 38814 3834
rect 38826 3782 38878 3834
rect 43570 3782 43622 3834
rect 43634 3782 43686 3834
rect 43698 3782 43750 3834
rect 43762 3782 43814 3834
rect 43826 3782 43878 3834
rect 4620 3680 4672 3732
rect 5724 3680 5776 3732
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 6460 3680 6512 3732
rect 7932 3680 7984 3732
rect 9036 3680 9088 3732
rect 11244 3680 11296 3732
rect 12164 3680 12216 3732
rect 13268 3680 13320 3732
rect 14832 3723 14884 3732
rect 14832 3689 14841 3723
rect 14841 3689 14875 3723
rect 14875 3689 14884 3723
rect 14832 3680 14884 3689
rect 1584 3612 1636 3664
rect 9680 3612 9732 3664
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 9312 3544 9364 3596
rect 10600 3544 10652 3596
rect 10968 3544 11020 3596
rect 19064 3680 19116 3732
rect 19248 3680 19300 3732
rect 21732 3680 21784 3732
rect 21824 3680 21876 3732
rect 23388 3680 23440 3732
rect 16304 3612 16356 3664
rect 14004 3544 14056 3596
rect 16672 3544 16724 3596
rect 18328 3612 18380 3664
rect 1492 3476 1544 3528
rect 2596 3476 2648 3528
rect 4712 3476 4764 3528
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 6644 3408 6696 3460
rect 4436 3340 4488 3392
rect 6460 3340 6512 3392
rect 7196 3476 7248 3528
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 8576 3451 8628 3460
rect 8576 3417 8585 3451
rect 8585 3417 8619 3451
rect 8619 3417 8628 3451
rect 8576 3408 8628 3417
rect 10140 3408 10192 3460
rect 12900 3476 12952 3528
rect 13912 3519 13964 3528
rect 13912 3485 13921 3519
rect 13921 3485 13955 3519
rect 13955 3485 13964 3519
rect 13912 3476 13964 3485
rect 14924 3476 14976 3528
rect 17040 3476 17092 3528
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 18328 3476 18380 3528
rect 11520 3408 11572 3460
rect 11888 3408 11940 3460
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 13176 3340 13228 3392
rect 14004 3383 14056 3392
rect 14004 3349 14013 3383
rect 14013 3349 14047 3383
rect 14047 3349 14056 3383
rect 14004 3340 14056 3349
rect 15292 3451 15344 3460
rect 15292 3417 15301 3451
rect 15301 3417 15335 3451
rect 15335 3417 15344 3451
rect 15292 3408 15344 3417
rect 16304 3340 16356 3392
rect 16580 3340 16632 3392
rect 16856 3383 16908 3392
rect 16856 3349 16865 3383
rect 16865 3349 16899 3383
rect 16899 3349 16908 3383
rect 16856 3340 16908 3349
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 19064 3519 19116 3528
rect 19064 3485 19073 3519
rect 19073 3485 19107 3519
rect 19107 3485 19116 3519
rect 19064 3476 19116 3485
rect 19248 3544 19300 3596
rect 20720 3544 20772 3596
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 22008 3544 22060 3596
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 18788 3408 18840 3460
rect 19156 3451 19208 3460
rect 19156 3417 19165 3451
rect 19165 3417 19199 3451
rect 19199 3417 19208 3451
rect 19156 3408 19208 3417
rect 21916 3476 21968 3528
rect 20536 3408 20588 3460
rect 20628 3451 20680 3460
rect 20628 3417 20637 3451
rect 20637 3417 20671 3451
rect 20671 3417 20680 3451
rect 20628 3408 20680 3417
rect 22376 3408 22428 3460
rect 23112 3476 23164 3528
rect 19892 3340 19944 3392
rect 20996 3340 21048 3392
rect 23940 3544 23992 3596
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 24032 3476 24084 3528
rect 24952 3544 25004 3596
rect 27252 3680 27304 3732
rect 28448 3680 28500 3732
rect 28540 3612 28592 3664
rect 29092 3612 29144 3664
rect 23020 3383 23072 3392
rect 23020 3349 23029 3383
rect 23029 3349 23063 3383
rect 23063 3349 23072 3383
rect 23020 3340 23072 3349
rect 23480 3340 23532 3392
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 24676 3383 24728 3392
rect 24676 3349 24685 3383
rect 24685 3349 24719 3383
rect 24719 3349 24728 3383
rect 24676 3340 24728 3349
rect 26332 3476 26384 3528
rect 26792 3544 26844 3596
rect 27344 3544 27396 3596
rect 25136 3408 25188 3460
rect 27344 3408 27396 3460
rect 27436 3451 27488 3460
rect 27436 3417 27477 3451
rect 27477 3417 27488 3451
rect 27896 3519 27948 3528
rect 27896 3485 27905 3519
rect 27905 3485 27939 3519
rect 27939 3485 27948 3519
rect 27896 3476 27948 3485
rect 28080 3544 28132 3596
rect 28172 3587 28224 3596
rect 28172 3553 28181 3587
rect 28181 3553 28215 3587
rect 28215 3553 28224 3587
rect 28172 3544 28224 3553
rect 29644 3680 29696 3732
rect 30012 3680 30064 3732
rect 31208 3680 31260 3732
rect 30840 3612 30892 3664
rect 28356 3476 28408 3528
rect 28448 3519 28500 3528
rect 28448 3485 28457 3519
rect 28457 3485 28491 3519
rect 28491 3485 28500 3519
rect 28448 3476 28500 3485
rect 29552 3544 29604 3596
rect 30656 3544 30708 3596
rect 31024 3544 31076 3596
rect 27436 3408 27488 3417
rect 27712 3408 27764 3460
rect 29000 3476 29052 3528
rect 29092 3519 29144 3528
rect 29092 3485 29101 3519
rect 29101 3485 29135 3519
rect 29135 3485 29144 3519
rect 29092 3476 29144 3485
rect 30840 3476 30892 3528
rect 31944 3680 31996 3732
rect 32404 3723 32456 3732
rect 32404 3689 32413 3723
rect 32413 3689 32447 3723
rect 32447 3689 32456 3723
rect 32404 3680 32456 3689
rect 32956 3680 33008 3732
rect 33232 3680 33284 3732
rect 34428 3680 34480 3732
rect 35900 3680 35952 3732
rect 38384 3680 38436 3732
rect 32680 3544 32732 3596
rect 32864 3587 32916 3596
rect 32864 3553 32873 3587
rect 32873 3553 32907 3587
rect 32907 3553 32916 3587
rect 32864 3544 32916 3553
rect 33140 3544 33192 3596
rect 31944 3476 31996 3528
rect 29368 3408 29420 3460
rect 29552 3408 29604 3460
rect 25228 3340 25280 3392
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 25688 3340 25740 3392
rect 25964 3340 26016 3392
rect 27068 3340 27120 3392
rect 27620 3383 27672 3392
rect 27620 3349 27629 3383
rect 27629 3349 27663 3383
rect 27663 3349 27672 3383
rect 27620 3340 27672 3349
rect 28264 3383 28316 3392
rect 28264 3349 28273 3383
rect 28273 3349 28307 3383
rect 28307 3349 28316 3383
rect 28264 3340 28316 3349
rect 28908 3340 28960 3392
rect 29276 3340 29328 3392
rect 29460 3340 29512 3392
rect 31392 3408 31444 3460
rect 31760 3451 31812 3460
rect 31760 3417 31769 3451
rect 31769 3417 31803 3451
rect 31803 3417 31812 3451
rect 31760 3408 31812 3417
rect 32312 3519 32364 3528
rect 32312 3485 32321 3519
rect 32321 3485 32355 3519
rect 32355 3485 32364 3519
rect 32312 3476 32364 3485
rect 33416 3519 33468 3528
rect 33416 3485 33425 3519
rect 33425 3485 33459 3519
rect 33459 3485 33468 3519
rect 33416 3476 33468 3485
rect 34612 3519 34664 3528
rect 34612 3485 34621 3519
rect 34621 3485 34655 3519
rect 34655 3485 34664 3519
rect 34612 3476 34664 3485
rect 32036 3383 32088 3392
rect 32036 3349 32045 3383
rect 32045 3349 32079 3383
rect 32079 3349 32088 3383
rect 32036 3340 32088 3349
rect 33140 3408 33192 3460
rect 33692 3451 33744 3460
rect 33692 3417 33701 3451
rect 33701 3417 33735 3451
rect 33735 3417 33744 3451
rect 33692 3408 33744 3417
rect 32772 3383 32824 3392
rect 32772 3349 32781 3383
rect 32781 3349 32815 3383
rect 32815 3349 32824 3383
rect 32772 3340 32824 3349
rect 33048 3340 33100 3392
rect 34428 3383 34480 3392
rect 34428 3349 34437 3383
rect 34437 3349 34471 3383
rect 34471 3349 34480 3383
rect 34428 3340 34480 3349
rect 35716 3587 35768 3596
rect 35716 3553 35725 3587
rect 35725 3553 35759 3587
rect 35759 3553 35768 3587
rect 35716 3544 35768 3553
rect 36544 3587 36596 3596
rect 36544 3553 36553 3587
rect 36553 3553 36587 3587
rect 36587 3553 36596 3587
rect 36544 3544 36596 3553
rect 35808 3476 35860 3528
rect 35900 3476 35952 3528
rect 37004 3476 37056 3528
rect 38200 3587 38252 3596
rect 38200 3553 38209 3587
rect 38209 3553 38243 3587
rect 38243 3553 38252 3587
rect 38200 3544 38252 3553
rect 39948 3680 40000 3732
rect 40960 3723 41012 3732
rect 40960 3689 40969 3723
rect 40969 3689 41003 3723
rect 41003 3689 41012 3723
rect 40960 3680 41012 3689
rect 41880 3680 41932 3732
rect 44548 3680 44600 3732
rect 44824 3680 44876 3732
rect 44916 3723 44968 3732
rect 44916 3689 44925 3723
rect 44925 3689 44959 3723
rect 44959 3689 44968 3723
rect 44916 3680 44968 3689
rect 40592 3612 40644 3664
rect 42248 3612 42300 3664
rect 40040 3544 40092 3596
rect 40224 3544 40276 3596
rect 42524 3612 42576 3664
rect 43352 3612 43404 3664
rect 44732 3612 44784 3664
rect 37188 3451 37240 3460
rect 37188 3417 37197 3451
rect 37197 3417 37231 3451
rect 37231 3417 37240 3451
rect 37188 3408 37240 3417
rect 38752 3408 38804 3460
rect 35992 3340 36044 3392
rect 36728 3340 36780 3392
rect 36820 3383 36872 3392
rect 36820 3349 36829 3383
rect 36829 3349 36863 3383
rect 36863 3349 36872 3383
rect 36820 3340 36872 3349
rect 37280 3383 37332 3392
rect 37280 3349 37289 3383
rect 37289 3349 37323 3383
rect 37323 3349 37332 3383
rect 37280 3340 37332 3349
rect 37648 3383 37700 3392
rect 37648 3349 37657 3383
rect 37657 3349 37691 3383
rect 37691 3349 37700 3383
rect 37648 3340 37700 3349
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 38108 3383 38160 3392
rect 38108 3349 38117 3383
rect 38117 3349 38151 3383
rect 38151 3349 38160 3383
rect 38108 3340 38160 3349
rect 6070 3238 6122 3290
rect 6134 3238 6186 3290
rect 6198 3238 6250 3290
rect 6262 3238 6314 3290
rect 6326 3238 6378 3290
rect 11070 3238 11122 3290
rect 11134 3238 11186 3290
rect 11198 3238 11250 3290
rect 11262 3238 11314 3290
rect 11326 3238 11378 3290
rect 16070 3238 16122 3290
rect 16134 3238 16186 3290
rect 16198 3238 16250 3290
rect 16262 3238 16314 3290
rect 16326 3238 16378 3290
rect 21070 3238 21122 3290
rect 21134 3238 21186 3290
rect 21198 3238 21250 3290
rect 21262 3238 21314 3290
rect 21326 3238 21378 3290
rect 26070 3238 26122 3290
rect 26134 3238 26186 3290
rect 26198 3238 26250 3290
rect 26262 3238 26314 3290
rect 26326 3238 26378 3290
rect 31070 3238 31122 3290
rect 31134 3238 31186 3290
rect 31198 3238 31250 3290
rect 31262 3238 31314 3290
rect 31326 3238 31378 3290
rect 36070 3238 36122 3290
rect 36134 3238 36186 3290
rect 36198 3238 36250 3290
rect 36262 3238 36314 3290
rect 36326 3238 36378 3290
rect 41070 3238 41122 3290
rect 41134 3238 41186 3290
rect 41198 3238 41250 3290
rect 41262 3238 41314 3290
rect 41326 3238 41378 3290
rect 1308 3136 1360 3188
rect 1584 3136 1636 3188
rect 2596 3136 2648 3188
rect 756 3043 808 3052
rect 756 3009 765 3043
rect 765 3009 799 3043
rect 799 3009 808 3043
rect 756 3000 808 3009
rect 4160 3136 4212 3188
rect 4436 3179 4488 3188
rect 4436 3145 4445 3179
rect 4445 3145 4479 3179
rect 4479 3145 4488 3179
rect 4436 3136 4488 3145
rect 5724 3136 5776 3188
rect 6460 3136 6512 3188
rect 7196 3136 7248 3188
rect 8576 3136 8628 3188
rect 10600 3136 10652 3188
rect 13176 3136 13228 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 15292 3136 15344 3188
rect 16856 3136 16908 3188
rect 4068 3068 4120 3120
rect 6644 3068 6696 3120
rect 11796 3068 11848 3120
rect 18236 3136 18288 3188
rect 18328 3136 18380 3188
rect 19340 3136 19392 3188
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 8300 3000 8352 3052
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 9956 3000 10008 3052
rect 11336 3043 11388 3052
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 14096 3000 14148 3052
rect 17776 3068 17828 3120
rect 19432 3068 19484 3120
rect 19892 3136 19944 3188
rect 20536 3136 20588 3188
rect 20628 3136 20680 3188
rect 23020 3136 23072 3188
rect 21548 3068 21600 3120
rect 21916 3068 21968 3120
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 3976 2932 4028 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9312 2932 9364 2984
rect 2412 2796 2464 2848
rect 8300 2907 8352 2916
rect 8300 2873 8309 2907
rect 8309 2873 8343 2907
rect 8343 2873 8352 2907
rect 8300 2864 8352 2873
rect 10968 2932 11020 2984
rect 11888 2932 11940 2984
rect 12348 2932 12400 2984
rect 13360 2932 13412 2984
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 16672 3000 16724 3052
rect 16764 3000 16816 3052
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 18788 3000 18840 3052
rect 20536 3000 20588 3052
rect 23480 3068 23532 3120
rect 24308 3068 24360 3120
rect 24676 3136 24728 3188
rect 24768 3136 24820 3188
rect 25688 3136 25740 3188
rect 25964 3136 26016 3188
rect 26608 3136 26660 3188
rect 27528 3136 27580 3188
rect 29736 3179 29788 3188
rect 29736 3145 29745 3179
rect 29745 3145 29779 3179
rect 29779 3145 29788 3179
rect 29736 3136 29788 3145
rect 2964 2796 3016 2848
rect 3332 2796 3384 2848
rect 11428 2796 11480 2848
rect 12348 2839 12400 2848
rect 12348 2805 12357 2839
rect 12357 2805 12391 2839
rect 12391 2805 12400 2839
rect 12348 2796 12400 2805
rect 12440 2839 12492 2848
rect 12440 2805 12449 2839
rect 12449 2805 12483 2839
rect 12483 2805 12492 2839
rect 12440 2796 12492 2805
rect 14832 2839 14884 2848
rect 14832 2805 14841 2839
rect 14841 2805 14875 2839
rect 14875 2805 14884 2839
rect 14832 2796 14884 2805
rect 14924 2796 14976 2848
rect 19156 2932 19208 2984
rect 19892 2932 19944 2984
rect 20444 2932 20496 2984
rect 21088 2932 21140 2984
rect 20720 2864 20772 2916
rect 22744 2932 22796 2984
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 25412 3000 25464 3052
rect 25872 3000 25924 3052
rect 26424 3000 26476 3052
rect 26884 3068 26936 3120
rect 30564 3136 30616 3188
rect 32036 3136 32088 3188
rect 32680 3136 32732 3188
rect 34612 3136 34664 3188
rect 35808 3136 35860 3188
rect 32956 3068 33008 3120
rect 35256 3068 35308 3120
rect 28172 3000 28224 3052
rect 29276 3000 29328 3052
rect 25596 2932 25648 2984
rect 21180 2796 21232 2848
rect 21916 2796 21968 2848
rect 22008 2796 22060 2848
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 26332 2839 26384 2848
rect 26332 2805 26341 2839
rect 26341 2805 26375 2839
rect 26375 2805 26384 2839
rect 26332 2796 26384 2805
rect 27436 2932 27488 2984
rect 28264 2932 28316 2984
rect 28540 2932 28592 2984
rect 29552 3000 29604 3052
rect 30104 3043 30156 3052
rect 30104 3009 30113 3043
rect 30113 3009 30147 3043
rect 30147 3009 30156 3043
rect 30104 3000 30156 3009
rect 30288 3000 30340 3052
rect 30380 3043 30432 3052
rect 30380 3009 30389 3043
rect 30389 3009 30423 3043
rect 30423 3009 30432 3043
rect 30380 3000 30432 3009
rect 30472 3000 30524 3052
rect 31484 3000 31536 3052
rect 33508 3043 33560 3052
rect 33508 3009 33517 3043
rect 33517 3009 33551 3043
rect 33551 3009 33560 3043
rect 33508 3000 33560 3009
rect 35992 3136 36044 3188
rect 36820 3136 36872 3188
rect 37004 3136 37056 3188
rect 37464 3068 37516 3120
rect 27896 2864 27948 2916
rect 27988 2796 28040 2848
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 29184 2796 29236 2848
rect 29460 2796 29512 2848
rect 29644 2796 29696 2848
rect 30104 2864 30156 2916
rect 31300 2932 31352 2984
rect 31484 2864 31536 2916
rect 34520 2932 34572 2984
rect 35900 2932 35952 2984
rect 30840 2796 30892 2848
rect 31668 2796 31720 2848
rect 33784 2864 33836 2916
rect 38292 3000 38344 3052
rect 38752 3068 38804 3120
rect 39028 3068 39080 3120
rect 39396 3068 39448 3120
rect 40316 3136 40368 3188
rect 41880 3136 41932 3188
rect 44732 3179 44784 3188
rect 44732 3145 44741 3179
rect 44741 3145 44775 3179
rect 44775 3145 44784 3179
rect 44732 3136 44784 3145
rect 40592 3068 40644 3120
rect 42248 3068 42300 3120
rect 40132 3000 40184 3052
rect 41420 3000 41472 3052
rect 44640 3000 44692 3052
rect 36360 2932 36412 2984
rect 37280 2932 37332 2984
rect 38752 2975 38804 2984
rect 38752 2941 38761 2975
rect 38761 2941 38795 2975
rect 38795 2941 38804 2975
rect 38752 2932 38804 2941
rect 40500 2932 40552 2984
rect 40868 2975 40920 2984
rect 40868 2941 40877 2975
rect 40877 2941 40911 2975
rect 40911 2941 40920 2975
rect 40868 2932 40920 2941
rect 34060 2796 34112 2848
rect 35808 2839 35860 2848
rect 35808 2805 35817 2839
rect 35817 2805 35851 2839
rect 35851 2805 35860 2839
rect 35808 2796 35860 2805
rect 35992 2796 36044 2848
rect 38292 2796 38344 2848
rect 39396 2796 39448 2848
rect 3570 2694 3622 2746
rect 3634 2694 3686 2746
rect 3698 2694 3750 2746
rect 3762 2694 3814 2746
rect 3826 2694 3878 2746
rect 8570 2694 8622 2746
rect 8634 2694 8686 2746
rect 8698 2694 8750 2746
rect 8762 2694 8814 2746
rect 8826 2694 8878 2746
rect 13570 2694 13622 2746
rect 13634 2694 13686 2746
rect 13698 2694 13750 2746
rect 13762 2694 13814 2746
rect 13826 2694 13878 2746
rect 18570 2694 18622 2746
rect 18634 2694 18686 2746
rect 18698 2694 18750 2746
rect 18762 2694 18814 2746
rect 18826 2694 18878 2746
rect 23570 2694 23622 2746
rect 23634 2694 23686 2746
rect 23698 2694 23750 2746
rect 23762 2694 23814 2746
rect 23826 2694 23878 2746
rect 28570 2694 28622 2746
rect 28634 2694 28686 2746
rect 28698 2694 28750 2746
rect 28762 2694 28814 2746
rect 28826 2694 28878 2746
rect 33570 2694 33622 2746
rect 33634 2694 33686 2746
rect 33698 2694 33750 2746
rect 33762 2694 33814 2746
rect 33826 2694 33878 2746
rect 38570 2694 38622 2746
rect 38634 2694 38686 2746
rect 38698 2694 38750 2746
rect 38762 2694 38814 2746
rect 38826 2694 38878 2746
rect 43570 2694 43622 2746
rect 43634 2694 43686 2746
rect 43698 2694 43750 2746
rect 43762 2694 43814 2746
rect 43826 2694 43878 2746
rect 1492 2635 1544 2644
rect 1492 2601 1501 2635
rect 1501 2601 1535 2635
rect 1535 2601 1544 2635
rect 1492 2592 1544 2601
rect 1768 2592 1820 2644
rect 2780 2592 2832 2644
rect 8484 2592 8536 2644
rect 1308 2524 1360 2576
rect 7012 2567 7064 2576
rect 7012 2533 7021 2567
rect 7021 2533 7055 2567
rect 7055 2533 7064 2567
rect 7012 2524 7064 2533
rect 2412 2456 2464 2508
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 11796 2635 11848 2644
rect 11796 2601 11805 2635
rect 11805 2601 11839 2635
rect 11839 2601 11848 2635
rect 11796 2592 11848 2601
rect 11888 2592 11940 2644
rect 12624 2524 12676 2576
rect 14096 2524 14148 2576
rect 15936 2592 15988 2644
rect 16488 2592 16540 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20352 2592 20404 2644
rect 22284 2592 22336 2644
rect 22560 2592 22612 2644
rect 24216 2592 24268 2644
rect 25688 2592 25740 2644
rect 1676 2252 1728 2304
rect 2504 2388 2556 2440
rect 2964 2388 3016 2440
rect 4712 2388 4764 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 9864 2456 9916 2508
rect 3424 2363 3476 2372
rect 3424 2329 3433 2363
rect 3433 2329 3467 2363
rect 3467 2329 3476 2363
rect 3424 2320 3476 2329
rect 4068 2252 4120 2304
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6000 2252 6052 2304
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 14188 2456 14240 2508
rect 14924 2456 14976 2508
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 18512 2456 18564 2508
rect 19248 2499 19300 2508
rect 19248 2465 19257 2499
rect 19257 2465 19291 2499
rect 19291 2465 19300 2499
rect 19248 2456 19300 2465
rect 19708 2456 19760 2508
rect 19800 2456 19852 2508
rect 21180 2456 21232 2508
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 11888 2388 11940 2440
rect 14004 2388 14056 2440
rect 24124 2456 24176 2508
rect 25596 2499 25648 2508
rect 25596 2465 25605 2499
rect 25605 2465 25639 2499
rect 25639 2465 25648 2499
rect 25596 2456 25648 2465
rect 26332 2456 26384 2508
rect 27252 2592 27304 2644
rect 27528 2635 27580 2644
rect 27528 2601 27537 2635
rect 27537 2601 27571 2635
rect 27571 2601 27580 2635
rect 27528 2592 27580 2601
rect 27160 2524 27212 2576
rect 29000 2592 29052 2644
rect 33232 2592 33284 2644
rect 21548 2388 21600 2440
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 26884 2388 26936 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 27712 2499 27764 2508
rect 27712 2465 27721 2499
rect 27721 2465 27755 2499
rect 27755 2465 27764 2499
rect 27712 2456 27764 2465
rect 29368 2567 29420 2576
rect 29368 2533 29377 2567
rect 29377 2533 29411 2567
rect 29411 2533 29420 2567
rect 29368 2524 29420 2533
rect 30104 2567 30156 2576
rect 30104 2533 30113 2567
rect 30113 2533 30147 2567
rect 30147 2533 30156 2567
rect 30104 2524 30156 2533
rect 30196 2524 30248 2576
rect 28724 2499 28776 2508
rect 28724 2465 28733 2499
rect 28733 2465 28767 2499
rect 28767 2465 28776 2499
rect 28724 2456 28776 2465
rect 28080 2388 28132 2440
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 28448 2388 28500 2397
rect 28540 2388 28592 2440
rect 29460 2388 29512 2440
rect 31300 2524 31352 2576
rect 10324 2363 10376 2372
rect 10324 2329 10333 2363
rect 10333 2329 10367 2363
rect 10367 2329 10376 2363
rect 10324 2320 10376 2329
rect 14188 2320 14240 2372
rect 14280 2320 14332 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 15844 2320 15896 2372
rect 16948 2363 17000 2372
rect 16948 2329 16957 2363
rect 16957 2329 16991 2363
rect 16991 2329 17000 2363
rect 16948 2320 17000 2329
rect 17684 2320 17736 2372
rect 11336 2252 11388 2304
rect 12348 2252 12400 2304
rect 13452 2252 13504 2304
rect 19064 2320 19116 2372
rect 20168 2363 20220 2372
rect 20168 2329 20177 2363
rect 20177 2329 20211 2363
rect 20211 2329 20220 2363
rect 20168 2320 20220 2329
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 21640 2295 21692 2304
rect 21640 2261 21649 2295
rect 21649 2261 21683 2295
rect 21683 2261 21692 2295
rect 21640 2252 21692 2261
rect 22100 2363 22152 2372
rect 22100 2329 22109 2363
rect 22109 2329 22143 2363
rect 22143 2329 22152 2363
rect 22100 2320 22152 2329
rect 24032 2363 24084 2372
rect 24032 2329 24041 2363
rect 24041 2329 24075 2363
rect 24075 2329 24084 2363
rect 24032 2320 24084 2329
rect 24768 2320 24820 2372
rect 27528 2320 27580 2372
rect 30564 2456 30616 2508
rect 31208 2499 31260 2508
rect 31208 2465 31217 2499
rect 31217 2465 31251 2499
rect 31251 2465 31260 2499
rect 31208 2456 31260 2465
rect 30288 2388 30340 2440
rect 30656 2388 30708 2440
rect 30012 2320 30064 2372
rect 31392 2320 31444 2372
rect 32864 2456 32916 2508
rect 32956 2388 33008 2440
rect 33140 2388 33192 2440
rect 33784 2388 33836 2440
rect 34152 2592 34204 2644
rect 34336 2499 34388 2508
rect 34336 2465 34345 2499
rect 34345 2465 34379 2499
rect 34379 2465 34388 2499
rect 34336 2456 34388 2465
rect 35900 2592 35952 2644
rect 37280 2592 37332 2644
rect 37648 2635 37700 2644
rect 37648 2601 37657 2635
rect 37657 2601 37691 2635
rect 37691 2601 37700 2635
rect 37648 2592 37700 2601
rect 38936 2592 38988 2644
rect 35808 2456 35860 2508
rect 36912 2456 36964 2508
rect 38108 2456 38160 2508
rect 38292 2499 38344 2508
rect 38292 2465 38301 2499
rect 38301 2465 38335 2499
rect 38335 2465 38344 2499
rect 38292 2456 38344 2465
rect 31944 2320 31996 2372
rect 25412 2252 25464 2304
rect 27436 2252 27488 2304
rect 29092 2252 29144 2304
rect 29184 2252 29236 2304
rect 31484 2252 31536 2304
rect 33232 2252 33284 2304
rect 33508 2295 33560 2304
rect 33508 2261 33517 2295
rect 33517 2261 33551 2295
rect 33551 2261 33560 2295
rect 33508 2252 33560 2261
rect 35256 2252 35308 2304
rect 35716 2252 35768 2304
rect 36452 2320 36504 2372
rect 37464 2320 37516 2372
rect 37648 2320 37700 2372
rect 38384 2388 38436 2440
rect 40408 2592 40460 2644
rect 41880 2592 41932 2644
rect 42432 2592 42484 2644
rect 43352 2635 43404 2644
rect 43352 2601 43361 2635
rect 43361 2601 43395 2635
rect 43395 2601 43404 2635
rect 43352 2592 43404 2601
rect 39580 2524 39632 2576
rect 39764 2499 39816 2508
rect 39764 2465 39773 2499
rect 39773 2465 39807 2499
rect 39807 2465 39816 2499
rect 39764 2456 39816 2465
rect 40316 2456 40368 2508
rect 42248 2524 42300 2576
rect 40868 2456 40920 2508
rect 44180 2635 44232 2644
rect 44180 2601 44189 2635
rect 44189 2601 44223 2635
rect 44223 2601 44232 2635
rect 44180 2592 44232 2601
rect 44732 2592 44784 2644
rect 43812 2456 43864 2508
rect 39396 2388 39448 2440
rect 39764 2320 39816 2372
rect 40132 2320 40184 2372
rect 35900 2252 35952 2304
rect 37832 2252 37884 2304
rect 40316 2252 40368 2304
rect 40868 2295 40920 2304
rect 40868 2261 40877 2295
rect 40877 2261 40911 2295
rect 40911 2261 40920 2295
rect 40868 2252 40920 2261
rect 40960 2252 41012 2304
rect 6070 2150 6122 2202
rect 6134 2150 6186 2202
rect 6198 2150 6250 2202
rect 6262 2150 6314 2202
rect 6326 2150 6378 2202
rect 11070 2150 11122 2202
rect 11134 2150 11186 2202
rect 11198 2150 11250 2202
rect 11262 2150 11314 2202
rect 11326 2150 11378 2202
rect 16070 2150 16122 2202
rect 16134 2150 16186 2202
rect 16198 2150 16250 2202
rect 16262 2150 16314 2202
rect 16326 2150 16378 2202
rect 21070 2150 21122 2202
rect 21134 2150 21186 2202
rect 21198 2150 21250 2202
rect 21262 2150 21314 2202
rect 21326 2150 21378 2202
rect 26070 2150 26122 2202
rect 26134 2150 26186 2202
rect 26198 2150 26250 2202
rect 26262 2150 26314 2202
rect 26326 2150 26378 2202
rect 31070 2150 31122 2202
rect 31134 2150 31186 2202
rect 31198 2150 31250 2202
rect 31262 2150 31314 2202
rect 31326 2150 31378 2202
rect 36070 2150 36122 2202
rect 36134 2150 36186 2202
rect 36198 2150 36250 2202
rect 36262 2150 36314 2202
rect 36326 2150 36378 2202
rect 41070 2150 41122 2202
rect 41134 2150 41186 2202
rect 41198 2150 41250 2202
rect 41262 2150 41314 2202
rect 41326 2150 41378 2202
rect 1676 2091 1728 2100
rect 1676 2057 1685 2091
rect 1685 2057 1719 2091
rect 1719 2057 1728 2091
rect 1676 2048 1728 2057
rect 2228 2048 2280 2100
rect 2964 2048 3016 2100
rect 3424 2048 3476 2100
rect 4068 2048 4120 2100
rect 4712 2048 4764 2100
rect 9864 2048 9916 2100
rect 10048 2048 10100 2100
rect 10324 2048 10376 2100
rect 11796 2048 11848 2100
rect 11888 2091 11940 2100
rect 11888 2057 11897 2091
rect 11897 2057 11931 2091
rect 11931 2057 11940 2091
rect 11888 2048 11940 2057
rect 12440 2048 12492 2100
rect 2320 1955 2372 1964
rect 2320 1921 2329 1955
rect 2329 1921 2363 1955
rect 2363 1921 2372 1955
rect 2320 1912 2372 1921
rect 3516 1955 3568 1964
rect 3516 1921 3525 1955
rect 3525 1921 3559 1955
rect 3559 1921 3568 1955
rect 3516 1912 3568 1921
rect 4712 1955 4764 1964
rect 4712 1921 4721 1955
rect 4721 1921 4755 1955
rect 4755 1921 4764 1955
rect 4712 1912 4764 1921
rect 5356 1955 5408 1964
rect 5356 1921 5365 1955
rect 5365 1921 5399 1955
rect 5399 1921 5408 1955
rect 5356 1912 5408 1921
rect 6736 1912 6788 1964
rect 8300 1912 8352 1964
rect 10416 1912 10468 1964
rect 10508 1955 10560 1964
rect 10508 1921 10517 1955
rect 10517 1921 10551 1955
rect 10551 1921 10560 1955
rect 10508 1912 10560 1921
rect 11428 1980 11480 2032
rect 3148 1844 3200 1896
rect 6000 1844 6052 1896
rect 8576 1844 8628 1896
rect 9220 1844 9272 1896
rect 8116 1776 8168 1828
rect 9956 1776 10008 1828
rect 14280 2091 14332 2100
rect 14280 2057 14289 2091
rect 14289 2057 14323 2091
rect 14323 2057 14332 2091
rect 14280 2048 14332 2057
rect 15936 2048 15988 2100
rect 16948 2048 17000 2100
rect 18604 2048 18656 2100
rect 19156 2048 19208 2100
rect 19248 2091 19300 2100
rect 19248 2057 19257 2091
rect 19257 2057 19291 2091
rect 19291 2057 19300 2091
rect 19248 2048 19300 2057
rect 19800 2048 19852 2100
rect 20168 2048 20220 2100
rect 12164 1955 12216 1964
rect 12164 1921 12173 1955
rect 12173 1921 12207 1955
rect 12207 1921 12216 1955
rect 12164 1912 12216 1921
rect 12348 1912 12400 1964
rect 12440 1955 12492 1964
rect 12440 1921 12449 1955
rect 12449 1921 12483 1955
rect 12483 1921 12492 1955
rect 12440 1912 12492 1921
rect 14096 1980 14148 2032
rect 14556 1955 14608 1964
rect 14556 1921 14565 1955
rect 14565 1921 14599 1955
rect 14599 1921 14608 1955
rect 14556 1912 14608 1921
rect 17040 1980 17092 2032
rect 17684 1980 17736 2032
rect 16580 1912 16632 1964
rect 16672 1912 16724 1964
rect 14924 1844 14976 1896
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 21640 2091 21692 2100
rect 21640 2057 21649 2091
rect 21649 2057 21683 2091
rect 21683 2057 21692 2091
rect 21640 2048 21692 2057
rect 22100 2048 22152 2100
rect 19892 1955 19944 1964
rect 19892 1921 19901 1955
rect 19901 1921 19935 1955
rect 19935 1921 19944 1955
rect 19892 1912 19944 1921
rect 20996 1955 21048 1964
rect 20996 1921 21005 1955
rect 21005 1921 21039 1955
rect 21039 1921 21048 1955
rect 20996 1912 21048 1921
rect 21548 1955 21600 1964
rect 21548 1921 21557 1955
rect 21557 1921 21591 1955
rect 21591 1921 21600 1955
rect 21548 1912 21600 1921
rect 22560 1912 22612 1964
rect 23756 2048 23808 2100
rect 24032 2048 24084 2100
rect 23020 2023 23072 2032
rect 23020 1989 23029 2023
rect 23029 1989 23063 2023
rect 23063 1989 23072 2023
rect 23020 1980 23072 1989
rect 24768 1980 24820 2032
rect 21916 1844 21968 1896
rect 24492 1912 24544 1964
rect 27620 2048 27672 2100
rect 28080 2048 28132 2100
rect 25688 1980 25740 2032
rect 25412 1955 25464 1964
rect 25412 1921 25421 1955
rect 25421 1921 25455 1955
rect 25455 1921 25464 1955
rect 25412 1912 25464 1921
rect 25596 1955 25648 1964
rect 25596 1921 25605 1955
rect 25605 1921 25639 1955
rect 25639 1921 25648 1955
rect 25596 1912 25648 1921
rect 26884 1980 26936 2032
rect 30012 2048 30064 2100
rect 30932 2048 30984 2100
rect 31852 2048 31904 2100
rect 33508 2048 33560 2100
rect 23664 1844 23716 1896
rect 1216 1751 1268 1760
rect 1216 1717 1225 1751
rect 1225 1717 1259 1751
rect 1259 1717 1268 1751
rect 1216 1708 1268 1717
rect 2136 1751 2188 1760
rect 2136 1717 2145 1751
rect 2145 1717 2179 1751
rect 2179 1717 2188 1751
rect 2136 1708 2188 1717
rect 2964 1708 3016 1760
rect 3976 1708 4028 1760
rect 4528 1751 4580 1760
rect 4528 1717 4537 1751
rect 4537 1717 4571 1751
rect 4571 1717 4580 1751
rect 4528 1708 4580 1717
rect 5172 1751 5224 1760
rect 5172 1717 5181 1751
rect 5181 1717 5215 1751
rect 5215 1717 5224 1751
rect 5172 1708 5224 1717
rect 6184 1751 6236 1760
rect 6184 1717 6193 1751
rect 6193 1717 6227 1751
rect 6227 1717 6236 1751
rect 6184 1708 6236 1717
rect 7748 1751 7800 1760
rect 7748 1717 7757 1751
rect 7757 1717 7791 1751
rect 7791 1717 7800 1751
rect 7748 1708 7800 1717
rect 8944 1751 8996 1760
rect 8944 1717 8953 1751
rect 8953 1717 8987 1751
rect 8987 1717 8996 1751
rect 8944 1708 8996 1717
rect 9680 1751 9732 1760
rect 9680 1717 9689 1751
rect 9689 1717 9723 1751
rect 9723 1717 9732 1751
rect 9680 1708 9732 1717
rect 10324 1751 10376 1760
rect 10324 1717 10333 1751
rect 10333 1717 10367 1751
rect 10367 1717 10376 1751
rect 10324 1708 10376 1717
rect 11152 1751 11204 1760
rect 11152 1717 11161 1751
rect 11161 1717 11195 1751
rect 11195 1717 11204 1751
rect 11152 1708 11204 1717
rect 11980 1751 12032 1760
rect 11980 1717 11989 1751
rect 11989 1717 12023 1751
rect 12023 1717 12032 1751
rect 11980 1708 12032 1717
rect 12256 1751 12308 1760
rect 12256 1717 12265 1751
rect 12265 1717 12299 1751
rect 12299 1717 12308 1751
rect 12256 1708 12308 1717
rect 14372 1751 14424 1760
rect 14372 1717 14381 1751
rect 14381 1717 14415 1751
rect 14415 1717 14424 1751
rect 14372 1708 14424 1717
rect 15384 1751 15436 1760
rect 15384 1717 15393 1751
rect 15393 1717 15427 1751
rect 15427 1717 15436 1751
rect 15384 1708 15436 1717
rect 16212 1751 16264 1760
rect 16212 1717 16221 1751
rect 16221 1717 16255 1751
rect 16255 1717 16264 1751
rect 16212 1708 16264 1717
rect 17592 1751 17644 1760
rect 17592 1717 17601 1751
rect 17601 1717 17635 1751
rect 17635 1717 17644 1751
rect 17592 1708 17644 1717
rect 18328 1751 18380 1760
rect 18328 1717 18337 1751
rect 18337 1717 18371 1751
rect 18371 1717 18380 1751
rect 18328 1708 18380 1717
rect 18420 1708 18472 1760
rect 19708 1751 19760 1760
rect 19708 1717 19717 1751
rect 19717 1717 19751 1751
rect 19751 1717 19760 1751
rect 19708 1708 19760 1717
rect 20168 1751 20220 1760
rect 20168 1717 20177 1751
rect 20177 1717 20211 1751
rect 20211 1717 20220 1751
rect 20168 1708 20220 1717
rect 20812 1751 20864 1760
rect 20812 1717 20821 1751
rect 20821 1717 20855 1751
rect 20855 1717 20864 1751
rect 20812 1708 20864 1717
rect 24308 1776 24360 1828
rect 24400 1776 24452 1828
rect 25136 1776 25188 1828
rect 22192 1751 22244 1760
rect 22192 1717 22201 1751
rect 22201 1717 22235 1751
rect 22235 1717 22244 1751
rect 22192 1708 22244 1717
rect 22376 1708 22428 1760
rect 27988 1912 28040 1964
rect 27896 1844 27948 1896
rect 29552 1912 29604 1964
rect 29736 1912 29788 1964
rect 32312 1980 32364 2032
rect 26240 1708 26292 1760
rect 28080 1751 28132 1760
rect 28080 1717 28089 1751
rect 28089 1717 28123 1751
rect 28123 1717 28132 1751
rect 28080 1708 28132 1717
rect 28172 1708 28224 1760
rect 28540 1844 28592 1896
rect 29920 1844 29972 1896
rect 31852 1912 31904 1964
rect 31944 1955 31996 1964
rect 31944 1921 31953 1955
rect 31953 1921 31987 1955
rect 31987 1921 31996 1955
rect 31944 1912 31996 1921
rect 30564 1776 30616 1828
rect 30012 1708 30064 1760
rect 30472 1751 30524 1760
rect 30472 1717 30481 1751
rect 30481 1717 30515 1751
rect 30515 1717 30524 1751
rect 30472 1708 30524 1717
rect 31576 1776 31628 1828
rect 30840 1708 30892 1760
rect 32220 1887 32272 1896
rect 32220 1853 32229 1887
rect 32229 1853 32263 1887
rect 32263 1853 32272 1887
rect 32220 1844 32272 1853
rect 32956 1844 33008 1896
rect 34152 2023 34204 2032
rect 34152 1989 34161 2023
rect 34161 1989 34195 2023
rect 34195 1989 34204 2023
rect 34152 1980 34204 1989
rect 35532 2048 35584 2100
rect 35900 2048 35952 2100
rect 37464 1980 37516 2032
rect 39028 2048 39080 2100
rect 39488 2048 39540 2100
rect 40040 2048 40092 2100
rect 40500 2048 40552 2100
rect 40684 2091 40736 2100
rect 40684 2057 40693 2091
rect 40693 2057 40727 2091
rect 40727 2057 40736 2091
rect 40684 2048 40736 2057
rect 42248 2048 42300 2100
rect 42984 2048 43036 2100
rect 43812 2091 43864 2100
rect 43812 2057 43821 2091
rect 43821 2057 43855 2091
rect 43855 2057 43864 2091
rect 43812 2048 43864 2057
rect 44548 2091 44600 2100
rect 44548 2057 44557 2091
rect 44557 2057 44591 2091
rect 44591 2057 44600 2091
rect 44548 2048 44600 2057
rect 44732 2048 44784 2100
rect 33784 1912 33836 1964
rect 36452 1912 36504 1964
rect 38200 1912 38252 1964
rect 34244 1844 34296 1896
rect 34888 1844 34940 1896
rect 35624 1887 35676 1896
rect 35624 1853 35633 1887
rect 35633 1853 35667 1887
rect 35667 1853 35676 1887
rect 35624 1844 35676 1853
rect 36544 1844 36596 1896
rect 40408 1980 40460 2032
rect 40592 1912 40644 1964
rect 41512 2023 41564 2032
rect 41512 1989 41521 2023
rect 41521 1989 41555 2023
rect 41555 1989 41564 2023
rect 41512 1980 41564 1989
rect 42432 2023 42484 2032
rect 42432 1989 42441 2023
rect 42441 1989 42475 2023
rect 42475 1989 42484 2023
rect 42432 1980 42484 1989
rect 38108 1776 38160 1828
rect 33324 1708 33376 1760
rect 38844 1708 38896 1760
rect 40224 1708 40276 1760
rect 3570 1606 3622 1658
rect 3634 1606 3686 1658
rect 3698 1606 3750 1658
rect 3762 1606 3814 1658
rect 3826 1606 3878 1658
rect 8570 1606 8622 1658
rect 8634 1606 8686 1658
rect 8698 1606 8750 1658
rect 8762 1606 8814 1658
rect 8826 1606 8878 1658
rect 13570 1606 13622 1658
rect 13634 1606 13686 1658
rect 13698 1606 13750 1658
rect 13762 1606 13814 1658
rect 13826 1606 13878 1658
rect 18570 1606 18622 1658
rect 18634 1606 18686 1658
rect 18698 1606 18750 1658
rect 18762 1606 18814 1658
rect 18826 1606 18878 1658
rect 23570 1606 23622 1658
rect 23634 1606 23686 1658
rect 23698 1606 23750 1658
rect 23762 1606 23814 1658
rect 23826 1606 23878 1658
rect 28570 1606 28622 1658
rect 28634 1606 28686 1658
rect 28698 1606 28750 1658
rect 28762 1606 28814 1658
rect 28826 1606 28878 1658
rect 33570 1606 33622 1658
rect 33634 1606 33686 1658
rect 33698 1606 33750 1658
rect 33762 1606 33814 1658
rect 33826 1606 33878 1658
rect 38570 1606 38622 1658
rect 38634 1606 38686 1658
rect 38698 1606 38750 1658
rect 38762 1606 38814 1658
rect 38826 1606 38878 1658
rect 43570 1606 43622 1658
rect 43634 1606 43686 1658
rect 43698 1606 43750 1658
rect 43762 1606 43814 1658
rect 43826 1606 43878 1658
rect 2872 1504 2924 1556
rect 6000 1547 6052 1556
rect 6000 1513 6009 1547
rect 6009 1513 6043 1547
rect 6043 1513 6052 1547
rect 6000 1504 6052 1513
rect 6920 1547 6972 1556
rect 6920 1513 6929 1547
rect 6929 1513 6963 1547
rect 6963 1513 6972 1547
rect 6920 1504 6972 1513
rect 8116 1504 8168 1556
rect 9220 1547 9272 1556
rect 9220 1513 9229 1547
rect 9229 1513 9263 1547
rect 9263 1513 9272 1547
rect 9220 1504 9272 1513
rect 10048 1504 10100 1556
rect 11060 1547 11112 1556
rect 11060 1513 11069 1547
rect 11069 1513 11103 1547
rect 11103 1513 11112 1547
rect 11060 1504 11112 1513
rect 15200 1547 15252 1556
rect 15200 1513 15209 1547
rect 15209 1513 15243 1547
rect 15243 1513 15252 1547
rect 15200 1504 15252 1513
rect 16672 1547 16724 1556
rect 16672 1513 16681 1547
rect 16681 1513 16715 1547
rect 16715 1513 16724 1547
rect 16672 1504 16724 1513
rect 17684 1547 17736 1556
rect 17684 1513 17693 1547
rect 17693 1513 17727 1547
rect 17727 1513 17736 1547
rect 17684 1504 17736 1513
rect 19340 1547 19392 1556
rect 19340 1513 19349 1547
rect 19349 1513 19383 1547
rect 19383 1513 19392 1547
rect 19340 1504 19392 1513
rect 24216 1504 24268 1556
rect 25596 1504 25648 1556
rect 1216 1436 1268 1488
rect 3148 1436 3200 1488
rect 12348 1436 12400 1488
rect 15844 1479 15896 1488
rect 15844 1445 15853 1479
rect 15853 1445 15887 1479
rect 15887 1445 15896 1479
rect 15844 1436 15896 1445
rect 1308 1300 1360 1352
rect 2136 1300 2188 1352
rect 2964 1300 3016 1352
rect 3976 1300 4028 1352
rect 4528 1300 4580 1352
rect 5172 1300 5224 1352
rect 6184 1300 6236 1352
rect 7012 1300 7064 1352
rect 7748 1343 7800 1352
rect 7748 1309 7757 1343
rect 7757 1309 7791 1343
rect 7791 1309 7800 1343
rect 7748 1300 7800 1309
rect 8944 1300 8996 1352
rect 9680 1300 9732 1352
rect 10324 1300 10376 1352
rect 11152 1300 11204 1352
rect 11980 1300 12032 1352
rect 12256 1300 12308 1352
rect 13452 1300 13504 1352
rect 14372 1343 14424 1352
rect 14372 1309 14381 1343
rect 14381 1309 14415 1343
rect 14415 1309 14424 1343
rect 14372 1300 14424 1309
rect 15384 1300 15436 1352
rect 16212 1300 16264 1352
rect 18328 1300 18380 1352
rect 18420 1300 18472 1352
rect 19708 1300 19760 1352
rect 20168 1343 20220 1352
rect 20168 1309 20177 1343
rect 20177 1309 20211 1343
rect 20211 1309 20220 1343
rect 20168 1300 20220 1309
rect 20812 1300 20864 1352
rect 2228 1232 2280 1284
rect 5724 1232 5776 1284
rect 14096 1232 14148 1284
rect 1308 1207 1360 1216
rect 1308 1173 1317 1207
rect 1317 1173 1351 1207
rect 1351 1173 1360 1207
rect 1308 1164 1360 1173
rect 1860 1164 1912 1216
rect 3516 1164 3568 1216
rect 4620 1207 4672 1216
rect 4620 1173 4629 1207
rect 4629 1173 4663 1207
rect 4663 1173 4672 1207
rect 4620 1164 4672 1173
rect 5448 1207 5500 1216
rect 5448 1173 5457 1207
rect 5457 1173 5491 1207
rect 5491 1173 5500 1207
rect 5448 1164 5500 1173
rect 6000 1164 6052 1216
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9588 1207 9640 1216
rect 9588 1173 9597 1207
rect 9597 1173 9631 1207
rect 9631 1173 9640 1207
rect 9588 1164 9640 1173
rect 10416 1207 10468 1216
rect 10416 1173 10425 1207
rect 10425 1173 10459 1207
rect 10459 1173 10468 1207
rect 10416 1164 10468 1173
rect 12072 1207 12124 1216
rect 12072 1173 12081 1207
rect 12081 1173 12115 1207
rect 12115 1173 12124 1207
rect 12072 1164 12124 1173
rect 12900 1207 12952 1216
rect 12900 1173 12909 1207
rect 12909 1173 12943 1207
rect 12943 1173 12952 1207
rect 12900 1164 12952 1173
rect 13728 1207 13780 1216
rect 13728 1173 13737 1207
rect 13737 1173 13771 1207
rect 13771 1173 13780 1207
rect 13728 1164 13780 1173
rect 14188 1207 14240 1216
rect 14188 1173 14197 1207
rect 14197 1173 14231 1207
rect 14231 1173 14240 1207
rect 14188 1164 14240 1173
rect 14280 1164 14332 1216
rect 15936 1164 15988 1216
rect 17040 1207 17092 1216
rect 17040 1173 17049 1207
rect 17049 1173 17083 1207
rect 17083 1173 17092 1207
rect 17040 1164 17092 1173
rect 19524 1232 19576 1284
rect 21732 1343 21784 1352
rect 21732 1309 21741 1343
rect 21741 1309 21775 1343
rect 21775 1309 21784 1343
rect 21732 1300 21784 1309
rect 22192 1300 22244 1352
rect 22560 1343 22612 1352
rect 22560 1309 22569 1343
rect 22569 1309 22603 1343
rect 22603 1309 22612 1343
rect 22560 1300 22612 1309
rect 25504 1436 25556 1488
rect 23020 1300 23072 1352
rect 25136 1368 25188 1420
rect 26148 1368 26200 1420
rect 27620 1504 27672 1556
rect 29092 1504 29144 1556
rect 29276 1504 29328 1556
rect 29644 1547 29696 1556
rect 29644 1513 29653 1547
rect 29653 1513 29687 1547
rect 29687 1513 29696 1547
rect 29644 1504 29696 1513
rect 29920 1547 29972 1556
rect 29920 1513 29929 1547
rect 29929 1513 29963 1547
rect 29963 1513 29972 1547
rect 29920 1504 29972 1513
rect 30012 1504 30064 1556
rect 28264 1436 28316 1488
rect 28356 1368 28408 1420
rect 18420 1164 18472 1216
rect 20076 1207 20128 1216
rect 20076 1173 20085 1207
rect 20085 1173 20119 1207
rect 20119 1173 20128 1207
rect 20076 1164 20128 1173
rect 20352 1207 20404 1216
rect 20352 1173 20361 1207
rect 20361 1173 20395 1207
rect 20395 1173 20404 1207
rect 20352 1164 20404 1173
rect 20996 1164 21048 1216
rect 21732 1164 21784 1216
rect 24124 1300 24176 1352
rect 26240 1300 26292 1352
rect 27160 1300 27212 1352
rect 28080 1300 28132 1352
rect 22560 1164 22612 1216
rect 23296 1207 23348 1216
rect 23296 1173 23305 1207
rect 23305 1173 23339 1207
rect 23339 1173 23348 1207
rect 23296 1164 23348 1173
rect 24492 1232 24544 1284
rect 24768 1232 24820 1284
rect 28448 1300 28500 1352
rect 29276 1368 29328 1420
rect 27068 1164 27120 1216
rect 31668 1504 31720 1556
rect 32036 1479 32088 1488
rect 32036 1445 32045 1479
rect 32045 1445 32079 1479
rect 32079 1445 32088 1479
rect 32036 1436 32088 1445
rect 32220 1504 32272 1556
rect 34980 1504 35032 1556
rect 38200 1504 38252 1556
rect 38936 1504 38988 1556
rect 40224 1504 40276 1556
rect 40960 1504 41012 1556
rect 42984 1547 43036 1556
rect 42984 1513 42993 1547
rect 42993 1513 43027 1547
rect 43027 1513 43036 1547
rect 42984 1504 43036 1513
rect 43904 1547 43956 1556
rect 43904 1513 43913 1547
rect 43913 1513 43947 1547
rect 43947 1513 43956 1547
rect 43904 1504 43956 1513
rect 33324 1436 33376 1488
rect 35256 1436 35308 1488
rect 32312 1368 32364 1420
rect 29276 1232 29328 1284
rect 29736 1232 29788 1284
rect 30288 1275 30340 1284
rect 30288 1241 30297 1275
rect 30297 1241 30331 1275
rect 30331 1241 30340 1275
rect 30288 1232 30340 1241
rect 31392 1300 31444 1352
rect 31484 1300 31536 1352
rect 32036 1300 32088 1352
rect 32496 1343 32548 1352
rect 32496 1309 32505 1343
rect 32505 1309 32539 1343
rect 32539 1309 32548 1343
rect 32496 1300 32548 1309
rect 29092 1164 29144 1216
rect 30380 1164 30432 1216
rect 32128 1164 32180 1216
rect 32404 1275 32456 1284
rect 32404 1241 32413 1275
rect 32413 1241 32447 1275
rect 32447 1241 32456 1275
rect 32404 1232 32456 1241
rect 32864 1275 32916 1284
rect 32864 1241 32889 1275
rect 32889 1241 32916 1275
rect 32864 1232 32916 1241
rect 33968 1368 34020 1420
rect 35624 1368 35676 1420
rect 33048 1300 33100 1352
rect 33232 1300 33284 1352
rect 33876 1343 33928 1352
rect 33876 1309 33885 1343
rect 33885 1309 33919 1343
rect 33919 1309 33928 1343
rect 33876 1300 33928 1309
rect 34244 1343 34296 1352
rect 34244 1309 34253 1343
rect 34253 1309 34287 1343
rect 34287 1309 34296 1343
rect 34244 1300 34296 1309
rect 34704 1300 34756 1352
rect 35164 1343 35216 1352
rect 35164 1309 35173 1343
rect 35173 1309 35207 1343
rect 35207 1309 35216 1343
rect 35164 1300 35216 1309
rect 35716 1300 35768 1352
rect 33048 1164 33100 1216
rect 33416 1164 33468 1216
rect 34336 1207 34388 1216
rect 34336 1173 34345 1207
rect 34345 1173 34379 1207
rect 34379 1173 34388 1207
rect 34336 1164 34388 1173
rect 35624 1207 35676 1216
rect 35624 1173 35633 1207
rect 35633 1173 35667 1207
rect 35667 1173 35676 1207
rect 35624 1164 35676 1173
rect 36452 1436 36504 1488
rect 36084 1343 36136 1352
rect 36084 1309 36093 1343
rect 36093 1309 36127 1343
rect 36127 1309 36136 1343
rect 36084 1300 36136 1309
rect 36176 1300 36228 1352
rect 36360 1343 36412 1352
rect 36360 1309 36369 1343
rect 36369 1309 36403 1343
rect 36403 1309 36412 1343
rect 36360 1300 36412 1309
rect 36820 1343 36872 1352
rect 36820 1309 36829 1343
rect 36829 1309 36863 1343
rect 36863 1309 36872 1343
rect 36820 1300 36872 1309
rect 37096 1343 37148 1352
rect 37096 1309 37105 1343
rect 37105 1309 37139 1343
rect 37139 1309 37148 1343
rect 37096 1300 37148 1309
rect 39488 1300 39540 1352
rect 39580 1343 39632 1352
rect 39580 1309 39589 1343
rect 39589 1309 39623 1343
rect 39623 1309 39632 1343
rect 39580 1300 39632 1309
rect 39672 1343 39724 1352
rect 39672 1309 39681 1343
rect 39681 1309 39715 1343
rect 39715 1309 39724 1343
rect 39672 1300 39724 1309
rect 39764 1300 39816 1352
rect 35992 1164 36044 1216
rect 37832 1232 37884 1284
rect 40316 1300 40368 1352
rect 40776 1343 40828 1352
rect 40776 1309 40785 1343
rect 40785 1309 40819 1343
rect 40819 1309 40828 1343
rect 40776 1300 40828 1309
rect 40868 1300 40920 1352
rect 41328 1343 41380 1352
rect 41328 1309 41337 1343
rect 41337 1309 41371 1343
rect 41371 1309 41380 1343
rect 41328 1300 41380 1309
rect 39948 1232 40000 1284
rect 41972 1343 42024 1352
rect 41972 1309 41981 1343
rect 41981 1309 42015 1343
rect 42015 1309 42024 1343
rect 41972 1300 42024 1309
rect 41696 1232 41748 1284
rect 42708 1343 42760 1352
rect 42708 1309 42717 1343
rect 42717 1309 42751 1343
rect 42751 1309 42760 1343
rect 42708 1300 42760 1309
rect 43260 1300 43312 1352
rect 43536 1343 43588 1352
rect 43536 1309 43545 1343
rect 43545 1309 43579 1343
rect 43579 1309 43588 1343
rect 43536 1300 43588 1309
rect 44364 1300 44416 1352
rect 44548 1343 44600 1352
rect 44548 1309 44557 1343
rect 44557 1309 44591 1343
rect 44591 1309 44600 1343
rect 44548 1300 44600 1309
rect 44824 1343 44876 1352
rect 44824 1309 44833 1343
rect 44833 1309 44867 1343
rect 44867 1309 44876 1343
rect 44824 1300 44876 1309
rect 45008 1300 45060 1352
rect 45192 1343 45244 1352
rect 45192 1309 45201 1343
rect 45201 1309 45235 1343
rect 45235 1309 45244 1343
rect 45192 1300 45244 1309
rect 39028 1207 39080 1216
rect 39028 1173 39037 1207
rect 39037 1173 39071 1207
rect 39071 1173 39080 1207
rect 39028 1164 39080 1173
rect 40408 1164 40460 1216
rect 40684 1164 40736 1216
rect 41420 1207 41472 1216
rect 41420 1173 41429 1207
rect 41429 1173 41463 1207
rect 41463 1173 41472 1207
rect 41420 1164 41472 1173
rect 41788 1207 41840 1216
rect 41788 1173 41797 1207
rect 41797 1173 41831 1207
rect 41831 1173 41840 1207
rect 41788 1164 41840 1173
rect 42064 1207 42116 1216
rect 42064 1173 42073 1207
rect 42073 1173 42107 1207
rect 42107 1173 42116 1207
rect 42064 1164 42116 1173
rect 42524 1207 42576 1216
rect 42524 1173 42533 1207
rect 42533 1173 42567 1207
rect 42567 1173 42576 1207
rect 42524 1164 42576 1173
rect 6070 1062 6122 1114
rect 6134 1062 6186 1114
rect 6198 1062 6250 1114
rect 6262 1062 6314 1114
rect 6326 1062 6378 1114
rect 11070 1062 11122 1114
rect 11134 1062 11186 1114
rect 11198 1062 11250 1114
rect 11262 1062 11314 1114
rect 11326 1062 11378 1114
rect 16070 1062 16122 1114
rect 16134 1062 16186 1114
rect 16198 1062 16250 1114
rect 16262 1062 16314 1114
rect 16326 1062 16378 1114
rect 21070 1062 21122 1114
rect 21134 1062 21186 1114
rect 21198 1062 21250 1114
rect 21262 1062 21314 1114
rect 21326 1062 21378 1114
rect 26070 1062 26122 1114
rect 26134 1062 26186 1114
rect 26198 1062 26250 1114
rect 26262 1062 26314 1114
rect 26326 1062 26378 1114
rect 31070 1062 31122 1114
rect 31134 1062 31186 1114
rect 31198 1062 31250 1114
rect 31262 1062 31314 1114
rect 31326 1062 31378 1114
rect 36070 1062 36122 1114
rect 36134 1062 36186 1114
rect 36198 1062 36250 1114
rect 36262 1062 36314 1114
rect 36326 1062 36378 1114
rect 41070 1062 41122 1114
rect 41134 1062 41186 1114
rect 41198 1062 41250 1114
rect 41262 1062 41314 1114
rect 41326 1062 41378 1114
rect 14096 960 14148 1012
rect 14188 960 14240 1012
rect 20076 960 20128 1012
rect 24584 960 24636 1012
rect 30288 960 30340 1012
rect 32864 960 32916 1012
rect 35624 960 35676 1012
rect 38292 960 38344 1012
rect 40868 960 40920 1012
rect 25228 892 25280 944
rect 34336 892 34388 944
rect 39028 892 39080 944
rect 40132 892 40184 944
rect 21548 824 21600 876
rect 27252 824 27304 876
rect 31484 824 31536 876
rect 38476 824 38528 876
rect 42524 824 42576 876
rect 32680 756 32732 808
rect 36452 756 36504 808
rect 39396 756 39448 808
rect 40960 756 41012 808
rect 34428 688 34480 740
rect 37096 688 37148 740
rect 37832 688 37884 740
rect 40776 688 40828 740
rect 28908 620 28960 672
rect 30380 620 30432 672
rect 33508 620 33560 672
rect 36820 620 36872 672
rect 40960 620 41012 672
rect 41972 620 42024 672
<< metal2 >>
rect 846 23840 902 24300
rect 1766 23840 1822 24300
rect 2686 23840 2742 24300
rect 3606 23840 3662 24300
rect 4526 23840 4582 24300
rect 5446 23840 5502 24300
rect 6366 23840 6422 24300
rect 7286 23840 7342 24300
rect 8206 23840 8262 24300
rect 9126 23840 9182 24300
rect 10046 23840 10102 24300
rect 10966 23840 11022 24300
rect 11886 23840 11942 24300
rect 12806 23840 12862 24300
rect 13726 23840 13782 24300
rect 14646 23840 14702 24300
rect 15566 23840 15622 24300
rect 16486 23840 16542 24300
rect 17406 23840 17462 24300
rect 18326 23840 18382 24300
rect 19246 23840 19302 24300
rect 20166 23840 20222 24300
rect 21086 23840 21142 24300
rect 22006 23840 22062 24300
rect 22926 23840 22982 24300
rect 23846 23840 23902 24300
rect 24766 23840 24822 24300
rect 25686 23840 25742 24300
rect 26606 23840 26662 24300
rect 27526 23840 27582 24300
rect 28446 23840 28502 24300
rect 29366 23840 29422 24300
rect 29472 23854 29776 23882
rect 860 22778 888 23840
rect 1780 22778 1808 23840
rect 848 22772 900 22778
rect 848 22714 900 22720
rect 1768 22772 1820 22778
rect 2700 22760 2728 23840
rect 3620 22778 3648 23840
rect 4540 22778 4568 23840
rect 5460 22778 5488 23840
rect 6380 23066 6408 23840
rect 6000 23044 6052 23050
rect 6380 23038 6500 23066
rect 6000 22986 6052 22992
rect 2780 22772 2832 22778
rect 2700 22732 2780 22760
rect 1768 22714 1820 22720
rect 2780 22714 2832 22720
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 940 22636 992 22642
rect 940 22578 992 22584
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 952 22234 980 22578
rect 1872 22234 1900 22578
rect 940 22228 992 22234
rect 940 22170 992 22176
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 1964 22030 1992 22646
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 3068 22030 3096 22510
rect 3252 22234 3280 22578
rect 3570 22332 3878 22341
rect 3570 22330 3576 22332
rect 3632 22330 3656 22332
rect 3712 22330 3736 22332
rect 3792 22330 3816 22332
rect 3872 22330 3878 22332
rect 3632 22278 3634 22330
rect 3814 22278 3816 22330
rect 3570 22276 3576 22278
rect 3632 22276 3656 22278
rect 3712 22276 3736 22278
rect 3792 22276 3816 22278
rect 3872 22276 3878 22278
rect 3570 22267 3878 22276
rect 3988 22234 4016 22578
rect 4632 22234 4660 22578
rect 5828 22234 5856 22578
rect 6012 22234 6040 22986
rect 6070 22876 6378 22885
rect 6070 22874 6076 22876
rect 6132 22874 6156 22876
rect 6212 22874 6236 22876
rect 6292 22874 6316 22876
rect 6372 22874 6378 22876
rect 6132 22822 6134 22874
rect 6314 22822 6316 22874
rect 6070 22820 6076 22822
rect 6132 22820 6156 22822
rect 6212 22820 6236 22822
rect 6292 22820 6316 22822
rect 6372 22820 6378 22822
rect 6070 22811 6378 22820
rect 6472 22778 6500 23038
rect 7300 22778 7328 23840
rect 8220 22778 8248 23840
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 6460 22772 6512 22778
rect 6460 22714 6512 22720
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8312 22642 8340 22918
rect 9140 22778 9168 23840
rect 10060 22778 10088 23840
rect 10980 22778 11008 23840
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11070 22876 11378 22885
rect 11070 22874 11076 22876
rect 11132 22874 11156 22876
rect 11212 22874 11236 22876
rect 11292 22874 11316 22876
rect 11372 22874 11378 22876
rect 11132 22822 11134 22874
rect 11314 22822 11316 22874
rect 11070 22820 11076 22822
rect 11132 22820 11156 22822
rect 11212 22820 11236 22822
rect 11292 22820 11316 22822
rect 11372 22820 11378 22822
rect 11070 22811 11378 22820
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 11716 22642 11744 23258
rect 11900 22778 11928 23840
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 6472 22234 6500 22578
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 5078 22128 5134 22137
rect 4724 22072 5078 22094
rect 7208 22094 7236 22374
rect 7392 22234 7420 22578
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 4724 22066 5134 22072
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 3056 22024 3108 22030
rect 4436 22024 4488 22030
rect 3056 21966 3108 21972
rect 4434 21992 4436 22001
rect 4488 21992 4490 22001
rect 940 20936 992 20942
rect 940 20878 992 20884
rect 756 20800 808 20806
rect 952 20777 980 20878
rect 756 20742 808 20748
rect 938 20768 994 20777
rect 768 20534 796 20742
rect 938 20703 994 20712
rect 756 20528 808 20534
rect 756 20470 808 20476
rect 940 15020 992 15026
rect 940 14962 992 14968
rect 756 14816 808 14822
rect 952 14793 980 14962
rect 756 14758 808 14764
rect 938 14784 994 14793
rect 768 13802 796 14758
rect 938 14719 994 14728
rect 756 13796 808 13802
rect 756 13738 808 13744
rect 940 8832 992 8838
rect 938 8800 940 8809
rect 992 8800 994 8809
rect 938 8735 994 8744
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 940 4480 992 4486
rect 940 4422 992 4428
rect 952 4010 980 4422
rect 940 4004 992 4010
rect 940 3946 992 3952
rect 1320 3194 1348 6258
rect 3068 5914 3096 21966
rect 4434 21927 4490 21936
rect 3570 21244 3878 21253
rect 3570 21242 3576 21244
rect 3632 21242 3656 21244
rect 3712 21242 3736 21244
rect 3792 21242 3816 21244
rect 3872 21242 3878 21244
rect 3632 21190 3634 21242
rect 3814 21190 3816 21242
rect 3570 21188 3576 21190
rect 3632 21188 3656 21190
rect 3712 21188 3736 21190
rect 3792 21188 3816 21190
rect 3872 21188 3878 21190
rect 3570 21179 3878 21188
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3160 20398 3188 20742
rect 3804 20398 3832 20742
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3792 20392 3844 20398
rect 3844 20340 4016 20346
rect 3792 20334 4016 20340
rect 3344 20058 3372 20334
rect 3804 20318 4016 20334
rect 3570 20156 3878 20165
rect 3570 20154 3576 20156
rect 3632 20154 3656 20156
rect 3712 20154 3736 20156
rect 3792 20154 3816 20156
rect 3872 20154 3878 20156
rect 3632 20102 3634 20154
rect 3814 20102 3816 20154
rect 3570 20100 3576 20102
rect 3632 20100 3656 20102
rect 3712 20100 3736 20102
rect 3792 20100 3816 20102
rect 3872 20100 3878 20102
rect 3570 20091 3878 20100
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3988 19922 4016 20318
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3436 17542 3464 19654
rect 3570 19068 3878 19077
rect 3570 19066 3576 19068
rect 3632 19066 3656 19068
rect 3712 19066 3736 19068
rect 3792 19066 3816 19068
rect 3872 19066 3878 19068
rect 3632 19014 3634 19066
rect 3814 19014 3816 19066
rect 3570 19012 3576 19014
rect 3632 19012 3656 19014
rect 3712 19012 3736 19014
rect 3792 19012 3816 19014
rect 3872 19012 3878 19014
rect 3570 19003 3878 19012
rect 3792 18284 3844 18290
rect 3988 18272 4016 19858
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 3844 18244 4016 18272
rect 3792 18226 3844 18232
rect 3570 17980 3878 17989
rect 3570 17978 3576 17980
rect 3632 17978 3656 17980
rect 3712 17978 3736 17980
rect 3792 17978 3816 17980
rect 3872 17978 3878 17980
rect 3632 17926 3634 17978
rect 3814 17926 3816 17978
rect 3570 17924 3576 17926
rect 3632 17924 3656 17926
rect 3712 17924 3736 17926
rect 3792 17924 3816 17926
rect 3872 17924 3878 17926
rect 3570 17915 3878 17924
rect 4448 17882 4476 18770
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3344 16454 3372 17070
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3344 16046 3372 16390
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3344 15348 3372 15982
rect 3436 15910 3464 17478
rect 3988 17354 4016 17478
rect 3988 17326 4108 17354
rect 4080 17134 4108 17326
rect 4172 17134 4200 17546
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3570 16892 3878 16901
rect 3570 16890 3576 16892
rect 3632 16890 3656 16892
rect 3712 16890 3736 16892
rect 3792 16890 3816 16892
rect 3872 16890 3878 16892
rect 3632 16838 3634 16890
rect 3814 16838 3816 16890
rect 3570 16836 3576 16838
rect 3632 16836 3656 16838
rect 3712 16836 3736 16838
rect 3792 16836 3816 16838
rect 3872 16836 3878 16838
rect 3570 16827 3878 16836
rect 4448 16590 4476 17614
rect 4632 17270 4660 18294
rect 4528 17264 4580 17270
rect 4620 17264 4672 17270
rect 4580 17212 4620 17218
rect 4528 17206 4672 17212
rect 4540 17190 4660 17206
rect 4632 16658 4660 17190
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4632 16250 4660 16594
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3570 15804 3878 15813
rect 3570 15802 3576 15804
rect 3632 15802 3656 15804
rect 3712 15802 3736 15804
rect 3792 15802 3816 15804
rect 3872 15802 3878 15804
rect 3632 15750 3634 15802
rect 3814 15750 3816 15802
rect 3570 15748 3576 15750
rect 3632 15748 3656 15750
rect 3712 15748 3736 15750
rect 3792 15748 3816 15750
rect 3872 15748 3878 15750
rect 3570 15739 3878 15748
rect 3424 15360 3476 15366
rect 3344 15320 3424 15348
rect 3424 15302 3476 15308
rect 3436 13870 3464 15302
rect 3570 14716 3878 14725
rect 3570 14714 3576 14716
rect 3632 14714 3656 14716
rect 3712 14714 3736 14716
rect 3792 14714 3816 14716
rect 3872 14714 3878 14716
rect 3632 14662 3634 14714
rect 3814 14662 3816 14714
rect 3570 14660 3576 14662
rect 3632 14660 3656 14662
rect 3712 14660 3736 14662
rect 3792 14660 3816 14662
rect 3872 14660 3878 14662
rect 3570 14651 3878 14660
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 13870 3832 14214
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3436 13190 3464 13806
rect 3570 13628 3878 13637
rect 3570 13626 3576 13628
rect 3632 13626 3656 13628
rect 3712 13626 3736 13628
rect 3792 13626 3816 13628
rect 3872 13626 3878 13628
rect 3632 13574 3634 13626
rect 3814 13574 3816 13626
rect 3570 13572 3576 13574
rect 3632 13572 3656 13574
rect 3712 13572 3736 13574
rect 3792 13572 3816 13574
rect 3872 13572 3878 13574
rect 3570 13563 3878 13572
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10266 3372 10542
rect 3436 10470 3464 13126
rect 3570 12540 3878 12549
rect 3570 12538 3576 12540
rect 3632 12538 3656 12540
rect 3712 12538 3736 12540
rect 3792 12538 3816 12540
rect 3872 12538 3878 12540
rect 3632 12486 3634 12538
rect 3814 12486 3816 12538
rect 3570 12484 3576 12486
rect 3632 12484 3656 12486
rect 3712 12484 3736 12486
rect 3792 12484 3816 12486
rect 3872 12484 3878 12486
rect 3570 12475 3878 12484
rect 4080 11898 4108 15846
rect 4356 15706 4384 16186
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4356 15162 4384 15642
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4356 14618 4384 15098
rect 4540 15026 4568 15506
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4356 14006 4384 14554
rect 4632 14482 4660 14758
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4252 13728 4304 13734
rect 4356 13716 4384 13942
rect 4304 13688 4384 13716
rect 4252 13670 4304 13676
rect 4264 13530 4292 13670
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4724 12434 4752 22066
rect 5078 22063 5134 22066
rect 7116 22066 7236 22094
rect 8312 22094 8340 22578
rect 8404 22234 8432 22578
rect 8570 22332 8878 22341
rect 8570 22330 8576 22332
rect 8632 22330 8656 22332
rect 8712 22330 8736 22332
rect 8792 22330 8816 22332
rect 8872 22330 8878 22332
rect 8632 22278 8634 22330
rect 8814 22278 8816 22330
rect 8570 22276 8576 22278
rect 8632 22276 8656 22278
rect 8712 22276 8736 22278
rect 8792 22276 8816 22278
rect 8872 22276 8878 22278
rect 8570 22267 8878 22276
rect 9232 22234 9260 22578
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 8312 22066 8524 22094
rect 5092 22030 5120 22063
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5354 21992 5410 22001
rect 5354 21927 5410 21936
rect 5448 21956 5500 21962
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5184 20058 5212 20402
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4908 18426 4936 18566
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 5092 16250 5120 16458
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4816 14618 4844 14894
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4908 14482 4936 14962
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4908 12850 4936 14418
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 5276 12782 5304 13398
rect 5368 12866 5396 21927
rect 5448 21898 5500 21904
rect 5460 19961 5488 21898
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6070 21788 6378 21797
rect 6070 21786 6076 21788
rect 6132 21786 6156 21788
rect 6212 21786 6236 21788
rect 6292 21786 6316 21788
rect 6372 21786 6378 21788
rect 6132 21734 6134 21786
rect 6314 21734 6316 21786
rect 6070 21732 6076 21734
rect 6132 21732 6156 21734
rect 6212 21732 6236 21734
rect 6292 21732 6316 21734
rect 6372 21732 6378 21734
rect 6070 21723 6378 21732
rect 6472 21593 6500 21830
rect 6458 21584 6514 21593
rect 6458 21519 6514 21528
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 20806 5948 21286
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5446 19952 5502 19961
rect 5446 19887 5502 19896
rect 5552 19446 5580 20742
rect 5644 20262 5672 20742
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19922 5672 20198
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5540 19440 5592 19446
rect 5540 19382 5592 19388
rect 5644 19378 5672 19858
rect 5920 19718 5948 20742
rect 6070 20700 6378 20709
rect 6070 20698 6076 20700
rect 6132 20698 6156 20700
rect 6212 20698 6236 20700
rect 6292 20698 6316 20700
rect 6372 20698 6378 20700
rect 6132 20646 6134 20698
rect 6314 20646 6316 20698
rect 6070 20644 6076 20646
rect 6132 20644 6156 20646
rect 6212 20644 6236 20646
rect 6292 20644 6316 20646
rect 6372 20644 6378 20646
rect 6070 20635 6378 20644
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 6070 19612 6378 19621
rect 6070 19610 6076 19612
rect 6132 19610 6156 19612
rect 6212 19610 6236 19612
rect 6292 19610 6316 19612
rect 6372 19610 6378 19612
rect 6132 19558 6134 19610
rect 6314 19558 6316 19610
rect 6070 19556 6076 19558
rect 6132 19556 6156 19558
rect 6212 19556 6236 19558
rect 6292 19556 6316 19558
rect 6372 19556 6378 19558
rect 6070 19547 6378 19556
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18902 6040 19110
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5460 18426 5488 18702
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5552 17746 5580 18566
rect 5644 18426 5672 18702
rect 6070 18524 6378 18533
rect 6070 18522 6076 18524
rect 6132 18522 6156 18524
rect 6212 18522 6236 18524
rect 6292 18522 6316 18524
rect 6372 18522 6378 18524
rect 6132 18470 6134 18522
rect 6314 18470 6316 18522
rect 6070 18468 6076 18470
rect 6132 18468 6156 18470
rect 6212 18468 6236 18470
rect 6292 18468 6316 18470
rect 6372 18468 6378 18470
rect 6070 18459 6378 18468
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5644 17542 5672 18226
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5644 17338 5672 17478
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5460 16250 5488 17138
rect 5736 16998 5764 18022
rect 5828 17542 5856 18158
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 17134 5856 17478
rect 6012 17218 6040 18022
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6380 17678 6408 17818
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6070 17436 6378 17445
rect 6070 17434 6076 17436
rect 6132 17434 6156 17436
rect 6212 17434 6236 17436
rect 6292 17434 6316 17436
rect 6372 17434 6378 17436
rect 6132 17382 6134 17434
rect 6314 17382 6316 17434
rect 6070 17380 6076 17382
rect 6132 17380 6156 17382
rect 6212 17380 6236 17382
rect 6292 17380 6316 17382
rect 6372 17380 6378 17382
rect 6070 17371 6378 17380
rect 5920 17202 6040 17218
rect 5908 17196 6040 17202
rect 5960 17190 6040 17196
rect 5908 17138 5960 17144
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 6070 16348 6378 16357
rect 6070 16346 6076 16348
rect 6132 16346 6156 16348
rect 6212 16346 6236 16348
rect 6292 16346 6316 16348
rect 6372 16346 6378 16348
rect 6132 16294 6134 16346
rect 6314 16294 6316 16346
rect 6070 16292 6076 16294
rect 6132 16292 6156 16294
rect 6212 16292 6236 16294
rect 6292 16292 6316 16294
rect 6372 16292 6378 16294
rect 6070 16283 6378 16292
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5460 16114 5488 16186
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 15570 5488 15914
rect 5828 15706 5856 15982
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 14822 5488 15506
rect 6070 15260 6378 15269
rect 6070 15258 6076 15260
rect 6132 15258 6156 15260
rect 6212 15258 6236 15260
rect 6292 15258 6316 15260
rect 6372 15258 6378 15260
rect 6132 15206 6134 15258
rect 6314 15206 6316 15258
rect 6070 15204 6076 15206
rect 6132 15204 6156 15206
rect 6212 15204 6236 15206
rect 6292 15204 6316 15206
rect 6372 15204 6378 15206
rect 6070 15195 6378 15204
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5644 14618 5672 14894
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5736 14482 5764 14894
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 6070 14172 6378 14181
rect 6070 14170 6076 14172
rect 6132 14170 6156 14172
rect 6212 14170 6236 14172
rect 6292 14170 6316 14172
rect 6372 14170 6378 14172
rect 6132 14118 6134 14170
rect 6314 14118 6316 14170
rect 6070 14116 6076 14118
rect 6132 14116 6156 14118
rect 6212 14116 6236 14118
rect 6292 14116 6316 14118
rect 6372 14116 6378 14118
rect 6070 14107 6378 14116
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 5552 13326 5580 13670
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5644 13326 5672 13466
rect 6196 13326 6224 13670
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5368 12838 5488 12866
rect 5644 12850 5672 13262
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 12986 5948 13126
rect 6070 13084 6378 13093
rect 6070 13082 6076 13084
rect 6132 13082 6156 13084
rect 6212 13082 6236 13084
rect 6292 13082 6316 13084
rect 6372 13082 6378 13084
rect 6132 13030 6134 13082
rect 6314 13030 6316 13082
rect 6070 13028 6076 13030
rect 6132 13028 6156 13030
rect 6212 13028 6236 13030
rect 6292 13028 6316 13030
rect 6372 13028 6378 13030
rect 6070 13019 6378 13028
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 4632 12406 4752 12434
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3570 11452 3878 11461
rect 3570 11450 3576 11452
rect 3632 11450 3656 11452
rect 3712 11450 3736 11452
rect 3792 11450 3816 11452
rect 3872 11450 3878 11452
rect 3632 11398 3634 11450
rect 3814 11398 3816 11450
rect 3570 11396 3576 11398
rect 3632 11396 3656 11398
rect 3712 11396 3736 11398
rect 3792 11396 3816 11398
rect 3872 11396 3878 11398
rect 3570 11387 3878 11396
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3436 9722 3464 10406
rect 3570 10364 3878 10373
rect 3570 10362 3576 10364
rect 3632 10362 3656 10364
rect 3712 10362 3736 10364
rect 3792 10362 3816 10364
rect 3872 10362 3878 10364
rect 3632 10310 3634 10362
rect 3814 10310 3816 10362
rect 3570 10308 3576 10310
rect 3632 10308 3656 10310
rect 3712 10308 3736 10310
rect 3792 10308 3816 10310
rect 3872 10308 3878 10310
rect 3570 10299 3878 10308
rect 3988 10248 4016 10406
rect 3896 10220 4016 10248
rect 3896 10062 3924 10220
rect 4172 10146 4200 11018
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10266 4384 10950
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4080 10118 4200 10146
rect 4080 10062 4108 10118
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3570 9276 3878 9285
rect 3570 9274 3576 9276
rect 3632 9274 3656 9276
rect 3712 9274 3736 9276
rect 3792 9274 3816 9276
rect 3872 9274 3878 9276
rect 3632 9222 3634 9274
rect 3814 9222 3816 9274
rect 3570 9220 3576 9222
rect 3632 9220 3656 9222
rect 3712 9220 3736 9222
rect 3792 9220 3816 9222
rect 3872 9220 3878 9222
rect 3570 9211 3878 9220
rect 4172 8974 4200 9862
rect 4356 9722 4384 9998
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9722 4476 9862
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4356 8974 4384 9658
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 3570 8188 3878 8197
rect 3570 8186 3576 8188
rect 3632 8186 3656 8188
rect 3712 8186 3736 8188
rect 3792 8186 3816 8188
rect 3872 8186 3878 8188
rect 3632 8134 3634 8186
rect 3814 8134 3816 8186
rect 3570 8132 3576 8134
rect 3632 8132 3656 8134
rect 3712 8132 3736 8134
rect 3792 8132 3816 8134
rect 3872 8132 3878 8134
rect 3570 8123 3878 8132
rect 3570 7100 3878 7109
rect 3570 7098 3576 7100
rect 3632 7098 3656 7100
rect 3712 7098 3736 7100
rect 3792 7098 3816 7100
rect 3872 7098 3878 7100
rect 3632 7046 3634 7098
rect 3814 7046 3816 7098
rect 3570 7044 3576 7046
rect 3632 7044 3656 7046
rect 3712 7044 3736 7046
rect 3792 7044 3816 7046
rect 3872 7044 3878 7046
rect 3570 7035 3878 7044
rect 3570 6012 3878 6021
rect 3570 6010 3576 6012
rect 3632 6010 3656 6012
rect 3712 6010 3736 6012
rect 3792 6010 3816 6012
rect 3872 6010 3878 6012
rect 3632 5958 3634 6010
rect 3814 5958 3816 6010
rect 3570 5956 3576 5958
rect 3632 5956 3656 5958
rect 3712 5956 3736 5958
rect 3792 5956 3816 5958
rect 3872 5956 3878 5958
rect 3570 5947 3878 5956
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1504 4554 1532 4966
rect 1596 4690 1624 4966
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1504 4214 1532 4490
rect 2332 4486 2360 4966
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1504 3754 1532 4150
rect 1504 3726 1624 3754
rect 1596 3670 1624 3726
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 756 3052 808 3058
rect 756 2994 808 3000
rect 768 2825 796 2994
rect 754 2816 810 2825
rect 754 2751 810 2760
rect 1504 2650 1532 3470
rect 1596 3194 1624 3606
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 2650 1808 2926
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1216 1760 1268 1766
rect 1216 1702 1268 1708
rect 1228 1494 1256 1702
rect 1216 1488 1268 1494
rect 1216 1430 1268 1436
rect 1320 1358 1348 2518
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 1688 2106 1716 2246
rect 2240 2106 2268 3334
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 2228 2100 2280 2106
rect 2228 2042 2280 2048
rect 2136 1760 2188 1766
rect 2136 1702 2188 1708
rect 2148 1358 2176 1702
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 2136 1352 2188 1358
rect 2136 1294 2188 1300
rect 2240 1290 2268 2042
rect 2332 1970 2360 4422
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2424 2514 2452 2790
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2516 2446 2544 5850
rect 3422 5672 3478 5681
rect 3422 5607 3478 5616
rect 2596 5568 2648 5574
rect 2872 5568 2924 5574
rect 2596 5510 2648 5516
rect 2700 5516 2872 5522
rect 2700 5510 2924 5516
rect 2608 5166 2636 5510
rect 2700 5494 2912 5510
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2700 4978 2728 5494
rect 3436 5370 3464 5607
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 2608 4950 2728 4978
rect 2608 4622 2636 4950
rect 3570 4924 3878 4933
rect 3570 4922 3576 4924
rect 3632 4922 3656 4924
rect 3712 4922 3736 4924
rect 3792 4922 3816 4924
rect 3872 4922 3878 4924
rect 3632 4870 3634 4922
rect 3814 4870 3816 4922
rect 3570 4868 3576 4870
rect 3632 4868 3656 4870
rect 3712 4868 3736 4870
rect 3792 4868 3816 4870
rect 3872 4868 3878 4870
rect 3570 4859 3878 4868
rect 3988 4622 4016 5510
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4690 4108 4966
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 2596 4616 2648 4622
rect 3516 4616 3568 4622
rect 2596 4558 2648 4564
rect 3514 4584 3516 4593
rect 3976 4616 4028 4622
rect 3568 4584 3570 4593
rect 2608 4146 2636 4558
rect 2780 4548 2832 4554
rect 3976 4558 4028 4564
rect 3514 4519 3570 4528
rect 2780 4490 2832 4496
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2608 3534 2636 4082
rect 2792 3942 2820 4490
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2608 3194 2636 3470
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2792 2650 2820 3878
rect 3344 3602 3372 3946
rect 3570 3836 3878 3845
rect 3570 3834 3576 3836
rect 3632 3834 3656 3836
rect 3712 3834 3736 3836
rect 3792 3834 3816 3836
rect 3872 3834 3878 3836
rect 3632 3782 3634 3834
rect 3814 3782 3816 3834
rect 3570 3780 3576 3782
rect 3632 3780 3656 3782
rect 3712 3780 3736 3782
rect 3792 3780 3816 3782
rect 3872 3780 3878 3782
rect 3570 3771 3878 3780
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 4080 3210 4108 4626
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3988 3182 4108 3210
rect 4172 3194 4200 4422
rect 4160 3188 4212 3194
rect 3988 2990 4016 3182
rect 4160 3130 4212 3136
rect 4068 3120 4120 3126
rect 4264 3074 4292 5850
rect 4632 5370 4660 12406
rect 5092 12374 5120 12718
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5184 12186 5212 12582
rect 5276 12442 5304 12718
rect 5264 12436 5316 12442
rect 5316 12396 5396 12424
rect 5264 12378 5316 12384
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 5080 12164 5132 12170
rect 5184 12158 5304 12186
rect 5080 12106 5132 12112
rect 5000 11937 5028 12106
rect 4986 11928 5042 11937
rect 5092 11898 5120 12106
rect 5276 12102 5304 12158
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 4986 11863 5042 11872
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5172 11824 5224 11830
rect 5170 11792 5172 11801
rect 5224 11792 5226 11801
rect 5170 11727 5226 11736
rect 5272 11756 5324 11762
rect 5368 11744 5396 12396
rect 5324 11716 5396 11744
rect 5272 11698 5324 11704
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5000 10452 5028 11086
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10606 5212 10950
rect 5368 10606 5396 11086
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5080 10464 5132 10470
rect 5000 10424 5080 10452
rect 5080 10406 5132 10412
rect 5092 9994 5120 10406
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5092 9382 5120 9930
rect 5184 9874 5212 10542
rect 5184 9846 5304 9874
rect 5276 9518 5304 9846
rect 5368 9518 5396 10542
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 5710 5028 6190
rect 5460 5914 5488 12838
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12300 5592 12306
rect 5644 12288 5672 12650
rect 6012 12306 6040 12718
rect 5592 12260 5672 12288
rect 5540 12242 5592 12248
rect 5538 11928 5594 11937
rect 5538 11863 5594 11872
rect 5552 11760 5580 11863
rect 5540 11754 5592 11760
rect 5540 11696 5592 11702
rect 5552 11626 5580 11696
rect 5644 11676 5672 12260
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6070 11996 6378 12005
rect 6070 11994 6076 11996
rect 6132 11994 6156 11996
rect 6212 11994 6236 11996
rect 6292 11994 6316 11996
rect 6372 11994 6378 11996
rect 6132 11942 6134 11994
rect 6314 11942 6316 11994
rect 6070 11940 6076 11942
rect 6132 11940 6156 11942
rect 6212 11940 6236 11942
rect 6292 11940 6316 11942
rect 6372 11940 6378 11942
rect 6070 11931 6378 11940
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5724 11824 5776 11830
rect 5722 11792 5724 11801
rect 5776 11792 5778 11801
rect 5722 11727 5778 11736
rect 5724 11688 5776 11694
rect 5644 11648 5724 11676
rect 5724 11630 5776 11636
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5736 11014 5764 11630
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5552 10266 5580 10950
rect 5920 10674 5948 11834
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10266 5856 10406
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9654 5764 9862
rect 5920 9722 5948 10610
rect 6012 10538 6040 10950
rect 6070 10908 6378 10917
rect 6070 10906 6076 10908
rect 6132 10906 6156 10908
rect 6212 10906 6236 10908
rect 6292 10906 6316 10908
rect 6372 10906 6378 10908
rect 6132 10854 6134 10906
rect 6314 10854 6316 10906
rect 6070 10852 6076 10854
rect 6132 10852 6156 10854
rect 6212 10852 6236 10854
rect 6292 10852 6316 10854
rect 6372 10852 6378 10854
rect 6070 10843 6378 10852
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6012 10130 6040 10474
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6196 9926 6224 10610
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6070 9820 6378 9829
rect 6070 9818 6076 9820
rect 6132 9818 6156 9820
rect 6212 9818 6236 9820
rect 6292 9818 6316 9820
rect 6372 9818 6378 9820
rect 6132 9766 6134 9818
rect 6314 9766 6316 9818
rect 6070 9764 6076 9766
rect 6132 9764 6156 9766
rect 6212 9764 6236 9766
rect 6292 9764 6316 9766
rect 6372 9764 6378 9766
rect 6070 9755 6378 9764
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 9178 6132 9318
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8634 6040 8842
rect 6070 8732 6378 8741
rect 6070 8730 6076 8732
rect 6132 8730 6156 8732
rect 6212 8730 6236 8732
rect 6292 8730 6316 8732
rect 6372 8730 6378 8732
rect 6132 8678 6134 8730
rect 6314 8678 6316 8730
rect 6070 8676 6076 8678
rect 6132 8676 6156 8678
rect 6212 8676 6236 8678
rect 6292 8676 6316 8678
rect 6372 8676 6378 8678
rect 6070 8667 6378 8676
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6070 7644 6378 7653
rect 6070 7642 6076 7644
rect 6132 7642 6156 7644
rect 6212 7642 6236 7644
rect 6292 7642 6316 7644
rect 6372 7642 6378 7644
rect 6132 7590 6134 7642
rect 6314 7590 6316 7642
rect 6070 7588 6076 7590
rect 6132 7588 6156 7590
rect 6212 7588 6236 7590
rect 6292 7588 6316 7590
rect 6372 7588 6378 7590
rect 6070 7579 6378 7588
rect 6070 6556 6378 6565
rect 6070 6554 6076 6556
rect 6132 6554 6156 6556
rect 6212 6554 6236 6556
rect 6292 6554 6316 6556
rect 6372 6554 6378 6556
rect 6132 6502 6134 6554
rect 6314 6502 6316 6554
rect 6070 6500 6076 6502
rect 6132 6500 6156 6502
rect 6212 6500 6236 6502
rect 6292 6500 6316 6502
rect 6372 6500 6378 6502
rect 6070 6491 6378 6500
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 4214 4384 4966
rect 4632 4622 4660 5306
rect 5000 4622 5028 5646
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5370 5488 5510
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5276 4690 5304 5102
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4988 4616 5040 4622
rect 5040 4576 5120 4604
rect 4988 4558 5040 4564
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4632 3738 4660 4422
rect 4724 4282 4752 4490
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3194 4476 3334
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4120 3068 4292 3074
rect 4068 3062 4292 3068
rect 4080 3046 4292 3062
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2976 2446 3004 2790
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2976 2106 3004 2382
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 3160 1902 3188 2450
rect 3344 1952 3372 2790
rect 3570 2748 3878 2757
rect 3570 2746 3576 2748
rect 3632 2746 3656 2748
rect 3712 2746 3736 2748
rect 3792 2746 3816 2748
rect 3872 2746 3878 2748
rect 3632 2694 3634 2746
rect 3814 2694 3816 2746
rect 3570 2692 3576 2694
rect 3632 2692 3656 2694
rect 3712 2692 3736 2694
rect 3792 2692 3816 2694
rect 3872 2692 3878 2694
rect 3570 2683 3878 2692
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3436 2106 3464 2314
rect 4080 2310 4108 2926
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 2106 4108 2246
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 3516 1964 3568 1970
rect 3344 1924 3516 1952
rect 4632 1952 4660 3674
rect 4724 3534 4752 4218
rect 5092 4146 5120 4576
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5368 4078 5396 5170
rect 5460 4729 5488 5306
rect 5446 4720 5502 4729
rect 5446 4655 5502 4664
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4282 5580 4490
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 2446 4752 3470
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4724 2106 4752 2382
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 5368 1970 5396 4014
rect 5736 3738 5764 5782
rect 6070 5468 6378 5477
rect 6070 5466 6076 5468
rect 6132 5466 6156 5468
rect 6212 5466 6236 5468
rect 6292 5466 6316 5468
rect 6372 5466 6378 5468
rect 6132 5414 6134 5466
rect 6314 5414 6316 5466
rect 6070 5412 6076 5414
rect 6132 5412 6156 5414
rect 6212 5412 6236 5414
rect 6292 5412 6316 5414
rect 6372 5412 6378 5414
rect 6070 5403 6378 5412
rect 6472 5370 6500 21519
rect 7116 21486 7144 22066
rect 8496 22030 8524 22066
rect 9600 22030 9628 22374
rect 10152 22234 10180 22578
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 6644 20868 6696 20874
rect 6644 20810 6696 20816
rect 6656 20602 6684 20810
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6748 19718 6776 21422
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6840 20398 6868 21286
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 20262 6868 20334
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 20058 6868 20198
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6748 19310 6776 19654
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6736 19304 6788 19310
rect 6734 19272 6736 19281
rect 6788 19272 6790 19281
rect 6644 19236 6696 19242
rect 6734 19207 6790 19216
rect 6644 19178 6696 19184
rect 6656 18970 6684 19178
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6564 18290 6592 18566
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6564 17542 6592 18226
rect 6736 18216 6788 18222
rect 6840 18204 6868 19314
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6788 18176 6868 18204
rect 6736 18158 6788 18164
rect 6840 17882 6868 18176
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6564 17338 6592 17478
rect 6656 17338 6684 17546
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6840 16998 6868 17818
rect 6932 17202 6960 18566
rect 7024 18086 7052 18838
rect 7116 18222 7144 18906
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7024 17134 7052 18022
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6564 16046 6592 16390
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6656 15502 6684 16526
rect 6840 16454 6868 16934
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6656 15094 6684 15438
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6656 14550 6684 15030
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6656 14074 6684 14486
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 13258 6684 14010
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 12918 6684 13194
rect 6932 12986 6960 13330
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6656 12782 6684 12854
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 7024 12442 7052 13466
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6840 11898 6868 12106
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7116 11762 7144 12242
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11354 7144 11698
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7116 10810 7144 11290
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6552 9920 6604 9926
rect 6604 9880 6684 9908
rect 6552 9862 6604 9868
rect 6656 9654 6684 9880
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6656 9178 6684 9590
rect 6932 9178 6960 9930
rect 7024 9382 7052 10066
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6656 8634 6684 9114
rect 7024 8838 7052 9318
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 7208 5914 7236 21830
rect 7300 21350 7328 21830
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 20262 7328 21286
rect 7932 20868 7984 20874
rect 7932 20810 7984 20816
rect 7944 20262 7972 20810
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7300 19786 7328 20198
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 8404 19718 8432 20198
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19514 8432 19654
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18426 7420 18566
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7576 17338 7604 19314
rect 7760 18902 7788 19314
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7760 17882 7788 18838
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7852 18426 7880 18634
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7852 17338 7880 18362
rect 8128 18290 8156 19314
rect 8116 18284 8168 18290
rect 8036 18244 8116 18272
rect 8036 17678 8064 18244
rect 8116 18226 8168 18232
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8128 17746 8156 18022
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8036 17338 8064 17614
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8036 16794 8064 17274
rect 8220 17105 8248 19382
rect 8312 18358 8340 19450
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8404 18766 8432 19246
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8404 17882 8432 18362
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8496 17762 8524 21966
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8570 21244 8878 21253
rect 8570 21242 8576 21244
rect 8632 21242 8656 21244
rect 8712 21242 8736 21244
rect 8792 21242 8816 21244
rect 8872 21242 8878 21244
rect 8632 21190 8634 21242
rect 8814 21190 8816 21242
rect 8570 21188 8576 21190
rect 8632 21188 8656 21190
rect 8712 21188 8736 21190
rect 8792 21188 8816 21190
rect 8872 21188 8878 21190
rect 8570 21179 8878 21188
rect 8956 20777 8984 21830
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9324 20874 9352 21354
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 8942 20768 8998 20777
rect 8942 20703 8998 20712
rect 9324 20602 9352 20810
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8570 20156 8878 20165
rect 8570 20154 8576 20156
rect 8632 20154 8656 20156
rect 8712 20154 8736 20156
rect 8792 20154 8816 20156
rect 8872 20154 8878 20156
rect 8632 20102 8634 20154
rect 8814 20102 8816 20154
rect 8570 20100 8576 20102
rect 8632 20100 8656 20102
rect 8712 20100 8736 20102
rect 8792 20100 8816 20102
rect 8872 20100 8878 20102
rect 8570 20091 8878 20100
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8588 19378 8616 19994
rect 9600 19922 9628 21966
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21690 10088 21830
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 20874 10272 21286
rect 10232 20868 10284 20874
rect 10232 20810 10284 20816
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9692 19854 9720 20538
rect 10244 20262 10272 20810
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10244 20074 10272 20198
rect 10152 20058 10272 20074
rect 10140 20052 10272 20058
rect 10192 20046 10272 20052
rect 10140 19994 10192 20000
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9232 19514 9260 19654
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8570 19068 8878 19077
rect 8570 19066 8576 19068
rect 8632 19066 8656 19068
rect 8712 19066 8736 19068
rect 8792 19066 8816 19068
rect 8872 19066 8878 19068
rect 8632 19014 8634 19066
rect 8814 19014 8816 19066
rect 8570 19012 8576 19014
rect 8632 19012 8656 19014
rect 8712 19012 8736 19014
rect 8792 19012 8816 19014
rect 8872 19012 8878 19014
rect 8570 19003 8878 19012
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 18290 8616 18566
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8570 17980 8878 17989
rect 8570 17978 8576 17980
rect 8632 17978 8656 17980
rect 8712 17978 8736 17980
rect 8792 17978 8816 17980
rect 8872 17978 8878 17980
rect 8632 17926 8634 17978
rect 8814 17926 8816 17978
rect 8570 17924 8576 17926
rect 8632 17924 8656 17926
rect 8712 17924 8736 17926
rect 8792 17924 8816 17926
rect 8872 17924 8878 17926
rect 8570 17915 8878 17924
rect 8404 17734 8524 17762
rect 8206 17096 8262 17105
rect 8206 17031 8262 17040
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7392 16250 7420 16730
rect 8128 16454 8156 16934
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8300 16448 8352 16454
rect 8404 16436 8432 17734
rect 9140 17678 9168 18770
rect 9324 17882 9352 19790
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9600 17882 9628 19450
rect 9876 19378 9904 19722
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 17882 9904 19314
rect 10152 18766 10180 19382
rect 10244 18970 10272 19722
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10428 18766 10456 19110
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10152 18358 10180 18702
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17338 8892 17478
rect 9784 17338 9812 17546
rect 9968 17542 9996 18022
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 8576 16992 8628 16998
rect 8496 16952 8576 16980
rect 8496 16590 8524 16952
rect 8576 16934 8628 16940
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8570 16892 8878 16901
rect 8570 16890 8576 16892
rect 8632 16890 8656 16892
rect 8712 16890 8736 16892
rect 8792 16890 8816 16892
rect 8872 16890 8878 16892
rect 8632 16838 8634 16890
rect 8814 16838 8816 16890
rect 8570 16836 8576 16838
rect 8632 16836 8656 16838
rect 8712 16836 8736 16838
rect 8792 16836 8816 16838
rect 8872 16836 8878 16838
rect 8570 16827 8878 16836
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8576 16448 8628 16454
rect 8404 16408 8524 16436
rect 8300 16390 8352 16396
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 8128 16182 8156 16390
rect 8116 16176 8168 16182
rect 8168 16124 8248 16130
rect 8116 16118 8248 16124
rect 8128 16102 8248 16118
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14550 7788 14894
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 8036 13870 8064 15506
rect 8220 15502 8248 16102
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8128 14958 8156 15438
rect 8116 14952 8168 14958
rect 8220 14940 8248 15438
rect 8312 15094 8340 16390
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8220 14912 8340 14940
rect 8116 14894 8168 14900
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14482 8248 14758
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8312 14414 8340 14912
rect 8116 14408 8168 14414
rect 8300 14408 8352 14414
rect 8116 14350 8168 14356
rect 8220 14356 8300 14362
rect 8220 14350 8352 14356
rect 8128 14074 8156 14350
rect 8220 14334 8340 14350
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 13938 8248 14334
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 14006 8432 14214
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7300 12306 7328 12922
rect 8220 12850 8248 13874
rect 8496 13818 8524 16408
rect 8576 16390 8628 16396
rect 8588 16250 8616 16390
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8570 15804 8878 15813
rect 8570 15802 8576 15804
rect 8632 15802 8656 15804
rect 8712 15802 8736 15804
rect 8792 15802 8816 15804
rect 8872 15802 8878 15804
rect 8632 15750 8634 15802
rect 8814 15750 8816 15802
rect 8570 15748 8576 15750
rect 8632 15748 8656 15750
rect 8712 15748 8736 15750
rect 8792 15748 8816 15750
rect 8872 15748 8878 15750
rect 8570 15739 8878 15748
rect 9048 14958 9076 16934
rect 9692 16726 9720 17138
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16250 9260 16390
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9600 15638 9628 16526
rect 9692 15910 9720 16662
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8570 14716 8878 14725
rect 8570 14714 8576 14716
rect 8632 14714 8656 14716
rect 8712 14714 8736 14716
rect 8792 14714 8816 14716
rect 8872 14714 8878 14716
rect 8632 14662 8634 14714
rect 8814 14662 8816 14714
rect 8570 14660 8576 14662
rect 8632 14660 8656 14662
rect 8712 14660 8736 14662
rect 8792 14660 8816 14662
rect 8872 14660 8878 14662
rect 8570 14651 8878 14660
rect 9692 14618 9720 15846
rect 9784 15570 9812 17274
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16794 9996 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 16658 10088 16934
rect 10152 16794 10180 17682
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10152 15910 10180 16730
rect 10336 16250 10364 17138
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16658 10456 16730
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10152 15706 10180 15846
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9784 15162 9812 15506
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 15162 9996 15302
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9784 14482 9812 15098
rect 10152 14958 10180 15642
rect 10428 15638 10456 15846
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14482 10088 14758
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 13938 9628 14350
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9876 13954 9904 14282
rect 10060 14278 10088 14418
rect 10152 14278 10180 14894
rect 10336 14414 10364 15098
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10140 14272 10192 14278
rect 10192 14232 10364 14260
rect 10140 14214 10192 14220
rect 10060 14074 10088 14214
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9692 13926 9904 13954
rect 10140 13932 10192 13938
rect 8404 13790 8524 13818
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11694 7420 12174
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7852 11558 7880 12582
rect 8036 12442 8064 12718
rect 8220 12646 8248 12786
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8024 12436 8076 12442
rect 8404 12434 8432 13790
rect 8570 13628 8878 13637
rect 8570 13626 8576 13628
rect 8632 13626 8656 13628
rect 8712 13626 8736 13628
rect 8792 13626 8816 13628
rect 8872 13626 8878 13628
rect 8632 13574 8634 13626
rect 8814 13574 8816 13626
rect 8570 13572 8576 13574
rect 8632 13572 8656 13574
rect 8712 13572 8736 13574
rect 8792 13572 8816 13574
rect 8872 13572 8878 13574
rect 8570 13563 8878 13572
rect 9588 13456 9640 13462
rect 9692 13410 9720 13926
rect 10140 13874 10192 13880
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9640 13404 9720 13410
rect 9588 13398 9720 13404
rect 9600 13382 9720 13398
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8496 12986 8524 13126
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 9140 12782 9168 13126
rect 9402 12880 9458 12889
rect 9402 12815 9458 12824
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9416 12646 9444 12815
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 8570 12540 8878 12549
rect 8570 12538 8576 12540
rect 8632 12538 8656 12540
rect 8712 12538 8736 12540
rect 8792 12538 8816 12540
rect 8872 12538 8878 12540
rect 8632 12486 8634 12538
rect 8814 12486 8816 12538
rect 8570 12484 8576 12486
rect 8632 12484 8656 12486
rect 8712 12484 8736 12486
rect 8792 12484 8816 12486
rect 8872 12484 8878 12486
rect 8570 12475 8878 12484
rect 8024 12378 8076 12384
rect 8312 12406 8432 12434
rect 8036 11898 8064 12378
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7668 8634 7696 11494
rect 7852 10538 7880 11494
rect 8312 10554 8340 12406
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11558 9076 12038
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8570 11452 8878 11461
rect 8570 11450 8576 11452
rect 8632 11450 8656 11452
rect 8712 11450 8736 11452
rect 8792 11450 8816 11452
rect 8872 11450 8878 11452
rect 8632 11398 8634 11450
rect 8814 11398 8816 11450
rect 8570 11396 8576 11398
rect 8632 11396 8656 11398
rect 8712 11396 8736 11398
rect 8792 11396 8816 11398
rect 8872 11396 8878 11398
rect 8570 11387 8878 11396
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 8220 10526 8340 10554
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7760 9654 7788 9998
rect 8036 9722 8064 9998
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 8220 9602 8248 10526
rect 8404 10470 8432 11018
rect 9048 10742 9076 11018
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10810 9352 10950
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9036 10736 9088 10742
rect 9088 10696 9168 10724
rect 9036 10678 9088 10684
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8496 10470 8524 10610
rect 8668 10600 8720 10606
rect 8720 10560 9076 10588
rect 8668 10542 8720 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8312 9722 8340 10406
rect 8404 9926 8432 10406
rect 8570 10364 8878 10373
rect 8570 10362 8576 10364
rect 8632 10362 8656 10364
rect 8712 10362 8736 10364
rect 8792 10362 8816 10364
rect 8872 10362 8878 10364
rect 8632 10310 8634 10362
rect 8814 10310 8816 10362
rect 8570 10308 8576 10310
rect 8632 10308 8656 10310
rect 8712 10308 8736 10310
rect 8792 10308 8816 10310
rect 8872 10308 8878 10310
rect 8570 10299 8878 10308
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 7760 9178 7788 9590
rect 8220 9574 8340 9602
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 9178 8248 9454
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 8634 8248 9114
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 7668 7546 7696 8570
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7546 7788 7686
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7668 7002 7696 7482
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7668 6662 7696 6938
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6390 7696 6598
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7668 6186 7696 6326
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4282 5948 4966
rect 6748 4486 6776 5102
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6070 4380 6378 4389
rect 6070 4378 6076 4380
rect 6132 4378 6156 4380
rect 6212 4378 6236 4380
rect 6292 4378 6316 4380
rect 6372 4378 6378 4380
rect 6132 4326 6134 4378
rect 6314 4326 6316 4378
rect 6070 4324 6076 4326
rect 6132 4324 6156 4326
rect 6212 4324 6236 4326
rect 6292 4324 6316 4326
rect 6372 4324 6378 4326
rect 6070 4315 6378 4324
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6472 3738 6500 4082
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 5736 3194 5764 3674
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2310 5764 3130
rect 5920 3058 5948 3674
rect 6656 3466 6684 3878
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6070 3292 6378 3301
rect 6070 3290 6076 3292
rect 6132 3290 6156 3292
rect 6212 3290 6236 3292
rect 6292 3290 6316 3292
rect 6372 3290 6378 3292
rect 6132 3238 6134 3290
rect 6314 3238 6316 3290
rect 6070 3236 6076 3238
rect 6132 3236 6156 3238
rect 6212 3236 6236 3238
rect 6292 3236 6316 3238
rect 6372 3236 6378 3238
rect 6070 3227 6378 3236
rect 6472 3194 6500 3334
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6656 3126 6684 3402
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5920 2774 5948 2994
rect 5920 2746 6040 2774
rect 6012 2310 6040 2746
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 4712 1964 4764 1970
rect 4632 1924 4712 1952
rect 3516 1906 3568 1912
rect 4712 1906 4764 1912
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 3148 1896 3200 1902
rect 3148 1838 3200 1844
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2872 1556 2924 1562
rect 2700 1516 2872 1544
rect 2228 1284 2280 1290
rect 2228 1226 2280 1232
rect 1308 1216 1360 1222
rect 1308 1158 1360 1164
rect 1860 1216 1912 1222
rect 1860 1158 1912 1164
rect 1030 82 1086 160
rect 1320 82 1348 1158
rect 1872 160 1900 1158
rect 2700 160 2728 1516
rect 2872 1498 2924 1504
rect 2976 1358 3004 1702
rect 3160 1494 3188 1838
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 4528 1760 4580 1766
rect 4528 1702 4580 1708
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 3570 1660 3878 1669
rect 3570 1658 3576 1660
rect 3632 1658 3656 1660
rect 3712 1658 3736 1660
rect 3792 1658 3816 1660
rect 3872 1658 3878 1660
rect 3632 1606 3634 1658
rect 3814 1606 3816 1658
rect 3570 1604 3576 1606
rect 3632 1604 3656 1606
rect 3712 1604 3736 1606
rect 3792 1604 3816 1606
rect 3872 1604 3878 1606
rect 3570 1595 3878 1604
rect 3148 1488 3200 1494
rect 3148 1430 3200 1436
rect 3988 1358 4016 1702
rect 4540 1358 4568 1702
rect 5184 1358 5212 1702
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 4528 1352 4580 1358
rect 4528 1294 4580 1300
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5736 1290 5764 2246
rect 6012 1902 6040 2246
rect 6070 2204 6378 2213
rect 6070 2202 6076 2204
rect 6132 2202 6156 2204
rect 6212 2202 6236 2204
rect 6292 2202 6316 2204
rect 6372 2202 6378 2204
rect 6132 2150 6134 2202
rect 6314 2150 6316 2202
rect 6070 2148 6076 2150
rect 6132 2148 6156 2150
rect 6212 2148 6236 2150
rect 6292 2148 6316 2150
rect 6372 2148 6378 2150
rect 6070 2139 6378 2148
rect 6748 1970 6776 4422
rect 6932 4078 6960 4422
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 7208 3534 7236 5850
rect 7300 5778 7328 6054
rect 7668 5914 7696 6122
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7300 5098 7328 5714
rect 7760 5574 7788 7482
rect 8312 5914 8340 9574
rect 8404 9058 8432 9862
rect 8496 9178 8524 9930
rect 8570 9276 8878 9285
rect 8570 9274 8576 9276
rect 8632 9274 8656 9276
rect 8712 9274 8736 9276
rect 8792 9274 8816 9276
rect 8872 9274 8878 9276
rect 8632 9222 8634 9274
rect 8814 9222 8816 9274
rect 8570 9220 8576 9222
rect 8632 9220 8656 9222
rect 8712 9220 8736 9222
rect 8792 9220 8816 9222
rect 8872 9220 8878 9222
rect 8570 9211 8878 9220
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8404 9030 8524 9058
rect 8496 8956 8524 9030
rect 8956 8974 8984 10406
rect 9048 10130 9076 10560
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9140 9722 9168 10696
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9048 8974 9076 9114
rect 8760 8968 8812 8974
rect 8496 8928 8760 8956
rect 8760 8910 8812 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9324 8906 9352 10746
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 8404 7886 8432 8842
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8430 8524 8774
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8496 8090 8524 8366
rect 8570 8188 8878 8197
rect 8570 8186 8576 8188
rect 8632 8186 8656 8188
rect 8712 8186 8736 8188
rect 8792 8186 8816 8188
rect 8872 8186 8878 8188
rect 8632 8134 8634 8186
rect 8814 8134 8816 8186
rect 8570 8132 8576 8134
rect 8632 8132 8656 8134
rect 8712 8132 8736 8134
rect 8792 8132 8816 8134
rect 8872 8132 8878 8134
rect 8570 8123 8878 8132
rect 8956 8090 8984 8502
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 9232 7546 9260 8230
rect 9324 8022 9352 8366
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 8496 6798 8524 7482
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8570 7100 8878 7109
rect 8570 7098 8576 7100
rect 8632 7098 8656 7100
rect 8712 7098 8736 7100
rect 8792 7098 8816 7100
rect 8872 7098 8878 7100
rect 8632 7046 8634 7098
rect 8814 7046 8816 7098
rect 8570 7044 8576 7046
rect 8632 7044 8656 7046
rect 8712 7044 8736 7046
rect 8792 7044 8816 7046
rect 8872 7044 8878 7046
rect 8570 7035 8878 7044
rect 8956 6934 8984 7346
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 9218 6896 9274 6905
rect 9416 6866 9444 12582
rect 9508 11898 9536 13262
rect 9600 12238 9628 13262
rect 9784 12866 9812 13806
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12986 9996 13194
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9692 12838 9812 12866
rect 9692 12646 9720 12838
rect 9772 12776 9824 12782
rect 9824 12724 9904 12730
rect 9772 12718 9904 12724
rect 9784 12702 9904 12718
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9692 11898 9720 12582
rect 9876 12434 9904 12702
rect 9784 12406 9904 12434
rect 9784 11898 9812 12406
rect 10060 12322 10088 13670
rect 10152 13258 10180 13874
rect 10244 13530 10272 13874
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 12850 10180 13194
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9876 12306 10088 12322
rect 9864 12300 10088 12306
rect 9916 12294 10088 12300
rect 9864 12242 9916 12248
rect 10152 12170 10180 12786
rect 10336 12434 10364 14232
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13394 10548 13670
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10244 12406 10364 12434
rect 10612 12434 10640 22442
rect 11164 22234 11192 22578
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11070 21788 11378 21797
rect 11070 21786 11076 21788
rect 11132 21786 11156 21788
rect 11212 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11378 21788
rect 11132 21734 11134 21786
rect 11314 21734 11316 21786
rect 11070 21732 11076 21734
rect 11132 21732 11156 21734
rect 11212 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11378 21734
rect 11070 21723 11378 21732
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20942 11100 21286
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11070 20700 11378 20709
rect 11070 20698 11076 20700
rect 11132 20698 11156 20700
rect 11212 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11378 20700
rect 11132 20646 11134 20698
rect 11314 20646 11316 20698
rect 11070 20644 11076 20646
rect 11132 20644 11156 20646
rect 11212 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11378 20646
rect 11070 20635 11378 20644
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10980 19854 11008 20198
rect 11440 20058 11468 20742
rect 11624 20369 11652 21830
rect 11716 21457 11744 21830
rect 11702 21448 11758 21457
rect 11702 21383 11758 21392
rect 11900 20942 11928 22374
rect 11992 22234 12020 22578
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12728 22030 12756 23054
rect 12820 22778 12848 23840
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13648 22778 13676 22986
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13740 22658 13768 23840
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14568 22778 14596 23190
rect 14660 22778 14688 23840
rect 14924 23384 14976 23390
rect 14924 23326 14976 23332
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 13832 22658 13860 22714
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 13452 22636 13504 22642
rect 13740 22630 13860 22658
rect 14740 22636 14792 22642
rect 13452 22578 13504 22584
rect 14740 22578 14792 22584
rect 12808 22568 12860 22574
rect 12806 22536 12808 22545
rect 12860 22536 12862 22545
rect 12806 22471 12862 22480
rect 12912 22234 12940 22578
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 13372 22094 13400 22374
rect 13464 22234 13492 22578
rect 13570 22332 13878 22341
rect 13570 22330 13576 22332
rect 13632 22330 13656 22332
rect 13712 22330 13736 22332
rect 13792 22330 13816 22332
rect 13872 22330 13878 22332
rect 13632 22278 13634 22330
rect 13814 22278 13816 22330
rect 13570 22276 13576 22278
rect 13632 22276 13656 22278
rect 13712 22276 13736 22278
rect 13792 22276 13816 22278
rect 13872 22276 13878 22278
rect 13570 22267 13878 22276
rect 14752 22234 14780 22578
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14016 22094 14044 22170
rect 14936 22094 14964 23326
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15120 22778 15148 23258
rect 15580 22778 15608 23840
rect 16070 22876 16378 22885
rect 16070 22874 16076 22876
rect 16132 22874 16156 22876
rect 16212 22874 16236 22876
rect 16292 22874 16316 22876
rect 16372 22874 16378 22876
rect 16132 22822 16134 22874
rect 16314 22822 16316 22874
rect 16070 22820 16076 22822
rect 16132 22820 16156 22822
rect 16212 22820 16236 22822
rect 16292 22820 16316 22822
rect 16372 22820 16378 22822
rect 16070 22811 16378 22820
rect 16500 22778 16528 23840
rect 17420 22778 17448 23840
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 15396 22506 15424 22578
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 13372 22066 13492 22094
rect 14016 22066 14964 22094
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 12084 21486 12112 21966
rect 13096 21554 13124 21966
rect 13464 21894 13492 22066
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11610 20360 11666 20369
rect 11610 20295 11666 20304
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19446 10916 19654
rect 10980 19514 11008 19790
rect 11070 19612 11378 19621
rect 11070 19610 11076 19612
rect 11132 19610 11156 19612
rect 11212 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11378 19612
rect 11132 19558 11134 19610
rect 11314 19558 11316 19610
rect 11070 19556 11076 19558
rect 11132 19556 11156 19558
rect 11212 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11378 19558
rect 11070 19547 11378 19556
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10704 18766 10732 19246
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10796 18630 10824 19246
rect 10888 18766 10916 19382
rect 11440 18970 11468 19858
rect 12084 19825 12112 21422
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12636 21049 12664 21286
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12622 21040 12678 21049
rect 12622 20975 12678 20984
rect 12728 20806 12756 21082
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12164 19848 12216 19854
rect 12070 19816 12126 19825
rect 12164 19790 12216 19796
rect 12070 19751 12126 19760
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11624 19174 11652 19654
rect 12176 19514 12204 19790
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18222 10824 18566
rect 11070 18524 11378 18533
rect 11070 18522 11076 18524
rect 11132 18522 11156 18524
rect 11212 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11378 18524
rect 11132 18470 11134 18522
rect 11314 18470 11316 18522
rect 11070 18468 11076 18470
rect 11132 18468 11156 18470
rect 11212 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11378 18470
rect 11070 18459 11378 18468
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 11440 18170 11468 18906
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11624 18426 11652 18634
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11900 18290 11928 18906
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11612 18216 11664 18222
rect 10796 17954 10824 18158
rect 11440 18142 11560 18170
rect 11992 18170 12020 18226
rect 11664 18164 12020 18170
rect 11612 18158 12020 18164
rect 11624 18142 12020 18158
rect 11532 18086 11560 18142
rect 12084 18086 12112 18566
rect 12176 18290 12204 19450
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 10796 17926 10916 17954
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10796 17202 10824 17478
rect 10888 17202 10916 17926
rect 11348 17814 11376 18022
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11070 17436 11378 17445
rect 11070 17434 11076 17436
rect 11132 17434 11156 17436
rect 11212 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11378 17436
rect 11132 17382 11134 17434
rect 11314 17382 11316 17434
rect 11070 17380 11076 17382
rect 11132 17380 11156 17382
rect 11212 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11378 17382
rect 11070 17371 11378 17380
rect 12268 17202 12296 17682
rect 12360 17678 12388 19994
rect 12544 19990 12572 20538
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 17746 12572 18226
rect 12728 17882 12756 20742
rect 12808 19304 12860 19310
rect 12860 19264 13032 19292
rect 12808 19246 12860 19252
rect 13004 18766 13032 19264
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13004 18426 13032 18702
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13004 17882 13032 18362
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 10704 16794 10732 17138
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10796 15434 10824 16934
rect 12268 16674 12296 17138
rect 12452 16998 12480 17478
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 11900 16658 12296 16674
rect 11888 16652 12296 16658
rect 11940 16646 12296 16652
rect 11888 16594 11940 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11070 16348 11378 16357
rect 11070 16346 11076 16348
rect 11132 16346 11156 16348
rect 11212 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11378 16348
rect 11132 16294 11134 16346
rect 11314 16294 11316 16346
rect 11070 16292 11076 16294
rect 11132 16292 11156 16294
rect 11212 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11378 16294
rect 11070 16283 11378 16292
rect 11440 16182 11468 16526
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15434 11192 15982
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11070 15260 11378 15269
rect 11070 15258 11076 15260
rect 11132 15258 11156 15260
rect 11212 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11378 15260
rect 11132 15206 11134 15258
rect 11314 15206 11316 15258
rect 11070 15204 11076 15206
rect 11132 15204 11156 15206
rect 11212 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11378 15206
rect 11070 15195 11378 15204
rect 11440 15026 11468 16118
rect 11532 15706 11560 16390
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11624 15162 11652 16458
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 15366 11836 16390
rect 12176 15910 12204 16526
rect 12268 16114 12296 16646
rect 12452 16454 12480 16934
rect 12440 16448 12492 16454
rect 12360 16408 12440 16436
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12268 15502 12296 16050
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11808 15026 11836 15302
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12360 14958 12388 16408
rect 12440 16390 12492 16396
rect 12728 15978 12756 17818
rect 13004 17610 13032 17818
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12820 17338 12848 17478
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 13004 16794 13032 17546
rect 13096 17241 13124 21490
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13372 21078 13400 21286
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13372 19922 13400 20470
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 18086 13216 18634
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13372 17882 13400 18226
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17338 13400 17614
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13082 17232 13138 17241
rect 13082 17167 13138 17176
rect 12992 16788 13044 16794
rect 12912 16748 12992 16776
rect 12912 16114 12940 16748
rect 12992 16730 13044 16736
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15706 12664 15846
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12728 15042 12756 15914
rect 13372 15502 13400 16390
rect 12808 15496 12860 15502
rect 13360 15496 13412 15502
rect 12808 15438 12860 15444
rect 12820 15094 12848 15438
rect 13004 15422 13216 15450
rect 13360 15438 13412 15444
rect 13004 15366 13032 15422
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12636 15014 12756 15042
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 13096 15026 13124 15302
rect 13188 15026 13216 15422
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13280 15162 13308 15370
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13084 15020 13136 15026
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14346 11928 14758
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 10704 14074 10732 14214
rect 11070 14172 11378 14181
rect 11070 14170 11076 14172
rect 11132 14170 11156 14172
rect 11212 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11378 14172
rect 11132 14118 11134 14170
rect 11314 14118 11316 14170
rect 11070 14116 11076 14118
rect 11132 14116 11156 14118
rect 11212 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11378 14118
rect 11070 14107 11378 14116
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11348 13326 11376 13806
rect 11440 13530 11468 14214
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11070 13084 11378 13093
rect 11070 13082 11076 13084
rect 11132 13082 11156 13084
rect 11212 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11378 13084
rect 11132 13030 11134 13082
rect 11314 13030 11316 13082
rect 11070 13028 11076 13030
rect 11132 13028 11156 13030
rect 11212 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11378 13030
rect 11070 13019 11378 13028
rect 11440 12986 11468 13466
rect 11532 13190 11560 14214
rect 12268 13530 12296 14214
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11336 12844 11388 12850
rect 11532 12832 11560 13126
rect 11388 12804 11560 12832
rect 11336 12786 11388 12792
rect 11348 12442 11376 12786
rect 11624 12764 11652 13126
rect 11532 12736 11652 12764
rect 11336 12436 11388 12442
rect 10612 12406 10732 12434
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 11898 10180 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10152 11354 10180 11834
rect 10244 11694 10272 12406
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 8974 9536 11018
rect 9692 10266 9720 11086
rect 10048 10668 10100 10674
rect 10152 10656 10180 11290
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10742 10272 10950
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10100 10628 10180 10656
rect 10048 10610 10100 10616
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 9586 9628 9862
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9692 9382 9720 10202
rect 10060 10062 10088 10610
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10060 9518 10088 9998
rect 10152 9722 10180 9998
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 8974 9720 9318
rect 10060 9110 10088 9454
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8430 9628 8774
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9600 6934 9628 7890
rect 9968 7342 9996 9046
rect 10152 8922 10180 9658
rect 10428 9586 10456 10406
rect 10520 10266 10548 11086
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10612 9654 10640 11086
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9178 10548 9522
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10060 8894 10180 8922
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10060 8022 10088 8894
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8634 10180 8774
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8090 10180 8570
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7546 10088 7958
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10060 7002 10088 7482
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9218 6831 9274 6840
rect 9404 6860 9456 6866
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 6322 8524 6734
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8570 6012 8878 6021
rect 8570 6010 8576 6012
rect 8632 6010 8656 6012
rect 8712 6010 8736 6012
rect 8792 6010 8816 6012
rect 8872 6010 8878 6012
rect 8632 5958 8634 6010
rect 8814 5958 8816 6010
rect 8570 5956 8576 5958
rect 8632 5956 8656 5958
rect 8712 5956 8736 5958
rect 8792 5956 8816 5958
rect 8872 5956 8878 5958
rect 8570 5947 8878 5956
rect 8300 5908 8352 5914
rect 8352 5868 8432 5896
rect 8300 5850 8352 5856
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5370 7788 5510
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 8404 5302 8432 5868
rect 9140 5574 9168 6258
rect 9232 5914 9260 6831
rect 9404 6802 9456 6808
rect 9416 6390 9444 6802
rect 10244 6662 10272 8910
rect 10336 8498 10364 9046
rect 10324 8492 10376 8498
rect 10376 8452 10640 8480
rect 10324 8434 10376 8440
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 7750 10456 8298
rect 10508 8084 10560 8090
rect 10612 8072 10640 8452
rect 10560 8044 10640 8072
rect 10508 8026 10560 8032
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7342 10456 7686
rect 10520 7410 10548 8026
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10612 7546 10640 7754
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10428 6730 10456 7278
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10520 6390 10548 7346
rect 10612 7206 10640 7482
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 7002 10640 7142
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10612 6118 10640 6598
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 10336 5710 10364 6054
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 9140 5302 9168 5510
rect 9968 5370 9996 5510
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4690 8340 4966
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4146 7972 4422
rect 8312 4214 8340 4626
rect 8404 4622 8432 5238
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4690 8524 4966
rect 8570 4924 8878 4933
rect 8570 4922 8576 4924
rect 8632 4922 8656 4924
rect 8712 4922 8736 4924
rect 8792 4922 8816 4924
rect 8872 4922 8878 4924
rect 8632 4870 8634 4922
rect 8814 4870 8816 4922
rect 8570 4868 8576 4870
rect 8632 4868 8656 4870
rect 8712 4868 8736 4870
rect 8792 4868 8816 4870
rect 8872 4868 8878 4870
rect 8570 4859 8878 4868
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7944 3738 7972 4082
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3194 7236 3334
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 6012 1562 6040 1838
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 6196 1358 6224 1702
rect 6920 1556 6972 1562
rect 6840 1516 6920 1544
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 5724 1284 5776 1290
rect 5724 1226 5776 1232
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 6000 1216 6052 1222
rect 6000 1158 6052 1164
rect 3528 160 3556 1158
rect 1030 54 1348 82
rect 1030 -300 1086 54
rect 1858 -300 1914 160
rect 2686 -300 2742 160
rect 3514 -300 3570 160
rect 4342 82 4398 160
rect 4632 82 4660 1158
rect 4342 54 4660 82
rect 5170 82 5226 160
rect 5460 82 5488 1158
rect 6012 160 6040 1158
rect 6070 1116 6378 1125
rect 6070 1114 6076 1116
rect 6132 1114 6156 1116
rect 6212 1114 6236 1116
rect 6292 1114 6316 1116
rect 6372 1114 6378 1116
rect 6132 1062 6134 1114
rect 6314 1062 6316 1114
rect 6070 1060 6076 1062
rect 6132 1060 6156 1062
rect 6212 1060 6236 1062
rect 6292 1060 6316 1062
rect 6372 1060 6378 1062
rect 6070 1051 6378 1060
rect 6840 160 6868 1516
rect 6920 1498 6972 1504
rect 7024 1358 7052 2518
rect 7208 2446 7236 3130
rect 7944 2774 7972 3674
rect 8312 3534 8340 4150
rect 8404 3942 8432 4422
rect 9140 4282 9168 5238
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 3058 8340 3470
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8298 2952 8354 2961
rect 8298 2887 8300 2896
rect 8352 2887 8354 2896
rect 8300 2858 8352 2864
rect 8404 2774 8432 3878
rect 8570 3836 8878 3845
rect 8570 3834 8576 3836
rect 8632 3834 8656 3836
rect 8712 3834 8736 3836
rect 8792 3834 8816 3836
rect 8872 3834 8878 3836
rect 8632 3782 8634 3834
rect 8814 3782 8816 3834
rect 8570 3780 8576 3782
rect 8632 3780 8656 3782
rect 8712 3780 8736 3782
rect 8792 3780 8816 3782
rect 8872 3780 8878 3782
rect 8570 3771 8878 3780
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8588 3194 8616 3402
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2938 8616 2994
rect 8956 2990 8984 3878
rect 9048 3738 9076 3878
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9324 3602 9352 4626
rect 10428 4486 10456 5510
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 9600 4282 9628 4422
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9324 2990 9352 3538
rect 7944 2746 8156 2774
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8128 2310 8156 2746
rect 8312 2746 8432 2774
rect 8496 2910 8616 2938
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8128 1834 8156 2246
rect 8312 1970 8340 2746
rect 8496 2650 8524 2910
rect 8570 2748 8878 2757
rect 8570 2746 8576 2748
rect 8632 2746 8656 2748
rect 8712 2746 8736 2748
rect 8792 2746 8816 2748
rect 8872 2746 8878 2748
rect 8632 2694 8634 2746
rect 8814 2694 8816 2746
rect 8570 2692 8576 2694
rect 8632 2692 8656 2694
rect 8712 2692 8736 2694
rect 8792 2692 8816 2694
rect 8872 2692 8878 2694
rect 8570 2683 8878 2692
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 9692 2514 9720 3606
rect 10140 3460 10192 3466
rect 10244 3448 10272 4082
rect 10428 3641 10456 4422
rect 10414 3632 10470 3641
rect 10414 3567 10470 3576
rect 10520 3534 10548 5850
rect 10704 5166 10732 12406
rect 11336 12378 11388 12384
rect 11070 11996 11378 12005
rect 11070 11994 11076 11996
rect 11132 11994 11156 11996
rect 11212 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11378 11996
rect 11132 11942 11134 11994
rect 11314 11942 11316 11994
rect 11070 11940 11076 11942
rect 11132 11940 11156 11942
rect 11212 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11378 11942
rect 11070 11931 11378 11940
rect 11532 11626 11560 12736
rect 11716 12442 11744 13194
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12238 11836 12582
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 12176 12102 12204 13194
rect 12360 12782 12388 14418
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12442 12480 13670
rect 12440 12436 12492 12442
rect 12544 12434 12572 14214
rect 12636 12850 12664 15014
rect 13084 14962 13136 14968
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13096 14618 13124 14962
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 13530 12940 14214
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12912 12986 12940 13466
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13188 12918 13216 14962
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 12912 13228 12918
rect 12714 12880 12770 12889
rect 12624 12844 12676 12850
rect 13176 12854 13228 12860
rect 13280 12850 13308 14758
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13372 12918 13400 14010
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 12714 12815 12716 12824
rect 12624 12786 12676 12792
rect 12768 12815 12770 12824
rect 13268 12844 13320 12850
rect 12716 12786 12768 12792
rect 13268 12786 13320 12792
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12544 12406 12664 12434
rect 12440 12378 12492 12384
rect 12636 12238 12664 12406
rect 13004 12238 13032 12718
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12176 11898 12204 12038
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 11144 11480 11150
rect 11480 11092 11560 11098
rect 11428 11086 11560 11092
rect 11440 11070 11560 11086
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11070 10908 11378 10917
rect 11070 10906 11076 10908
rect 11132 10906 11156 10908
rect 11212 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11378 10908
rect 11132 10854 11134 10906
rect 11314 10854 11316 10906
rect 11070 10852 11076 10854
rect 11132 10852 11156 10854
rect 11212 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11378 10854
rect 11070 10843 11378 10852
rect 11440 10742 11468 10950
rect 11532 10810 11560 11070
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11624 10606 11652 11630
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 10796 9994 10824 10542
rect 11716 10266 11744 10950
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11808 10606 11836 10746
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10266 11836 10542
rect 11900 10470 11928 11698
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11888 10464 11940 10470
rect 11940 10424 12020 10452
rect 11888 10406 11940 10412
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11070 9820 11378 9829
rect 11070 9818 11076 9820
rect 11132 9818 11156 9820
rect 11212 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11378 9820
rect 11132 9766 11134 9818
rect 11314 9766 11316 9818
rect 11070 9764 11076 9766
rect 11132 9764 11156 9766
rect 11212 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11378 9766
rect 11070 9755 11378 9764
rect 11532 9586 11560 9862
rect 11808 9586 11836 10202
rect 11992 10062 12020 10424
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11992 9382 12020 9998
rect 12084 9654 12112 11086
rect 12176 10742 12204 11834
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11354 12572 11630
rect 12636 11558 12664 12038
rect 12992 11824 13044 11830
rect 13044 11784 13124 11812
rect 12992 11766 13044 11772
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12636 11286 12664 11494
rect 13096 11286 13124 11784
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10198 12204 10678
rect 12360 10266 12388 11086
rect 13004 10674 13032 11222
rect 13096 10810 13124 11222
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12360 9518 12388 10202
rect 12728 9926 12756 10406
rect 12820 10266 12848 10406
rect 13096 10282 13124 10746
rect 13280 10577 13308 12786
rect 13360 10600 13412 10606
rect 13266 10568 13322 10577
rect 13360 10542 13412 10548
rect 13266 10503 13322 10512
rect 12808 10260 12860 10266
rect 13096 10254 13308 10282
rect 13372 10266 13400 10542
rect 12808 10202 12860 10208
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13280 10146 13308 10254
rect 13360 10260 13412 10266
rect 13464 10248 13492 21830
rect 13924 21622 13952 21898
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13570 21244 13878 21253
rect 13570 21242 13576 21244
rect 13632 21242 13656 21244
rect 13712 21242 13736 21244
rect 13792 21242 13816 21244
rect 13872 21242 13878 21244
rect 13632 21190 13634 21242
rect 13814 21190 13816 21242
rect 13570 21188 13576 21190
rect 13632 21188 13656 21190
rect 13712 21188 13736 21190
rect 13792 21188 13816 21190
rect 13872 21188 13878 21190
rect 13570 21179 13878 21188
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13556 20602 13584 20810
rect 13832 20602 13860 21014
rect 13924 20924 13952 21558
rect 14002 21176 14058 21185
rect 14002 21111 14004 21120
rect 14056 21111 14058 21120
rect 14004 21082 14056 21088
rect 13924 20896 14044 20924
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13570 20156 13878 20165
rect 13570 20154 13576 20156
rect 13632 20154 13656 20156
rect 13712 20154 13736 20156
rect 13792 20154 13816 20156
rect 13872 20154 13878 20156
rect 13632 20102 13634 20154
rect 13814 20102 13816 20154
rect 13570 20100 13576 20102
rect 13632 20100 13656 20102
rect 13712 20100 13736 20102
rect 13792 20100 13816 20102
rect 13872 20100 13878 20102
rect 13570 20091 13878 20100
rect 13924 19718 13952 20198
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 19446 13952 19654
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 13570 19068 13878 19077
rect 13570 19066 13576 19068
rect 13632 19066 13656 19068
rect 13712 19066 13736 19068
rect 13792 19066 13816 19068
rect 13872 19066 13878 19068
rect 13632 19014 13634 19066
rect 13814 19014 13816 19066
rect 13570 19012 13576 19014
rect 13632 19012 13656 19014
rect 13712 19012 13736 19014
rect 13792 19012 13816 19014
rect 13872 19012 13878 19014
rect 13570 19003 13878 19012
rect 14016 18873 14044 20896
rect 14002 18864 14058 18873
rect 14002 18799 14058 18808
rect 13570 17980 13878 17989
rect 13570 17978 13576 17980
rect 13632 17978 13656 17980
rect 13712 17978 13736 17980
rect 13792 17978 13816 17980
rect 13872 17978 13878 17980
rect 13632 17926 13634 17978
rect 13814 17926 13816 17978
rect 13570 17924 13576 17926
rect 13632 17924 13656 17926
rect 13712 17924 13736 17926
rect 13792 17924 13816 17926
rect 13872 17924 13878 17926
rect 13570 17915 13878 17924
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13570 16892 13878 16901
rect 13570 16890 13576 16892
rect 13632 16890 13656 16892
rect 13712 16890 13736 16892
rect 13792 16890 13816 16892
rect 13872 16890 13878 16892
rect 13632 16838 13634 16890
rect 13814 16838 13816 16890
rect 13570 16836 13576 16838
rect 13632 16836 13656 16838
rect 13712 16836 13736 16838
rect 13792 16836 13816 16838
rect 13872 16836 13878 16838
rect 13570 16827 13878 16836
rect 13570 15804 13878 15813
rect 13570 15802 13576 15804
rect 13632 15802 13656 15804
rect 13712 15802 13736 15804
rect 13792 15802 13816 15804
rect 13872 15802 13878 15804
rect 13632 15750 13634 15802
rect 13814 15750 13816 15802
rect 13570 15748 13576 15750
rect 13632 15748 13656 15750
rect 13712 15748 13736 15750
rect 13792 15748 13816 15750
rect 13872 15748 13878 15750
rect 13570 15739 13878 15748
rect 13924 15434 13952 17614
rect 14108 15586 14136 21830
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 20346 14228 21422
rect 14292 21321 14320 21626
rect 14476 21486 14504 21966
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14278 21312 14334 21321
rect 14278 21247 14334 21256
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14292 20505 14320 20538
rect 14278 20496 14334 20505
rect 14384 20466 14412 20878
rect 14476 20874 14504 21422
rect 14568 21146 14596 21422
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14464 20528 14516 20534
rect 14462 20496 14464 20505
rect 14516 20496 14518 20505
rect 14278 20431 14334 20440
rect 14372 20460 14424 20466
rect 14462 20431 14518 20440
rect 14372 20402 14424 20408
rect 14200 20330 14412 20346
rect 14200 20324 14424 20330
rect 14200 20318 14372 20324
rect 14372 20266 14424 20272
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 20097 14228 20198
rect 14186 20088 14242 20097
rect 14186 20023 14242 20032
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 18834 14412 19654
rect 14372 18828 14424 18834
rect 14476 18816 14504 19722
rect 14568 18970 14596 19790
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14556 18828 14608 18834
rect 14476 18788 14556 18816
rect 14372 18770 14424 18776
rect 14556 18770 14608 18776
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17202 14320 17478
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14292 16454 14320 17138
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16114 14320 16390
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15706 14228 15982
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14108 15558 14228 15586
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 14200 15026 14228 15558
rect 14292 15502 14320 15846
rect 14568 15706 14596 16594
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14568 15162 14596 15642
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 13570 14716 13878 14725
rect 13570 14714 13576 14716
rect 13632 14714 13656 14716
rect 13712 14714 13736 14716
rect 13792 14714 13816 14716
rect 13872 14714 13878 14716
rect 13632 14662 13634 14714
rect 13814 14662 13816 14714
rect 13570 14660 13576 14662
rect 13632 14660 13656 14662
rect 13712 14660 13736 14662
rect 13792 14660 13816 14662
rect 13872 14660 13878 14662
rect 13570 14651 13878 14660
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13556 14278 13584 14554
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13556 14074 13584 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13648 13841 13676 13942
rect 13924 13870 13952 14214
rect 14016 14074 14044 14282
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 13864 13964 13870
rect 13634 13832 13690 13841
rect 13912 13806 13964 13812
rect 13634 13767 13690 13776
rect 13570 13628 13878 13637
rect 13570 13626 13576 13628
rect 13632 13626 13656 13628
rect 13712 13626 13736 13628
rect 13792 13626 13816 13628
rect 13872 13626 13878 13628
rect 13632 13574 13634 13626
rect 13814 13574 13816 13626
rect 13570 13572 13576 13574
rect 13632 13572 13656 13574
rect 13712 13572 13736 13574
rect 13792 13572 13816 13574
rect 13872 13572 13878 13574
rect 13570 13563 13878 13572
rect 13924 12986 13952 13806
rect 14016 13258 14044 14010
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14016 12986 14044 13194
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13570 12540 13878 12549
rect 13570 12538 13576 12540
rect 13632 12538 13656 12540
rect 13712 12538 13736 12540
rect 13792 12538 13816 12540
rect 13872 12538 13878 12540
rect 13632 12486 13634 12538
rect 13814 12486 13816 12538
rect 13570 12484 13576 12486
rect 13632 12484 13656 12486
rect 13712 12484 13736 12486
rect 13792 12484 13816 12486
rect 13872 12484 13878 12486
rect 13570 12475 13878 12484
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11898 13860 12038
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14016 11694 14044 12718
rect 14108 12646 14136 14962
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13734 14228 14214
rect 14278 13832 14334 13841
rect 14384 13818 14412 14758
rect 14568 14278 14596 15098
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14334 13790 14412 13818
rect 14278 13767 14334 13776
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12782 14320 13330
rect 14384 13258 14412 13790
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14384 12918 14412 13194
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14292 12238 14320 12718
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14384 11812 14412 12854
rect 14464 11824 14516 11830
rect 14384 11784 14464 11812
rect 14464 11766 14516 11772
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13570 11452 13878 11461
rect 13570 11450 13576 11452
rect 13632 11450 13656 11452
rect 13712 11450 13736 11452
rect 13792 11450 13816 11452
rect 13872 11450 13878 11452
rect 13632 11398 13634 11450
rect 13814 11398 13816 11450
rect 13570 11396 13576 11398
rect 13632 11396 13656 11398
rect 13712 11396 13736 11398
rect 13792 11396 13816 11398
rect 13872 11396 13878 11398
rect 13570 11387 13878 11396
rect 13820 11212 13872 11218
rect 13924 11200 13952 11494
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 13872 11172 13952 11200
rect 13820 11154 13872 11160
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 14004 11144 14056 11150
rect 14056 11104 14228 11132
rect 14004 11086 14056 11092
rect 13636 11008 13688 11014
rect 13740 10985 13768 11086
rect 13912 11008 13964 11014
rect 13636 10950 13688 10956
rect 13726 10976 13782 10985
rect 13648 10606 13676 10950
rect 13912 10950 13964 10956
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13726 10911 13782 10920
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13570 10364 13878 10373
rect 13570 10362 13576 10364
rect 13632 10362 13656 10364
rect 13712 10362 13736 10364
rect 13792 10362 13816 10364
rect 13872 10362 13878 10364
rect 13632 10310 13634 10362
rect 13814 10310 13816 10362
rect 13570 10308 13576 10310
rect 13632 10308 13656 10310
rect 13712 10308 13736 10310
rect 13792 10308 13816 10310
rect 13872 10308 13878 10310
rect 13570 10299 13878 10308
rect 13464 10220 13676 10248
rect 13360 10202 13412 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11256 9217 11284 9318
rect 11242 9208 11298 9217
rect 11060 9172 11112 9178
rect 11242 9143 11298 9152
rect 11060 9114 11112 9120
rect 11072 8820 11100 9114
rect 10796 8792 11100 8820
rect 10796 8294 10824 8792
rect 11070 8732 11378 8741
rect 11070 8730 11076 8732
rect 11132 8730 11156 8732
rect 11212 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11378 8732
rect 11132 8678 11134 8730
rect 11314 8678 11316 8730
rect 11070 8676 11076 8678
rect 11132 8676 11156 8678
rect 11212 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11378 8678
rect 11070 8667 11378 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11256 8514 11284 8570
rect 11532 8514 11560 9318
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 8945 12020 9114
rect 11978 8936 12034 8945
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11888 8900 11940 8906
rect 11978 8871 12034 8880
rect 11888 8842 11940 8848
rect 11256 8486 11560 8514
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7954 10916 8230
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 11070 7644 11378 7653
rect 11070 7642 11076 7644
rect 11132 7642 11156 7644
rect 11212 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11378 7644
rect 11132 7590 11134 7642
rect 11314 7590 11316 7642
rect 11070 7588 11076 7590
rect 11132 7588 11156 7590
rect 11212 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11378 7590
rect 11070 7579 11378 7588
rect 11440 7546 11468 8486
rect 11716 8430 11744 8842
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11808 7750 11836 8502
rect 11900 8294 11928 8842
rect 12084 8634 12112 9318
rect 12440 8832 12492 8838
rect 12544 8820 12572 9590
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12492 8792 12572 8820
rect 12440 8774 12492 8780
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 8090 11928 8230
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11808 7410 11836 7686
rect 11900 7546 11928 8026
rect 12452 7886 12480 8434
rect 12544 8430 12572 8792
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12544 7750 12572 8366
rect 12636 7886 12664 9318
rect 12728 9178 12756 9522
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8650 12756 8842
rect 12820 8838 12848 9522
rect 12912 9382 12940 9522
rect 12900 9376 12952 9382
rect 13004 9364 13032 9998
rect 13096 9602 13124 10134
rect 13188 10062 13216 10134
rect 13280 10118 13492 10146
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9722 13308 9998
rect 13464 9722 13492 10118
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9722 13584 9862
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13360 9648 13412 9654
rect 13096 9596 13360 9602
rect 13096 9590 13412 9596
rect 13096 9574 13400 9590
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13004 9336 13124 9364
rect 12900 9318 12952 9324
rect 12992 9104 13044 9110
rect 13096 9081 13124 9336
rect 13266 9208 13322 9217
rect 13372 9178 13400 9454
rect 13266 9143 13322 9152
rect 13360 9172 13412 9178
rect 12992 9046 13044 9052
rect 13082 9072 13138 9081
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12728 8622 12848 8650
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 8022 12756 8434
rect 12820 8362 12848 8622
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12912 8090 12940 8910
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 13004 7750 13032 9046
rect 13082 9007 13138 9016
rect 13096 8906 13124 9007
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13084 8560 13136 8566
rect 13188 8548 13216 8842
rect 13280 8634 13308 9143
rect 13464 9160 13492 9658
rect 13648 9364 13676 10220
rect 13924 9926 13952 10950
rect 14016 10470 14044 10950
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14108 9994 14136 10202
rect 14200 9994 14228 11104
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10810 14320 10950
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14292 10062 14320 10746
rect 14384 10130 14412 11222
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14476 10266 14504 11086
rect 14660 10656 14688 22066
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21690 14780 21966
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 15488 21418 15516 22578
rect 15672 22030 15700 22578
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15672 21418 15700 21830
rect 15856 21622 15884 22374
rect 16776 22234 16804 22578
rect 17132 22568 17184 22574
rect 17130 22536 17132 22545
rect 17184 22536 17186 22545
rect 17130 22471 17186 22480
rect 17512 22234 17540 22578
rect 17972 22545 18000 23462
rect 18340 22778 18368 23840
rect 19260 22778 19288 23840
rect 20180 22778 20208 23840
rect 21100 23066 21128 23840
rect 21008 23038 21128 23066
rect 21008 22778 21036 23038
rect 21070 22876 21378 22885
rect 21070 22874 21076 22876
rect 21132 22874 21156 22876
rect 21212 22874 21236 22876
rect 21292 22874 21316 22876
rect 21372 22874 21378 22876
rect 21132 22822 21134 22874
rect 21314 22822 21316 22874
rect 21070 22820 21076 22822
rect 21132 22820 21156 22822
rect 21212 22820 21236 22822
rect 21292 22820 21316 22822
rect 21372 22820 21378 22822
rect 21070 22811 21378 22820
rect 22020 22778 22048 23840
rect 22836 23452 22888 23458
rect 22836 23394 22888 23400
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 17958 22536 18014 22545
rect 17958 22471 18014 22480
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17696 22234 17724 22374
rect 18248 22234 18276 22578
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 18570 22332 18878 22341
rect 18570 22330 18576 22332
rect 18632 22330 18656 22332
rect 18712 22330 18736 22332
rect 18792 22330 18816 22332
rect 18872 22330 18878 22332
rect 18632 22278 18634 22330
rect 18814 22278 18816 22330
rect 18570 22276 18576 22278
rect 18632 22276 18656 22278
rect 18712 22276 18736 22278
rect 18792 22276 18816 22278
rect 18872 22276 18878 22278
rect 18570 22267 18878 22276
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15948 21554 15976 21898
rect 16316 21876 16344 22102
rect 16396 22024 16448 22030
rect 17316 22024 17368 22030
rect 16448 21984 16712 22012
rect 16396 21966 16448 21972
rect 16316 21848 16436 21876
rect 16070 21788 16378 21797
rect 16070 21786 16076 21788
rect 16132 21786 16156 21788
rect 16212 21786 16236 21788
rect 16292 21786 16316 21788
rect 16372 21786 16378 21788
rect 16132 21734 16134 21786
rect 16314 21734 16316 21786
rect 16070 21732 16076 21734
rect 16132 21732 16156 21734
rect 16212 21732 16236 21734
rect 16292 21732 16316 21734
rect 16372 21732 16378 21734
rect 16070 21723 16378 21732
rect 16408 21622 16436 21848
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15476 21412 15528 21418
rect 15476 21354 15528 21360
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15488 21146 15516 21354
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 14740 20936 14792 20942
rect 15290 20904 15346 20913
rect 14740 20878 14792 20884
rect 14752 20398 14780 20878
rect 15212 20862 15290 20890
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15120 20602 15148 20742
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15212 20534 15240 20862
rect 15290 20839 15346 20848
rect 15384 20868 15436 20874
rect 15580 20856 15608 21082
rect 15436 20828 15608 20856
rect 15384 20810 15436 20816
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 20262 14780 20334
rect 14740 20256 14792 20262
rect 14922 20224 14978 20233
rect 14792 20204 14922 20210
rect 14740 20198 14922 20204
rect 14752 20182 14922 20198
rect 14922 20159 14978 20168
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19514 14872 19790
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14752 18970 14780 19450
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14844 18834 14872 19110
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14752 18086 14780 18634
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14752 17542 14780 18022
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14844 17270 14872 18770
rect 15028 18630 15056 19382
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 18834 15240 19246
rect 15304 19242 15332 20470
rect 15672 20330 15700 21354
rect 15948 20924 15976 21490
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16120 20936 16172 20942
rect 15856 20896 16120 20924
rect 15750 20496 15806 20505
rect 15750 20431 15806 20440
rect 15764 20398 15792 20431
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15396 19310 15424 19790
rect 15488 19718 15516 20266
rect 15856 19786 15884 20896
rect 16316 20913 16344 21422
rect 16120 20878 16172 20884
rect 16302 20904 16358 20913
rect 16302 20839 16358 20848
rect 16408 20806 16436 21558
rect 16684 21554 16712 21984
rect 17316 21966 17368 21972
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 16764 21956 16816 21962
rect 16816 21916 16896 21944
rect 16764 21898 16816 21904
rect 16868 21554 16896 21916
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16488 20936 16540 20942
rect 16486 20904 16488 20913
rect 16540 20904 16542 20913
rect 16486 20839 16542 20848
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 15948 20602 15976 20742
rect 16070 20700 16378 20709
rect 16070 20698 16076 20700
rect 16132 20698 16156 20700
rect 16212 20698 16236 20700
rect 16292 20698 16316 20700
rect 16372 20698 16378 20700
rect 16132 20646 16134 20698
rect 16314 20646 16316 20698
rect 16070 20644 16076 20646
rect 16132 20644 16156 20646
rect 16212 20644 16236 20646
rect 16292 20644 16316 20646
rect 16372 20644 16378 20646
rect 16070 20635 16378 20644
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15948 20466 15976 20538
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16040 19922 16068 20538
rect 16592 20505 16620 20742
rect 16868 20602 16896 20810
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16578 20496 16634 20505
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16488 20460 16540 20466
rect 16946 20496 17002 20505
rect 16578 20431 16634 20440
rect 16672 20460 16724 20466
rect 16488 20402 16540 20408
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15936 19712 15988 19718
rect 16132 19700 16160 20402
rect 16316 20262 16344 20402
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16132 19672 16436 19700
rect 15936 19654 15988 19660
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18290 15056 18566
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15028 16998 15056 18226
rect 15304 18193 15332 18702
rect 15290 18184 15346 18193
rect 15108 18148 15160 18154
rect 15290 18119 15346 18128
rect 15108 18090 15160 18096
rect 15120 17746 15148 18090
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15212 17338 15240 17750
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15304 17066 15332 18119
rect 15488 17954 15516 19654
rect 15948 19514 15976 19654
rect 16070 19612 16378 19621
rect 16070 19610 16076 19612
rect 16132 19610 16156 19612
rect 16212 19610 16236 19612
rect 16292 19610 16316 19612
rect 16372 19610 16378 19612
rect 16132 19558 16134 19610
rect 16314 19558 16316 19610
rect 16070 19556 16076 19558
rect 16132 19556 16156 19558
rect 16212 19556 16236 19558
rect 16292 19556 16316 19558
rect 16372 19556 16378 19558
rect 16070 19547 16378 19556
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15580 18834 15608 19314
rect 15764 19174 15792 19314
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18834 15792 19110
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 16224 18766 16252 19246
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 15660 18624 15712 18630
rect 16028 18624 16080 18630
rect 15660 18566 15712 18572
rect 15948 18584 16028 18612
rect 15672 18306 15700 18566
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15856 18306 15884 18362
rect 15948 18358 15976 18584
rect 16028 18566 16080 18572
rect 16070 18524 16378 18533
rect 16070 18522 16076 18524
rect 16132 18522 16156 18524
rect 16212 18522 16236 18524
rect 16292 18522 16316 18524
rect 16372 18522 16378 18524
rect 16132 18470 16134 18522
rect 16314 18470 16316 18522
rect 16070 18468 16076 18470
rect 16132 18468 16156 18470
rect 16212 18468 16236 18470
rect 16292 18468 16316 18470
rect 16372 18468 16378 18470
rect 16070 18459 16378 18468
rect 15672 18278 15884 18306
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15488 17926 15608 17954
rect 15580 17202 15608 17926
rect 15856 17746 15884 18158
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17746 16068 18022
rect 16316 17882 16344 18226
rect 16408 17921 16436 19672
rect 16500 18766 16528 20402
rect 16592 19922 16620 20431
rect 16724 20420 16804 20448
rect 16946 20431 16948 20440
rect 16672 20402 16724 20408
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16684 20097 16712 20266
rect 16670 20088 16726 20097
rect 16670 20023 16726 20032
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19514 16620 19858
rect 16776 19718 16804 20420
rect 17000 20431 17002 20440
rect 16948 20402 17000 20408
rect 16960 19854 16988 20402
rect 17052 20233 17080 21830
rect 17328 21457 17356 21966
rect 17314 21448 17370 21457
rect 17314 21383 17370 21392
rect 17130 20768 17186 20777
rect 17328 20754 17356 21383
rect 17512 21321 17540 21966
rect 17696 21554 17724 22170
rect 19536 22166 19564 22374
rect 19720 22234 19748 22578
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 19524 22160 19576 22166
rect 19524 22102 19576 22108
rect 17868 22024 17920 22030
rect 18696 22024 18748 22030
rect 17868 21966 17920 21972
rect 18326 21992 18382 22001
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17498 21312 17554 21321
rect 17498 21247 17554 21256
rect 17406 20904 17462 20913
rect 17406 20839 17408 20848
rect 17460 20839 17462 20848
rect 17408 20810 17460 20816
rect 17512 20777 17540 21247
rect 17696 21146 17724 21490
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17880 21049 17908 21966
rect 18696 21966 18748 21972
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19156 22024 19208 22030
rect 19156 21966 19208 21972
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18326 21927 18328 21936
rect 18380 21927 18382 21936
rect 18328 21898 18380 21904
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18052 21480 18104 21486
rect 18156 21457 18184 21830
rect 18248 21622 18276 21830
rect 18708 21690 18736 21966
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18800 21690 18828 21898
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18972 21480 19024 21486
rect 18052 21422 18104 21428
rect 18142 21448 18198 21457
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17866 21040 17922 21049
rect 17866 20975 17922 20984
rect 17776 20800 17828 20806
rect 17186 20726 17356 20754
rect 17498 20768 17554 20777
rect 17130 20703 17186 20712
rect 17776 20742 17828 20748
rect 17498 20703 17554 20712
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17038 20224 17094 20233
rect 17038 20159 17094 20168
rect 16948 19848 17000 19854
rect 16868 19808 16948 19836
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16776 19446 16804 19654
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18426 16528 18702
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16684 18358 16712 19110
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18358 16804 18566
rect 16580 18352 16632 18358
rect 16486 18320 16542 18329
rect 16580 18294 16632 18300
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16486 18255 16488 18264
rect 16540 18255 16542 18264
rect 16488 18226 16540 18232
rect 16592 18057 16620 18294
rect 16578 18048 16634 18057
rect 16578 17983 16634 17992
rect 16394 17912 16450 17921
rect 16304 17876 16356 17882
rect 16394 17847 16450 17856
rect 16304 17818 16356 17824
rect 16394 17776 16450 17785
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 16028 17740 16080 17746
rect 16592 17762 16620 17983
rect 16764 17808 16816 17814
rect 16592 17734 16712 17762
rect 16764 17750 16816 17756
rect 16394 17711 16450 17720
rect 16028 17682 16080 17688
rect 16408 17678 16436 17711
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16070 17436 16378 17445
rect 16070 17434 16076 17436
rect 16132 17434 16156 17436
rect 16212 17434 16236 17436
rect 16292 17434 16316 17436
rect 16372 17434 16378 17436
rect 16132 17382 16134 17434
rect 16314 17382 16316 17434
rect 16070 17380 16076 17382
rect 16132 17380 16156 17382
rect 16212 17380 16236 17382
rect 16292 17380 16316 17382
rect 16372 17380 16378 17382
rect 16070 17371 16378 17380
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15580 17066 15608 17138
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15304 16250 15332 16594
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15488 16114 15516 16934
rect 15580 16114 15608 17002
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15570 14780 15982
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14752 15473 14780 15506
rect 14832 15496 14884 15502
rect 14738 15464 14794 15473
rect 14832 15438 14884 15444
rect 15198 15464 15254 15473
rect 14738 15399 14794 15408
rect 14844 15162 14872 15438
rect 14924 15428 14976 15434
rect 15198 15399 15254 15408
rect 15660 15428 15712 15434
rect 14924 15370 14976 15376
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14936 14822 14964 15370
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14752 14006 14780 14282
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14844 13870 14872 14418
rect 15120 14006 15148 14486
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 12434 14872 13806
rect 14752 12406 14872 12434
rect 14752 12306 14780 12406
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15028 11694 15056 12106
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 15028 11150 15056 11630
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14660 10628 14780 10656
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14568 10062 14596 10406
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 14200 9722 14228 9930
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14004 9376 14056 9382
rect 13648 9336 13952 9364
rect 13570 9276 13878 9285
rect 13570 9274 13576 9276
rect 13632 9274 13656 9276
rect 13712 9274 13736 9276
rect 13792 9274 13816 9276
rect 13872 9274 13878 9276
rect 13632 9222 13634 9274
rect 13814 9222 13816 9274
rect 13570 9220 13576 9222
rect 13632 9220 13656 9222
rect 13712 9220 13736 9222
rect 13792 9220 13816 9222
rect 13872 9220 13878 9222
rect 13570 9211 13878 9220
rect 13924 9160 13952 9336
rect 14004 9318 14056 9324
rect 13464 9132 13676 9160
rect 13360 9114 13412 9120
rect 13542 9072 13598 9081
rect 13452 9036 13504 9042
rect 13542 9007 13598 9016
rect 13452 8978 13504 8984
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13136 8520 13216 8548
rect 13084 8502 13136 8508
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7954 13216 8230
rect 13372 8090 13400 8910
rect 13464 8566 13492 8978
rect 13556 8906 13584 9007
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13648 8566 13676 9132
rect 13740 9132 13952 9160
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13648 8430 13676 8502
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13740 8276 13768 9132
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8945 13860 8978
rect 14016 8974 14044 9318
rect 14200 9110 14228 9658
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14004 8968 14056 8974
rect 13818 8936 13874 8945
rect 14004 8910 14056 8916
rect 13818 8871 13874 8880
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14188 8424 14240 8430
rect 14476 8412 14504 8774
rect 14240 8384 14504 8412
rect 14188 8366 14240 8372
rect 13464 8248 13768 8276
rect 14280 8288 14332 8294
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11900 7002 11928 7482
rect 12544 7206 12572 7686
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 12544 6730 12572 7142
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 13096 6662 13124 7210
rect 13188 7206 13216 7754
rect 13464 7290 13492 8248
rect 14280 8230 14332 8236
rect 13570 8188 13878 8197
rect 13570 8186 13576 8188
rect 13632 8186 13656 8188
rect 13712 8186 13736 8188
rect 13792 8186 13816 8188
rect 13872 8186 13878 8188
rect 13632 8134 13634 8186
rect 13814 8134 13816 8186
rect 13570 8132 13576 8134
rect 13632 8132 13656 8134
rect 13712 8132 13736 8134
rect 13792 8132 13816 8134
rect 13872 8132 13878 8134
rect 13570 8123 13878 8132
rect 14292 7954 14320 8230
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14476 7818 14504 8384
rect 14752 8362 14780 10628
rect 15028 10044 15056 11086
rect 15106 10976 15162 10985
rect 15106 10911 15162 10920
rect 15120 10742 15148 10911
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15120 10266 15148 10678
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15108 10056 15160 10062
rect 15028 10016 15108 10044
rect 15108 9998 15160 10004
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15028 9450 15056 9862
rect 15120 9722 15148 9998
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 9178 15056 9386
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 8838 15056 9114
rect 15212 9042 15240 15399
rect 15660 15370 15712 15376
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15396 14482 15424 15302
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15672 14346 15700 15370
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15764 14618 15792 14894
rect 15856 14822 15884 17138
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16114 15976 16934
rect 16316 16794 16344 17070
rect 16408 17066 16436 17614
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16500 16794 16528 17478
rect 16592 17202 16620 17614
rect 16684 17338 16712 17734
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16304 16788 16356 16794
rect 16488 16788 16540 16794
rect 16356 16748 16436 16776
rect 16304 16730 16356 16736
rect 16070 16348 16378 16357
rect 16070 16346 16076 16348
rect 16132 16346 16156 16348
rect 16212 16346 16236 16348
rect 16292 16346 16316 16348
rect 16372 16346 16378 16348
rect 16132 16294 16134 16346
rect 16314 16294 16316 16346
rect 16070 16292 16076 16294
rect 16132 16292 16156 16294
rect 16212 16292 16236 16294
rect 16292 16292 16316 16294
rect 16372 16292 16378 16294
rect 16070 16283 16378 16292
rect 16408 16250 16436 16748
rect 16488 16730 16540 16736
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16210 16144 16266 16153
rect 16132 16114 16210 16130
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 16120 16108 16210 16114
rect 16172 16102 16210 16108
rect 16210 16079 16266 16088
rect 16304 16108 16356 16114
rect 16120 16050 16172 16056
rect 16356 16068 16436 16096
rect 16304 16050 16356 16056
rect 16070 15260 16378 15269
rect 16070 15258 16076 15260
rect 16132 15258 16156 15260
rect 16212 15258 16236 15260
rect 16292 15258 16316 15260
rect 16372 15258 16378 15260
rect 16132 15206 16134 15258
rect 16314 15206 16316 15258
rect 16070 15204 16076 15206
rect 16132 15204 16156 15206
rect 16212 15204 16236 15206
rect 16292 15204 16316 15206
rect 16372 15204 16378 15206
rect 16070 15195 16378 15204
rect 16302 15056 16358 15065
rect 16224 15026 16302 15042
rect 16212 15020 16302 15026
rect 16264 15014 16302 15020
rect 16302 14991 16358 15000
rect 16212 14962 16264 14968
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 16408 14550 16436 16068
rect 16500 16046 16528 16730
rect 16592 16114 16620 17138
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16684 15978 16712 17274
rect 16776 17134 16804 17750
rect 16868 17746 16896 19808
rect 16948 19790 17000 19796
rect 17052 19446 17080 20159
rect 17222 19952 17278 19961
rect 17222 19887 17278 19896
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16960 18834 16988 19314
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17144 18714 17172 19790
rect 17236 19417 17264 19887
rect 17420 19514 17448 20402
rect 17788 20398 17816 20742
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17590 19952 17646 19961
rect 17590 19887 17592 19896
rect 17644 19887 17646 19896
rect 17592 19858 17644 19864
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17696 19446 17724 20334
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17592 19440 17644 19446
rect 17222 19408 17278 19417
rect 17592 19382 17644 19388
rect 17684 19440 17736 19446
rect 17684 19382 17736 19388
rect 17222 19343 17278 19352
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18766 17264 19246
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 16960 18686 17172 18714
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 16960 17814 16988 18686
rect 17328 18358 17356 19110
rect 17512 18766 17540 19314
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17132 18352 17184 18358
rect 17038 18320 17094 18329
rect 17132 18294 17184 18300
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17038 18255 17094 18264
rect 17052 18154 17080 18255
rect 17144 18193 17172 18294
rect 17130 18184 17186 18193
rect 17040 18148 17092 18154
rect 17130 18119 17186 18128
rect 17040 18090 17092 18096
rect 17132 18080 17184 18086
rect 17316 18080 17368 18086
rect 17132 18022 17184 18028
rect 17314 18048 17316 18057
rect 17368 18048 17370 18057
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17144 17678 17172 18022
rect 17314 17983 17370 17992
rect 17328 17746 17356 17983
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16776 15978 16804 17070
rect 16868 16250 16896 17546
rect 17052 17338 17080 17546
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16960 16182 16988 17138
rect 17052 16794 17080 17138
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17144 16232 17172 17002
rect 17224 16244 17276 16250
rect 17144 16204 17224 16232
rect 17224 16186 17276 16192
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16684 15688 16712 15914
rect 16764 15700 16816 15706
rect 16684 15660 16764 15688
rect 16764 15642 16816 15648
rect 16868 15638 16896 16050
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15026 16528 15302
rect 16868 15094 16896 15574
rect 16856 15088 16908 15094
rect 16856 15030 16908 15036
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12646 15332 13262
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12238 15332 12582
rect 15488 12238 15516 12718
rect 15580 12238 15608 13670
rect 15672 13462 15700 14282
rect 16070 14172 16378 14181
rect 16070 14170 16076 14172
rect 16132 14170 16156 14172
rect 16212 14170 16236 14172
rect 16292 14170 16316 14172
rect 16372 14170 16378 14172
rect 16132 14118 16134 14170
rect 16314 14118 16316 14170
rect 16070 14116 16076 14118
rect 16132 14116 16156 14118
rect 16212 14116 16236 14118
rect 16292 14116 16316 14118
rect 16372 14116 16378 14118
rect 16070 14107 16378 14116
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15764 11898 15792 13874
rect 16684 13870 16712 14758
rect 16868 14482 16896 14894
rect 16960 14618 16988 15846
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17052 14822 17080 15642
rect 17236 15366 17264 16186
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17132 15088 17184 15094
rect 17236 15076 17264 15302
rect 17184 15048 17264 15076
rect 17132 15030 17184 15036
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 14346 16896 14418
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 17328 13938 17356 17478
rect 17420 17184 17448 18566
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 18193 17540 18226
rect 17498 18184 17554 18193
rect 17498 18119 17554 18128
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17512 17678 17540 18022
rect 17604 17678 17632 19382
rect 17696 19310 17724 19382
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17788 19174 17816 19790
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17880 19122 17908 20975
rect 17972 19242 18000 21286
rect 18064 20913 18092 21422
rect 18972 21422 19024 21428
rect 18142 21383 18198 21392
rect 18570 21244 18878 21253
rect 18570 21242 18576 21244
rect 18632 21242 18656 21244
rect 18712 21242 18736 21244
rect 18792 21242 18816 21244
rect 18872 21242 18878 21244
rect 18632 21190 18634 21242
rect 18814 21190 18816 21242
rect 18570 21188 18576 21190
rect 18632 21188 18656 21190
rect 18712 21188 18736 21190
rect 18792 21188 18816 21190
rect 18872 21188 18878 21190
rect 18234 21176 18290 21185
rect 18570 21179 18878 21188
rect 18984 21185 19012 21422
rect 18234 21111 18290 21120
rect 18970 21176 19026 21185
rect 18970 21111 19026 21120
rect 18248 20913 18276 21111
rect 19076 21049 19104 21966
rect 19062 21040 19118 21049
rect 19062 20975 19118 20984
rect 18972 20936 19024 20942
rect 18050 20904 18106 20913
rect 18050 20839 18106 20848
rect 18234 20904 18290 20913
rect 18972 20878 19024 20884
rect 18234 20839 18290 20848
rect 18328 20800 18380 20806
rect 18064 20760 18328 20788
rect 18064 20058 18092 20760
rect 18328 20742 18380 20748
rect 18788 20596 18840 20602
rect 18156 20556 18644 20584
rect 18156 20466 18184 20556
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18328 20460 18380 20466
rect 18512 20460 18564 20466
rect 18328 20402 18380 20408
rect 18432 20420 18512 20448
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18064 19844 18092 19994
rect 18052 19838 18104 19844
rect 18052 19780 18104 19786
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17880 19094 18000 19122
rect 17868 18760 17920 18766
rect 17972 18737 18000 19094
rect 18064 18766 18092 19780
rect 18156 19718 18184 20198
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18248 19514 18276 20402
rect 18340 19922 18368 20402
rect 18432 20058 18460 20420
rect 18512 20402 18564 20408
rect 18616 20262 18644 20556
rect 18984 20584 19012 20878
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 19076 20602 19104 20742
rect 19168 20602 19196 21966
rect 18840 20556 19012 20584
rect 19064 20596 19116 20602
rect 18788 20538 18840 20544
rect 19064 20538 19116 20544
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19260 20482 19288 21966
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19076 20454 19288 20482
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18570 20156 18878 20165
rect 18570 20154 18576 20156
rect 18632 20154 18656 20156
rect 18712 20154 18736 20156
rect 18792 20154 18816 20156
rect 18872 20154 18878 20156
rect 18632 20102 18634 20154
rect 18814 20102 18816 20154
rect 18570 20100 18576 20102
rect 18632 20100 18656 20102
rect 18712 20100 18736 20102
rect 18792 20100 18816 20102
rect 18872 20100 18878 20102
rect 18570 20091 18878 20100
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18340 19689 18368 19722
rect 18326 19680 18382 19689
rect 18326 19615 18382 19624
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18236 18896 18288 18902
rect 18236 18838 18288 18844
rect 18052 18760 18104 18766
rect 17868 18702 17920 18708
rect 17958 18728 18014 18737
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17696 17746 17724 18226
rect 17774 18184 17830 18193
rect 17880 18154 17908 18702
rect 18052 18702 18104 18708
rect 17958 18663 18014 18672
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18426 18000 18566
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17958 18320 18014 18329
rect 17958 18255 17960 18264
rect 18012 18255 18014 18264
rect 17960 18226 18012 18232
rect 17774 18119 17830 18128
rect 17868 18148 17920 18154
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17500 17196 17552 17202
rect 17420 17156 17500 17184
rect 17788 17184 17816 18119
rect 17868 18090 17920 18096
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17958 17912 18014 17921
rect 17958 17847 17960 17856
rect 18012 17847 18014 17856
rect 17960 17818 18012 17824
rect 18156 17678 18184 18022
rect 18248 17785 18276 18838
rect 18340 18834 18368 19110
rect 18432 18970 18460 19994
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 19446 18736 19858
rect 18984 19786 19012 20402
rect 19076 20262 19104 20454
rect 19352 20398 19380 21830
rect 19444 21690 19472 21830
rect 19536 21729 19564 22102
rect 20088 22094 20116 22442
rect 20272 22234 20300 22578
rect 21548 22500 21600 22506
rect 21548 22442 21600 22448
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20088 22066 20208 22094
rect 20180 22030 20208 22066
rect 21560 22030 21588 22442
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21652 22030 21680 22374
rect 20168 22024 20220 22030
rect 19798 21992 19854 22001
rect 20168 21966 20220 21972
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 19798 21927 19854 21936
rect 19812 21894 19840 21927
rect 20548 21916 21036 21944
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19892 21888 19944 21894
rect 20444 21888 20496 21894
rect 19892 21830 19944 21836
rect 20258 21856 20314 21865
rect 19522 21720 19578 21729
rect 19432 21684 19484 21690
rect 19522 21655 19578 21664
rect 19432 21626 19484 21632
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19076 20058 19104 20198
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 19064 19780 19116 19786
rect 19064 19722 19116 19728
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18984 19378 19012 19722
rect 19076 19689 19104 19722
rect 19062 19680 19118 19689
rect 19062 19615 19118 19624
rect 19168 19514 19196 20266
rect 19444 19961 19472 21626
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19524 21072 19576 21078
rect 19522 21040 19524 21049
rect 19576 21040 19578 21049
rect 19522 20975 19578 20984
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19536 20398 19564 20878
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19430 19952 19486 19961
rect 19536 19922 19564 20334
rect 19430 19887 19486 19896
rect 19524 19916 19576 19922
rect 19444 19854 19472 19887
rect 19524 19858 19576 19864
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19536 19514 19564 19654
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 18570 19068 18878 19077
rect 18570 19066 18576 19068
rect 18632 19066 18656 19068
rect 18712 19066 18736 19068
rect 18792 19066 18816 19068
rect 18872 19066 18878 19068
rect 18632 19014 18634 19066
rect 18814 19014 18816 19066
rect 18570 19012 18576 19014
rect 18632 19012 18656 19014
rect 18712 19012 18736 19014
rect 18792 19012 18816 19014
rect 18872 19012 18878 19014
rect 18570 19003 18878 19012
rect 19444 18970 19472 19246
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19062 18728 19118 18737
rect 18570 17980 18878 17989
rect 18570 17978 18576 17980
rect 18632 17978 18656 17980
rect 18712 17978 18736 17980
rect 18792 17978 18816 17980
rect 18872 17978 18878 17980
rect 18632 17926 18634 17978
rect 18814 17926 18816 17978
rect 18570 17924 18576 17926
rect 18632 17924 18656 17926
rect 18712 17924 18736 17926
rect 18792 17924 18816 17926
rect 18872 17924 18878 17926
rect 18570 17915 18878 17924
rect 18234 17776 18290 17785
rect 18234 17711 18290 17720
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17868 17196 17920 17202
rect 17788 17156 17868 17184
rect 17500 17138 17552 17144
rect 17868 17138 17920 17144
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16658 17448 16934
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17512 15094 17540 17138
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16658 17724 16934
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17604 16114 17632 16186
rect 17696 16114 17724 16594
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17604 15978 17632 16050
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17788 15502 17816 16050
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 13297 16068 13330
rect 16500 13326 16528 13670
rect 16488 13320 16540 13326
rect 16026 13288 16082 13297
rect 16488 13262 16540 13268
rect 16026 13223 16082 13232
rect 16070 13084 16378 13093
rect 16070 13082 16076 13084
rect 16132 13082 16156 13084
rect 16212 13082 16236 13084
rect 16292 13082 16316 13084
rect 16372 13082 16378 13084
rect 16132 13030 16134 13082
rect 16314 13030 16316 13082
rect 16070 13028 16076 13030
rect 16132 13028 16156 13030
rect 16212 13028 16236 13030
rect 16292 13028 16316 13030
rect 16372 13028 16378 13030
rect 16070 13019 16378 13028
rect 16500 12850 16528 13262
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16592 12434 16620 13806
rect 16960 12986 16988 13806
rect 17052 13530 17080 13806
rect 17604 13734 17632 14758
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17604 12850 17632 13670
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17132 12436 17184 12442
rect 16592 12406 16712 12434
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16070 11996 16378 12005
rect 16070 11994 16076 11996
rect 16132 11994 16156 11996
rect 16212 11994 16236 11996
rect 16292 11994 16316 11996
rect 16372 11994 16378 11996
rect 16132 11942 16134 11994
rect 16314 11942 16316 11994
rect 16070 11940 16076 11942
rect 16132 11940 16156 11942
rect 16212 11940 16236 11942
rect 16292 11940 16316 11942
rect 16372 11940 16378 11942
rect 16070 11931 16378 11940
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 11082 15700 11494
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15672 10538 15700 11018
rect 15764 10674 15792 11698
rect 16592 11694 16620 12038
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 15856 11082 15884 11630
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15856 10470 15884 11018
rect 15948 10742 15976 11494
rect 16070 10908 16378 10917
rect 16070 10906 16076 10908
rect 16132 10906 16156 10908
rect 16212 10906 16236 10908
rect 16292 10906 16316 10908
rect 16372 10906 16378 10908
rect 16132 10854 16134 10906
rect 16314 10854 16316 10906
rect 16070 10852 16076 10854
rect 16132 10852 16156 10854
rect 16212 10852 16236 10854
rect 16292 10852 16316 10854
rect 16372 10852 16378 10854
rect 16070 10843 16378 10852
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 15856 9994 15884 10406
rect 16592 10266 16620 10406
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16684 10062 16712 12406
rect 17132 12378 17184 12384
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16868 11898 16896 12310
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16960 11354 16988 11698
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16868 10742 16896 10950
rect 17144 10810 17172 12378
rect 17408 12368 17460 12374
rect 17406 12336 17408 12345
rect 17460 12336 17462 12345
rect 17696 12306 17724 14350
rect 17788 14278 17816 14554
rect 17880 14346 17908 17138
rect 18156 16590 18184 17614
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17338 18920 17478
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16046 18184 16526
rect 18248 16153 18276 17138
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16454 18368 16934
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18432 16182 18460 17002
rect 18570 16892 18878 16901
rect 18570 16890 18576 16892
rect 18632 16890 18656 16892
rect 18712 16890 18736 16892
rect 18792 16890 18816 16892
rect 18872 16890 18878 16892
rect 18632 16838 18634 16890
rect 18814 16838 18816 16890
rect 18570 16836 18576 16838
rect 18632 16836 18656 16838
rect 18712 16836 18736 16838
rect 18792 16836 18816 16838
rect 18872 16836 18878 16838
rect 18570 16827 18878 16836
rect 18984 16561 19012 18702
rect 19352 18714 19380 18906
rect 19430 18728 19486 18737
rect 19352 18686 19430 18714
rect 19062 18663 19118 18672
rect 19430 18663 19486 18672
rect 18970 16552 19026 16561
rect 18970 16487 19026 16496
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16182 18552 16390
rect 18420 16176 18472 16182
rect 18234 16144 18290 16153
rect 18420 16118 18472 16124
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18234 16079 18290 16088
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 14958 18000 15438
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18156 14822 18184 15982
rect 18248 15910 18276 16079
rect 18524 16028 18552 16118
rect 18432 16000 18552 16028
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18248 15162 18276 15846
rect 18432 15366 18460 16000
rect 18570 15804 18878 15813
rect 18570 15802 18576 15804
rect 18632 15802 18656 15804
rect 18712 15802 18736 15804
rect 18792 15802 18816 15804
rect 18872 15802 18878 15804
rect 18632 15750 18634 15802
rect 18814 15750 18816 15802
rect 18570 15748 18576 15750
rect 18632 15748 18656 15750
rect 18712 15748 18736 15750
rect 18792 15748 18816 15750
rect 18872 15748 18878 15750
rect 18570 15739 18878 15748
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18432 14890 18460 15302
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18432 14618 18460 14826
rect 18800 14822 18828 15302
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18570 14716 18878 14725
rect 18570 14714 18576 14716
rect 18632 14714 18656 14716
rect 18712 14714 18736 14716
rect 18792 14714 18816 14716
rect 18872 14714 18878 14716
rect 18632 14662 18634 14714
rect 18814 14662 18816 14714
rect 18570 14660 18576 14662
rect 18632 14660 18656 14662
rect 18712 14660 18736 14662
rect 18792 14660 18816 14662
rect 18872 14660 18878 14662
rect 18570 14651 18878 14660
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18708 14414 18736 14554
rect 18970 14512 19026 14521
rect 19076 14498 19104 18663
rect 19628 18426 19656 21422
rect 19720 20534 19748 21830
rect 19812 20777 19840 21830
rect 19904 21690 19932 21830
rect 20444 21830 20496 21836
rect 20258 21791 20314 21800
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19798 20768 19854 20777
rect 19798 20703 19854 20712
rect 19904 20602 19932 21490
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19996 21350 20024 21422
rect 20180 21418 20208 21626
rect 20272 21457 20300 21791
rect 20456 21486 20484 21830
rect 20548 21554 20576 21916
rect 20640 21814 20944 21842
rect 20640 21690 20668 21814
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20444 21480 20496 21486
rect 20258 21448 20314 21457
rect 20168 21412 20220 21418
rect 20444 21422 20496 21428
rect 20258 21383 20314 21392
rect 20168 21354 20220 21360
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 19996 21078 20024 21286
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 20076 20868 20128 20874
rect 20076 20810 20128 20816
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19720 19689 19748 20470
rect 19996 20398 20024 20742
rect 20088 20505 20116 20810
rect 20074 20496 20130 20505
rect 20180 20466 20208 20810
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20074 20431 20130 20440
rect 20168 20460 20220 20466
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20088 20330 20116 20431
rect 20168 20402 20220 20408
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 19984 20256 20036 20262
rect 19904 20216 19984 20244
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19706 19680 19762 19689
rect 19706 19615 19762 19624
rect 19720 19378 19748 19615
rect 19812 19378 19840 19790
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19904 19242 19932 20216
rect 19984 20198 20036 20204
rect 20074 19952 20130 19961
rect 20074 19887 20130 19896
rect 20088 19786 20116 19887
rect 20272 19854 20300 20742
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19984 19372 20036 19378
rect 20088 19360 20116 19722
rect 20180 19514 20208 19722
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20272 19394 20300 19654
rect 20036 19332 20116 19360
rect 20180 19366 20300 19394
rect 19984 19314 20036 19320
rect 19892 19236 19944 19242
rect 19892 19178 19944 19184
rect 19892 18692 19944 18698
rect 19996 18680 20024 19314
rect 20180 18902 20208 19366
rect 20258 19000 20314 19009
rect 20258 18935 20314 18944
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20272 18766 20300 18935
rect 20364 18766 20392 21286
rect 20548 20806 20576 21286
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 19718 20484 20402
rect 20548 20398 20576 20742
rect 20640 20602 20668 21490
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20732 20398 20760 21558
rect 20824 20398 20852 21626
rect 20916 20806 20944 21814
rect 21008 21672 21036 21916
rect 21070 21788 21378 21797
rect 21070 21786 21076 21788
rect 21132 21786 21156 21788
rect 21212 21786 21236 21788
rect 21292 21786 21316 21788
rect 21372 21786 21378 21788
rect 21132 21734 21134 21786
rect 21314 21734 21316 21786
rect 21070 21732 21076 21734
rect 21132 21732 21156 21734
rect 21212 21732 21236 21734
rect 21292 21732 21316 21734
rect 21372 21732 21378 21734
rect 21070 21723 21378 21732
rect 21008 21644 21128 21672
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21008 20874 21036 21422
rect 21100 21418 21128 21644
rect 21560 21554 21588 21966
rect 21652 21622 21680 21966
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21178 21176 21234 21185
rect 21178 21111 21234 21120
rect 21192 20874 21220 21111
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 21070 20700 21378 20709
rect 21070 20698 21076 20700
rect 21132 20698 21156 20700
rect 21212 20698 21236 20700
rect 21292 20698 21316 20700
rect 21372 20698 21378 20700
rect 21132 20646 21134 20698
rect 21314 20646 21316 20698
rect 21070 20644 21076 20646
rect 21132 20644 21156 20646
rect 21212 20644 21236 20646
rect 21292 20644 21316 20646
rect 21372 20644 21378 20646
rect 21070 20635 21378 20644
rect 21468 20534 21496 21490
rect 21560 20924 21588 21490
rect 21652 21185 21680 21558
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21638 21176 21694 21185
rect 21638 21111 21694 21120
rect 21744 21078 21772 21286
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 21732 20936 21784 20942
rect 21560 20896 21732 20924
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20444 19712 20496 19718
rect 20548 19689 20576 19926
rect 20640 19922 20668 20198
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20628 19712 20680 19718
rect 20444 19654 20496 19660
rect 20534 19680 20590 19689
rect 20628 19654 20680 19660
rect 20534 19615 20590 19624
rect 20536 19304 20588 19310
rect 20456 19264 20536 19292
rect 20456 18970 20484 19264
rect 20536 19246 20588 19252
rect 20640 19174 20668 19654
rect 20732 19514 20760 19790
rect 20824 19718 20852 20334
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 19944 18652 20024 18680
rect 20168 18692 20220 18698
rect 19892 18634 19944 18640
rect 20168 18634 20220 18640
rect 20180 18426 20208 18634
rect 19616 18420 19668 18426
rect 19444 18380 19616 18408
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19352 17954 19380 18294
rect 19260 17926 19380 17954
rect 19260 16504 19288 17926
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19352 17066 19380 17546
rect 19444 17542 19472 18380
rect 19616 18362 19668 18368
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 20168 18420 20220 18426
rect 20364 18408 20392 18702
rect 20640 18426 20668 19110
rect 20168 18362 20220 18368
rect 20272 18380 20392 18408
rect 20628 18420 20680 18426
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19536 17338 19564 17478
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19352 16969 19380 17002
rect 19338 16960 19394 16969
rect 19338 16895 19394 16904
rect 19340 16516 19392 16522
rect 19260 16476 19340 16504
rect 19340 16458 19392 16464
rect 19444 15706 19472 17206
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16658 19564 16934
rect 19628 16794 19656 17818
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19720 17377 19748 17682
rect 19798 17640 19854 17649
rect 19798 17575 19854 17584
rect 19706 17368 19762 17377
rect 19706 17303 19762 17312
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19720 16250 19748 17138
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19026 14470 19104 14498
rect 18970 14447 19026 14456
rect 19260 14414 19288 14554
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 18248 14006 18276 14350
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 13530 18000 13806
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12442 17816 12718
rect 17880 12442 17908 12922
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17406 12271 17462 12280
rect 17684 12300 17736 12306
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 17132 10600 17184 10606
rect 17236 10588 17264 11494
rect 17184 10560 17264 10588
rect 17132 10542 17184 10548
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16070 9820 16378 9829
rect 16070 9818 16076 9820
rect 16132 9818 16156 9820
rect 16212 9818 16236 9820
rect 16292 9818 16316 9820
rect 16372 9818 16378 9820
rect 16132 9766 16134 9818
rect 16314 9766 16316 9818
rect 16070 9764 16076 9766
rect 16132 9764 16156 9766
rect 16212 9764 16236 9766
rect 16292 9764 16316 9766
rect 16372 9764 16378 9766
rect 16070 9755 16378 9764
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15396 8838 15424 9454
rect 16592 8974 16620 9658
rect 16868 9586 16896 9862
rect 16960 9654 16988 9862
rect 17144 9722 17172 10542
rect 17420 10266 17448 12271
rect 17684 12242 17736 12248
rect 17696 12209 17724 12242
rect 17880 12238 17908 12378
rect 17868 12232 17920 12238
rect 17682 12200 17738 12209
rect 17868 12174 17920 12180
rect 17682 12135 17738 12144
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17512 10266 17540 10542
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16580 8968 16632 8974
rect 15842 8936 15898 8945
rect 16580 8910 16632 8916
rect 15842 8871 15898 8880
rect 15856 8838 15884 8871
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15120 8634 15148 8774
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14936 8090 14964 8230
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 7546 14504 7754
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13280 7262 13492 7290
rect 14648 7268 14700 7274
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 11070 6556 11378 6565
rect 11070 6554 11076 6556
rect 11132 6554 11156 6556
rect 11212 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11378 6556
rect 11132 6502 11134 6554
rect 11314 6502 11316 6554
rect 11070 6500 11076 6502
rect 11132 6500 11156 6502
rect 11212 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11378 6502
rect 11070 6491 11378 6500
rect 12636 6118 12664 6598
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 11808 5574 11836 6054
rect 13188 5914 13216 6122
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11070 5468 11378 5477
rect 11070 5466 11076 5468
rect 11132 5466 11156 5468
rect 11212 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11378 5468
rect 11132 5414 11134 5466
rect 11314 5414 11316 5466
rect 11070 5412 11076 5414
rect 11132 5412 11156 5414
rect 11212 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11378 5414
rect 11070 5403 11378 5412
rect 11532 5302 11560 5510
rect 11808 5370 11836 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 3602 10640 4626
rect 11532 4486 11560 5238
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11624 4554 11652 4966
rect 11808 4826 11836 5306
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 10704 3942 10732 4422
rect 11070 4380 11378 4389
rect 11070 4378 11076 4380
rect 11132 4378 11156 4380
rect 11212 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11378 4380
rect 11132 4326 11134 4378
rect 11314 4326 11316 4378
rect 11070 4324 11076 4326
rect 11132 4324 11156 4326
rect 11212 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11378 4326
rect 11070 4315 11378 4324
rect 11532 4078 11560 4422
rect 11716 4282 11744 4422
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 12084 4214 12112 4966
rect 12268 4826 12296 5170
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10192 3420 10272 3448
rect 10140 3402 10192 3408
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3176 10088 3334
rect 9876 3148 10088 3176
rect 9876 2514 9904 3148
rect 9956 3052 10008 3058
rect 10152 3040 10180 3402
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3194 10640 3334
rect 10600 3188 10652 3194
rect 10008 3012 10180 3040
rect 10428 3148 10600 3176
rect 9956 2994 10008 3000
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8588 1902 8616 2246
rect 9876 2106 9904 2450
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 8576 1896 8628 1902
rect 8576 1838 8628 1844
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 8116 1828 8168 1834
rect 8116 1770 8168 1776
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7760 1358 7788 1702
rect 8128 1562 8156 1770
rect 8944 1760 8996 1766
rect 8944 1702 8996 1708
rect 8570 1660 8878 1669
rect 8570 1658 8576 1660
rect 8632 1658 8656 1660
rect 8712 1658 8736 1660
rect 8792 1658 8816 1660
rect 8872 1658 8878 1660
rect 8632 1606 8634 1658
rect 8814 1606 8816 1658
rect 8570 1604 8576 1606
rect 8632 1604 8656 1606
rect 8712 1604 8736 1606
rect 8792 1604 8816 1606
rect 8872 1604 8878 1606
rect 8570 1595 8878 1604
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8956 1358 8984 1702
rect 9232 1562 9260 1838
rect 9968 1834 9996 2994
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10060 2106 10088 2382
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10336 2106 10364 2314
rect 10048 2100 10100 2106
rect 10048 2042 10100 2048
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9692 1358 9720 1702
rect 10060 1562 10088 2042
rect 10428 1970 10456 3148
rect 10600 3130 10652 3136
rect 10704 2774 10732 3878
rect 11256 3738 11284 3878
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 2990 11008 3538
rect 11532 3466 11560 4014
rect 12176 3738 12204 4422
rect 12544 4282 12572 5102
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11070 3292 11378 3301
rect 11070 3290 11076 3292
rect 11132 3290 11156 3292
rect 11212 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11378 3292
rect 11132 3238 11134 3290
rect 11314 3238 11316 3290
rect 11070 3236 11076 3238
rect 11132 3236 11156 3238
rect 11212 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11378 3238
rect 11070 3227 11378 3236
rect 11796 3120 11848 3126
rect 11334 3088 11390 3097
rect 11796 3062 11848 3068
rect 11334 3023 11336 3032
rect 11388 3023 11390 3032
rect 11336 2994 11388 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10520 2746 10732 2774
rect 10520 1970 10548 2746
rect 11348 2310 11376 2994
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11070 2204 11378 2213
rect 11070 2202 11076 2204
rect 11132 2202 11156 2204
rect 11212 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11378 2204
rect 11132 2150 11134 2202
rect 11314 2150 11316 2202
rect 11070 2148 11076 2150
rect 11132 2148 11156 2150
rect 11212 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11378 2150
rect 11070 2139 11378 2148
rect 11440 2038 11468 2790
rect 11808 2650 11836 3062
rect 11900 2990 11928 3402
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11808 2106 11836 2586
rect 11900 2446 11928 2586
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11900 2106 11928 2382
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 12176 1970 12204 3674
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 2854 12388 2926
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12360 2310 12388 2790
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 1970 12388 2246
rect 12452 2106 12480 2790
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 12164 1964 12216 1970
rect 12164 1906 12216 1912
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12440 1964 12492 1970
rect 12544 1952 12572 3878
rect 12636 2582 12664 5102
rect 12820 4486 12848 5782
rect 13188 5370 13216 5850
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13188 4622 13216 5306
rect 13280 5234 13308 7262
rect 14648 7210 14700 7216
rect 13570 7100 13878 7109
rect 13570 7098 13576 7100
rect 13632 7098 13656 7100
rect 13712 7098 13736 7100
rect 13792 7098 13816 7100
rect 13872 7098 13878 7100
rect 13632 7046 13634 7098
rect 13814 7046 13816 7098
rect 13570 7044 13576 7046
rect 13632 7044 13656 7046
rect 13712 7044 13736 7046
rect 13792 7044 13816 7046
rect 13872 7044 13878 7046
rect 13570 7035 13878 7044
rect 14660 6730 14688 7210
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 15028 6458 15056 8366
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15212 7410 15240 7754
rect 15304 7410 15332 8434
rect 15396 8294 15424 8774
rect 15948 8430 15976 8774
rect 16070 8732 16378 8741
rect 16070 8730 16076 8732
rect 16132 8730 16156 8732
rect 16212 8730 16236 8732
rect 16292 8730 16316 8732
rect 16372 8730 16378 8732
rect 16132 8678 16134 8730
rect 16314 8678 16316 8730
rect 16070 8676 16076 8678
rect 16132 8676 16156 8678
rect 16212 8676 16236 8678
rect 16292 8676 16316 8678
rect 16372 8676 16378 8678
rect 16070 8667 16378 8676
rect 16592 8566 16620 8910
rect 16868 8906 16896 9522
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 17236 8634 17264 9998
rect 17420 9382 17448 10066
rect 17696 9654 17724 11222
rect 17788 10810 17816 11222
rect 17880 11150 17908 12174
rect 17972 12102 18000 12922
rect 18156 12764 18184 13874
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 12918 18276 13670
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18236 12776 18288 12782
rect 18156 12736 18236 12764
rect 18236 12718 18288 12724
rect 18248 12238 18276 12718
rect 18340 12238 18368 14214
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 13410 18460 14010
rect 18708 14006 18736 14214
rect 18800 14074 18828 14350
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18570 13628 18878 13637
rect 18570 13626 18576 13628
rect 18632 13626 18656 13628
rect 18712 13626 18736 13628
rect 18792 13626 18816 13628
rect 18872 13626 18878 13628
rect 18632 13574 18634 13626
rect 18814 13574 18816 13626
rect 18570 13572 18576 13574
rect 18632 13572 18656 13574
rect 18712 13572 18736 13574
rect 18792 13572 18816 13574
rect 18872 13572 18878 13574
rect 18570 13563 18878 13572
rect 18696 13524 18748 13530
rect 18748 13484 18920 13512
rect 18696 13466 18748 13472
rect 18432 13394 18552 13410
rect 18432 13388 18564 13394
rect 18432 13382 18512 13388
rect 18512 13330 18564 13336
rect 18892 13326 18920 13484
rect 18984 13326 19012 14350
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18708 13190 18736 13262
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18696 13184 18748 13190
rect 18984 13172 19012 13262
rect 18696 13126 18748 13132
rect 18892 13144 19012 13172
rect 18432 12306 18460 13126
rect 18892 12782 18920 13144
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18570 12540 18878 12549
rect 18570 12538 18576 12540
rect 18632 12538 18656 12540
rect 18712 12538 18736 12540
rect 18792 12538 18816 12540
rect 18872 12538 18878 12540
rect 18632 12486 18634 12538
rect 18814 12486 18816 12538
rect 18570 12484 18576 12486
rect 18632 12484 18656 12486
rect 18712 12484 18736 12486
rect 18792 12484 18816 12486
rect 18872 12484 18878 12486
rect 18570 12475 18878 12484
rect 18880 12436 18932 12442
rect 18984 12424 19012 12718
rect 19076 12458 19104 14350
rect 19444 14346 19472 14758
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19168 13258 19196 13942
rect 19352 13546 19380 14282
rect 19352 13530 19472 13546
rect 19352 13524 19484 13530
rect 19352 13518 19432 13524
rect 19432 13466 19484 13472
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19168 12986 19196 13194
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19260 12782 19288 13194
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19076 12442 19109 12458
rect 18932 12396 19012 12424
rect 18880 12378 18932 12384
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18984 12238 19012 12396
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19352 12322 19380 13194
rect 19536 12696 19564 13262
rect 19628 12986 19656 14486
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 13802 19748 14350
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19616 12708 19668 12714
rect 19536 12668 19616 12696
rect 19616 12650 19668 12656
rect 19628 12458 19656 12650
rect 19720 12646 19748 13738
rect 19812 13297 19840 17575
rect 19904 17236 19932 18362
rect 20272 18290 20300 18380
rect 20628 18362 20680 18368
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20444 18284 20496 18290
rect 20496 18244 20576 18272
rect 20444 18226 20496 18232
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17882 20024 18022
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19996 17338 20024 17546
rect 20272 17338 20300 18226
rect 20364 17882 20392 18226
rect 20548 18170 20576 18244
rect 20732 18170 20760 19450
rect 20444 18148 20496 18154
rect 20548 18142 20760 18170
rect 20444 18090 20496 18096
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20456 17678 20484 18090
rect 20732 17864 20760 18142
rect 20824 18086 20852 19450
rect 20916 19310 20944 20198
rect 21284 20058 21312 20266
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21456 20052 21508 20058
rect 21560 20040 21588 20896
rect 21732 20878 21784 20884
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21744 20466 21772 20742
rect 21732 20460 21784 20466
rect 21732 20402 21784 20408
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21652 20058 21680 20198
rect 21508 20012 21588 20040
rect 21640 20052 21692 20058
rect 21456 19994 21508 20000
rect 21640 19994 21692 20000
rect 20994 19952 21050 19961
rect 20994 19887 20996 19896
rect 21048 19887 21050 19896
rect 20996 19858 21048 19864
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20916 18086 20944 19246
rect 21008 18358 21036 19858
rect 21744 19854 21772 20402
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21070 19612 21378 19621
rect 21070 19610 21076 19612
rect 21132 19610 21156 19612
rect 21212 19610 21236 19612
rect 21292 19610 21316 19612
rect 21372 19610 21378 19612
rect 21132 19558 21134 19610
rect 21314 19558 21316 19610
rect 21070 19556 21076 19558
rect 21132 19556 21156 19558
rect 21212 19556 21236 19558
rect 21292 19556 21316 19558
rect 21372 19556 21378 19558
rect 21070 19547 21378 19556
rect 21744 19446 21772 19790
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 19009 21220 19110
rect 21178 19000 21234 19009
rect 21178 18935 21234 18944
rect 21070 18524 21378 18533
rect 21070 18522 21076 18524
rect 21132 18522 21156 18524
rect 21212 18522 21236 18524
rect 21292 18522 21316 18524
rect 21372 18522 21378 18524
rect 21132 18470 21134 18522
rect 21314 18470 21316 18522
rect 21070 18468 21076 18470
rect 21132 18468 21156 18470
rect 21212 18468 21236 18470
rect 21292 18468 21316 18470
rect 21372 18468 21378 18470
rect 21070 18459 21378 18468
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21364 18284 21416 18290
rect 21468 18272 21496 19314
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21560 18630 21588 19110
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21560 18358 21588 18566
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21416 18244 21496 18272
rect 21364 18226 21416 18232
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20812 17876 20864 17882
rect 20732 17836 20812 17864
rect 20812 17818 20864 17824
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 21008 17678 21036 17750
rect 21192 17746 21220 18226
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19892 17230 19944 17236
rect 20364 17202 20392 17478
rect 20442 17368 20498 17377
rect 20640 17338 20668 17546
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20442 17303 20444 17312
rect 20496 17303 20498 17312
rect 20628 17332 20680 17338
rect 20444 17274 20496 17280
rect 20628 17274 20680 17280
rect 20352 17196 20404 17202
rect 19892 17172 19944 17178
rect 20272 17156 20352 17184
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19890 16960 19946 16969
rect 19890 16895 19946 16904
rect 19904 15978 19932 16895
rect 20180 16794 20208 17070
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20180 16114 20208 16390
rect 20272 16182 20300 17156
rect 20352 17138 20404 17144
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16522 20392 17002
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20456 16114 20484 17274
rect 21008 17202 21036 17478
rect 21070 17436 21378 17445
rect 21070 17434 21076 17436
rect 21132 17434 21156 17436
rect 21212 17434 21236 17436
rect 21292 17434 21316 17436
rect 21372 17434 21378 17436
rect 21132 17382 21134 17434
rect 21314 17382 21316 17434
rect 21070 17380 21076 17382
rect 21132 17380 21156 17382
rect 21212 17380 21236 17382
rect 21292 17380 21316 17382
rect 21372 17380 21378 17382
rect 21070 17371 21378 17380
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20902 17096 20958 17105
rect 20548 16969 20576 17070
rect 20902 17031 20904 17040
rect 20956 17031 20958 17040
rect 20904 17002 20956 17008
rect 20534 16960 20590 16969
rect 20534 16895 20590 16904
rect 20916 16674 20944 17002
rect 21008 16794 21036 17138
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20916 16646 21036 16674
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20824 16114 20852 16526
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19904 15502 19932 15914
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 20168 15428 20220 15434
rect 20220 15388 20300 15416
rect 20168 15370 20220 15376
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14550 19932 14758
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19904 14278 19932 14486
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19798 13288 19854 13297
rect 19798 13223 19854 13232
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19812 12850 19840 13126
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19628 12430 19748 12458
rect 19260 12294 19380 12322
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19260 12238 19288 12294
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 19064 12232 19116 12238
rect 19248 12232 19300 12238
rect 19064 12174 19116 12180
rect 19154 12200 19210 12209
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 18064 10266 18092 12106
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18420 12096 18472 12102
rect 18696 12096 18748 12102
rect 18420 12038 18472 12044
rect 18694 12064 18696 12073
rect 18748 12064 18750 12073
rect 18248 11830 18276 12038
rect 18432 11898 18460 12038
rect 18694 11999 18750 12008
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18248 10742 18276 11766
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18570 11452 18878 11461
rect 18570 11450 18576 11452
rect 18632 11450 18656 11452
rect 18712 11450 18736 11452
rect 18792 11450 18816 11452
rect 18872 11450 18878 11452
rect 18632 11398 18634 11450
rect 18814 11398 18816 11450
rect 18570 11396 18576 11398
rect 18632 11396 18656 11398
rect 18712 11396 18736 11398
rect 18792 11396 18816 11398
rect 18872 11396 18878 11398
rect 18570 11387 18878 11396
rect 18984 11014 19012 11494
rect 19076 11354 19104 12174
rect 19248 12174 19300 12180
rect 19154 12135 19156 12144
rect 19208 12135 19210 12144
rect 19156 12106 19208 12112
rect 19168 11898 19196 12106
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19444 11801 19472 12038
rect 19430 11792 19486 11801
rect 19430 11727 19486 11736
rect 19536 11694 19564 12310
rect 19720 12170 19748 12430
rect 19812 12434 19840 12786
rect 19904 12646 19932 14214
rect 19996 14074 20024 14962
rect 20088 14618 20116 14962
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20180 14414 20208 14758
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19996 12850 20024 13466
rect 20166 13424 20222 13433
rect 20166 13359 20222 13368
rect 20180 12889 20208 13359
rect 20166 12880 20222 12889
rect 19984 12844 20036 12850
rect 20166 12815 20168 12824
rect 19984 12786 20036 12792
rect 20220 12815 20222 12824
rect 20168 12786 20220 12792
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 20180 12481 20208 12786
rect 20166 12472 20222 12481
rect 19892 12436 19944 12442
rect 19812 12406 19856 12434
rect 19828 12356 19856 12406
rect 20166 12407 20222 12416
rect 19892 12378 19944 12384
rect 19812 12328 19856 12356
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19628 11812 19656 12106
rect 19708 11824 19760 11830
rect 19628 11784 19708 11812
rect 19708 11766 19760 11772
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19720 11370 19748 11766
rect 19812 11762 19840 12328
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19904 11744 19932 12378
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 11762 20208 12174
rect 19984 11756 20036 11762
rect 19904 11716 19984 11744
rect 19904 11626 19932 11716
rect 19984 11698 20036 11704
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 19982 11656 20038 11665
rect 19892 11620 19944 11626
rect 19982 11591 19984 11600
rect 19892 11562 19944 11568
rect 20036 11591 20038 11600
rect 19984 11562 20036 11568
rect 20180 11370 20208 11698
rect 20272 11626 20300 15388
rect 20456 15366 20484 16050
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15638 20852 15846
rect 20916 15706 20944 16526
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20732 15026 20760 15438
rect 20720 15020 20772 15026
rect 20824 15008 20852 15574
rect 21008 15434 21036 16646
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21284 16454 21312 16526
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21070 16348 21378 16357
rect 21070 16346 21076 16348
rect 21132 16346 21156 16348
rect 21212 16346 21236 16348
rect 21292 16346 21316 16348
rect 21372 16346 21378 16348
rect 21132 16294 21134 16346
rect 21314 16294 21316 16346
rect 21070 16292 21076 16294
rect 21132 16292 21156 16294
rect 21212 16292 21236 16294
rect 21292 16292 21316 16294
rect 21372 16292 21378 16294
rect 21070 16283 21378 16292
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15706 21128 15914
rect 21468 15706 21496 16526
rect 21560 16250 21588 18158
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21652 16998 21680 17478
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 20904 15020 20956 15026
rect 20824 14980 20904 15008
rect 20720 14962 20772 14968
rect 20904 14962 20956 14968
rect 21008 14906 21036 15370
rect 21070 15260 21378 15269
rect 21070 15258 21076 15260
rect 21132 15258 21156 15260
rect 21212 15258 21236 15260
rect 21292 15258 21316 15260
rect 21372 15258 21378 15260
rect 21132 15206 21134 15258
rect 21314 15206 21316 15258
rect 21070 15204 21076 15206
rect 21132 15204 21156 15206
rect 21212 15204 21236 15206
rect 21292 15204 21316 15206
rect 21372 15204 21378 15206
rect 21070 15195 21378 15204
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 20824 14878 21036 14906
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14618 20484 14758
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 13190 20392 14214
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20456 13002 20484 13670
rect 20364 12974 20484 13002
rect 20364 12442 20392 12974
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20364 12306 20392 12378
rect 20456 12345 20484 12854
rect 20442 12336 20498 12345
rect 20352 12300 20404 12306
rect 20442 12271 20498 12280
rect 20352 12242 20404 12248
rect 20352 11892 20404 11898
rect 20456 11880 20484 12271
rect 20404 11852 20484 11880
rect 20352 11834 20404 11840
rect 20548 11762 20576 13806
rect 20824 13433 20852 14878
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14006 21036 14758
rect 21192 14414 21220 14894
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21284 14346 21312 14554
rect 21468 14550 21496 14962
rect 21560 14618 21588 14962
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21468 14414 21496 14486
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21272 14340 21324 14346
rect 21324 14300 21404 14328
rect 21272 14282 21324 14288
rect 21376 14260 21404 14300
rect 21652 14260 21680 16934
rect 21730 16688 21786 16697
rect 21730 16623 21786 16632
rect 21744 16522 21772 16623
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21744 16182 21772 16458
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21376 14232 21680 14260
rect 21070 14172 21378 14181
rect 21070 14170 21076 14172
rect 21132 14170 21156 14172
rect 21212 14170 21236 14172
rect 21292 14170 21316 14172
rect 21372 14170 21378 14172
rect 21132 14118 21134 14170
rect 21314 14118 21316 14170
rect 21070 14116 21076 14118
rect 21132 14116 21156 14118
rect 21212 14116 21236 14118
rect 21292 14116 21316 14118
rect 21372 14116 21378 14118
rect 21070 14107 21378 14116
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20810 13424 20866 13433
rect 20810 13359 20866 13368
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20824 12782 20852 13126
rect 20916 12986 20944 13466
rect 21468 13240 21496 14232
rect 21546 13968 21602 13977
rect 21546 13903 21602 13912
rect 21560 13870 21588 13903
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21548 13252 21600 13258
rect 21468 13212 21548 13240
rect 21548 13194 21600 13200
rect 21070 13084 21378 13093
rect 21070 13082 21076 13084
rect 21132 13082 21156 13084
rect 21212 13082 21236 13084
rect 21292 13082 21316 13084
rect 21372 13082 21378 13084
rect 21132 13030 21134 13082
rect 21314 13030 21316 13082
rect 21070 13028 21076 13030
rect 21132 13028 21156 13030
rect 21212 13028 21236 13030
rect 21292 13028 21316 13030
rect 21372 13028 21378 13030
rect 21070 13019 21378 13028
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21560 12782 21588 13194
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 12238 20668 12582
rect 20824 12434 20852 12718
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20732 12406 20852 12434
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20628 12096 20680 12102
rect 20626 12064 20628 12073
rect 20680 12064 20682 12073
rect 20626 11999 20682 12008
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 19064 11348 19116 11354
rect 19720 11342 20208 11370
rect 19064 11290 19116 11296
rect 19062 11248 19118 11257
rect 19062 11183 19118 11192
rect 19340 11212 19392 11218
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18984 10810 19012 10950
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18570 10364 18878 10373
rect 18570 10362 18576 10364
rect 18632 10362 18656 10364
rect 18712 10362 18736 10364
rect 18792 10362 18816 10364
rect 18872 10362 18878 10364
rect 18632 10310 18634 10362
rect 18814 10310 18816 10362
rect 18570 10308 18576 10310
rect 18632 10308 18656 10310
rect 18712 10308 18736 10310
rect 18792 10308 18816 10310
rect 18872 10308 18878 10310
rect 18570 10299 18878 10308
rect 18052 10260 18104 10266
rect 18984 10248 19012 10746
rect 18052 10202 18104 10208
rect 18892 10220 19012 10248
rect 18892 10062 18920 10220
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 17776 10056 17828 10062
rect 18420 10056 18472 10062
rect 17828 10004 18092 10010
rect 17776 9998 18092 10004
rect 18420 9998 18472 10004
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 17788 9982 18092 9998
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15396 7886 15424 8230
rect 16040 7886 16068 8230
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 7206 15332 7346
rect 15396 7324 15424 7822
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15672 7342 15700 7686
rect 15856 7478 15884 7686
rect 16070 7644 16378 7653
rect 16070 7642 16076 7644
rect 16132 7642 16156 7644
rect 16212 7642 16236 7644
rect 16292 7642 16316 7644
rect 16372 7642 16378 7644
rect 16132 7590 16134 7642
rect 16314 7590 16316 7642
rect 16070 7588 16076 7590
rect 16132 7588 16156 7590
rect 16212 7588 16236 7590
rect 16292 7588 16316 7590
rect 16372 7588 16378 7590
rect 16070 7579 16378 7588
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 15568 7336 15620 7342
rect 15396 7296 15568 7324
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15120 7002 15148 7142
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15396 6730 15424 7296
rect 15568 7278 15620 7284
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15672 6730 15700 7278
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 13358 6352 13414 6361
rect 13358 6287 13414 6296
rect 15660 6316 15712 6322
rect 13372 5846 13400 6287
rect 15660 6258 15712 6264
rect 15568 6248 15620 6254
rect 13634 6216 13690 6225
rect 15568 6190 15620 6196
rect 13634 6151 13636 6160
rect 13688 6151 13690 6160
rect 13636 6122 13688 6128
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 13570 6012 13878 6021
rect 13570 6010 13576 6012
rect 13632 6010 13656 6012
rect 13712 6010 13736 6012
rect 13792 6010 13816 6012
rect 13872 6010 13878 6012
rect 13632 5958 13634 6010
rect 13814 5958 13816 6010
rect 13570 5956 13576 5958
rect 13632 5956 13656 5958
rect 13712 5956 13736 5958
rect 13792 5956 13816 5958
rect 13872 5956 13878 5958
rect 13570 5947 13878 5956
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13726 5264 13782 5273
rect 13268 5228 13320 5234
rect 13726 5199 13728 5208
rect 13268 5170 13320 5176
rect 13780 5199 13782 5208
rect 13728 5170 13780 5176
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12912 3534 12940 4082
rect 13004 3942 13032 4422
rect 13280 4078 13308 5170
rect 14002 5128 14058 5137
rect 14002 5063 14004 5072
rect 14056 5063 14058 5072
rect 14004 5034 14056 5040
rect 13570 4924 13878 4933
rect 13570 4922 13576 4924
rect 13632 4922 13656 4924
rect 13712 4922 13736 4924
rect 13792 4922 13816 4924
rect 13872 4922 13878 4924
rect 13632 4870 13634 4922
rect 13814 4870 13816 4922
rect 13570 4868 13576 4870
rect 13632 4868 13656 4870
rect 13712 4868 13736 4870
rect 13792 4868 13816 4870
rect 13872 4868 13878 4870
rect 13570 4859 13878 4868
rect 14108 4826 14136 6054
rect 14462 5944 14518 5953
rect 14372 5908 14424 5914
rect 14462 5879 14518 5888
rect 15200 5908 15252 5914
rect 14372 5850 14424 5856
rect 14278 5808 14334 5817
rect 14278 5743 14334 5752
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13280 3738 13308 4014
rect 13924 4010 13952 4694
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 4078 14044 4626
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 3194 13216 3334
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13372 2990 13400 3878
rect 13570 3836 13878 3845
rect 13570 3834 13576 3836
rect 13632 3834 13656 3836
rect 13712 3834 13736 3836
rect 13792 3834 13816 3836
rect 13872 3834 13878 3836
rect 13632 3782 13634 3834
rect 13814 3782 13816 3834
rect 13570 3780 13576 3782
rect 13632 3780 13656 3782
rect 13712 3780 13736 3782
rect 13792 3780 13816 3782
rect 13872 3780 13878 3782
rect 13570 3771 13878 3780
rect 13924 3534 13952 3946
rect 14016 3602 14044 4014
rect 14096 3936 14148 3942
rect 14200 3924 14228 5510
rect 14292 4282 14320 5743
rect 14384 5302 14412 5850
rect 14476 5846 14504 5879
rect 15200 5850 15252 5856
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14462 5672 14518 5681
rect 15212 5642 15240 5850
rect 15580 5778 15608 6190
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 14462 5607 14464 5616
rect 14516 5607 14518 5616
rect 14648 5636 14700 5642
rect 14464 5578 14516 5584
rect 14648 5578 14700 5584
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14660 5148 14688 5578
rect 14924 5568 14976 5574
rect 14844 5528 14924 5556
rect 14740 5160 14792 5166
rect 14660 5120 14740 5148
rect 14740 5102 14792 5108
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14384 4282 14412 4490
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14844 4185 14872 5528
rect 14924 5510 14976 5516
rect 15120 5370 15148 5578
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 14830 4176 14886 4185
rect 14464 4140 14516 4146
rect 15212 4146 15240 5578
rect 15580 5166 15608 5714
rect 15672 5234 15700 6258
rect 15764 5302 15792 6802
rect 15856 6662 15884 7142
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15948 6458 15976 7210
rect 16500 6798 16528 7754
rect 16684 7546 16712 8434
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7954 16804 8230
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16592 7002 16620 7414
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16776 6866 16804 7686
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 7002 17080 7142
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16070 6556 16378 6565
rect 16070 6554 16076 6556
rect 16132 6554 16156 6556
rect 16212 6554 16236 6556
rect 16292 6554 16316 6556
rect 16372 6554 16378 6556
rect 16132 6502 16134 6554
rect 16314 6502 16316 6554
rect 16070 6500 16076 6502
rect 16132 6500 16156 6502
rect 16212 6500 16236 6502
rect 16292 6500 16316 6502
rect 16372 6500 16378 6502
rect 16070 6491 16378 6500
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16500 6322 16528 6734
rect 16776 6730 16804 6802
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 17236 6662 17264 8434
rect 17328 7868 17356 8434
rect 17512 7886 17540 8842
rect 17972 8566 18000 9862
rect 18064 9654 18092 9982
rect 18432 9722 18460 9998
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18064 8634 18092 9590
rect 18984 9382 19012 10066
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18570 9276 18878 9285
rect 18570 9274 18576 9276
rect 18632 9274 18656 9276
rect 18712 9274 18736 9276
rect 18792 9274 18816 9276
rect 18872 9274 18878 9276
rect 18632 9222 18634 9274
rect 18814 9222 18816 9274
rect 18570 9220 18576 9222
rect 18632 9220 18656 9222
rect 18712 9220 18736 9222
rect 18792 9220 18816 9222
rect 18872 9220 18878 9222
rect 18570 9211 18878 9220
rect 18984 9042 19012 9318
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 18248 8090 18276 8978
rect 18512 8832 18564 8838
rect 18432 8792 18512 8820
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18432 7886 18460 8792
rect 18512 8774 18564 8780
rect 18570 8188 18878 8197
rect 18570 8186 18576 8188
rect 18632 8186 18656 8188
rect 18712 8186 18736 8188
rect 18792 8186 18816 8188
rect 18872 8186 18878 8188
rect 18632 8134 18634 8186
rect 18814 8134 18816 8186
rect 18570 8132 18576 8134
rect 18632 8132 18656 8134
rect 18712 8132 18736 8134
rect 18792 8132 18816 8134
rect 18872 8132 18878 8134
rect 18570 8123 18878 8132
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 17408 7880 17460 7886
rect 17328 7840 17408 7868
rect 17328 7002 17356 7840
rect 17408 7822 17460 7828
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17420 7410 17448 7686
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17420 6662 17448 7346
rect 17604 6798 17632 7482
rect 18064 7410 18092 7686
rect 18616 7478 18644 7890
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18892 7546 18920 7754
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 17684 7404 17736 7410
rect 17960 7404 18012 7410
rect 17684 7346 17736 7352
rect 17880 7364 17960 7392
rect 17696 6866 17724 7346
rect 17880 6934 17908 7364
rect 17960 7346 18012 7352
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 16580 6452 16632 6458
rect 16948 6452 17000 6458
rect 16580 6394 16632 6400
rect 16776 6412 16948 6440
rect 16592 6322 16620 6394
rect 16776 6322 16804 6412
rect 16948 6394 17000 6400
rect 17880 6390 17908 6870
rect 17972 6458 18000 6938
rect 18340 6798 18368 7142
rect 18570 7100 18878 7109
rect 18570 7098 18576 7100
rect 18632 7098 18656 7100
rect 18712 7098 18736 7100
rect 18792 7098 18816 7100
rect 18872 7098 18878 7100
rect 18632 7046 18634 7098
rect 18814 7046 18816 7098
rect 18570 7044 18576 7046
rect 18632 7044 18656 7046
rect 18712 7044 18736 7046
rect 18792 7044 18816 7046
rect 18872 7044 18878 7046
rect 18570 7035 18878 7044
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 16040 5914 16068 6258
rect 16120 6248 16172 6254
rect 16304 6248 16356 6254
rect 16120 6190 16172 6196
rect 16224 6208 16304 6236
rect 16132 6089 16160 6190
rect 16224 6118 16252 6208
rect 16304 6190 16356 6196
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16212 6112 16264 6118
rect 16118 6080 16174 6089
rect 16212 6054 16264 6060
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16118 6015 16174 6024
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16684 5710 16712 6054
rect 16776 5778 16804 6122
rect 16868 6089 16896 6258
rect 16854 6080 16910 6089
rect 16854 6015 16910 6024
rect 16960 5914 16988 6258
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15672 4554 15700 5170
rect 15856 4826 15884 5578
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16070 5468 16378 5477
rect 16070 5466 16076 5468
rect 16132 5466 16156 5468
rect 16212 5466 16236 5468
rect 16292 5466 16316 5468
rect 16372 5466 16378 5468
rect 16132 5414 16134 5466
rect 16314 5414 16316 5466
rect 16070 5412 16076 5414
rect 16132 5412 16156 5414
rect 16212 5412 16236 5414
rect 16292 5412 16316 5414
rect 16372 5412 16378 5414
rect 16070 5403 16378 5412
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15764 4282 15792 4558
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 14830 4111 14886 4120
rect 15200 4140 15252 4146
rect 14464 4082 14516 4088
rect 14148 3896 14228 3924
rect 14096 3878 14148 3884
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13570 2748 13878 2757
rect 13570 2746 13576 2748
rect 13632 2746 13656 2748
rect 13712 2746 13736 2748
rect 13792 2746 13816 2748
rect 13872 2746 13878 2748
rect 13632 2694 13634 2746
rect 13814 2694 13816 2746
rect 13570 2692 13576 2694
rect 13632 2692 13656 2694
rect 13712 2692 13736 2694
rect 13792 2692 13816 2694
rect 13872 2692 13878 2694
rect 13570 2683 13878 2692
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 14016 2446 14044 3334
rect 14108 3058 14136 3878
rect 14476 3194 14504 4082
rect 14844 3738 14872 4111
rect 15200 4082 15252 4088
rect 15856 3942 15884 4490
rect 15948 4214 15976 4694
rect 16040 4554 16068 5238
rect 16408 4826 16436 5510
rect 16500 5370 16528 5510
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16592 5302 16620 5510
rect 16776 5302 16804 5714
rect 17144 5658 17172 5850
rect 17512 5710 17540 6054
rect 17696 5914 17724 6258
rect 17774 5944 17830 5953
rect 17684 5908 17736 5914
rect 17774 5879 17776 5888
rect 17684 5850 17736 5856
rect 17828 5879 17830 5888
rect 17776 5850 17828 5856
rect 16868 5630 17172 5658
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 16868 5574 16896 5630
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 17222 5536 17278 5545
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16856 5160 16908 5166
rect 16776 5120 16856 5148
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16486 4720 16542 4729
rect 16486 4655 16542 4664
rect 16394 4584 16450 4593
rect 16028 4548 16080 4554
rect 16394 4519 16450 4528
rect 16028 4490 16080 4496
rect 16070 4380 16378 4389
rect 16070 4378 16076 4380
rect 16132 4378 16156 4380
rect 16212 4378 16236 4380
rect 16292 4378 16316 4380
rect 16372 4378 16378 4380
rect 16132 4326 16134 4378
rect 16314 4326 16316 4378
rect 16070 4324 16076 4326
rect 16132 4324 16156 4326
rect 16212 4324 16236 4326
rect 16292 4324 16316 4326
rect 16372 4324 16378 4326
rect 16070 4315 16378 4324
rect 15936 4208 15988 4214
rect 16408 4162 16436 4519
rect 15936 4150 15988 4156
rect 16224 4146 16436 4162
rect 16212 4140 16436 4146
rect 16264 4134 16436 4140
rect 16212 4082 16264 4088
rect 16304 4072 16356 4078
rect 16500 4026 16528 4655
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 4214 16620 4490
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16684 4078 16712 4966
rect 16776 4214 16804 5120
rect 16856 5102 16908 5108
rect 16960 4554 16988 5510
rect 17222 5471 17278 5480
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 16948 4548 17000 4554
rect 17052 4536 17080 5238
rect 17144 4826 17172 5238
rect 17236 5030 17264 5471
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17132 4548 17184 4554
rect 17052 4508 17132 4536
rect 16948 4490 17000 4496
rect 17132 4490 17184 4496
rect 17144 4214 17172 4490
rect 16764 4208 16816 4214
rect 17132 4208 17184 4214
rect 16764 4150 16816 4156
rect 17052 4168 17132 4196
rect 16356 4020 16528 4026
rect 16304 4014 16528 4020
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16316 3998 16528 4014
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14108 2582 14136 2994
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 12492 1924 12572 1952
rect 12440 1906 12492 1912
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 12256 1760 12308 1766
rect 12256 1702 12308 1708
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10336 1358 10364 1702
rect 11060 1556 11112 1562
rect 10980 1516 11060 1544
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 8944 1352 8996 1358
rect 8944 1294 8996 1300
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 10416 1216 10468 1222
rect 10416 1158 10468 1164
rect 5170 54 5488 82
rect 4342 -300 4398 54
rect 5170 -300 5226 54
rect 5998 -300 6054 160
rect 6826 -300 6882 160
rect 7654 82 7710 160
rect 7944 82 7972 1158
rect 7654 54 7972 82
rect 8482 82 8538 160
rect 8772 82 8800 1158
rect 8482 54 8800 82
rect 9310 82 9366 160
rect 9600 82 9628 1158
rect 9310 54 9628 82
rect 10138 82 10194 160
rect 10428 82 10456 1158
rect 10980 160 11008 1516
rect 11060 1498 11112 1504
rect 11164 1358 11192 1702
rect 11992 1358 12020 1702
rect 12268 1358 12296 1702
rect 12360 1494 12388 1906
rect 12348 1488 12400 1494
rect 12348 1430 12400 1436
rect 13464 1358 13492 2246
rect 14108 2038 14136 2518
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14200 2378 14228 2450
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14292 2106 14320 2314
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 14476 1952 14504 3130
rect 14936 2854 14964 3470
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 15304 3194 15332 3402
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 14832 2848 14884 2854
rect 14660 2796 14832 2802
rect 14660 2790 14884 2796
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14660 2774 14872 2790
rect 14556 2372 14608 2378
rect 14660 2360 14688 2774
rect 14936 2514 14964 2790
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 14608 2332 14688 2360
rect 14556 2314 14608 2320
rect 14556 1964 14608 1970
rect 14476 1924 14556 1952
rect 14556 1906 14608 1912
rect 14936 1902 14964 2450
rect 15856 2378 15884 3878
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16316 3398 16344 3606
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16070 3292 16378 3301
rect 16070 3290 16076 3292
rect 16132 3290 16156 3292
rect 16212 3290 16236 3292
rect 16292 3290 16316 3292
rect 16372 3290 16378 3292
rect 16132 3238 16134 3290
rect 16314 3238 16316 3290
rect 16070 3236 16076 3238
rect 16132 3236 16156 3238
rect 16212 3236 16236 3238
rect 16292 3236 16316 3238
rect 16372 3236 16378 3238
rect 16070 3227 16378 3236
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16408 2961 16436 2994
rect 16488 2984 16540 2990
rect 16394 2952 16450 2961
rect 16488 2926 16540 2932
rect 16394 2887 16450 2896
rect 16500 2650 16528 2926
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14372 1760 14424 1766
rect 14372 1702 14424 1708
rect 15384 1760 15436 1766
rect 15384 1702 15436 1708
rect 13570 1660 13878 1669
rect 13570 1658 13576 1660
rect 13632 1658 13656 1660
rect 13712 1658 13736 1660
rect 13792 1658 13816 1660
rect 13872 1658 13878 1660
rect 13632 1606 13634 1658
rect 13814 1606 13816 1658
rect 13570 1604 13576 1606
rect 13632 1604 13656 1606
rect 13712 1604 13736 1606
rect 13792 1604 13816 1606
rect 13872 1604 13878 1606
rect 13570 1595 13878 1604
rect 14384 1358 14412 1702
rect 15200 1556 15252 1562
rect 15200 1498 15252 1504
rect 15212 1442 15240 1498
rect 15120 1414 15240 1442
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 12256 1352 12308 1358
rect 12256 1294 12308 1300
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14096 1284 14148 1290
rect 14096 1226 14148 1232
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 13728 1216 13780 1222
rect 13728 1158 13780 1164
rect 11070 1116 11378 1125
rect 11070 1114 11076 1116
rect 11132 1114 11156 1116
rect 11212 1114 11236 1116
rect 11292 1114 11316 1116
rect 11372 1114 11378 1116
rect 11132 1062 11134 1114
rect 11314 1062 11316 1114
rect 11070 1060 11076 1062
rect 11132 1060 11156 1062
rect 11212 1060 11236 1062
rect 11292 1060 11316 1062
rect 11372 1060 11378 1062
rect 11070 1051 11378 1060
rect 10138 54 10456 82
rect 7654 -300 7710 54
rect 8482 -300 8538 54
rect 9310 -300 9366 54
rect 10138 -300 10194 54
rect 10966 -300 11022 160
rect 11794 82 11850 160
rect 12084 82 12112 1158
rect 11794 54 12112 82
rect 12622 82 12678 160
rect 12912 82 12940 1158
rect 12622 54 12940 82
rect 13450 82 13506 160
rect 13740 82 13768 1158
rect 14108 1018 14136 1226
rect 14188 1216 14240 1222
rect 14188 1158 14240 1164
rect 14280 1216 14332 1222
rect 14280 1158 14332 1164
rect 14200 1018 14228 1158
rect 14096 1012 14148 1018
rect 14096 954 14148 960
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 14292 160 14320 1158
rect 15120 160 15148 1414
rect 15396 1358 15424 1702
rect 15856 1494 15884 2314
rect 15948 2106 15976 2586
rect 16070 2204 16378 2213
rect 16070 2202 16076 2204
rect 16132 2202 16156 2204
rect 16212 2202 16236 2204
rect 16292 2202 16316 2204
rect 16372 2202 16378 2204
rect 16132 2150 16134 2202
rect 16314 2150 16316 2202
rect 16070 2148 16076 2150
rect 16132 2148 16156 2150
rect 16212 2148 16236 2150
rect 16292 2148 16316 2150
rect 16372 2148 16378 2150
rect 16070 2139 16378 2148
rect 15936 2100 15988 2106
rect 15936 2042 15988 2048
rect 16592 1970 16620 3334
rect 16684 3058 16712 3538
rect 16776 3058 16804 4150
rect 17052 3534 17080 4168
rect 17132 4150 17184 4156
rect 17236 3534 17264 4966
rect 17696 4078 17724 5850
rect 17880 5642 17908 6326
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17972 4758 18000 5782
rect 18064 5710 18092 6190
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18064 4758 18092 5646
rect 18340 5642 18368 6734
rect 18432 6730 18460 6938
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18432 5896 18460 6666
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6458 18552 6598
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18570 6012 18878 6021
rect 18570 6010 18576 6012
rect 18632 6010 18656 6012
rect 18712 6010 18736 6012
rect 18792 6010 18816 6012
rect 18872 6010 18878 6012
rect 18632 5958 18634 6010
rect 18814 5958 18816 6010
rect 18570 5956 18576 5958
rect 18632 5956 18656 5958
rect 18712 5956 18736 5958
rect 18792 5956 18816 5958
rect 18872 5956 18878 5958
rect 18570 5947 18878 5956
rect 18432 5868 18552 5896
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5370 18184 5510
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18432 4622 18460 5714
rect 18524 5642 18552 5868
rect 18984 5710 19012 6190
rect 19076 6089 19104 11183
rect 19340 11154 19392 11160
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10810 19288 11086
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19260 10266 19288 10746
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19168 8634 19196 9590
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9178 19288 9454
rect 19352 9450 19380 11154
rect 19536 10674 19564 11154
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19996 10470 20024 11086
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19444 8974 19472 9862
rect 19628 9110 19656 10134
rect 20180 10130 20208 11342
rect 20272 11218 20300 11562
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20272 10742 20300 10950
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19536 8294 19564 8502
rect 19628 8498 19656 9046
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19168 6854 19472 6882
rect 19168 6662 19196 6854
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19062 6080 19118 6089
rect 19062 6015 19118 6024
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18708 5234 18736 5578
rect 19076 5556 19104 6015
rect 19168 5710 19196 6394
rect 19260 6118 19288 6598
rect 19352 6254 19380 6734
rect 19444 6662 19472 6854
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5778 19288 6054
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 18984 5528 19104 5556
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18570 4924 18878 4933
rect 18570 4922 18576 4924
rect 18632 4922 18656 4924
rect 18712 4922 18736 4924
rect 18792 4922 18816 4924
rect 18872 4922 18878 4924
rect 18632 4870 18634 4922
rect 18814 4870 18816 4922
rect 18570 4868 18576 4870
rect 18632 4868 18656 4870
rect 18712 4868 18736 4870
rect 18792 4868 18816 4870
rect 18872 4868 18878 4870
rect 18570 4859 18878 4868
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 18570 3836 18878 3845
rect 18570 3834 18576 3836
rect 18632 3834 18656 3836
rect 18712 3834 18736 3836
rect 18792 3834 18816 3836
rect 18872 3834 18878 3836
rect 18632 3782 18634 3834
rect 18814 3782 18816 3834
rect 18570 3780 18576 3782
rect 18632 3780 18656 3782
rect 18712 3780 18736 3782
rect 18792 3780 18816 3782
rect 18872 3780 18878 3782
rect 18570 3771 18878 3780
rect 18984 3720 19012 5528
rect 19352 5302 19380 5646
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 5114 19472 6598
rect 19536 5778 19564 6802
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19352 5086 19472 5114
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 4622 19104 4966
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 19076 3738 19104 4150
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19156 4072 19208 4078
rect 19154 4040 19156 4049
rect 19208 4040 19210 4049
rect 19154 3975 19210 3984
rect 19260 3738 19288 4082
rect 18892 3692 19012 3720
rect 19064 3732 19116 3738
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18340 3534 18368 3606
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3194 16896 3334
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16672 2508 16724 2514
rect 16776 2496 16804 2994
rect 16724 2468 16804 2496
rect 16672 2450 16724 2456
rect 16684 1970 16712 2450
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 16960 2106 16988 2314
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 17052 2038 17080 3470
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18248 3194 18276 3334
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17776 3120 17828 3126
rect 17696 3080 17776 3108
rect 17696 2378 17724 3080
rect 17828 3080 18184 3108
rect 17776 3062 17828 3068
rect 18156 3074 18184 3080
rect 18340 3074 18368 3130
rect 18156 3046 18368 3074
rect 18800 3058 18828 3402
rect 18892 3380 18920 3692
rect 19064 3674 19116 3680
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19076 3534 19104 3674
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18892 3352 19104 3380
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18570 2748 18878 2757
rect 18570 2746 18576 2748
rect 18632 2746 18656 2748
rect 18712 2746 18736 2748
rect 18792 2746 18816 2748
rect 18872 2746 18878 2748
rect 18632 2694 18634 2746
rect 18814 2694 18816 2746
rect 18570 2692 18576 2694
rect 18632 2692 18656 2694
rect 18712 2692 18736 2694
rect 18792 2692 18816 2694
rect 18872 2692 18878 2694
rect 18570 2683 18878 2692
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17696 2038 17724 2314
rect 17040 2032 17092 2038
rect 17040 1974 17092 1980
rect 17684 2032 17736 2038
rect 17684 1974 17736 1980
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 16672 1964 16724 1970
rect 16672 1906 16724 1912
rect 16212 1760 16264 1766
rect 16212 1702 16264 1708
rect 15844 1488 15896 1494
rect 15844 1430 15896 1436
rect 16224 1358 16252 1702
rect 16684 1562 16712 1906
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 16672 1556 16724 1562
rect 16672 1498 16724 1504
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 16212 1352 16264 1358
rect 16212 1294 16264 1300
rect 15936 1216 15988 1222
rect 15936 1158 15988 1164
rect 17040 1216 17092 1222
rect 17040 1158 17092 1164
rect 15948 160 15976 1158
rect 16070 1116 16378 1125
rect 16070 1114 16076 1116
rect 16132 1114 16156 1116
rect 16212 1114 16236 1116
rect 16292 1114 16316 1116
rect 16372 1114 16378 1116
rect 16132 1062 16134 1114
rect 16314 1062 16316 1114
rect 16070 1060 16076 1062
rect 16132 1060 16156 1062
rect 16212 1060 16236 1062
rect 16292 1060 16316 1062
rect 16372 1060 16378 1062
rect 16070 1051 16378 1060
rect 13450 54 13768 82
rect 11794 -300 11850 54
rect 12622 -300 12678 54
rect 13450 -300 13506 54
rect 14278 -300 14334 160
rect 15106 -300 15162 160
rect 15934 -300 15990 160
rect 16762 82 16818 160
rect 17052 82 17080 1158
rect 17604 160 17632 1702
rect 17696 1562 17724 1974
rect 18524 1970 18552 2450
rect 19076 2378 19104 3352
rect 19168 2990 19196 3402
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 2106 18644 2246
rect 19168 2106 19196 2926
rect 19260 2514 19288 3538
rect 19352 3194 19380 5086
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 4826 19472 4966
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19444 3233 19472 4762
rect 19536 4758 19564 5510
rect 19628 4865 19656 8298
rect 19812 7342 19840 8910
rect 19904 8430 19932 9454
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19996 8566 20024 9386
rect 20180 8906 20208 9930
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20180 8430 20208 8842
rect 20272 8634 20300 10678
rect 20364 9654 20392 11086
rect 20640 10266 20668 11698
rect 20732 11626 20760 12406
rect 20824 12238 20852 12406
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20916 11898 20944 12650
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21070 11996 21378 12005
rect 21070 11994 21076 11996
rect 21132 11994 21156 11996
rect 21212 11994 21236 11996
rect 21292 11994 21316 11996
rect 21372 11994 21378 11996
rect 21132 11942 21134 11994
rect 21314 11942 21316 11994
rect 21070 11940 21076 11942
rect 21132 11940 21156 11942
rect 21212 11940 21236 11942
rect 21292 11940 21316 11942
rect 21372 11940 21378 11942
rect 21070 11931 21378 11940
rect 21468 11898 21496 12106
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20732 11354 20760 11562
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11354 20944 11494
rect 21376 11354 21404 11698
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20352 9648 20404 9654
rect 20640 9636 20668 9998
rect 20824 9722 20852 10406
rect 20916 10266 20944 11086
rect 21560 11014 21588 11494
rect 21652 11286 21680 11698
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21652 11014 21680 11222
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21070 10908 21378 10917
rect 21070 10906 21076 10908
rect 21132 10906 21156 10908
rect 21212 10906 21236 10908
rect 21292 10906 21316 10908
rect 21372 10906 21378 10908
rect 21132 10854 21134 10906
rect 21314 10854 21316 10906
rect 21070 10852 21076 10854
rect 21132 10852 21156 10854
rect 21212 10852 21236 10854
rect 21292 10852 21316 10854
rect 21372 10852 21378 10854
rect 21070 10843 21378 10852
rect 21640 10736 21692 10742
rect 21640 10678 21692 10684
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21088 10124 21140 10130
rect 21008 10084 21088 10112
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20352 9590 20404 9596
rect 20456 9608 20668 9636
rect 20456 9382 20484 9608
rect 20824 9586 20852 9658
rect 21008 9602 21036 10084
rect 21088 10066 21140 10072
rect 21192 10062 21220 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21070 9820 21378 9829
rect 21070 9818 21076 9820
rect 21132 9818 21156 9820
rect 21212 9818 21236 9820
rect 21292 9818 21316 9820
rect 21372 9818 21378 9820
rect 21132 9766 21134 9818
rect 21314 9766 21316 9818
rect 21070 9764 21076 9766
rect 21132 9764 21156 9766
rect 21212 9764 21236 9766
rect 21292 9764 21316 9766
rect 21372 9764 21378 9766
rect 21070 9755 21378 9764
rect 20916 9586 21036 9602
rect 21272 9648 21324 9654
rect 21468 9636 21496 9998
rect 21560 9994 21588 10406
rect 21652 10130 21680 10678
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21836 10010 21864 22442
rect 22204 22234 22232 22578
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22296 22094 22324 23054
rect 22112 22066 22324 22094
rect 22008 21480 22060 21486
rect 22008 21422 22060 21428
rect 22020 21146 22048 21422
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22020 20466 22048 20946
rect 22112 20505 22140 22066
rect 22388 22030 22416 23190
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22098 20496 22154 20505
rect 22008 20460 22060 20466
rect 22204 20466 22232 21830
rect 22296 21622 22324 21830
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22388 20777 22416 21966
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22480 20806 22508 20878
rect 22468 20800 22520 20806
rect 22374 20768 22430 20777
rect 22468 20742 22520 20748
rect 22374 20703 22430 20712
rect 22098 20431 22154 20440
rect 22192 20460 22244 20466
rect 22008 20402 22060 20408
rect 22244 20420 22324 20448
rect 22192 20402 22244 20408
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 21928 19990 21956 20266
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 22020 19718 22048 19994
rect 22204 19786 22232 20266
rect 22296 19922 22324 20420
rect 22572 20058 22600 20878
rect 22848 20398 22876 23394
rect 22940 22778 22968 23840
rect 23480 23384 23532 23390
rect 23480 23326 23532 23332
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23032 22234 23060 22578
rect 23124 22234 23152 22578
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23216 21486 23244 21830
rect 23308 21593 23336 23122
rect 23492 22094 23520 23326
rect 23860 22778 23888 23840
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23570 22332 23878 22341
rect 23570 22330 23576 22332
rect 23632 22330 23656 22332
rect 23712 22330 23736 22332
rect 23792 22330 23816 22332
rect 23872 22330 23878 22332
rect 23632 22278 23634 22330
rect 23814 22278 23816 22330
rect 23570 22276 23576 22278
rect 23632 22276 23656 22278
rect 23712 22276 23736 22278
rect 23792 22276 23816 22278
rect 23872 22276 23878 22278
rect 23570 22267 23878 22276
rect 24044 22094 24072 23258
rect 24780 22778 24808 23840
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 23492 22066 23704 22094
rect 24044 22066 24256 22094
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23294 21584 23350 21593
rect 23294 21519 23350 21528
rect 23204 21480 23256 21486
rect 23018 21448 23074 21457
rect 23204 21422 23256 21428
rect 23018 21383 23074 21392
rect 23032 20913 23060 21383
rect 23112 20936 23164 20942
rect 23018 20904 23074 20913
rect 23112 20878 23164 20884
rect 23018 20839 23074 20848
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23032 20534 23060 20742
rect 23124 20602 23152 20878
rect 23216 20874 23244 21422
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23308 20777 23336 21519
rect 23400 21457 23428 21966
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23386 21448 23442 21457
rect 23386 21383 23442 21392
rect 23492 21010 23520 21830
rect 23584 21690 23612 21966
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23676 21593 23704 22066
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23662 21584 23718 21593
rect 23662 21519 23718 21528
rect 23860 21350 23888 21830
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23570 21244 23878 21253
rect 23570 21242 23576 21244
rect 23632 21242 23656 21244
rect 23712 21242 23736 21244
rect 23792 21242 23816 21244
rect 23872 21242 23878 21244
rect 23632 21190 23634 21242
rect 23814 21190 23816 21242
rect 23570 21188 23576 21190
rect 23632 21188 23656 21190
rect 23712 21188 23736 21190
rect 23792 21188 23816 21190
rect 23872 21188 23878 21190
rect 23570 21179 23878 21188
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23294 20768 23350 20777
rect 23294 20703 23350 20712
rect 23400 20602 23428 20878
rect 23952 20602 23980 21422
rect 24136 20806 24164 21558
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23020 20528 23072 20534
rect 23020 20470 23072 20476
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 24228 20330 24256 22066
rect 24320 20874 24348 22374
rect 24780 22234 24808 22578
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24872 22094 24900 22986
rect 25700 22778 25728 23840
rect 26070 22876 26378 22885
rect 26070 22874 26076 22876
rect 26132 22874 26156 22876
rect 26212 22874 26236 22876
rect 26292 22874 26316 22876
rect 26372 22874 26378 22876
rect 26132 22822 26134 22874
rect 26314 22822 26316 22874
rect 26070 22820 26076 22822
rect 26132 22820 26156 22822
rect 26212 22820 26236 22822
rect 26292 22820 26316 22822
rect 26372 22820 26378 22822
rect 26070 22811 26378 22820
rect 26620 22778 26648 23840
rect 27436 23248 27488 23254
rect 27436 23190 27488 23196
rect 27540 23202 27568 23840
rect 28460 23202 28488 23840
rect 29380 23746 29408 23840
rect 29472 23746 29500 23854
rect 29380 23718 29500 23746
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 27448 22710 27476 23190
rect 27540 23174 27660 23202
rect 27632 22710 27660 23174
rect 28172 23180 28224 23186
rect 28460 23174 28672 23202
rect 28172 23122 28224 23128
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 27896 23044 27948 23050
rect 27896 22986 27948 22992
rect 27908 22778 27936 22986
rect 27896 22772 27948 22778
rect 27896 22714 27948 22720
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 24872 22066 25176 22094
rect 24492 21956 24544 21962
rect 24492 21898 24544 21904
rect 24504 21486 24532 21898
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24780 21010 24808 22034
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24308 20868 24360 20874
rect 24308 20810 24360 20816
rect 24780 20602 24808 20946
rect 24872 20777 24900 22066
rect 25148 22030 25176 22066
rect 25332 22030 25360 22374
rect 25608 22137 25636 22578
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25594 22128 25650 22137
rect 25594 22063 25650 22072
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25320 22024 25372 22030
rect 25372 21984 25452 22012
rect 25320 21966 25372 21972
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21622 25360 21830
rect 25320 21616 25372 21622
rect 25424 21604 25452 21984
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25504 21616 25556 21622
rect 25424 21576 25504 21604
rect 25320 21558 25372 21564
rect 25504 21558 25556 21564
rect 25332 20942 25360 21558
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 24858 20768 24914 20777
rect 24858 20703 24914 20712
rect 25608 20602 25636 21898
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25686 21720 25742 21729
rect 25792 21690 25820 21830
rect 25884 21690 25912 22510
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25686 21655 25742 21664
rect 25780 21684 25832 21690
rect 25700 21185 25728 21655
rect 25780 21626 25832 21632
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25686 21176 25742 21185
rect 25884 21146 25912 21626
rect 25686 21111 25742 21120
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 25976 21026 26004 21830
rect 26070 21788 26378 21797
rect 26070 21786 26076 21788
rect 26132 21786 26156 21788
rect 26212 21786 26236 21788
rect 26292 21786 26316 21788
rect 26372 21786 26378 21788
rect 26132 21734 26134 21786
rect 26314 21734 26316 21786
rect 26070 21732 26076 21734
rect 26132 21732 26156 21734
rect 26212 21732 26236 21734
rect 26292 21732 26316 21734
rect 26372 21732 26378 21734
rect 26070 21723 26378 21732
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 25884 20998 26004 21026
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20602 25728 20742
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 24584 20460 24636 20466
rect 24636 20420 24900 20448
rect 24584 20402 24636 20408
rect 24216 20324 24268 20330
rect 24216 20266 24268 20272
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 23570 20156 23878 20165
rect 23570 20154 23576 20156
rect 23632 20154 23656 20156
rect 23712 20154 23736 20156
rect 23792 20154 23816 20156
rect 23872 20154 23878 20156
rect 23632 20102 23634 20154
rect 23814 20102 23816 20154
rect 23570 20100 23576 20102
rect 23632 20100 23656 20102
rect 23712 20100 23736 20102
rect 23792 20100 23816 20102
rect 23872 20100 23878 20102
rect 23570 20091 23878 20100
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22296 19378 22324 19858
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21928 18834 21956 19110
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21928 17882 21956 18770
rect 22388 17954 22416 19654
rect 23308 19514 23336 19790
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23940 19780 23992 19786
rect 23940 19722 23992 19728
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22480 18698 22508 19110
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22480 18426 22508 18634
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22572 18426 22600 18566
rect 22756 18426 22784 18702
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22848 18290 22876 19246
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22296 17926 22416 17954
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 16114 21956 17478
rect 22020 16454 22048 17682
rect 22296 17066 22324 17926
rect 22756 17882 22784 18226
rect 23124 18222 23152 19246
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23216 18465 23244 18566
rect 23202 18456 23258 18465
rect 23202 18391 23258 18400
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22388 17338 22416 17818
rect 23308 17746 23336 19450
rect 23492 18970 23520 19722
rect 23570 19068 23878 19077
rect 23570 19066 23576 19068
rect 23632 19066 23656 19068
rect 23712 19066 23736 19068
rect 23792 19066 23816 19068
rect 23872 19066 23878 19068
rect 23632 19014 23634 19066
rect 23814 19014 23816 19066
rect 23570 19012 23576 19014
rect 23632 19012 23656 19014
rect 23712 19012 23736 19014
rect 23792 19012 23816 19014
rect 23872 19012 23878 19014
rect 23570 19003 23878 19012
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23952 18465 23980 19722
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 24044 18970 24072 19654
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23938 18456 23994 18465
rect 23938 18391 23994 18400
rect 23570 17980 23878 17989
rect 23570 17978 23576 17980
rect 23632 17978 23656 17980
rect 23712 17978 23736 17980
rect 23792 17978 23816 17980
rect 23872 17978 23878 17980
rect 23632 17926 23634 17978
rect 23814 17926 23816 17978
rect 23570 17924 23576 17926
rect 23632 17924 23656 17926
rect 23712 17924 23736 17926
rect 23792 17924 23816 17926
rect 23872 17924 23878 17926
rect 23570 17915 23878 17924
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 22572 17338 22600 17478
rect 22376 17332 22428 17338
rect 22560 17332 22612 17338
rect 22428 17292 22508 17320
rect 22376 17274 22428 17280
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15910 21956 16050
rect 22296 16046 22324 16526
rect 22388 16454 22416 16934
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21928 15706 21956 15846
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 22112 15502 22140 15982
rect 22296 15570 22324 15982
rect 22480 15910 22508 17292
rect 22560 17274 22612 17280
rect 23216 16794 23244 17478
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22652 16040 22704 16046
rect 22558 16008 22614 16017
rect 22652 15982 22704 15988
rect 22558 15943 22614 15952
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22572 15706 22600 15943
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21928 14414 21956 14826
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 22020 14278 22048 15370
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 21928 13530 21956 14214
rect 22112 13938 22140 15438
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22204 14482 22232 14962
rect 22388 14770 22416 15370
rect 22480 14890 22508 15506
rect 22572 15042 22600 15642
rect 22664 15162 22692 15982
rect 23032 15706 23060 16390
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22572 15014 22692 15042
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22572 14770 22600 14894
rect 22388 14742 22600 14770
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22204 13802 22232 14418
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22296 13682 22324 14214
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22204 13654 22324 13682
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21914 13424 21970 13433
rect 21914 13359 21916 13368
rect 21968 13359 21970 13368
rect 21916 13330 21968 13336
rect 22204 13326 22232 13654
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 11898 22232 13262
rect 22296 13025 22324 13398
rect 22480 13190 22508 13874
rect 22572 13462 22600 14742
rect 22664 14414 22692 15014
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22664 13938 22692 14350
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22282 13016 22338 13025
rect 22282 12951 22338 12960
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 22020 11354 22048 11630
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22296 11150 22324 12951
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12238 22508 12786
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22480 11830 22508 12174
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22664 11218 22692 13874
rect 22756 12986 22784 14486
rect 22848 13326 22876 14758
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22940 13870 22968 14350
rect 23032 13920 23060 15642
rect 23216 14618 23244 16730
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 15570 23336 16390
rect 23400 15570 23428 17682
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23400 15162 23428 15506
rect 23492 15366 23520 17478
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23570 16892 23878 16901
rect 23570 16890 23576 16892
rect 23632 16890 23656 16892
rect 23712 16890 23736 16892
rect 23792 16890 23816 16892
rect 23872 16890 23878 16892
rect 23632 16838 23634 16890
rect 23814 16838 23816 16890
rect 23570 16836 23576 16838
rect 23632 16836 23656 16838
rect 23712 16836 23736 16838
rect 23792 16836 23816 16838
rect 23872 16836 23878 16838
rect 23570 16827 23878 16836
rect 23754 16552 23810 16561
rect 23754 16487 23810 16496
rect 23768 16454 23796 16487
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23570 15804 23878 15813
rect 23570 15802 23576 15804
rect 23632 15802 23656 15804
rect 23712 15802 23736 15804
rect 23792 15802 23816 15804
rect 23872 15802 23878 15804
rect 23632 15750 23634 15802
rect 23814 15750 23816 15802
rect 23570 15748 23576 15750
rect 23632 15748 23656 15750
rect 23712 15748 23736 15750
rect 23792 15748 23816 15750
rect 23872 15748 23878 15750
rect 23570 15739 23878 15748
rect 23664 15632 23716 15638
rect 23952 15609 23980 16934
rect 24044 16590 24072 18770
rect 24136 18766 24164 19926
rect 24308 19916 24360 19922
rect 24308 19858 24360 19864
rect 24320 18834 24348 19858
rect 24412 19310 24440 20198
rect 24872 19961 24900 20420
rect 25884 20330 25912 20998
rect 26068 20924 26096 21558
rect 26528 21146 26556 22578
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26620 21622 26648 22374
rect 27448 22094 27476 22646
rect 28092 22574 28120 23054
rect 28184 22642 28212 23122
rect 28644 22778 28672 23174
rect 29748 22778 29776 23854
rect 30286 23840 30342 24300
rect 31206 23840 31262 24300
rect 32126 23840 32182 24300
rect 32232 23854 32628 23882
rect 28632 22772 28684 22778
rect 28632 22714 28684 22720
rect 29736 22772 29788 22778
rect 29736 22714 29788 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27264 22066 27476 22094
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 26608 21616 26660 21622
rect 26608 21558 26660 21564
rect 26698 21448 26754 21457
rect 26698 21383 26754 21392
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 25976 20896 26096 20924
rect 25872 20324 25924 20330
rect 25872 20266 25924 20272
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 24858 19952 24914 19961
rect 24858 19887 24914 19896
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 24872 19514 24900 19654
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24228 17270 24256 18226
rect 24320 17610 24348 18566
rect 24412 18290 24440 19246
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24492 18760 24544 18766
rect 24544 18720 24716 18748
rect 24492 18702 24544 18708
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 24320 17338 24348 17546
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24044 16250 24072 16526
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23664 15574 23716 15580
rect 23938 15600 23994 15609
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23400 14521 23428 14962
rect 23386 14512 23442 14521
rect 23308 14470 23386 14498
rect 23308 14278 23336 14470
rect 23386 14447 23442 14456
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23112 13932 23164 13938
rect 23032 13892 23112 13920
rect 23112 13874 23164 13880
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 23124 13530 23152 13874
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22756 12238 22784 12922
rect 22940 12442 22968 13262
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22848 12238 22876 12310
rect 23124 12238 23152 13466
rect 23216 13258 23244 13874
rect 23308 13326 23336 14214
rect 23492 14056 23520 15302
rect 23676 15162 23704 15574
rect 23938 15535 23994 15544
rect 23952 15162 23980 15535
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 24044 15162 24072 15370
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24136 14890 24164 16390
rect 24228 16182 24256 17206
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 16658 24440 17138
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24216 16176 24268 16182
rect 24216 16118 24268 16124
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24214 15056 24270 15065
rect 24412 15026 24440 15098
rect 24214 14991 24270 15000
rect 24400 15020 24452 15026
rect 24228 14958 24256 14991
rect 24400 14962 24452 14968
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23570 14716 23878 14725
rect 23570 14714 23576 14716
rect 23632 14714 23656 14716
rect 23712 14714 23736 14716
rect 23792 14714 23816 14716
rect 23872 14714 23878 14716
rect 23632 14662 23634 14714
rect 23814 14662 23816 14714
rect 23570 14660 23576 14662
rect 23632 14660 23656 14662
rect 23712 14660 23736 14662
rect 23792 14660 23816 14662
rect 23872 14660 23878 14662
rect 23570 14651 23878 14660
rect 23952 14550 23980 14758
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23940 14544 23992 14550
rect 24228 14498 24256 14894
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 23940 14486 23992 14492
rect 23400 14028 23520 14056
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23216 12714 23244 13194
rect 23294 13016 23350 13025
rect 23400 13002 23428 14028
rect 23768 14006 23796 14486
rect 24136 14470 24256 14498
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23952 13938 23980 14350
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23492 13190 23520 13874
rect 23570 13628 23878 13637
rect 23570 13626 23576 13628
rect 23632 13626 23656 13628
rect 23712 13626 23736 13628
rect 23792 13626 23816 13628
rect 23872 13626 23878 13628
rect 23632 13574 23634 13626
rect 23814 13574 23816 13626
rect 23570 13572 23576 13574
rect 23632 13572 23656 13574
rect 23712 13572 23736 13574
rect 23792 13572 23816 13574
rect 23872 13572 23878 13574
rect 23570 13563 23878 13572
rect 23848 13320 23900 13326
rect 23846 13288 23848 13297
rect 23900 13288 23902 13297
rect 23846 13223 23902 13232
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23400 12974 23520 13002
rect 23294 12951 23350 12960
rect 23308 12850 23336 12951
rect 23492 12866 23520 12974
rect 23846 12880 23902 12889
rect 23296 12844 23348 12850
rect 23492 12844 23846 12866
rect 23492 12838 23756 12844
rect 23296 12786 23348 12792
rect 23808 12838 23846 12844
rect 23846 12815 23902 12824
rect 23756 12786 23808 12792
rect 23204 12708 23256 12714
rect 23204 12650 23256 12656
rect 23296 12708 23348 12714
rect 23296 12650 23348 12656
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21928 10674 21956 10950
rect 22204 10810 22232 11086
rect 22480 10810 22508 11154
rect 22756 11150 22784 12174
rect 22848 11898 22876 12174
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22848 11218 22876 11834
rect 23124 11558 23152 12174
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23308 11354 23336 12650
rect 23570 12540 23878 12549
rect 23570 12538 23576 12540
rect 23632 12538 23656 12540
rect 23712 12538 23736 12540
rect 23792 12538 23816 12540
rect 23872 12538 23878 12540
rect 23632 12486 23634 12538
rect 23814 12486 23816 12538
rect 23570 12484 23576 12486
rect 23632 12484 23656 12486
rect 23712 12484 23736 12486
rect 23792 12484 23816 12486
rect 23872 12484 23878 12486
rect 23570 12475 23878 12484
rect 23952 12442 23980 13874
rect 24044 13530 24072 14214
rect 24136 14074 24164 14470
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24044 13190 24072 13466
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12782 24072 13126
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24136 12646 24164 13738
rect 24124 12640 24176 12646
rect 24044 12600 24124 12628
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23400 12238 23428 12378
rect 24044 12238 24072 12600
rect 24124 12582 24176 12588
rect 24228 12442 24256 14350
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24412 12968 24440 13466
rect 24504 13326 24532 14758
rect 24582 14648 24638 14657
rect 24582 14583 24584 14592
rect 24636 14583 24638 14592
rect 24584 14554 24636 14560
rect 24688 14226 24716 18720
rect 24780 18426 24808 19110
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24872 18426 24900 18634
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 24858 18320 24914 18329
rect 24858 18255 24860 18264
rect 24912 18255 24914 18264
rect 24952 18284 25004 18290
rect 24860 18226 24912 18232
rect 24952 18226 25004 18232
rect 24964 18086 24992 18226
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24872 17746 24900 18022
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24964 17338 24992 17614
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24780 16182 24808 16934
rect 24964 16794 24992 17138
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24964 16046 24992 16390
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24872 15366 24900 15982
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24596 14198 24716 14226
rect 24596 13394 24624 14198
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24688 13870 24716 14010
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13462 24716 13806
rect 24780 13734 24808 14894
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24872 14618 24900 14758
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24320 12940 24440 12968
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24320 12238 24348 12940
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12238 24440 12786
rect 24504 12442 24532 13262
rect 24676 13184 24728 13190
rect 24582 13152 24638 13161
rect 24676 13126 24728 13132
rect 24582 13087 24638 13096
rect 24596 12986 24624 13087
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 23570 11452 23878 11461
rect 23570 11450 23576 11452
rect 23632 11450 23656 11452
rect 23712 11450 23736 11452
rect 23792 11450 23816 11452
rect 23872 11450 23878 11452
rect 23632 11398 23634 11450
rect 23814 11398 23816 11450
rect 23570 11396 23576 11398
rect 23632 11396 23656 11398
rect 23712 11396 23736 11398
rect 23792 11396 23816 11398
rect 23872 11396 23878 11398
rect 23570 11387 23878 11396
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22020 10198 22048 10406
rect 22480 10266 22508 10610
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22008 10192 22060 10198
rect 22008 10134 22060 10140
rect 21548 9988 21600 9994
rect 21836 9982 21956 10010
rect 21548 9930 21600 9936
rect 21560 9874 21588 9930
rect 21732 9920 21784 9926
rect 21560 9846 21680 9874
rect 21732 9862 21784 9868
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21324 9608 21496 9636
rect 21272 9590 21324 9596
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20904 9580 21036 9586
rect 20956 9574 21036 9580
rect 20904 9522 20956 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19904 7342 19932 7754
rect 20180 7546 20208 8230
rect 20456 7818 20484 9318
rect 20732 8548 20760 9522
rect 21178 9480 21234 9489
rect 21178 9415 21180 9424
rect 21232 9415 21234 9424
rect 21548 9444 21600 9450
rect 21180 9386 21232 9392
rect 21548 9386 21600 9392
rect 21560 9178 21588 9386
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21652 9058 21680 9846
rect 21744 9602 21772 9862
rect 21836 9722 21864 9862
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21744 9574 21864 9602
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21468 9030 21680 9058
rect 21070 8732 21378 8741
rect 21070 8730 21076 8732
rect 21132 8730 21156 8732
rect 21212 8730 21236 8732
rect 21292 8730 21316 8732
rect 21372 8730 21378 8732
rect 21132 8678 21134 8730
rect 21314 8678 21316 8730
rect 21070 8676 21076 8678
rect 21132 8676 21156 8678
rect 21212 8676 21236 8678
rect 21292 8676 21316 8678
rect 21372 8676 21378 8678
rect 21070 8667 21378 8676
rect 20812 8560 20864 8566
rect 20732 8520 20812 8548
rect 20812 8502 20864 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20640 8090 20668 8434
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19798 6896 19854 6905
rect 19798 6831 19854 6840
rect 19812 5914 19840 6831
rect 19904 6662 19932 7278
rect 20548 6934 20576 7822
rect 20640 7002 20668 7890
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20536 6928 20588 6934
rect 20536 6870 20588 6876
rect 20732 6866 20760 8298
rect 20824 7546 20852 8502
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20916 7478 20944 7754
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 19904 6390 19932 6598
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19890 5536 19946 5545
rect 19614 4856 19670 4865
rect 19720 4826 19748 5510
rect 19812 5370 19840 5510
rect 19890 5471 19946 5480
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19614 4791 19670 4800
rect 19708 4820 19760 4826
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19628 4604 19656 4791
rect 19708 4762 19760 4768
rect 19812 4622 19840 5306
rect 19904 4729 19932 5471
rect 19890 4720 19946 4729
rect 19890 4655 19946 4664
rect 19536 4576 19656 4604
rect 19800 4616 19852 4622
rect 19430 3224 19486 3233
rect 19340 3188 19392 3194
rect 19430 3159 19486 3168
rect 19340 3130 19392 3136
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19444 2650 19472 3062
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19246 2408 19302 2417
rect 19246 2343 19302 2352
rect 19260 2106 19288 2343
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18328 1760 18380 1766
rect 18328 1702 18380 1708
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 17684 1556 17736 1562
rect 17684 1498 17736 1504
rect 18340 1358 18368 1702
rect 18432 1358 18460 1702
rect 18570 1660 18878 1669
rect 18570 1658 18576 1660
rect 18632 1658 18656 1660
rect 18712 1658 18736 1660
rect 18792 1658 18816 1660
rect 18872 1658 18878 1660
rect 18632 1606 18634 1658
rect 18814 1606 18816 1658
rect 18570 1604 18576 1606
rect 18632 1604 18656 1606
rect 18712 1604 18736 1606
rect 18792 1604 18816 1606
rect 18872 1604 18878 1606
rect 18570 1595 18878 1604
rect 19340 1556 19392 1562
rect 19340 1498 19392 1504
rect 19352 1442 19380 1498
rect 19260 1414 19380 1442
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 18420 1352 18472 1358
rect 18420 1294 18472 1300
rect 18420 1216 18472 1222
rect 18420 1158 18472 1164
rect 18432 160 18460 1158
rect 19260 160 19288 1414
rect 19536 1290 19564 4576
rect 19800 4558 19852 4564
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19720 2514 19748 3878
rect 19904 3534 19932 4655
rect 19996 4554 20024 6598
rect 20180 5778 20208 6598
rect 20364 6186 20392 6598
rect 20456 6322 20484 6802
rect 20916 6497 20944 6938
rect 21008 6730 21036 8298
rect 21468 7954 21496 9030
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21560 8634 21588 8910
rect 21744 8906 21772 9454
rect 21836 9382 21864 9574
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21560 8401 21588 8570
rect 21928 8480 21956 9982
rect 22020 9586 22048 10134
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 9722 22324 9862
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 22020 8974 22048 9007
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21744 8452 21956 8480
rect 21546 8392 21602 8401
rect 21546 8327 21602 8336
rect 21560 7970 21588 8327
rect 21456 7948 21508 7954
rect 21560 7942 21680 7970
rect 21456 7890 21508 7896
rect 21070 7644 21378 7653
rect 21070 7642 21076 7644
rect 21132 7642 21156 7644
rect 21212 7642 21236 7644
rect 21292 7642 21316 7644
rect 21372 7642 21378 7644
rect 21132 7590 21134 7642
rect 21314 7590 21316 7642
rect 21070 7588 21076 7590
rect 21132 7588 21156 7590
rect 21212 7588 21236 7590
rect 21292 7588 21316 7590
rect 21372 7588 21378 7590
rect 21070 7579 21378 7588
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20902 6488 20958 6497
rect 21008 6458 21036 6666
rect 21070 6556 21378 6565
rect 21070 6554 21076 6556
rect 21132 6554 21156 6556
rect 21212 6554 21236 6556
rect 21292 6554 21316 6556
rect 21372 6554 21378 6556
rect 21132 6502 21134 6554
rect 21314 6502 21316 6554
rect 21070 6500 21076 6502
rect 21132 6500 21156 6502
rect 21212 6500 21236 6502
rect 21292 6500 21316 6502
rect 21372 6500 21378 6502
rect 21070 6491 21378 6500
rect 20902 6423 20958 6432
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21468 6322 21496 7890
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6458 21588 6666
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 20456 5914 20484 6258
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20272 5778 20300 5850
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 20088 4146 20116 5306
rect 20456 4690 20484 5850
rect 20916 5760 20944 6258
rect 21652 6186 21680 7942
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 20996 5772 21048 5778
rect 20916 5732 20996 5760
rect 20810 5400 20866 5409
rect 20810 5335 20866 5344
rect 20824 5166 20852 5335
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20916 5030 20944 5732
rect 20996 5714 21048 5720
rect 21100 5710 21128 6054
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21192 5556 21220 6054
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21008 5528 21220 5556
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20916 4622 20944 4966
rect 21008 4826 21036 5528
rect 21070 5468 21378 5477
rect 21070 5466 21076 5468
rect 21132 5466 21156 5468
rect 21212 5466 21236 5468
rect 21292 5466 21316 5468
rect 21372 5466 21378 5468
rect 21132 5414 21134 5466
rect 21314 5414 21316 5466
rect 21070 5412 21076 5414
rect 21132 5412 21156 5414
rect 21212 5412 21236 5414
rect 21292 5412 21316 5414
rect 21372 5412 21378 5414
rect 21070 5403 21378 5412
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20364 4049 20392 4150
rect 21008 4146 21036 4626
rect 21468 4593 21496 5850
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21560 5098 21588 5578
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21454 4584 21510 4593
rect 21652 4554 21680 5714
rect 21454 4519 21510 4528
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21070 4380 21378 4389
rect 21070 4378 21076 4380
rect 21132 4378 21156 4380
rect 21212 4378 21236 4380
rect 21292 4378 21316 4380
rect 21372 4378 21378 4380
rect 21132 4326 21134 4378
rect 21314 4326 21316 4378
rect 21070 4324 21076 4326
rect 21132 4324 21156 4326
rect 21212 4324 21236 4326
rect 21292 4324 21316 4326
rect 21372 4324 21378 4326
rect 21070 4315 21378 4324
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20350 4040 20406 4049
rect 20350 3975 20406 3984
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19904 3194 19932 3334
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19812 2106 19840 2450
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19904 1970 19932 2926
rect 20364 2650 20392 3975
rect 20456 2990 20484 4082
rect 20548 3466 20576 4082
rect 21560 4078 21588 4422
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 21548 4072 21600 4078
rect 21744 4049 21772 8452
rect 22020 8430 22048 8910
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7478 21864 7686
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21928 6458 21956 8298
rect 22020 7478 22048 8366
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 22112 7410 22140 8502
rect 22204 8090 22232 9318
rect 22388 8974 22416 9454
rect 22572 8974 22600 9998
rect 22848 9897 22876 10066
rect 22940 10062 22968 10950
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23216 10266 23244 10542
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 22834 9888 22890 9897
rect 22834 9823 22890 9832
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22848 8974 22876 9318
rect 22940 9178 22968 9998
rect 23216 9674 23244 9998
rect 23308 9926 23336 10202
rect 23400 10130 23428 11222
rect 24044 11150 24072 12174
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11354 24164 11494
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23940 10600 23992 10606
rect 24044 10588 24072 11086
rect 23992 10560 24072 10588
rect 23940 10542 23992 10548
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23570 10364 23878 10373
rect 23570 10362 23576 10364
rect 23632 10362 23656 10364
rect 23712 10362 23736 10364
rect 23792 10362 23816 10364
rect 23872 10362 23878 10364
rect 23632 10310 23634 10362
rect 23814 10310 23816 10362
rect 23570 10308 23576 10310
rect 23632 10308 23656 10310
rect 23712 10308 23736 10310
rect 23792 10308 23816 10310
rect 23872 10308 23878 10310
rect 23570 10299 23878 10308
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23756 10056 23808 10062
rect 23952 10044 23980 10406
rect 24320 10130 24348 12174
rect 24412 11558 24440 12174
rect 24492 11824 24544 11830
rect 24596 11812 24624 12582
rect 24688 12442 24716 13126
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24780 12306 24808 13330
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24872 13190 24900 13262
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24964 12918 24992 13738
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24872 12481 24900 12650
rect 24858 12472 24914 12481
rect 25056 12434 25084 20198
rect 25332 19417 25360 20198
rect 25870 19952 25926 19961
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25792 19910 25870 19938
rect 25318 19408 25374 19417
rect 25318 19343 25374 19352
rect 25320 19304 25372 19310
rect 25240 19264 25320 19292
rect 25136 19236 25188 19242
rect 25136 19178 25188 19184
rect 25148 18630 25176 19178
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25148 18290 25176 18566
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25148 16658 25176 18022
rect 25240 17134 25268 19264
rect 25424 19292 25452 19858
rect 25372 19264 25452 19292
rect 25320 19246 25372 19252
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25608 18290 25636 18906
rect 25686 18456 25742 18465
rect 25686 18391 25688 18400
rect 25740 18391 25742 18400
rect 25688 18362 25740 18368
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25424 17338 25452 17478
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25240 16658 25268 17070
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25148 13734 25176 16594
rect 25240 15162 25268 16594
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25332 15366 25360 15438
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25240 14550 25268 15098
rect 25228 14544 25280 14550
rect 25228 14486 25280 14492
rect 25240 14278 25268 14486
rect 25332 14396 25360 15302
rect 25424 15162 25452 16390
rect 25516 15706 25544 16390
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25424 14822 25452 14894
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25412 14408 25464 14414
rect 25332 14368 25412 14396
rect 25412 14350 25464 14356
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25424 13734 25452 14350
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25136 13184 25188 13190
rect 25332 13161 25360 13670
rect 25424 13190 25452 13670
rect 25516 13530 25544 15302
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25516 13433 25544 13466
rect 25502 13424 25558 13433
rect 25502 13359 25558 13368
rect 25502 13288 25558 13297
rect 25608 13274 25636 18226
rect 25700 16776 25728 18362
rect 25792 17898 25820 19910
rect 25976 19922 26004 20896
rect 26070 20700 26378 20709
rect 26070 20698 26076 20700
rect 26132 20698 26156 20700
rect 26212 20698 26236 20700
rect 26292 20698 26316 20700
rect 26372 20698 26378 20700
rect 26132 20646 26134 20698
rect 26314 20646 26316 20698
rect 26070 20644 26076 20646
rect 26132 20644 26156 20646
rect 26212 20644 26236 20646
rect 26292 20644 26316 20646
rect 26372 20644 26378 20646
rect 26070 20635 26378 20644
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 25870 19887 25926 19896
rect 25964 19916 26016 19922
rect 25964 19858 26016 19864
rect 26160 19825 26188 20402
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26252 19922 26280 20334
rect 26240 19916 26292 19922
rect 26292 19876 26464 19904
rect 26240 19858 26292 19864
rect 26146 19816 26202 19825
rect 26146 19751 26202 19760
rect 26070 19612 26378 19621
rect 26070 19610 26076 19612
rect 26132 19610 26156 19612
rect 26212 19610 26236 19612
rect 26292 19610 26316 19612
rect 26372 19610 26378 19612
rect 26132 19558 26134 19610
rect 26314 19558 26316 19610
rect 26070 19556 26076 19558
rect 26132 19556 26156 19558
rect 26212 19556 26236 19558
rect 26292 19556 26316 19558
rect 26372 19556 26378 19558
rect 26070 19547 26378 19556
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26252 18970 26280 19450
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25976 18329 26004 18702
rect 26344 18630 26372 19314
rect 26436 19174 26464 19876
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 26528 19514 26556 19722
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26436 18766 26464 19110
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26070 18524 26378 18533
rect 26070 18522 26076 18524
rect 26132 18522 26156 18524
rect 26212 18522 26236 18524
rect 26292 18522 26316 18524
rect 26372 18522 26378 18524
rect 26132 18470 26134 18522
rect 26314 18470 26316 18522
rect 26070 18468 26076 18470
rect 26132 18468 26156 18470
rect 26212 18468 26236 18470
rect 26292 18468 26316 18470
rect 26372 18468 26378 18470
rect 26070 18459 26378 18468
rect 25962 18320 26018 18329
rect 25962 18255 26018 18264
rect 25976 18154 26004 18255
rect 25964 18148 26016 18154
rect 25964 18090 26016 18096
rect 26620 18086 26648 19110
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 25792 17870 25912 17898
rect 25700 16748 25820 16776
rect 25792 15366 25820 16748
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25700 14278 25728 14894
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25558 13246 25636 13274
rect 25502 13223 25558 13232
rect 25412 13184 25464 13190
rect 25136 13126 25188 13132
rect 25318 13152 25374 13161
rect 24858 12407 24914 12416
rect 24964 12406 25084 12434
rect 24768 12300 24820 12306
rect 24820 12260 24900 12288
rect 24768 12242 24820 12248
rect 24872 12209 24900 12260
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24544 11784 24624 11812
rect 24492 11766 24544 11772
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11150 24440 11494
rect 24584 11212 24636 11218
rect 24636 11172 24716 11200
rect 24584 11154 24636 11160
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24032 10056 24084 10062
rect 23952 10016 24032 10044
rect 23756 9998 23808 10004
rect 24032 9998 24084 10004
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23386 9888 23442 9897
rect 23386 9823 23442 9832
rect 23112 9648 23164 9654
rect 23216 9646 23336 9674
rect 23112 9590 23164 9596
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 23032 9178 23060 9454
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22388 8809 22416 8910
rect 22374 8800 22430 8809
rect 22374 8735 22430 8744
rect 22388 8430 22416 8735
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 7290 22140 7346
rect 22112 7262 22232 7290
rect 22204 7206 22232 7262
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22112 7018 22140 7142
rect 22296 7018 22324 7754
rect 22112 6990 22324 7018
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22020 6390 22048 6802
rect 22296 6780 22324 6990
rect 22388 6934 22416 8366
rect 22480 7546 22508 8502
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22572 7546 22600 7958
rect 22664 7818 22692 8910
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22480 7410 22692 7426
rect 22468 7404 22692 7410
rect 22520 7398 22692 7404
rect 22468 7346 22520 7352
rect 22560 7336 22612 7342
rect 22558 7304 22560 7313
rect 22612 7304 22614 7313
rect 22558 7239 22614 7248
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22376 6792 22428 6798
rect 22296 6752 22376 6780
rect 22428 6752 22508 6780
rect 22376 6734 22428 6740
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22008 6384 22060 6390
rect 22008 6326 22060 6332
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21836 5302 21864 5646
rect 21824 5296 21876 5302
rect 21824 5238 21876 5244
rect 21836 4826 21864 5238
rect 21928 5234 21956 6122
rect 22204 6118 22232 6598
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22388 5710 22416 6734
rect 22480 6633 22508 6752
rect 22466 6624 22522 6633
rect 22466 6559 22522 6568
rect 22572 6390 22600 7239
rect 22664 6798 22692 7398
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22756 6390 22784 8298
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22848 7002 22876 7822
rect 23032 7750 23060 9114
rect 23124 8566 23152 9590
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23216 8974 23244 9386
rect 23308 9110 23336 9646
rect 23296 9104 23348 9110
rect 23400 9092 23428 9823
rect 23768 9722 23796 9998
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23860 9654 23888 9862
rect 24044 9674 24072 9998
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24412 9722 24440 9862
rect 24400 9716 24452 9722
rect 23848 9648 23900 9654
rect 24044 9646 24164 9674
rect 24400 9658 24452 9664
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 23848 9590 23900 9596
rect 23940 9512 23992 9518
rect 23478 9480 23534 9489
rect 23940 9454 23992 9460
rect 23478 9415 23480 9424
rect 23532 9415 23534 9424
rect 23480 9386 23532 9392
rect 23952 9382 23980 9454
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23570 9276 23878 9285
rect 23570 9274 23576 9276
rect 23632 9274 23656 9276
rect 23712 9274 23736 9276
rect 23792 9274 23816 9276
rect 23872 9274 23878 9276
rect 23632 9222 23634 9274
rect 23814 9222 23816 9274
rect 23570 9220 23576 9222
rect 23632 9220 23656 9222
rect 23712 9220 23736 9222
rect 23792 9220 23816 9222
rect 23872 9220 23878 9222
rect 23570 9211 23878 9220
rect 23664 9172 23716 9178
rect 23584 9132 23664 9160
rect 23584 9092 23612 9132
rect 23664 9114 23716 9120
rect 23400 9064 23612 9092
rect 23296 9046 23348 9052
rect 23952 9042 23980 9318
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23388 8832 23440 8838
rect 23386 8800 23388 8809
rect 23440 8800 23442 8809
rect 23386 8735 23442 8744
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23018 7032 23074 7041
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 22940 6990 23018 7018
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22466 5944 22522 5953
rect 22466 5879 22522 5888
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22376 5568 22428 5574
rect 22296 5528 22376 5556
rect 22006 5400 22062 5409
rect 22006 5335 22062 5344
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 22020 5030 22048 5335
rect 22008 5024 22060 5030
rect 22296 5012 22324 5528
rect 22376 5510 22428 5516
rect 22480 5250 22508 5879
rect 22572 5302 22600 6326
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22848 5710 22876 6054
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22008 4966 22060 4972
rect 22112 4984 22324 5012
rect 22388 5222 22508 5250
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21548 4014 21600 4020
rect 21730 4040 21786 4049
rect 20732 3602 20760 4014
rect 21730 3975 21786 3984
rect 21730 3768 21786 3777
rect 21836 3738 21864 4762
rect 22112 4690 22140 4984
rect 22388 4842 22416 5222
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22480 5001 22508 5102
rect 22466 4992 22522 5001
rect 22466 4927 22522 4936
rect 22204 4814 22416 4842
rect 22572 4826 22600 5238
rect 22664 4826 22692 5646
rect 22940 5574 22968 6990
rect 23018 6967 23074 6976
rect 23216 6934 23244 7278
rect 23204 6928 23256 6934
rect 23018 6896 23074 6905
rect 23204 6870 23256 6876
rect 23308 6866 23336 8026
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23400 7206 23428 7890
rect 23492 7750 23520 8366
rect 24136 8294 24164 9646
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 24412 8566 24440 8774
rect 24400 8560 24452 8566
rect 24320 8520 24400 8548
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 23570 8188 23878 8197
rect 23570 8186 23576 8188
rect 23632 8186 23656 8188
rect 23712 8186 23736 8188
rect 23792 8186 23816 8188
rect 23872 8186 23878 8188
rect 23632 8134 23634 8186
rect 23814 8134 23816 8186
rect 23570 8132 23576 8134
rect 23632 8132 23656 8134
rect 23712 8132 23736 8134
rect 23792 8132 23816 8134
rect 23872 8132 23878 8134
rect 23570 8123 23878 8132
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 24044 7342 24072 8230
rect 24136 7954 24164 8230
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24032 7336 24084 7342
rect 24136 7313 24164 7890
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7478 24256 7686
rect 24320 7546 24348 8520
rect 24400 8502 24452 8508
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24412 7546 24440 8366
rect 24504 7954 24532 8842
rect 24492 7948 24544 7954
rect 24492 7890 24544 7896
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 24032 7278 24084 7284
rect 24122 7304 24178 7313
rect 24122 7239 24178 7248
rect 23388 7200 23440 7206
rect 24228 7154 24256 7414
rect 23388 7142 23440 7148
rect 23018 6831 23074 6840
rect 23296 6860 23348 6866
rect 23032 5778 23060 6831
rect 23296 6802 23348 6808
rect 23400 6458 23428 7142
rect 24136 7126 24256 7154
rect 23570 7100 23878 7109
rect 23570 7098 23576 7100
rect 23632 7098 23656 7100
rect 23712 7098 23736 7100
rect 23792 7098 23816 7100
rect 23872 7098 23878 7100
rect 23632 7046 23634 7098
rect 23814 7046 23816 7098
rect 23570 7044 23576 7046
rect 23632 7044 23656 7046
rect 23712 7044 23736 7046
rect 23792 7044 23816 7046
rect 23872 7044 23878 7046
rect 23570 7035 23878 7044
rect 24136 6633 24164 7126
rect 24320 7002 24348 7482
rect 24216 6996 24268 7002
rect 24216 6938 24268 6944
rect 24308 6996 24360 7002
rect 24308 6938 24360 6944
rect 24228 6662 24256 6938
rect 24306 6896 24362 6905
rect 24306 6831 24362 6840
rect 24216 6656 24268 6662
rect 24122 6624 24178 6633
rect 24216 6598 24268 6604
rect 24122 6559 24178 6568
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23110 6352 23166 6361
rect 23166 6310 23520 6338
rect 24136 6322 24164 6559
rect 23110 6287 23166 6296
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 22928 5568 22980 5574
rect 22928 5510 22980 5516
rect 23124 5234 23152 6190
rect 23492 6100 23520 6310
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24032 6180 24084 6186
rect 24032 6122 24084 6128
rect 23756 6112 23808 6118
rect 23492 6072 23756 6100
rect 23756 6054 23808 6060
rect 23570 6012 23878 6021
rect 23570 6010 23576 6012
rect 23632 6010 23656 6012
rect 23712 6010 23736 6012
rect 23792 6010 23816 6012
rect 23872 6010 23878 6012
rect 23632 5958 23634 6010
rect 23814 5958 23816 6010
rect 23570 5956 23576 5958
rect 23632 5956 23656 5958
rect 23712 5956 23736 5958
rect 23792 5956 23816 5958
rect 23872 5956 23878 5958
rect 23386 5944 23442 5953
rect 23570 5947 23878 5956
rect 23386 5879 23442 5888
rect 23400 5710 23428 5879
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23202 5536 23258 5545
rect 23202 5471 23258 5480
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 22756 4865 22784 5170
rect 22742 4856 22798 4865
rect 22560 4820 22612 4826
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 22204 3942 22232 4814
rect 22560 4762 22612 4768
rect 22652 4820 22704 4826
rect 22742 4791 22798 4800
rect 22652 4762 22704 4768
rect 22940 4729 22968 5170
rect 23216 5030 23244 5471
rect 23294 5264 23350 5273
rect 23294 5199 23296 5208
rect 23348 5199 23350 5208
rect 23296 5170 23348 5176
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 22926 4720 22982 4729
rect 22926 4655 22982 4664
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22282 4448 22338 4457
rect 22282 4383 22338 4392
rect 22296 4282 22324 4383
rect 22388 4282 22416 4490
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 21730 3703 21732 3712
rect 21784 3703 21786 3712
rect 21824 3732 21876 3738
rect 21732 3674 21784 3680
rect 21824 3674 21876 3680
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20640 3194 20668 3402
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20548 3058 20576 3130
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20732 2922 20760 3538
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20180 2106 20208 2314
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 21008 1970 21036 3334
rect 21070 3292 21378 3301
rect 21070 3290 21076 3292
rect 21132 3290 21156 3292
rect 21212 3290 21236 3292
rect 21292 3290 21316 3292
rect 21372 3290 21378 3292
rect 21132 3238 21134 3290
rect 21314 3238 21316 3290
rect 21070 3236 21076 3238
rect 21132 3236 21156 3238
rect 21212 3236 21236 3238
rect 21292 3236 21316 3238
rect 21372 3236 21378 3238
rect 21070 3227 21378 3236
rect 21928 3126 21956 3470
rect 21548 3120 21600 3126
rect 21178 3088 21234 3097
rect 21548 3062 21600 3068
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21178 3023 21234 3032
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 21100 2496 21128 2926
rect 21192 2854 21220 3023
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21180 2508 21232 2514
rect 21100 2468 21180 2496
rect 21180 2450 21232 2456
rect 21560 2446 21588 3062
rect 22020 2938 22048 3538
rect 21744 2910 22048 2938
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21070 2204 21378 2213
rect 21070 2202 21076 2204
rect 21132 2202 21156 2204
rect 21212 2202 21236 2204
rect 21292 2202 21316 2204
rect 21372 2202 21378 2204
rect 21132 2150 21134 2202
rect 21314 2150 21316 2202
rect 21070 2148 21076 2150
rect 21132 2148 21156 2150
rect 21212 2148 21236 2150
rect 21292 2148 21316 2150
rect 21372 2148 21378 2150
rect 21070 2139 21378 2148
rect 21652 2106 21680 2246
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 21546 2000 21602 2009
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 20996 1964 21048 1970
rect 21546 1935 21548 1944
rect 20996 1906 21048 1912
rect 21600 1935 21602 1944
rect 21548 1906 21600 1912
rect 19708 1760 19760 1766
rect 19708 1702 19760 1708
rect 20168 1760 20220 1766
rect 20168 1702 20220 1708
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 19720 1358 19748 1702
rect 20180 1358 20208 1702
rect 20824 1358 20852 1702
rect 19708 1352 19760 1358
rect 19708 1294 19760 1300
rect 20168 1352 20220 1358
rect 20168 1294 20220 1300
rect 20812 1352 20864 1358
rect 20812 1294 20864 1300
rect 19524 1284 19576 1290
rect 19524 1226 19576 1232
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 20352 1216 20404 1222
rect 20352 1158 20404 1164
rect 20996 1216 21048 1222
rect 20996 1158 21048 1164
rect 20088 1018 20116 1158
rect 20076 1012 20128 1018
rect 20076 954 20128 960
rect 16762 54 17080 82
rect 16762 -300 16818 54
rect 17590 -300 17646 160
rect 18418 -300 18474 160
rect 19246 -300 19302 160
rect 20074 82 20130 160
rect 20364 82 20392 1158
rect 20074 54 20392 82
rect 20902 82 20958 160
rect 21008 82 21036 1158
rect 21070 1116 21378 1125
rect 21070 1114 21076 1116
rect 21132 1114 21156 1116
rect 21212 1114 21236 1116
rect 21292 1114 21316 1116
rect 21372 1114 21378 1116
rect 21132 1062 21134 1114
rect 21314 1062 21316 1114
rect 21070 1060 21076 1062
rect 21132 1060 21156 1062
rect 21212 1060 21236 1062
rect 21292 1060 21316 1062
rect 21372 1060 21378 1062
rect 21070 1051 21378 1060
rect 21560 882 21588 1906
rect 21744 1358 21772 2910
rect 22020 2854 22048 2910
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21928 1902 21956 2790
rect 22296 2650 22324 3878
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 22112 2106 22140 2314
rect 22100 2100 22152 2106
rect 22100 2042 22152 2048
rect 21916 1896 21968 1902
rect 21916 1838 21968 1844
rect 22388 1766 22416 3402
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 22376 1760 22428 1766
rect 22376 1702 22428 1708
rect 22204 1358 22232 1702
rect 21732 1352 21784 1358
rect 21732 1294 21784 1300
rect 22192 1352 22244 1358
rect 22480 1340 22508 4422
rect 23124 4146 23152 4558
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 2990 22784 3538
rect 23124 3534 23152 3946
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 3194 23060 3334
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22572 1970 22600 2586
rect 23032 2038 23060 2790
rect 23216 2774 23244 4966
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23308 4593 23336 4626
rect 23294 4584 23350 4593
rect 23294 4519 23350 4528
rect 23492 4282 23520 4966
rect 23570 4924 23878 4933
rect 23570 4922 23576 4924
rect 23632 4922 23656 4924
rect 23712 4922 23736 4924
rect 23792 4922 23816 4924
rect 23872 4922 23878 4924
rect 23632 4870 23634 4922
rect 23814 4870 23816 4922
rect 23570 4868 23576 4870
rect 23632 4868 23656 4870
rect 23712 4868 23736 4870
rect 23792 4868 23816 4870
rect 23872 4868 23878 4870
rect 23570 4859 23878 4868
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23860 4185 23888 4762
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23846 4176 23902 4185
rect 23846 4111 23848 4120
rect 23900 4111 23902 4120
rect 23848 4082 23900 4088
rect 23952 4078 23980 4626
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23570 3836 23878 3845
rect 23570 3834 23576 3836
rect 23632 3834 23656 3836
rect 23712 3834 23736 3836
rect 23792 3834 23816 3836
rect 23872 3834 23878 3836
rect 23632 3782 23634 3834
rect 23814 3782 23816 3834
rect 23570 3780 23576 3782
rect 23632 3780 23656 3782
rect 23712 3780 23736 3782
rect 23792 3780 23816 3782
rect 23872 3780 23878 3782
rect 23386 3768 23442 3777
rect 23570 3771 23878 3780
rect 23386 3703 23388 3712
rect 23440 3703 23442 3712
rect 23388 3674 23440 3680
rect 23386 3632 23442 3641
rect 23952 3602 23980 4014
rect 23386 3567 23442 3576
rect 23940 3596 23992 3602
rect 23400 3516 23428 3567
rect 23940 3538 23992 3544
rect 24044 3534 24072 6122
rect 24214 6080 24270 6089
rect 24214 6015 24270 6024
rect 24228 5914 24256 6015
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24136 5137 24164 5170
rect 24122 5128 24178 5137
rect 24122 5063 24178 5072
rect 24124 4480 24176 4486
rect 24122 4448 24124 4457
rect 24176 4448 24178 4457
rect 24122 4383 24178 4392
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 23572 3528 23624 3534
rect 23400 3488 23572 3516
rect 23572 3470 23624 3476
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23756 3392 23808 3398
rect 23808 3352 23980 3380
rect 23756 3334 23808 3340
rect 23492 3126 23520 3334
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23124 2746 23244 2774
rect 23570 2748 23878 2757
rect 23570 2746 23576 2748
rect 23632 2746 23656 2748
rect 23712 2746 23736 2748
rect 23792 2746 23816 2748
rect 23872 2746 23878 2748
rect 23020 2032 23072 2038
rect 23020 1974 23072 1980
rect 22560 1964 22612 1970
rect 22560 1906 22612 1912
rect 22560 1352 22612 1358
rect 22480 1312 22560 1340
rect 22192 1294 22244 1300
rect 22560 1294 22612 1300
rect 23020 1352 23072 1358
rect 23124 1340 23152 2746
rect 23632 2694 23634 2746
rect 23814 2694 23816 2746
rect 23570 2692 23576 2694
rect 23632 2692 23656 2694
rect 23712 2692 23736 2694
rect 23792 2692 23816 2694
rect 23872 2692 23878 2694
rect 23570 2683 23878 2692
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23768 2106 23796 2382
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 23664 1896 23716 1902
rect 23952 1884 23980 3352
rect 24136 3058 24164 4218
rect 24228 3618 24256 5850
rect 24320 5710 24348 6831
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24412 5710 24440 6054
rect 24596 5914 24624 9658
rect 24688 6866 24716 11172
rect 24872 10810 24900 12135
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24872 10266 24900 10406
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24964 9722 24992 12406
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25056 11540 25084 12242
rect 25148 12238 25176 13126
rect 25412 13126 25464 13132
rect 25318 13087 25374 13096
rect 25320 12912 25372 12918
rect 25412 12912 25464 12918
rect 25320 12854 25372 12860
rect 25410 12880 25412 12889
rect 25464 12880 25466 12889
rect 25228 12776 25280 12782
rect 25226 12744 25228 12753
rect 25280 12744 25282 12753
rect 25226 12679 25282 12688
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25148 11694 25176 12174
rect 25136 11688 25188 11694
rect 25240 11676 25268 12679
rect 25332 11801 25360 12854
rect 25410 12815 25466 12824
rect 25608 12442 25636 13246
rect 25700 12782 25728 14214
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25792 12646 25820 15030
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25596 12436 25648 12442
rect 25516 12396 25596 12424
rect 25318 11792 25374 11801
rect 25318 11727 25374 11736
rect 25412 11688 25464 11694
rect 25240 11648 25412 11676
rect 25136 11630 25188 11636
rect 25412 11630 25464 11636
rect 25056 11512 25176 11540
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25056 9518 25084 10610
rect 25148 9926 25176 11512
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 24780 9178 24808 9454
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 25056 9081 25084 9318
rect 25136 9104 25188 9110
rect 25042 9072 25098 9081
rect 24860 9036 24912 9042
rect 25136 9046 25188 9052
rect 25240 9058 25268 9454
rect 25332 9178 25360 10746
rect 25412 10192 25464 10198
rect 25412 10134 25464 10140
rect 25424 9722 25452 10134
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25042 9007 25098 9016
rect 24860 8978 24912 8984
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24780 7410 24808 8366
rect 24872 8090 24900 8978
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24964 7546 24992 8774
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 25056 7342 25084 8230
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24766 6896 24822 6905
rect 24676 6860 24728 6866
rect 25042 6896 25098 6905
rect 24766 6831 24822 6840
rect 24964 6854 25042 6882
rect 24676 6802 24728 6808
rect 24780 6322 24808 6831
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24308 5704 24360 5710
rect 24306 5672 24308 5681
rect 24400 5704 24452 5710
rect 24360 5672 24362 5681
rect 24490 5672 24546 5681
rect 24452 5652 24490 5658
rect 24400 5646 24490 5652
rect 24412 5630 24490 5646
rect 24306 5607 24362 5616
rect 24490 5607 24546 5616
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24582 5536 24638 5545
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 24320 4146 24348 4966
rect 24412 4146 24440 5510
rect 24582 5471 24638 5480
rect 24490 5128 24546 5137
rect 24490 5063 24546 5072
rect 24504 5030 24532 5063
rect 24492 5024 24544 5030
rect 24596 5001 24624 5471
rect 24492 4966 24544 4972
rect 24582 4992 24638 5001
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24306 3632 24362 3641
rect 24228 3590 24306 3618
rect 24306 3567 24362 3576
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 24136 2514 24164 2994
rect 24228 2650 24256 3334
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24044 2106 24072 2314
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 23716 1856 23980 1884
rect 23664 1838 23716 1844
rect 23570 1660 23878 1669
rect 23570 1658 23576 1660
rect 23632 1658 23656 1660
rect 23712 1658 23736 1660
rect 23792 1658 23816 1660
rect 23872 1658 23878 1660
rect 23632 1606 23634 1658
rect 23814 1606 23816 1658
rect 23570 1604 23576 1606
rect 23632 1604 23656 1606
rect 23712 1604 23736 1606
rect 23792 1604 23816 1606
rect 23872 1604 23878 1606
rect 23570 1595 23878 1604
rect 24136 1358 24164 2450
rect 24228 1562 24256 2586
rect 24320 1834 24348 3062
rect 24504 2774 24532 4966
rect 24582 4927 24638 4936
rect 24596 4826 24624 4927
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 24688 4758 24716 6258
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24688 3482 24716 4694
rect 24780 4554 24808 6258
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24768 4548 24820 4554
rect 24768 4490 24820 4496
rect 24872 3942 24900 5510
rect 24964 4690 24992 6854
rect 25042 6831 25098 6840
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 5953 25084 6598
rect 25148 6458 25176 9046
rect 25240 9030 25360 9058
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8634 25268 8910
rect 25332 8838 25360 9030
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25228 7472 25280 7478
rect 25332 7460 25360 8774
rect 25424 7546 25452 9658
rect 25516 8906 25544 12396
rect 25596 12378 25648 12384
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25700 11762 25728 12106
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25700 11286 25728 11494
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 25608 10742 25636 10950
rect 25700 10810 25728 11222
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25596 10736 25648 10742
rect 25648 10684 25728 10690
rect 25596 10678 25728 10684
rect 25608 10662 25728 10678
rect 25596 10600 25648 10606
rect 25596 10542 25648 10548
rect 25608 9654 25636 10542
rect 25700 9994 25728 10662
rect 25792 10470 25820 11630
rect 25780 10464 25832 10470
rect 25780 10406 25832 10412
rect 25688 9988 25740 9994
rect 25688 9930 25740 9936
rect 25700 9654 25728 9930
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25700 9500 25728 9590
rect 25608 9472 25728 9500
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25516 8090 25544 8842
rect 25608 8401 25636 9472
rect 25792 9042 25820 10406
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25594 8392 25650 8401
rect 25594 8327 25650 8336
rect 25504 8084 25556 8090
rect 25504 8026 25556 8032
rect 25502 7848 25558 7857
rect 25502 7783 25558 7792
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25280 7432 25360 7460
rect 25228 7414 25280 7420
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25134 6352 25190 6361
rect 25134 6287 25190 6296
rect 25042 5944 25098 5953
rect 25148 5914 25176 6287
rect 25240 6118 25268 7278
rect 25332 6934 25360 7432
rect 25320 6928 25372 6934
rect 25320 6870 25372 6876
rect 25516 6610 25544 7783
rect 25608 6866 25636 8327
rect 25700 7886 25728 8434
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25778 7304 25834 7313
rect 25778 7239 25834 7248
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25594 6760 25650 6769
rect 25700 6746 25728 7142
rect 25650 6718 25728 6746
rect 25594 6695 25650 6704
rect 25332 6582 25544 6610
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25332 6390 25360 6582
rect 25410 6488 25466 6497
rect 25410 6423 25466 6432
rect 25504 6452 25556 6458
rect 25424 6390 25452 6423
rect 25504 6394 25556 6400
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25042 5879 25098 5888
rect 25136 5908 25188 5914
rect 25056 5710 25084 5879
rect 25136 5850 25188 5856
rect 25148 5817 25176 5850
rect 25134 5808 25190 5817
rect 25240 5778 25268 6054
rect 25134 5743 25190 5752
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25042 5400 25098 5409
rect 25042 5335 25098 5344
rect 25056 5166 25084 5335
rect 25134 5264 25190 5273
rect 25134 5199 25190 5208
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24964 3602 24992 4626
rect 25056 4593 25084 5102
rect 25148 4758 25176 5199
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25136 4752 25188 4758
rect 25136 4694 25188 4700
rect 25042 4584 25098 4593
rect 25042 4519 25098 4528
rect 25148 4214 25176 4694
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25240 4049 25268 4966
rect 25226 4040 25282 4049
rect 25226 3975 25282 3984
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24688 3454 24808 3482
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24688 3194 24716 3334
rect 24780 3194 24808 3454
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24504 2746 24624 2774
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24308 1828 24360 1834
rect 24308 1770 24360 1776
rect 24400 1828 24452 1834
rect 24400 1770 24452 1776
rect 24216 1556 24268 1562
rect 24216 1498 24268 1504
rect 23072 1312 23152 1340
rect 24124 1352 24176 1358
rect 23020 1294 23072 1300
rect 24124 1294 24176 1300
rect 21732 1216 21784 1222
rect 21732 1158 21784 1164
rect 22560 1216 22612 1222
rect 22560 1158 22612 1164
rect 23296 1216 23348 1222
rect 23296 1158 23348 1164
rect 21548 876 21600 882
rect 21548 818 21600 824
rect 21744 160 21772 1158
rect 22572 160 22600 1158
rect 20902 54 21036 82
rect 20074 -300 20130 54
rect 20902 -300 20958 54
rect 21730 -300 21786 160
rect 22558 -300 22614 160
rect 23308 82 23336 1158
rect 24412 898 24440 1770
rect 24504 1290 24532 1906
rect 24492 1284 24544 1290
rect 24492 1226 24544 1232
rect 24596 1018 24624 2746
rect 24780 2378 24808 3130
rect 25148 3097 25176 3402
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25134 3088 25190 3097
rect 25134 3023 25190 3032
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 24780 2038 24808 2314
rect 24768 2032 24820 2038
rect 24768 1974 24820 1980
rect 24780 1290 24808 1974
rect 25136 1828 25188 1834
rect 25136 1770 25188 1776
rect 25148 1426 25176 1770
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 24584 1012 24636 1018
rect 24584 954 24636 960
rect 25240 950 25268 3334
rect 25332 3074 25360 6326
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25424 3942 25452 5510
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25412 3392 25464 3398
rect 25516 3380 25544 6394
rect 25608 6225 25636 6598
rect 25594 6216 25650 6225
rect 25594 6151 25650 6160
rect 25608 5817 25636 6151
rect 25594 5808 25650 5817
rect 25594 5743 25650 5752
rect 25608 5642 25636 5743
rect 25596 5636 25648 5642
rect 25596 5578 25648 5584
rect 25700 5234 25728 6718
rect 25792 6458 25820 7239
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25884 6254 25912 17870
rect 26070 17436 26378 17445
rect 26070 17434 26076 17436
rect 26132 17434 26156 17436
rect 26212 17434 26236 17436
rect 26292 17434 26316 17436
rect 26372 17434 26378 17436
rect 26132 17382 26134 17434
rect 26314 17382 26316 17434
rect 26070 17380 26076 17382
rect 26132 17380 26156 17382
rect 26212 17380 26236 17382
rect 26292 17380 26316 17382
rect 26372 17380 26378 17382
rect 26070 17371 26378 17380
rect 26436 17270 26464 18022
rect 26620 17610 26648 18022
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26424 17264 26476 17270
rect 26424 17206 26476 17212
rect 26620 16658 26648 17546
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26070 16348 26378 16357
rect 26070 16346 26076 16348
rect 26132 16346 26156 16348
rect 26212 16346 26236 16348
rect 26292 16346 26316 16348
rect 26372 16346 26378 16348
rect 26132 16294 26134 16346
rect 26314 16294 26316 16346
rect 26070 16292 26076 16294
rect 26132 16292 26156 16294
rect 26212 16292 26236 16294
rect 26292 16292 26316 16294
rect 26372 16292 26378 16294
rect 26070 16283 26378 16292
rect 26332 16108 26384 16114
rect 26436 16096 26464 16594
rect 26712 16266 26740 21383
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 21010 27016 21286
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 27080 20874 27108 21830
rect 27160 21480 27212 21486
rect 27160 21422 27212 21428
rect 27172 21049 27200 21422
rect 27158 21040 27214 21049
rect 27158 20975 27160 20984
rect 27212 20975 27214 20984
rect 27160 20946 27212 20952
rect 27068 20868 27120 20874
rect 27068 20810 27120 20816
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 26882 18864 26938 18873
rect 26882 18799 26938 18808
rect 26792 18692 26844 18698
rect 26792 18634 26844 18640
rect 26804 17678 26832 18634
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26804 16998 26832 17614
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16436 26832 16934
rect 26896 16561 26924 18799
rect 27172 18698 27200 19110
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26988 18154 27016 18226
rect 26976 18148 27028 18154
rect 26976 18090 27028 18096
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27172 17678 27200 18022
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 26976 16584 27028 16590
rect 26882 16552 26938 16561
rect 26976 16526 27028 16532
rect 26882 16487 26938 16496
rect 26884 16448 26936 16454
rect 26804 16408 26884 16436
rect 26884 16390 26936 16396
rect 26712 16238 26832 16266
rect 26384 16068 26464 16096
rect 26332 16050 26384 16056
rect 26344 15434 26372 16050
rect 26514 16008 26570 16017
rect 26514 15943 26516 15952
rect 26568 15943 26570 15952
rect 26516 15914 26568 15920
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26332 15428 26384 15434
rect 26424 15428 26476 15434
rect 26384 15388 26424 15416
rect 26332 15370 26384 15376
rect 26424 15370 26476 15376
rect 26070 15260 26378 15269
rect 26070 15258 26076 15260
rect 26132 15258 26156 15260
rect 26212 15258 26236 15260
rect 26292 15258 26316 15260
rect 26372 15258 26378 15260
rect 26132 15206 26134 15258
rect 26314 15206 26316 15258
rect 26070 15204 26076 15206
rect 26132 15204 26156 15206
rect 26212 15204 26236 15206
rect 26292 15204 26316 15206
rect 26372 15204 26378 15206
rect 26070 15195 26378 15204
rect 26436 15042 26464 15370
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26528 15162 26556 15302
rect 26620 15162 26648 15506
rect 26804 15162 26832 16238
rect 26896 16046 26924 16390
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26792 15156 26844 15162
rect 26792 15098 26844 15104
rect 26240 15020 26292 15026
rect 26436 15014 26832 15042
rect 26240 14962 26292 14968
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25976 12306 26004 14758
rect 26252 14657 26280 14962
rect 26608 14952 26660 14958
rect 26528 14900 26608 14906
rect 26528 14894 26660 14900
rect 26528 14878 26648 14894
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26238 14648 26294 14657
rect 26238 14583 26294 14592
rect 26070 14172 26378 14181
rect 26070 14170 26076 14172
rect 26132 14170 26156 14172
rect 26212 14170 26236 14172
rect 26292 14170 26316 14172
rect 26372 14170 26378 14172
rect 26132 14118 26134 14170
rect 26314 14118 26316 14170
rect 26070 14116 26076 14118
rect 26132 14116 26156 14118
rect 26212 14116 26236 14118
rect 26292 14116 26316 14118
rect 26372 14116 26378 14118
rect 26070 14107 26378 14116
rect 26436 13394 26464 14758
rect 26528 13394 26556 14878
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26620 13530 26648 14214
rect 26712 14074 26740 14418
rect 26804 14414 26832 15014
rect 26896 14958 26924 15982
rect 26988 15638 27016 16526
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27080 15722 27108 16050
rect 27080 15706 27200 15722
rect 27080 15700 27212 15706
rect 27080 15694 27160 15700
rect 27160 15642 27212 15648
rect 26976 15632 27028 15638
rect 26976 15574 27028 15580
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26608 13524 26660 13530
rect 26804 13512 26832 14350
rect 26896 14074 26924 14758
rect 26988 14414 27016 15574
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 27172 15162 27200 15302
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27080 14618 27108 14962
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27172 14482 27200 14962
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27066 14376 27122 14385
rect 27066 14311 27122 14320
rect 27080 14090 27108 14311
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26988 14062 27108 14090
rect 27172 14074 27200 14418
rect 27160 14068 27212 14074
rect 26884 13524 26936 13530
rect 26804 13484 26884 13512
rect 26608 13466 26660 13472
rect 26884 13466 26936 13472
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26424 13252 26476 13258
rect 26424 13194 26476 13200
rect 26070 13084 26378 13093
rect 26070 13082 26076 13084
rect 26132 13082 26156 13084
rect 26212 13082 26236 13084
rect 26292 13082 26316 13084
rect 26372 13082 26378 13084
rect 26132 13030 26134 13082
rect 26314 13030 26316 13082
rect 26070 13028 26076 13030
rect 26132 13028 26156 13030
rect 26212 13028 26236 13030
rect 26292 13028 26316 13030
rect 26372 13028 26378 13030
rect 26070 13019 26378 13028
rect 26436 12918 26464 13194
rect 26424 12912 26476 12918
rect 26054 12880 26110 12889
rect 26424 12854 26476 12860
rect 26054 12815 26110 12824
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 26068 12084 26096 12815
rect 26620 12782 26648 13466
rect 26896 13326 26924 13466
rect 26988 13326 27016 14062
rect 27160 14010 27212 14016
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 27080 13530 27108 13874
rect 27158 13560 27214 13569
rect 27068 13524 27120 13530
rect 27158 13495 27160 13504
rect 27068 13466 27120 13472
rect 27212 13495 27214 13504
rect 27160 13466 27212 13472
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26804 12918 26832 13126
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26608 12776 26660 12782
rect 26608 12718 26660 12724
rect 26424 12708 26476 12714
rect 26424 12650 26476 12656
rect 26436 12345 26464 12650
rect 26528 12628 26556 12718
rect 26700 12640 26752 12646
rect 26528 12600 26648 12628
rect 26422 12336 26478 12345
rect 26422 12271 26478 12280
rect 25976 12056 26096 12084
rect 25976 11354 26004 12056
rect 26070 11996 26378 12005
rect 26070 11994 26076 11996
rect 26132 11994 26156 11996
rect 26212 11994 26236 11996
rect 26292 11994 26316 11996
rect 26372 11994 26378 11996
rect 26132 11942 26134 11994
rect 26314 11942 26316 11994
rect 26070 11940 26076 11942
rect 26132 11940 26156 11942
rect 26212 11940 26236 11942
rect 26292 11940 26316 11942
rect 26372 11940 26378 11942
rect 26070 11931 26378 11940
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26252 11354 26280 11630
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 25976 10674 26004 11154
rect 26070 10908 26378 10917
rect 26070 10906 26076 10908
rect 26132 10906 26156 10908
rect 26212 10906 26236 10908
rect 26292 10906 26316 10908
rect 26372 10906 26378 10908
rect 26132 10854 26134 10906
rect 26314 10854 26316 10906
rect 26070 10852 26076 10854
rect 26132 10852 26156 10854
rect 26212 10852 26236 10854
rect 26292 10852 26316 10854
rect 26372 10852 26378 10854
rect 26070 10843 26378 10852
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26160 10062 26188 10610
rect 26148 10056 26200 10062
rect 26148 9998 26200 10004
rect 26070 9820 26378 9829
rect 26070 9818 26076 9820
rect 26132 9818 26156 9820
rect 26212 9818 26236 9820
rect 26292 9818 26316 9820
rect 26372 9818 26378 9820
rect 26132 9766 26134 9818
rect 26314 9766 26316 9818
rect 26070 9764 26076 9766
rect 26132 9764 26156 9766
rect 26212 9764 26236 9766
rect 26292 9764 26316 9766
rect 26372 9764 26378 9766
rect 26070 9755 26378 9764
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25976 8838 26004 9114
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 26436 8786 26464 12271
rect 26516 12232 26568 12238
rect 26516 12174 26568 12180
rect 26528 11830 26556 12174
rect 26620 11830 26648 12600
rect 26700 12582 26752 12588
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26712 12238 26740 12582
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26712 9178 26740 9454
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26514 8936 26570 8945
rect 26514 8871 26516 8880
rect 26568 8871 26570 8880
rect 26516 8842 26568 8848
rect 25976 8430 26004 8774
rect 26436 8758 26556 8786
rect 26070 8732 26378 8741
rect 26070 8730 26076 8732
rect 26132 8730 26156 8732
rect 26212 8730 26236 8732
rect 26292 8730 26316 8732
rect 26372 8730 26378 8732
rect 26132 8678 26134 8730
rect 26314 8678 26316 8730
rect 26070 8676 26076 8678
rect 26132 8676 26156 8678
rect 26212 8676 26236 8678
rect 26292 8676 26316 8678
rect 26372 8676 26378 8678
rect 26070 8667 26378 8676
rect 26528 8634 26556 8758
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26804 8566 26832 12582
rect 26896 12306 26924 13262
rect 26974 12744 27030 12753
rect 26974 12679 26976 12688
rect 27028 12679 27030 12688
rect 26976 12650 27028 12656
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26882 11248 26938 11257
rect 26988 11218 27016 12038
rect 26882 11183 26938 11192
rect 26976 11212 27028 11218
rect 26896 8906 26924 11183
rect 26976 11154 27028 11160
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26792 8560 26844 8566
rect 26792 8502 26844 8508
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 26804 7993 26832 8502
rect 26988 8430 27016 8842
rect 26976 8424 27028 8430
rect 26976 8366 27028 8372
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26790 7984 26846 7993
rect 26790 7919 26846 7928
rect 26514 7848 26570 7857
rect 26514 7783 26570 7792
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 26070 7644 26378 7653
rect 26070 7642 26076 7644
rect 26132 7642 26156 7644
rect 26212 7642 26236 7644
rect 26292 7642 26316 7644
rect 26372 7642 26378 7644
rect 26132 7590 26134 7642
rect 26314 7590 26316 7642
rect 26070 7588 26076 7590
rect 26132 7588 26156 7590
rect 26212 7588 26236 7590
rect 26292 7588 26316 7590
rect 26372 7588 26378 7590
rect 26070 7579 26378 7588
rect 26436 7002 26464 7686
rect 26528 7546 26556 7783
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26620 7342 26648 7686
rect 26896 7546 26924 8230
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 26620 6934 26648 7278
rect 26608 6928 26660 6934
rect 26146 6896 26202 6905
rect 26608 6870 26660 6876
rect 26146 6831 26202 6840
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 25976 6458 26004 6734
rect 26160 6662 26188 6831
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 26070 6556 26378 6565
rect 26070 6554 26076 6556
rect 26132 6554 26156 6556
rect 26212 6554 26236 6556
rect 26292 6554 26316 6556
rect 26372 6554 26378 6556
rect 26132 6502 26134 6554
rect 26314 6502 26316 6554
rect 26070 6500 26076 6502
rect 26132 6500 26156 6502
rect 26212 6500 26236 6502
rect 26292 6500 26316 6502
rect 26372 6500 26378 6502
rect 26070 6491 26378 6500
rect 25964 6452 26016 6458
rect 26988 6440 27016 8366
rect 25964 6394 26016 6400
rect 26804 6412 27016 6440
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25792 5234 25820 5306
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25608 4282 25636 4490
rect 25688 4480 25740 4486
rect 25688 4422 25740 4428
rect 25596 4276 25648 4282
rect 25596 4218 25648 4224
rect 25464 3352 25544 3380
rect 25412 3334 25464 3340
rect 25332 3058 25452 3074
rect 25332 3052 25464 3058
rect 25332 3046 25412 3052
rect 25412 2994 25464 3000
rect 25608 2990 25636 4218
rect 25700 4146 25728 4422
rect 25792 4146 25820 4966
rect 25884 4214 25912 6054
rect 26056 5772 26108 5778
rect 25976 5732 26056 5760
rect 25976 5234 26004 5732
rect 26056 5714 26108 5720
rect 26070 5468 26378 5477
rect 26070 5466 26076 5468
rect 26132 5466 26156 5468
rect 26212 5466 26236 5468
rect 26292 5466 26316 5468
rect 26372 5466 26378 5468
rect 26132 5414 26134 5466
rect 26314 5414 26316 5466
rect 26070 5412 26076 5414
rect 26132 5412 26156 5414
rect 26212 5412 26236 5414
rect 26292 5412 26316 5414
rect 26372 5412 26378 5414
rect 26070 5403 26378 5412
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 26160 5030 26188 5306
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 26056 5024 26108 5030
rect 26056 4966 26108 4972
rect 26148 5024 26200 5030
rect 26148 4966 26200 4972
rect 26068 4865 26096 4966
rect 26054 4856 26110 4865
rect 26054 4791 26110 4800
rect 26344 4554 26372 5170
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 26332 4548 26384 4554
rect 26332 4490 26384 4496
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25976 4078 26004 4490
rect 26070 4380 26378 4389
rect 26070 4378 26076 4380
rect 26132 4378 26156 4380
rect 26212 4378 26236 4380
rect 26292 4378 26316 4380
rect 26372 4378 26378 4380
rect 26132 4326 26134 4378
rect 26314 4326 26316 4378
rect 26070 4324 26076 4326
rect 26132 4324 26156 4326
rect 26212 4324 26236 4326
rect 26292 4324 26316 4326
rect 26372 4324 26378 4326
rect 26070 4315 26378 4324
rect 26436 4282 26464 6190
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26608 6180 26660 6186
rect 26608 6122 26660 6128
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 25964 4072 26016 4078
rect 26528 4026 26556 6122
rect 25964 4014 26016 4020
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 26344 3998 26556 4026
rect 26620 4010 26648 6122
rect 26712 4282 26740 6258
rect 26804 5710 26832 6412
rect 27080 6338 27108 13330
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27172 12442 27200 12786
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 27264 9674 27292 22066
rect 27540 22030 27568 22374
rect 27632 22094 27660 22374
rect 28092 22098 28120 22510
rect 28570 22332 28878 22341
rect 28570 22330 28576 22332
rect 28632 22330 28656 22332
rect 28712 22330 28736 22332
rect 28792 22330 28816 22332
rect 28872 22330 28878 22332
rect 28632 22278 28634 22330
rect 28814 22278 28816 22330
rect 28570 22276 28576 22278
rect 28632 22276 28656 22278
rect 28712 22276 28736 22278
rect 28792 22276 28816 22278
rect 28872 22276 28878 22278
rect 28570 22267 28878 22276
rect 27632 22066 27752 22094
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27618 21992 27674 22001
rect 27618 21927 27674 21936
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27356 20602 27384 21014
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27540 20058 27568 21830
rect 27632 21690 27660 21927
rect 27724 21729 27752 22066
rect 27804 22092 27856 22098
rect 27804 22034 27856 22040
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 27710 21720 27766 21729
rect 27620 21684 27672 21690
rect 27710 21655 27766 21664
rect 27620 21626 27672 21632
rect 27816 21418 27844 22034
rect 28354 21992 28410 22001
rect 27896 21956 27948 21962
rect 28354 21927 28356 21936
rect 27896 21898 27948 21904
rect 28408 21927 28410 21936
rect 28356 21898 28408 21904
rect 27908 21486 27936 21898
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27804 21412 27856 21418
rect 27804 21354 27856 21360
rect 27816 21010 27844 21354
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 28000 20942 28028 21830
rect 28092 21350 28120 21830
rect 28264 21412 28316 21418
rect 28264 21354 28316 21360
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27632 20602 27660 20742
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27896 20528 27948 20534
rect 27710 20496 27766 20505
rect 27896 20470 27948 20476
rect 27710 20431 27766 20440
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19372 27488 19378
rect 27540 19360 27568 19994
rect 27632 19990 27660 20334
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27620 19372 27672 19378
rect 27540 19332 27620 19360
rect 27436 19314 27488 19320
rect 27620 19314 27672 19320
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27356 16658 27384 17478
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27356 15609 27384 16594
rect 27342 15600 27398 15609
rect 27342 15535 27398 15544
rect 27356 15026 27384 15535
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 13920 27384 14962
rect 27448 14906 27476 19314
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27540 17882 27568 18294
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27632 17542 27660 18294
rect 27724 17898 27752 20431
rect 27908 19854 27936 20470
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 28000 19854 28028 20334
rect 28092 20262 28120 20742
rect 28184 20534 28212 20878
rect 28276 20602 28304 21354
rect 28460 21128 28488 22034
rect 28908 22024 28960 22030
rect 28908 21966 28960 21972
rect 28920 21690 28948 21966
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28570 21244 28878 21253
rect 28570 21242 28576 21244
rect 28632 21242 28656 21244
rect 28712 21242 28736 21244
rect 28792 21242 28816 21244
rect 28872 21242 28878 21244
rect 28632 21190 28634 21242
rect 28814 21190 28816 21242
rect 28570 21188 28576 21190
rect 28632 21188 28656 21190
rect 28712 21188 28736 21190
rect 28792 21188 28816 21190
rect 28872 21188 28878 21190
rect 28570 21179 28878 21188
rect 28460 21100 28580 21128
rect 28356 21072 28408 21078
rect 28408 21032 28488 21060
rect 28356 21014 28408 21020
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28368 20602 28396 20810
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 28172 20392 28224 20398
rect 28172 20334 28224 20340
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28092 19718 28120 20198
rect 28184 20074 28212 20334
rect 28276 20262 28304 20538
rect 28460 20482 28488 21032
rect 28368 20454 28488 20482
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28368 20074 28396 20454
rect 28552 20380 28580 21100
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 28920 20942 28948 21014
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28724 20800 28776 20806
rect 28828 20788 28856 20878
rect 28828 20760 28948 20788
rect 28724 20742 28776 20748
rect 28736 20534 28764 20742
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 28184 20046 28396 20074
rect 28460 20352 28580 20380
rect 28184 19922 28212 20046
rect 28354 19952 28410 19961
rect 28172 19916 28224 19922
rect 28354 19887 28410 19896
rect 28172 19858 28224 19864
rect 28172 19780 28224 19786
rect 28172 19722 28224 19728
rect 28264 19780 28316 19786
rect 28264 19722 28316 19728
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 28080 19712 28132 19718
rect 28080 19654 28132 19660
rect 27816 18970 27844 19654
rect 28078 19544 28134 19553
rect 28078 19479 28134 19488
rect 28092 19378 28120 19479
rect 28184 19446 28212 19722
rect 28172 19440 28224 19446
rect 28276 19417 28304 19722
rect 28368 19514 28396 19887
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28172 19382 28224 19388
rect 28262 19408 28318 19417
rect 28080 19372 28132 19378
rect 28262 19343 28318 19352
rect 28080 19314 28132 19320
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27988 18896 28040 18902
rect 27988 18838 28040 18844
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27724 17870 27844 17898
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27632 16250 27660 16390
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27632 15570 27660 16186
rect 27724 16114 27752 16390
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27816 15722 27844 17870
rect 27908 17338 27936 18226
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27894 16688 27950 16697
rect 27894 16623 27950 16632
rect 27908 16590 27936 16623
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27724 15694 27844 15722
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27448 14878 27660 14906
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27434 14512 27490 14521
rect 27434 14447 27490 14456
rect 27448 14346 27476 14447
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27356 13892 27476 13920
rect 27344 13796 27396 13802
rect 27344 13738 27396 13744
rect 27356 13394 27384 13738
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27448 12646 27476 13892
rect 27540 12850 27568 14758
rect 27632 13190 27660 14878
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27618 13016 27674 13025
rect 27618 12951 27620 12960
rect 27672 12951 27674 12960
rect 27620 12922 27672 12928
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27724 12594 27752 15694
rect 27804 15564 27856 15570
rect 27804 15506 27856 15512
rect 27816 14482 27844 15506
rect 27908 15337 27936 16526
rect 27894 15328 27950 15337
rect 27894 15263 27950 15272
rect 27908 15026 27936 15263
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 27816 13870 27844 14418
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27816 12782 27844 13806
rect 27908 13190 27936 14962
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27896 12640 27948 12646
rect 27724 12566 27844 12594
rect 27896 12582 27948 12588
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27632 11354 27660 12038
rect 27724 11762 27752 12242
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27724 11082 27752 11698
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27172 9646 27292 9674
rect 27172 6905 27200 9646
rect 27632 9518 27660 10746
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27724 10062 27752 10610
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27724 9722 27752 9998
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27436 9036 27488 9042
rect 27436 8978 27488 8984
rect 27448 8430 27476 8978
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 27158 6896 27214 6905
rect 27158 6831 27214 6840
rect 27264 6780 27292 8230
rect 27448 7449 27476 8366
rect 27434 7440 27490 7449
rect 27434 7375 27490 7384
rect 26988 6310 27108 6338
rect 27172 6752 27292 6780
rect 27436 6792 27488 6798
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 26804 5370 26832 5646
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 26804 4690 26832 5306
rect 26988 5273 27016 6310
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 27080 5914 27108 6190
rect 27068 5908 27120 5914
rect 27068 5850 27120 5856
rect 27080 5710 27108 5850
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 26974 5264 27030 5273
rect 26974 5199 27030 5208
rect 27172 4865 27200 6752
rect 27540 6780 27568 9114
rect 27632 8838 27660 9454
rect 27620 8832 27672 8838
rect 27672 8792 27752 8820
rect 27620 8774 27672 8780
rect 27724 8498 27752 8792
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27632 8090 27660 8434
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27724 7002 27752 8434
rect 27712 6996 27764 7002
rect 27712 6938 27764 6944
rect 27816 6848 27844 12566
rect 27908 12306 27936 12582
rect 27896 12300 27948 12306
rect 27896 12242 27948 12248
rect 27896 12164 27948 12170
rect 27896 12106 27948 12112
rect 27908 11354 27936 12106
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 28000 10010 28028 18838
rect 28092 14385 28120 19314
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28172 18964 28224 18970
rect 28172 18906 28224 18912
rect 28184 16590 28212 18906
rect 28276 18766 28304 19110
rect 28460 18766 28488 20352
rect 28570 20156 28878 20165
rect 28570 20154 28576 20156
rect 28632 20154 28656 20156
rect 28712 20154 28736 20156
rect 28792 20154 28816 20156
rect 28872 20154 28878 20156
rect 28632 20102 28634 20154
rect 28814 20102 28816 20154
rect 28570 20100 28576 20102
rect 28632 20100 28656 20102
rect 28712 20100 28736 20102
rect 28792 20100 28816 20102
rect 28872 20100 28878 20102
rect 28570 20091 28878 20100
rect 28630 19952 28686 19961
rect 28630 19887 28686 19896
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28552 19378 28580 19654
rect 28644 19553 28672 19887
rect 28920 19718 28948 20760
rect 29012 20398 29040 22578
rect 29368 22568 29420 22574
rect 29368 22510 29420 22516
rect 29380 22234 29408 22510
rect 30300 22506 30328 23840
rect 31220 23338 31248 23840
rect 32140 23746 32168 23840
rect 32232 23746 32260 23854
rect 32140 23718 32260 23746
rect 31220 23310 31340 23338
rect 31312 23254 31340 23310
rect 31300 23248 31352 23254
rect 31300 23190 31352 23196
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 32404 22976 32456 22982
rect 32404 22918 32456 22924
rect 30668 22778 30696 22918
rect 31070 22876 31378 22885
rect 31070 22874 31076 22876
rect 31132 22874 31156 22876
rect 31212 22874 31236 22876
rect 31292 22874 31316 22876
rect 31372 22874 31378 22876
rect 31132 22822 31134 22874
rect 31314 22822 31316 22874
rect 31070 22820 31076 22822
rect 31132 22820 31156 22822
rect 31212 22820 31236 22822
rect 31292 22820 31316 22822
rect 31372 22820 31378 22822
rect 31070 22811 31378 22820
rect 30656 22772 30708 22778
rect 30656 22714 30708 22720
rect 32416 22710 32444 22918
rect 32404 22704 32456 22710
rect 32404 22646 32456 22652
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 30288 22500 30340 22506
rect 30288 22442 30340 22448
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 30024 21978 30052 22034
rect 30196 22024 30248 22030
rect 30024 21950 30144 21978
rect 30196 21966 30248 21972
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 29104 20777 29132 21830
rect 30024 21593 30052 21830
rect 30010 21584 30066 21593
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 29920 21548 29972 21554
rect 30010 21519 30066 21528
rect 29920 21490 29972 21496
rect 29184 20868 29236 20874
rect 29184 20810 29236 20816
rect 29090 20768 29146 20777
rect 29090 20703 29146 20712
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28630 19544 28686 19553
rect 28630 19479 28686 19488
rect 28540 19372 28592 19378
rect 28540 19314 28592 19320
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28570 19068 28878 19077
rect 28570 19066 28576 19068
rect 28632 19066 28656 19068
rect 28712 19066 28736 19068
rect 28792 19066 28816 19068
rect 28872 19066 28878 19068
rect 28632 19014 28634 19066
rect 28814 19014 28816 19066
rect 28570 19012 28576 19014
rect 28632 19012 28656 19014
rect 28712 19012 28736 19014
rect 28792 19012 28816 19014
rect 28872 19012 28878 19014
rect 28570 19003 28878 19012
rect 28920 18970 28948 19314
rect 28908 18964 28960 18970
rect 28908 18906 28960 18912
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28368 17270 28396 18566
rect 29104 18329 29132 20538
rect 29196 20505 29224 20810
rect 29380 20806 29408 21490
rect 29932 20913 29960 21490
rect 30116 21486 30144 21950
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30208 21418 30236 21966
rect 30196 21412 30248 21418
rect 30196 21354 30248 21360
rect 30300 20942 30328 21966
rect 30392 21690 30420 22578
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30378 21176 30434 21185
rect 30378 21111 30434 21120
rect 30288 20936 30340 20942
rect 29918 20904 29974 20913
rect 30288 20878 30340 20884
rect 29918 20839 29974 20848
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 29380 20602 29408 20742
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29182 20496 29238 20505
rect 29182 20431 29238 20440
rect 29184 20392 29236 20398
rect 29236 20352 29316 20380
rect 29184 20334 29236 20340
rect 29184 18896 29236 18902
rect 29184 18838 29236 18844
rect 29196 18426 29224 18838
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 29288 18358 29316 20352
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 29642 19544 29698 19553
rect 29642 19479 29698 19488
rect 29656 19446 29684 19479
rect 29644 19440 29696 19446
rect 29644 19382 29696 19388
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29736 19372 29788 19378
rect 29840 19360 29868 19654
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29788 19332 29868 19360
rect 29736 19314 29788 19320
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 29276 18352 29328 18358
rect 29090 18320 29146 18329
rect 29276 18294 29328 18300
rect 29090 18255 29146 18264
rect 28908 18216 28960 18222
rect 28908 18158 28960 18164
rect 28570 17980 28878 17989
rect 28570 17978 28576 17980
rect 28632 17978 28656 17980
rect 28712 17978 28736 17980
rect 28792 17978 28816 17980
rect 28872 17978 28878 17980
rect 28632 17926 28634 17978
rect 28814 17926 28816 17978
rect 28570 17924 28576 17926
rect 28632 17924 28656 17926
rect 28712 17924 28736 17926
rect 28792 17924 28816 17926
rect 28872 17924 28878 17926
rect 28570 17915 28878 17924
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28356 17264 28408 17270
rect 28356 17206 28408 17212
rect 28264 17196 28316 17202
rect 28264 17138 28316 17144
rect 28276 16794 28304 17138
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28356 16584 28408 16590
rect 28460 16574 28488 17750
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28552 17270 28580 17682
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28540 17264 28592 17270
rect 28540 17206 28592 17212
rect 28736 16998 28764 17478
rect 28724 16992 28776 16998
rect 28724 16934 28776 16940
rect 28570 16892 28878 16901
rect 28570 16890 28576 16892
rect 28632 16890 28656 16892
rect 28712 16890 28736 16892
rect 28792 16890 28816 16892
rect 28872 16890 28878 16892
rect 28632 16838 28634 16890
rect 28814 16838 28816 16890
rect 28570 16836 28576 16838
rect 28632 16836 28656 16838
rect 28712 16836 28736 16838
rect 28792 16836 28816 16838
rect 28872 16836 28878 16838
rect 28570 16827 28878 16836
rect 28408 16546 28488 16574
rect 28632 16584 28684 16590
rect 28356 16526 28408 16532
rect 28684 16544 28764 16572
rect 28632 16526 28684 16532
rect 28736 16250 28764 16544
rect 28920 16522 28948 18158
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17338 29040 18022
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 29012 16726 29040 16934
rect 29000 16720 29052 16726
rect 29000 16662 29052 16668
rect 28908 16516 28960 16522
rect 28908 16458 28960 16464
rect 28724 16244 28776 16250
rect 28724 16186 28776 16192
rect 28736 16114 28764 16186
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 28184 15502 28212 15574
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28276 15026 28304 16050
rect 28570 15804 28878 15813
rect 28570 15802 28576 15804
rect 28632 15802 28656 15804
rect 28712 15802 28736 15804
rect 28792 15802 28816 15804
rect 28872 15802 28878 15804
rect 28632 15750 28634 15802
rect 28814 15750 28816 15802
rect 28570 15748 28576 15750
rect 28632 15748 28656 15750
rect 28712 15748 28736 15750
rect 28792 15748 28816 15750
rect 28872 15748 28878 15750
rect 28570 15739 28878 15748
rect 28920 15706 28948 16458
rect 29104 16046 29132 18255
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29288 16998 29316 17138
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29472 16946 29500 19246
rect 29564 17338 29592 19314
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29656 18358 29684 19110
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29748 17762 29776 19314
rect 29826 18864 29882 18873
rect 29826 18799 29882 18808
rect 29840 18766 29868 18799
rect 29932 18766 29960 19450
rect 30024 19378 30052 19654
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29932 17882 29960 18702
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29748 17734 29868 17762
rect 29552 17332 29604 17338
rect 29552 17274 29604 17280
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29092 16040 29144 16046
rect 29090 16008 29092 16017
rect 29144 16008 29146 16017
rect 29090 15943 29146 15952
rect 29092 15904 29144 15910
rect 29092 15846 29144 15852
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28078 14376 28134 14385
rect 28078 14311 28134 14320
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 28092 13326 28120 14214
rect 28184 14074 28212 14758
rect 28276 14618 28304 14962
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14618 28396 14894
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28172 14068 28224 14074
rect 28172 14010 28224 14016
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12918 28120 13126
rect 28080 12912 28132 12918
rect 28080 12854 28132 12860
rect 28080 12096 28132 12102
rect 28080 12038 28132 12044
rect 28092 11898 28120 12038
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28092 10810 28120 11630
rect 28184 10810 28212 13738
rect 28276 13025 28304 14350
rect 28354 14104 28410 14113
rect 28460 14074 28488 15438
rect 28816 15360 28868 15366
rect 28868 15320 28948 15348
rect 28816 15302 28868 15308
rect 28570 14716 28878 14725
rect 28570 14714 28576 14716
rect 28632 14714 28656 14716
rect 28712 14714 28736 14716
rect 28792 14714 28816 14716
rect 28872 14714 28878 14716
rect 28632 14662 28634 14714
rect 28814 14662 28816 14714
rect 28570 14660 28576 14662
rect 28632 14660 28656 14662
rect 28712 14660 28736 14662
rect 28792 14660 28816 14662
rect 28872 14660 28878 14662
rect 28570 14651 28878 14660
rect 28920 14362 28948 15320
rect 29012 14414 29040 15574
rect 29104 15502 29132 15846
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29104 15337 29132 15438
rect 29090 15328 29146 15337
rect 29090 15263 29146 15272
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 28828 14334 28948 14362
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 28354 14039 28356 14048
rect 28408 14039 28410 14048
rect 28448 14068 28500 14074
rect 28356 14010 28408 14016
rect 28448 14010 28500 14016
rect 28368 13920 28396 14010
rect 28448 13932 28500 13938
rect 28368 13892 28448 13920
rect 28448 13874 28500 13880
rect 28828 13802 28856 14334
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28816 13796 28868 13802
rect 28816 13738 28868 13744
rect 28570 13628 28878 13637
rect 28570 13626 28576 13628
rect 28632 13626 28656 13628
rect 28712 13626 28736 13628
rect 28792 13626 28816 13628
rect 28872 13626 28878 13628
rect 28632 13574 28634 13626
rect 28814 13574 28816 13626
rect 28570 13572 28576 13574
rect 28632 13572 28656 13574
rect 28712 13572 28736 13574
rect 28792 13572 28816 13574
rect 28872 13572 28878 13574
rect 28570 13563 28878 13572
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28724 13524 28776 13530
rect 28724 13466 28776 13472
rect 28356 13456 28408 13462
rect 28356 13398 28408 13404
rect 28262 13016 28318 13025
rect 28368 12986 28396 13398
rect 28262 12951 28318 12960
rect 28356 12980 28408 12986
rect 28356 12922 28408 12928
rect 28368 12889 28396 12922
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 28460 12764 28488 13466
rect 28540 13388 28592 13394
rect 28540 13330 28592 13336
rect 28552 12850 28580 13330
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28736 13274 28764 13466
rect 28920 13394 28948 14214
rect 29012 14074 29040 14214
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 29104 13938 29132 14554
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29012 13818 29040 13874
rect 29090 13832 29146 13841
rect 29012 13790 29090 13818
rect 29090 13767 29146 13776
rect 28908 13388 28960 13394
rect 28908 13330 28960 13336
rect 28644 13190 28672 13262
rect 28736 13246 28948 13274
rect 28632 13184 28684 13190
rect 28632 13126 28684 13132
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28736 12968 28764 13126
rect 28644 12940 28764 12968
rect 28644 12850 28672 12940
rect 28920 12918 28948 13246
rect 29092 13252 29144 13258
rect 29092 13194 29144 13200
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 28540 12844 28592 12850
rect 28540 12786 28592 12792
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 29104 12764 29132 13194
rect 28276 12736 28488 12764
rect 28920 12736 29132 12764
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28276 10674 28304 12736
rect 28816 12708 28868 12714
rect 28460 12668 28816 12696
rect 28460 12306 28488 12668
rect 28816 12650 28868 12656
rect 28570 12540 28878 12549
rect 28570 12538 28576 12540
rect 28632 12538 28656 12540
rect 28712 12538 28736 12540
rect 28792 12538 28816 12540
rect 28872 12538 28878 12540
rect 28632 12486 28634 12538
rect 28814 12486 28816 12538
rect 28570 12484 28576 12486
rect 28632 12484 28656 12486
rect 28712 12484 28736 12486
rect 28792 12484 28816 12486
rect 28872 12484 28878 12486
rect 28570 12475 28878 12484
rect 28920 12442 28948 12736
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 28908 12436 28960 12442
rect 28908 12378 28960 12384
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28448 11824 28500 11830
rect 28448 11766 28500 11772
rect 28460 11354 28488 11766
rect 28570 11452 28878 11461
rect 28570 11450 28576 11452
rect 28632 11450 28656 11452
rect 28712 11450 28736 11452
rect 28792 11450 28816 11452
rect 28872 11450 28878 11452
rect 28632 11398 28634 11450
rect 28814 11398 28816 11450
rect 28570 11396 28576 11398
rect 28632 11396 28656 11398
rect 28712 11396 28736 11398
rect 28792 11396 28816 11398
rect 28872 11396 28878 11398
rect 28570 11387 28878 11396
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28276 10538 28304 10610
rect 28264 10532 28316 10538
rect 28264 10474 28316 10480
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 27908 9982 28028 10010
rect 27908 9178 27936 9982
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 28000 9586 28028 9862
rect 27988 9580 28040 9586
rect 27988 9522 28040 9528
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 28092 9042 28120 10406
rect 28368 10146 28396 10746
rect 28460 10266 28488 10950
rect 29104 10690 29132 12582
rect 29196 12209 29224 16390
rect 29288 16114 29316 16934
rect 29380 16590 29408 16934
rect 29472 16918 29684 16946
rect 29368 16584 29420 16590
rect 29368 16526 29420 16532
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29380 14929 29408 15098
rect 29366 14920 29422 14929
rect 29366 14855 29422 14864
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29288 13433 29316 14554
rect 29274 13424 29330 13433
rect 29274 13359 29330 13368
rect 29288 12782 29316 13359
rect 29368 13320 29420 13326
rect 29368 13262 29420 13268
rect 29380 12986 29408 13262
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29276 12776 29328 12782
rect 29276 12718 29328 12724
rect 29182 12200 29238 12209
rect 29472 12186 29500 16918
rect 29552 16516 29604 16522
rect 29552 16458 29604 16464
rect 29564 16250 29592 16458
rect 29552 16244 29604 16250
rect 29552 16186 29604 16192
rect 29564 15502 29592 16186
rect 29656 15502 29684 16918
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 29748 15706 29776 15982
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29736 15496 29788 15502
rect 29840 15484 29868 17734
rect 29918 17640 29974 17649
rect 29918 17575 29974 17584
rect 29932 17066 29960 17575
rect 29920 17060 29972 17066
rect 29920 17002 29972 17008
rect 29920 16584 29972 16590
rect 29920 16526 29972 16532
rect 29788 15456 29868 15484
rect 29736 15438 29788 15444
rect 29564 12986 29592 15438
rect 29748 15366 29776 15438
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29932 15026 29960 16526
rect 30024 15162 30052 18158
rect 30116 16250 30144 20742
rect 30300 20398 30328 20878
rect 30392 20534 30420 21111
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30300 19854 30328 20334
rect 30484 20330 30512 22578
rect 30944 22094 30972 22578
rect 30852 22066 30972 22094
rect 30564 21956 30616 21962
rect 30564 21898 30616 21904
rect 30576 21078 30604 21898
rect 30746 21584 30802 21593
rect 30656 21548 30708 21554
rect 30746 21519 30748 21528
rect 30656 21490 30708 21496
rect 30800 21519 30802 21528
rect 30748 21490 30800 21496
rect 30564 21072 30616 21078
rect 30564 21014 30616 21020
rect 30576 20534 30604 21014
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30472 20324 30524 20330
rect 30472 20266 30524 20272
rect 30564 20324 30616 20330
rect 30564 20266 30616 20272
rect 30378 20088 30434 20097
rect 30378 20023 30434 20032
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30196 19440 30248 19446
rect 30196 19382 30248 19388
rect 30208 18680 30236 19382
rect 30392 18834 30420 20023
rect 30470 19408 30526 19417
rect 30470 19343 30526 19352
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30208 18652 30328 18680
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 30208 17610 30236 18362
rect 30196 17604 30248 17610
rect 30196 17546 30248 17552
rect 30104 16244 30156 16250
rect 30104 16186 30156 16192
rect 30116 15502 30144 16186
rect 30208 16182 30236 17546
rect 30300 16454 30328 18652
rect 30484 17678 30512 19343
rect 30576 19258 30604 20266
rect 30668 19990 30696 21490
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 30760 21146 30788 21354
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30746 20632 30802 20641
rect 30746 20567 30802 20576
rect 30760 20233 30788 20567
rect 30852 20262 30880 22066
rect 30932 21956 30984 21962
rect 30932 21898 30984 21904
rect 30944 21350 30972 21898
rect 31070 21788 31378 21797
rect 31070 21786 31076 21788
rect 31132 21786 31156 21788
rect 31212 21786 31236 21788
rect 31292 21786 31316 21788
rect 31372 21786 31378 21788
rect 31132 21734 31134 21786
rect 31314 21734 31316 21786
rect 31070 21732 31076 21734
rect 31132 21732 31156 21734
rect 31212 21732 31236 21734
rect 31292 21732 31316 21734
rect 31372 21732 31378 21734
rect 31070 21723 31378 21732
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 31036 20788 31064 21490
rect 31392 21480 31444 21486
rect 31114 21448 31170 21457
rect 31444 21440 31524 21468
rect 31392 21422 31444 21428
rect 31114 21383 31170 21392
rect 31128 20942 31156 21383
rect 31496 21010 31524 21440
rect 31484 21004 31536 21010
rect 31484 20946 31536 20952
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 30944 20760 31064 20788
rect 30944 20584 30972 20760
rect 31070 20700 31378 20709
rect 31070 20698 31076 20700
rect 31132 20698 31156 20700
rect 31212 20698 31236 20700
rect 31292 20698 31316 20700
rect 31372 20698 31378 20700
rect 31132 20646 31134 20698
rect 31314 20646 31316 20698
rect 31070 20644 31076 20646
rect 31132 20644 31156 20646
rect 31212 20644 31236 20646
rect 31292 20644 31316 20646
rect 31372 20644 31378 20646
rect 31070 20635 31378 20644
rect 31496 20618 31524 20946
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 20806 31800 20878
rect 31864 20874 31892 22578
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 32128 22568 32180 22574
rect 32128 22510 32180 22516
rect 32048 22166 32076 22510
rect 32036 22160 32088 22166
rect 32036 22102 32088 22108
rect 32140 21350 32168 22510
rect 32416 22137 32444 22646
rect 32600 22574 32628 23854
rect 33046 23840 33102 24300
rect 33966 23840 34022 24300
rect 34886 23840 34942 24300
rect 35806 23840 35862 24300
rect 36726 23840 36782 24300
rect 37646 23840 37702 24300
rect 37752 23854 38056 23882
rect 32864 23112 32916 23118
rect 32864 23054 32916 23060
rect 32588 22568 32640 22574
rect 32588 22510 32640 22516
rect 32496 22160 32548 22166
rect 32402 22128 32458 22137
rect 32496 22102 32548 22108
rect 32680 22160 32732 22166
rect 32680 22102 32732 22108
rect 32402 22063 32458 22072
rect 32508 22030 32536 22102
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32692 21962 32720 22102
rect 32876 22098 32904 23054
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32968 22137 32996 22578
rect 32954 22128 33010 22137
rect 32864 22092 32916 22098
rect 32954 22063 33010 22072
rect 32864 22034 32916 22040
rect 32680 21956 32732 21962
rect 32680 21898 32732 21904
rect 32312 21888 32364 21894
rect 32312 21830 32364 21836
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32324 21486 32352 21830
rect 32600 21690 32628 21830
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32220 21480 32272 21486
rect 32220 21422 32272 21428
rect 32312 21480 32364 21486
rect 32364 21440 32444 21468
rect 32312 21422 32364 21428
rect 31944 21344 31996 21350
rect 31944 21286 31996 21292
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 31956 21146 31984 21286
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31760 20800 31812 20806
rect 31760 20742 31812 20748
rect 31404 20590 31524 20618
rect 30944 20556 31340 20584
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 30840 20256 30892 20262
rect 30746 20224 30802 20233
rect 30840 20198 30892 20204
rect 30746 20159 30802 20168
rect 31036 20097 31064 20334
rect 31022 20088 31078 20097
rect 31022 20023 31078 20032
rect 30656 19984 30708 19990
rect 31128 19938 31156 20402
rect 30656 19926 30708 19932
rect 30760 19910 31156 19938
rect 30760 19854 30788 19910
rect 30748 19848 30800 19854
rect 31116 19848 31168 19854
rect 30748 19790 30800 19796
rect 30852 19808 31116 19836
rect 30748 19712 30800 19718
rect 30748 19654 30800 19660
rect 30576 19230 30696 19258
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30576 17814 30604 19110
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30472 17672 30524 17678
rect 30472 17614 30524 17620
rect 30484 17513 30512 17614
rect 30564 17536 30616 17542
rect 30470 17504 30526 17513
rect 30564 17478 30616 17484
rect 30470 17439 30526 17448
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30472 17332 30524 17338
rect 30472 17274 30524 17280
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 30196 15428 30248 15434
rect 30196 15370 30248 15376
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 29656 13530 29684 14962
rect 30208 14958 30236 15370
rect 30392 15366 30420 17274
rect 30484 15434 30512 17274
rect 30576 17202 30604 17478
rect 30668 17320 30696 19230
rect 30760 19009 30788 19654
rect 30852 19514 30880 19808
rect 31116 19790 31168 19796
rect 31312 19700 31340 20556
rect 31404 20330 31432 20590
rect 31668 20460 31720 20466
rect 31588 20420 31668 20448
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 30944 19672 31340 19700
rect 31484 19712 31536 19718
rect 30944 19553 30972 19672
rect 31484 19654 31536 19660
rect 31070 19612 31378 19621
rect 31070 19610 31076 19612
rect 31132 19610 31156 19612
rect 31212 19610 31236 19612
rect 31292 19610 31316 19612
rect 31372 19610 31378 19612
rect 31132 19558 31134 19610
rect 31314 19558 31316 19610
rect 31070 19556 31076 19558
rect 31132 19556 31156 19558
rect 31212 19556 31236 19558
rect 31292 19556 31316 19558
rect 31372 19556 31378 19558
rect 30930 19544 30986 19553
rect 31070 19547 31378 19556
rect 30840 19508 30892 19514
rect 31496 19496 31524 19654
rect 30930 19479 30986 19488
rect 30840 19450 30892 19456
rect 30840 19304 30892 19310
rect 30840 19246 30892 19252
rect 30746 19000 30802 19009
rect 30746 18935 30802 18944
rect 30852 18834 30880 19246
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30760 18426 30788 18634
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30840 18352 30892 18358
rect 30840 18294 30892 18300
rect 30852 17610 30880 18294
rect 30944 18222 30972 19479
rect 31404 19468 31524 19496
rect 31404 19378 31432 19468
rect 31588 19428 31616 20420
rect 31668 20402 31720 20408
rect 31852 20460 31904 20466
rect 31852 20402 31904 20408
rect 31666 20224 31722 20233
rect 31666 20159 31722 20168
rect 31680 19514 31708 20159
rect 31864 19922 31892 20402
rect 31956 20380 31984 21082
rect 32140 21049 32168 21286
rect 32232 21146 32260 21422
rect 32220 21140 32272 21146
rect 32220 21082 32272 21088
rect 32126 21040 32182 21049
rect 32126 20975 32182 20984
rect 32036 20596 32088 20602
rect 32036 20538 32088 20544
rect 32048 20505 32076 20538
rect 32034 20496 32090 20505
rect 32034 20431 32090 20440
rect 31956 20352 32076 20380
rect 31852 19916 31904 19922
rect 31852 19858 31904 19864
rect 31944 19712 31996 19718
rect 31944 19654 31996 19660
rect 31668 19508 31720 19514
rect 31852 19508 31904 19514
rect 31668 19450 31720 19456
rect 31772 19468 31852 19496
rect 31496 19400 31616 19428
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 31116 19304 31168 19310
rect 31116 19246 31168 19252
rect 31128 18630 31156 19246
rect 31312 19174 31340 19314
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 31070 18524 31378 18533
rect 31070 18522 31076 18524
rect 31132 18522 31156 18524
rect 31212 18522 31236 18524
rect 31292 18522 31316 18524
rect 31372 18522 31378 18524
rect 31132 18470 31134 18522
rect 31314 18470 31316 18522
rect 31070 18468 31076 18470
rect 31132 18468 31156 18470
rect 31212 18468 31236 18470
rect 31292 18468 31316 18470
rect 31372 18468 31378 18470
rect 31070 18459 31378 18468
rect 31496 18290 31524 19400
rect 31772 19334 31800 19468
rect 31852 19450 31904 19456
rect 31588 19306 31800 19334
rect 31588 19242 31616 19306
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 31576 19236 31628 19242
rect 31576 19178 31628 19184
rect 31574 19000 31630 19009
rect 31574 18935 31630 18944
rect 31484 18284 31536 18290
rect 31484 18226 31536 18232
rect 30932 18216 30984 18222
rect 30932 18158 30984 18164
rect 31206 18184 31262 18193
rect 31206 18119 31262 18128
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 31128 17882 31156 18022
rect 31220 17882 31248 18119
rect 31588 17882 31616 18935
rect 31864 18902 31892 19246
rect 31956 18970 31984 19654
rect 31944 18964 31996 18970
rect 31944 18906 31996 18912
rect 31852 18896 31904 18902
rect 31852 18838 31904 18844
rect 31760 18828 31812 18834
rect 31680 18788 31760 18816
rect 31680 18290 31708 18788
rect 31760 18770 31812 18776
rect 31956 18442 31984 18906
rect 32048 18902 32076 20352
rect 32310 20360 32366 20369
rect 32310 20295 32312 20304
rect 32364 20295 32366 20304
rect 32312 20266 32364 20272
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32036 18896 32088 18902
rect 32036 18838 32088 18844
rect 31864 18414 31984 18442
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31760 18284 31812 18290
rect 31864 18272 31892 18414
rect 31812 18244 31892 18272
rect 31760 18226 31812 18232
rect 31116 17876 31168 17882
rect 31116 17818 31168 17824
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 31576 17876 31628 17882
rect 31576 17818 31628 17824
rect 31588 17649 31616 17818
rect 31680 17814 31708 18226
rect 32048 18222 32076 18838
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 32140 18358 32168 18566
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32036 18216 32088 18222
rect 32036 18158 32088 18164
rect 31668 17808 31720 17814
rect 31668 17750 31720 17756
rect 31852 17808 31904 17814
rect 31852 17750 31904 17756
rect 31574 17640 31630 17649
rect 30840 17604 30892 17610
rect 31574 17575 31630 17584
rect 30840 17546 30892 17552
rect 30852 17338 30880 17546
rect 31484 17536 31536 17542
rect 31484 17478 31536 17484
rect 31070 17436 31378 17445
rect 31070 17434 31076 17436
rect 31132 17434 31156 17436
rect 31212 17434 31236 17436
rect 31292 17434 31316 17436
rect 31372 17434 31378 17436
rect 31132 17382 31134 17434
rect 31314 17382 31316 17434
rect 31070 17380 31076 17382
rect 31132 17380 31156 17382
rect 31212 17380 31236 17382
rect 31292 17380 31316 17382
rect 31372 17380 31378 17382
rect 31070 17371 31378 17380
rect 30840 17332 30892 17338
rect 30668 17292 30788 17320
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30564 17060 30616 17066
rect 30564 17002 30616 17008
rect 30576 16590 30604 17002
rect 30668 16794 30696 17138
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30564 16584 30616 16590
rect 30564 16526 30616 16532
rect 30668 15706 30696 16594
rect 30656 15700 30708 15706
rect 30576 15660 30656 15688
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30484 15162 30512 15370
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 29734 14376 29790 14385
rect 29734 14311 29790 14320
rect 29748 14090 29776 14311
rect 30300 14278 30328 15030
rect 30576 14822 30604 15660
rect 30656 15642 30708 15648
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 30668 15162 30696 15506
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30656 14952 30708 14958
rect 30656 14894 30708 14900
rect 30564 14816 30616 14822
rect 30564 14758 30616 14764
rect 30668 14482 30696 14894
rect 30760 14618 30788 17292
rect 30840 17274 30892 17280
rect 31024 17196 31076 17202
rect 30852 17156 31024 17184
rect 30852 16454 30880 17156
rect 31024 17138 31076 17144
rect 31116 16992 31168 16998
rect 31116 16934 31168 16940
rect 31128 16794 31156 16934
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31496 16658 31524 17478
rect 31680 16794 31708 17750
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31772 17338 31800 17614
rect 31760 17332 31812 17338
rect 31760 17274 31812 17280
rect 31758 17232 31814 17241
rect 31864 17202 31892 17750
rect 32140 17542 32168 18294
rect 32232 17746 32260 19382
rect 32416 18766 32444 21440
rect 32864 21412 32916 21418
rect 32864 21354 32916 21360
rect 32876 21146 32904 21354
rect 32864 21140 32916 21146
rect 32864 21082 32916 21088
rect 32586 21040 32642 21049
rect 32586 20975 32642 20984
rect 32600 20874 32628 20975
rect 32588 20868 32640 20874
rect 32588 20810 32640 20816
rect 32968 20777 32996 22063
rect 33060 22030 33088 23840
rect 33600 23248 33652 23254
rect 33980 23236 34008 23840
rect 34060 23248 34112 23254
rect 33980 23208 34060 23236
rect 33600 23190 33652 23196
rect 34060 23190 34112 23196
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 33428 22778 33456 22986
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 33612 22642 33640 23190
rect 34612 23112 34664 23118
rect 34612 23054 34664 23060
rect 33600 22636 33652 22642
rect 33600 22578 33652 22584
rect 34624 22574 34652 23054
rect 34900 22710 34928 23840
rect 35072 23248 35124 23254
rect 35072 23190 35124 23196
rect 34888 22704 34940 22710
rect 34888 22646 34940 22652
rect 35084 22642 35112 23190
rect 35072 22636 35124 22642
rect 35820 22624 35848 23840
rect 36740 23236 36768 23840
rect 37660 23746 37688 23840
rect 37752 23746 37780 23854
rect 37660 23718 37780 23746
rect 36740 23208 36952 23236
rect 36070 22876 36378 22885
rect 36070 22874 36076 22876
rect 36132 22874 36156 22876
rect 36212 22874 36236 22876
rect 36292 22874 36316 22876
rect 36372 22874 36378 22876
rect 36132 22822 36134 22874
rect 36314 22822 36316 22874
rect 36070 22820 36076 22822
rect 36132 22820 36156 22822
rect 36212 22820 36236 22822
rect 36292 22820 36316 22822
rect 36372 22820 36378 22822
rect 36070 22811 36378 22820
rect 36924 22710 36952 23208
rect 36912 22704 36964 22710
rect 36912 22646 36964 22652
rect 38028 22658 38056 23854
rect 38566 23840 38622 24300
rect 39486 23840 39542 24300
rect 40406 23840 40462 24300
rect 41326 23840 41382 24300
rect 41432 23854 41644 23882
rect 38580 23236 38608 23840
rect 38580 23208 38700 23236
rect 38672 22710 38700 23208
rect 38292 22704 38344 22710
rect 38028 22652 38292 22658
rect 38028 22646 38344 22652
rect 38660 22704 38712 22710
rect 38660 22646 38712 22652
rect 35992 22636 36044 22642
rect 35820 22596 35992 22624
rect 35072 22578 35124 22584
rect 35992 22578 36044 22584
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37648 22636 37700 22642
rect 38028 22630 38332 22646
rect 39500 22642 39528 23840
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 38384 22636 38436 22642
rect 37648 22578 37700 22584
rect 38384 22578 38436 22584
rect 39488 22636 39540 22642
rect 39488 22578 39540 22584
rect 34060 22568 34112 22574
rect 34060 22510 34112 22516
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 37096 22568 37148 22574
rect 37096 22510 37148 22516
rect 33140 22432 33192 22438
rect 33508 22432 33560 22438
rect 33140 22374 33192 22380
rect 33428 22392 33508 22420
rect 33152 22234 33180 22374
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33336 21486 33364 22034
rect 33428 22001 33456 22392
rect 33508 22374 33560 22380
rect 33968 22432 34020 22438
rect 33968 22374 34020 22380
rect 33570 22332 33878 22341
rect 33570 22330 33576 22332
rect 33632 22330 33656 22332
rect 33712 22330 33736 22332
rect 33792 22330 33816 22332
rect 33872 22330 33878 22332
rect 33632 22278 33634 22330
rect 33814 22278 33816 22330
rect 33570 22276 33576 22278
rect 33632 22276 33656 22278
rect 33712 22276 33736 22278
rect 33792 22276 33816 22278
rect 33872 22276 33878 22278
rect 33570 22267 33878 22276
rect 33980 22234 34008 22374
rect 33968 22228 34020 22234
rect 33968 22170 34020 22176
rect 34072 22094 34100 22510
rect 33704 22066 34100 22094
rect 33414 21992 33470 22001
rect 33414 21927 33470 21936
rect 33140 21480 33192 21486
rect 33140 21422 33192 21428
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 33048 21344 33100 21350
rect 33048 21286 33100 21292
rect 33060 21146 33088 21286
rect 33048 21140 33100 21146
rect 33048 21082 33100 21088
rect 33152 21078 33180 21422
rect 33704 21350 33732 22066
rect 33876 22024 33928 22030
rect 33876 21966 33928 21972
rect 33888 21690 33916 21966
rect 33876 21684 33928 21690
rect 33876 21626 33928 21632
rect 34060 21616 34112 21622
rect 34060 21558 34112 21564
rect 34072 21486 34100 21558
rect 34060 21480 34112 21486
rect 34060 21422 34112 21428
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33692 21344 33744 21350
rect 33692 21286 33744 21292
rect 33140 21072 33192 21078
rect 33244 21049 33272 21286
rect 33140 21014 33192 21020
rect 33230 21040 33286 21049
rect 33428 21010 33456 21286
rect 33570 21244 33878 21253
rect 33570 21242 33576 21244
rect 33632 21242 33656 21244
rect 33712 21242 33736 21244
rect 33792 21242 33816 21244
rect 33872 21242 33878 21244
rect 33632 21190 33634 21242
rect 33814 21190 33816 21242
rect 33570 21188 33576 21190
rect 33632 21188 33656 21190
rect 33712 21188 33736 21190
rect 33792 21188 33816 21190
rect 33872 21188 33878 21190
rect 33570 21179 33878 21188
rect 34520 21140 34572 21146
rect 34520 21082 34572 21088
rect 33230 20975 33286 20984
rect 33324 21004 33376 21010
rect 33244 20806 33272 20975
rect 33324 20946 33376 20952
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33968 21004 34020 21010
rect 33968 20946 34020 20952
rect 33232 20800 33284 20806
rect 32954 20768 33010 20777
rect 33232 20742 33284 20748
rect 32954 20703 33010 20712
rect 32770 20632 32826 20641
rect 32770 20567 32826 20576
rect 33232 20596 33284 20602
rect 32494 19816 32550 19825
rect 32784 19786 32812 20567
rect 33232 20538 33284 20544
rect 32956 20528 33008 20534
rect 32954 20496 32956 20505
rect 33008 20496 33010 20505
rect 32954 20431 33010 20440
rect 33140 20392 33192 20398
rect 33244 20369 33272 20538
rect 33336 20398 33364 20946
rect 33416 20868 33468 20874
rect 33416 20810 33468 20816
rect 33428 20602 33456 20810
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33980 20534 34008 20946
rect 34060 20800 34112 20806
rect 34060 20742 34112 20748
rect 34072 20602 34100 20742
rect 34532 20602 34560 21082
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34520 20596 34572 20602
rect 34520 20538 34572 20544
rect 33968 20528 34020 20534
rect 33968 20470 34020 20476
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 33324 20392 33376 20398
rect 33140 20334 33192 20340
rect 33230 20360 33286 20369
rect 33152 20058 33180 20334
rect 33324 20334 33376 20340
rect 33230 20295 33286 20304
rect 33322 20088 33378 20097
rect 33140 20052 33192 20058
rect 33322 20023 33378 20032
rect 33140 19994 33192 20000
rect 33336 19786 33364 20023
rect 32494 19751 32550 19760
rect 32772 19780 32824 19786
rect 32508 19718 32536 19751
rect 32772 19722 32824 19728
rect 33324 19780 33376 19786
rect 33324 19722 33376 19728
rect 32496 19712 32548 19718
rect 32496 19654 32548 19660
rect 33140 19712 33192 19718
rect 33140 19654 33192 19660
rect 32956 19508 33008 19514
rect 32956 19450 33008 19456
rect 32968 19334 32996 19450
rect 33152 19334 33180 19654
rect 33428 19514 33456 20402
rect 34244 20392 34296 20398
rect 34244 20334 34296 20340
rect 34334 20360 34390 20369
rect 33570 20156 33878 20165
rect 33570 20154 33576 20156
rect 33632 20154 33656 20156
rect 33712 20154 33736 20156
rect 33792 20154 33816 20156
rect 33872 20154 33878 20156
rect 33632 20102 33634 20154
rect 33814 20102 33816 20154
rect 33570 20100 33576 20102
rect 33632 20100 33656 20102
rect 33712 20100 33736 20102
rect 33792 20100 33816 20102
rect 33872 20100 33878 20102
rect 33570 20091 33878 20100
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33520 19394 33548 19858
rect 34150 19816 34206 19825
rect 34150 19751 34152 19760
rect 34204 19751 34206 19760
rect 34152 19722 34204 19728
rect 32968 19306 33180 19334
rect 33232 19372 33284 19378
rect 33232 19314 33284 19320
rect 33428 19366 33548 19394
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 32324 18426 32352 18566
rect 32312 18420 32364 18426
rect 32312 18362 32364 18368
rect 32508 18358 32536 18634
rect 32496 18352 32548 18358
rect 32496 18294 32548 18300
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32680 18216 32732 18222
rect 32680 18158 32732 18164
rect 32220 17740 32272 17746
rect 32220 17682 32272 17688
rect 32324 17610 32352 18158
rect 32588 17740 32640 17746
rect 32588 17682 32640 17688
rect 32312 17604 32364 17610
rect 32312 17546 32364 17552
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31758 17167 31760 17176
rect 31812 17167 31814 17176
rect 31852 17196 31904 17202
rect 31760 17138 31812 17144
rect 31852 17138 31904 17144
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 31484 16652 31536 16658
rect 31484 16594 31536 16600
rect 30840 16448 30892 16454
rect 30840 16390 30892 16396
rect 30932 16448 30984 16454
rect 30932 16390 30984 16396
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30852 14498 30880 16390
rect 30944 16046 30972 16390
rect 31070 16348 31378 16357
rect 31070 16346 31076 16348
rect 31132 16346 31156 16348
rect 31212 16346 31236 16348
rect 31292 16346 31316 16348
rect 31372 16346 31378 16348
rect 31132 16294 31134 16346
rect 31314 16294 31316 16346
rect 31070 16292 31076 16294
rect 31132 16292 31156 16294
rect 31212 16292 31236 16294
rect 31292 16292 31316 16294
rect 31372 16292 31378 16294
rect 31070 16283 31378 16292
rect 32048 16250 32076 17274
rect 32140 16726 32168 17478
rect 32324 17338 32352 17546
rect 32404 17536 32456 17542
rect 32404 17478 32456 17484
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32324 16794 32352 17070
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32128 16720 32180 16726
rect 32128 16662 32180 16668
rect 32036 16244 32088 16250
rect 32088 16204 32168 16232
rect 32036 16186 32088 16192
rect 30932 16040 30984 16046
rect 30932 15982 30984 15988
rect 30944 15570 30972 15982
rect 30932 15564 30984 15570
rect 30932 15506 30984 15512
rect 31852 15360 31904 15366
rect 31852 15302 31904 15308
rect 31070 15260 31378 15269
rect 31070 15258 31076 15260
rect 31132 15258 31156 15260
rect 31212 15258 31236 15260
rect 31292 15258 31316 15260
rect 31372 15258 31378 15260
rect 31132 15206 31134 15258
rect 31314 15206 31316 15258
rect 31070 15204 31076 15206
rect 31132 15204 31156 15206
rect 31212 15204 31236 15206
rect 31292 15204 31316 15206
rect 31372 15204 31378 15206
rect 31070 15195 31378 15204
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30760 14470 30880 14498
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 29748 14062 29868 14090
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 29644 13524 29696 13530
rect 29644 13466 29696 13472
rect 29748 13326 29776 13942
rect 29840 13530 29868 14062
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 29828 13524 29880 13530
rect 29828 13466 29880 13472
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29840 12986 29868 13466
rect 29552 12980 29604 12986
rect 29552 12922 29604 12928
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 29932 12889 29960 13942
rect 30484 13546 30512 14010
rect 30576 13734 30604 14214
rect 30564 13728 30616 13734
rect 30564 13670 30616 13676
rect 30484 13518 30604 13546
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 30484 13326 30512 13398
rect 30576 13326 30604 13518
rect 30472 13320 30524 13326
rect 30102 13288 30158 13297
rect 30472 13262 30524 13268
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30102 13223 30158 13232
rect 30012 12912 30064 12918
rect 29918 12880 29974 12889
rect 29736 12844 29788 12850
rect 29736 12786 29788 12792
rect 29840 12838 29918 12866
rect 29644 12300 29696 12306
rect 29644 12242 29696 12248
rect 29182 12135 29238 12144
rect 29380 12158 29500 12186
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29196 10742 29224 11154
rect 29380 11082 29408 12158
rect 29552 11620 29604 11626
rect 29656 11608 29684 12242
rect 29748 11694 29776 12786
rect 29840 12646 29868 12838
rect 30012 12854 30064 12860
rect 29918 12815 29974 12824
rect 29828 12640 29880 12646
rect 29828 12582 29880 12588
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29828 12300 29880 12306
rect 29828 12242 29880 12248
rect 29840 11830 29868 12242
rect 29828 11824 29880 11830
rect 29828 11766 29880 11772
rect 29736 11688 29788 11694
rect 29736 11630 29788 11636
rect 29604 11580 29684 11608
rect 29552 11562 29604 11568
rect 29458 11384 29514 11393
rect 29656 11354 29684 11580
rect 29458 11319 29514 11328
rect 29644 11348 29696 11354
rect 29472 11286 29500 11319
rect 29644 11290 29696 11296
rect 29460 11280 29512 11286
rect 29460 11222 29512 11228
rect 29368 11076 29420 11082
rect 29288 11036 29368 11064
rect 29012 10662 29132 10690
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 29288 10674 29316 11036
rect 29368 11018 29420 11024
rect 29366 10976 29422 10985
rect 29366 10911 29422 10920
rect 29380 10810 29408 10911
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 29276 10668 29328 10674
rect 28570 10364 28878 10373
rect 28570 10362 28576 10364
rect 28632 10362 28656 10364
rect 28712 10362 28736 10364
rect 28792 10362 28816 10364
rect 28872 10362 28878 10364
rect 28632 10310 28634 10362
rect 28814 10310 28816 10362
rect 28570 10308 28576 10310
rect 28632 10308 28656 10310
rect 28712 10308 28736 10310
rect 28792 10308 28816 10310
rect 28872 10308 28878 10310
rect 28570 10299 28878 10308
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28368 10130 28580 10146
rect 28264 10124 28316 10130
rect 28368 10124 28592 10130
rect 28368 10118 28540 10124
rect 28264 10066 28316 10072
rect 28540 10066 28592 10072
rect 28170 9616 28226 9625
rect 28170 9551 28226 9560
rect 28184 9518 28212 9551
rect 28172 9512 28224 9518
rect 28172 9454 28224 9460
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 28000 8401 28028 8842
rect 27986 8392 28042 8401
rect 27986 8327 28042 8336
rect 28000 7886 28028 8327
rect 27988 7880 28040 7886
rect 28184 7834 28212 9454
rect 28276 8566 28304 10066
rect 28356 10056 28408 10062
rect 28408 10016 28488 10044
rect 28356 9998 28408 10004
rect 28460 8838 28488 10016
rect 29012 9994 29040 10662
rect 29276 10610 29328 10616
rect 29276 10532 29328 10538
rect 29276 10474 29328 10480
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 28570 9276 28878 9285
rect 28570 9274 28576 9276
rect 28632 9274 28656 9276
rect 28712 9274 28736 9276
rect 28792 9274 28816 9276
rect 28872 9274 28878 9276
rect 28632 9222 28634 9274
rect 28814 9222 28816 9274
rect 28570 9220 28576 9222
rect 28632 9220 28656 9222
rect 28712 9220 28736 9222
rect 28792 9220 28816 9222
rect 28872 9220 28878 9222
rect 28570 9211 28878 9220
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28264 8560 28316 8566
rect 28736 8537 28764 8774
rect 28264 8502 28316 8508
rect 28722 8528 28778 8537
rect 28722 8463 28778 8472
rect 28356 8424 28408 8430
rect 28540 8424 28592 8430
rect 28356 8366 28408 8372
rect 28538 8392 28540 8401
rect 28592 8392 28594 8401
rect 27988 7822 28040 7828
rect 28000 7410 28028 7822
rect 28092 7806 28212 7834
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 28000 7002 28028 7210
rect 27988 6996 28040 7002
rect 27988 6938 28040 6944
rect 27488 6752 27568 6780
rect 27724 6820 27844 6848
rect 27436 6734 27488 6740
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27448 6118 27476 6598
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27448 5710 27476 6054
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27252 5636 27304 5642
rect 27252 5578 27304 5584
rect 27158 4856 27214 4865
rect 27158 4791 27214 4800
rect 26792 4684 26844 4690
rect 26844 4644 26924 4672
rect 26792 4626 26844 4632
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 26608 4004 26660 4010
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25700 3194 25728 3334
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 25608 2514 25636 2926
rect 25700 2650 25728 3130
rect 25884 3058 25912 3946
rect 26344 3534 26372 3998
rect 26608 3946 26660 3952
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 25976 3194 26004 3334
rect 26070 3292 26378 3301
rect 26070 3290 26076 3292
rect 26132 3290 26156 3292
rect 26212 3290 26236 3292
rect 26292 3290 26316 3292
rect 26372 3290 26378 3292
rect 26132 3238 26134 3290
rect 26314 3238 26316 3290
rect 26070 3236 26076 3238
rect 26132 3236 26156 3238
rect 26212 3236 26236 3238
rect 26292 3236 26316 3238
rect 26372 3236 26378 3238
rect 26070 3227 26378 3236
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 26436 3058 26464 3878
rect 26608 3188 26660 3194
rect 26712 3176 26740 4082
rect 26804 3602 26832 4422
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26660 3148 26740 3176
rect 26608 3130 26660 3136
rect 26896 3126 26924 4644
rect 27264 4146 27292 5578
rect 27632 5370 27660 6326
rect 27724 6254 27752 6820
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27816 6458 27844 6666
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27908 5302 27936 6258
rect 28092 6066 28120 7806
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 28368 7698 28396 8366
rect 28538 8327 28594 8336
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 28460 8090 28488 8230
rect 28570 8188 28878 8197
rect 28570 8186 28576 8188
rect 28632 8186 28656 8188
rect 28712 8186 28736 8188
rect 28792 8186 28816 8188
rect 28872 8186 28878 8188
rect 28632 8134 28634 8186
rect 28814 8134 28816 8186
rect 28570 8132 28576 8134
rect 28632 8132 28656 8134
rect 28712 8132 28736 8134
rect 28792 8132 28816 8134
rect 28872 8132 28878 8134
rect 28570 8123 28878 8132
rect 28448 8084 28500 8090
rect 28448 8026 28500 8032
rect 28446 7984 28502 7993
rect 29104 7954 29132 10202
rect 29288 9994 29316 10474
rect 29380 10169 29408 10746
rect 29366 10160 29422 10169
rect 29366 10095 29422 10104
rect 29368 10056 29420 10062
rect 29472 10044 29500 11222
rect 29644 11212 29696 11218
rect 29644 11154 29696 11160
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 29564 10810 29592 11018
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29656 10742 29684 11154
rect 29748 11150 29776 11630
rect 29828 11552 29880 11558
rect 29826 11520 29828 11529
rect 29932 11540 29960 12582
rect 30024 12186 30052 12854
rect 30116 12782 30144 13223
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30104 12776 30156 12782
rect 30104 12718 30156 12724
rect 30024 12158 30144 12186
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 30024 11898 30052 12038
rect 30116 11898 30144 12158
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30208 11626 30236 12038
rect 30300 11778 30328 12786
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30392 11898 30420 12582
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30300 11750 30420 11778
rect 30196 11620 30248 11626
rect 30196 11562 30248 11568
rect 30012 11552 30064 11558
rect 29880 11520 29882 11529
rect 29932 11512 30012 11540
rect 30012 11494 30064 11500
rect 29826 11455 29882 11464
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29644 10736 29696 10742
rect 29644 10678 29696 10684
rect 29748 10674 29776 11086
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29828 10532 29880 10538
rect 29828 10474 29880 10480
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29420 10016 29500 10044
rect 29552 10056 29604 10062
rect 29368 9998 29420 10004
rect 29552 9998 29604 10004
rect 29276 9988 29328 9994
rect 29276 9930 29328 9936
rect 29380 9518 29408 9998
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 29184 9172 29236 9178
rect 29184 9114 29236 9120
rect 29196 8838 29224 9114
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29182 8392 29238 8401
rect 29182 8327 29238 8336
rect 29196 8022 29224 8327
rect 29380 8294 29408 9454
rect 29564 9178 29592 9998
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29550 9072 29606 9081
rect 29472 9030 29550 9058
rect 29368 8288 29420 8294
rect 29368 8230 29420 8236
rect 29184 8016 29236 8022
rect 29184 7958 29236 7964
rect 28446 7919 28502 7928
rect 28816 7948 28868 7954
rect 28460 7886 28488 7919
rect 28816 7890 28868 7896
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28184 7546 28212 7686
rect 28368 7670 28488 7698
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28368 6458 28396 7482
rect 28460 6780 28488 7670
rect 28632 7540 28684 7546
rect 28828 7528 28856 7890
rect 29104 7818 29132 7890
rect 29196 7868 29224 7958
rect 29276 7880 29328 7886
rect 29196 7840 29276 7868
rect 29276 7822 29328 7828
rect 29092 7812 29144 7818
rect 29092 7754 29144 7760
rect 28684 7500 28856 7528
rect 28632 7482 28684 7488
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28570 7100 28878 7109
rect 28570 7098 28576 7100
rect 28632 7098 28656 7100
rect 28712 7098 28736 7100
rect 28792 7098 28816 7100
rect 28872 7098 28878 7100
rect 28632 7046 28634 7098
rect 28814 7046 28816 7098
rect 28570 7044 28576 7046
rect 28632 7044 28656 7046
rect 28712 7044 28736 7046
rect 28792 7044 28816 7046
rect 28872 7044 28878 7046
rect 28570 7035 28878 7044
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 28736 6798 28764 6938
rect 28540 6792 28592 6798
rect 28460 6752 28540 6780
rect 28540 6734 28592 6740
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28356 6452 28408 6458
rect 28356 6394 28408 6400
rect 28736 6338 28764 6734
rect 28920 6458 28948 7142
rect 29472 6730 29500 9030
rect 29550 9007 29606 9016
rect 29656 7954 29684 10406
rect 29736 9716 29788 9722
rect 29736 9658 29788 9664
rect 29748 9382 29776 9658
rect 29840 9586 29868 10474
rect 29932 10130 29960 10678
rect 29920 10124 29972 10130
rect 29920 10066 29972 10072
rect 29932 9586 29960 10066
rect 30024 9674 30052 11494
rect 30208 10810 30236 11562
rect 30392 11370 30420 11750
rect 30300 11342 30420 11370
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30300 10606 30328 11342
rect 30484 10674 30512 12922
rect 30668 12442 30696 14418
rect 30760 12986 30788 14470
rect 31036 14346 31064 15030
rect 31758 14920 31814 14929
rect 31758 14855 31760 14864
rect 31812 14855 31814 14864
rect 31760 14826 31812 14832
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 14600 31248 14758
rect 31300 14612 31352 14618
rect 31220 14572 31300 14600
rect 31300 14554 31352 14560
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31116 14544 31168 14550
rect 31116 14486 31168 14492
rect 31484 14544 31536 14550
rect 31484 14486 31536 14492
rect 31128 14385 31156 14486
rect 31114 14376 31170 14385
rect 30840 14340 30892 14346
rect 30840 14282 30892 14288
rect 31024 14340 31076 14346
rect 31114 14311 31170 14320
rect 31024 14282 31076 14288
rect 30852 13938 30880 14282
rect 30932 14272 30984 14278
rect 30932 14214 30984 14220
rect 30840 13932 30892 13938
rect 30840 13874 30892 13880
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30748 12980 30800 12986
rect 30748 12922 30800 12928
rect 30852 12782 30880 13262
rect 30944 13190 30972 14214
rect 31070 14172 31378 14181
rect 31070 14170 31076 14172
rect 31132 14170 31156 14172
rect 31212 14170 31236 14172
rect 31292 14170 31316 14172
rect 31372 14170 31378 14172
rect 31132 14118 31134 14170
rect 31314 14118 31316 14170
rect 31070 14116 31076 14118
rect 31132 14116 31156 14118
rect 31212 14116 31236 14118
rect 31292 14116 31316 14118
rect 31372 14116 31378 14118
rect 31070 14107 31378 14116
rect 31392 14000 31444 14006
rect 31392 13942 31444 13948
rect 31404 13512 31432 13942
rect 31496 13938 31524 14486
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 31484 13524 31536 13530
rect 31404 13484 31484 13512
rect 31404 13258 31432 13484
rect 31484 13466 31536 13472
rect 31392 13252 31444 13258
rect 31392 13194 31444 13200
rect 30932 13184 30984 13190
rect 30932 13126 30984 13132
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31070 13084 31378 13093
rect 31070 13082 31076 13084
rect 31132 13082 31156 13084
rect 31212 13082 31236 13084
rect 31292 13082 31316 13084
rect 31372 13082 31378 13084
rect 31132 13030 31134 13082
rect 31314 13030 31316 13082
rect 31070 13028 31076 13030
rect 31132 13028 31156 13030
rect 31212 13028 31236 13030
rect 31292 13028 31316 13030
rect 31372 13028 31378 13030
rect 31070 13019 31378 13028
rect 31496 12918 31524 13126
rect 31484 12912 31536 12918
rect 31484 12854 31536 12860
rect 30840 12776 30892 12782
rect 30840 12718 30892 12724
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 30748 12640 30800 12646
rect 30748 12582 30800 12588
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30576 11642 30604 11834
rect 30668 11762 30696 12174
rect 30760 11898 30788 12582
rect 30840 12436 30892 12442
rect 30840 12378 30892 12384
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30852 11830 30880 12378
rect 31070 11996 31378 12005
rect 31070 11994 31076 11996
rect 31132 11994 31156 11996
rect 31212 11994 31236 11996
rect 31292 11994 31316 11996
rect 31372 11994 31378 11996
rect 31132 11942 31134 11994
rect 31314 11942 31316 11994
rect 31070 11940 31076 11942
rect 31132 11940 31156 11942
rect 31212 11940 31236 11942
rect 31292 11940 31316 11942
rect 31372 11940 31378 11942
rect 31070 11931 31378 11940
rect 30840 11824 30892 11830
rect 30840 11766 30892 11772
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30576 11614 30696 11642
rect 30668 11082 30696 11614
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30472 10668 30524 10674
rect 30472 10610 30524 10616
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30300 10130 30328 10542
rect 30760 10470 30788 11154
rect 30838 11112 30894 11121
rect 30894 11070 30972 11098
rect 30838 11047 30894 11056
rect 30944 10742 30972 11070
rect 31070 10908 31378 10917
rect 31070 10906 31076 10908
rect 31132 10906 31156 10908
rect 31212 10906 31236 10908
rect 31292 10906 31316 10908
rect 31372 10906 31378 10908
rect 31132 10854 31134 10906
rect 31314 10854 31316 10906
rect 31070 10852 31076 10854
rect 31132 10852 31156 10854
rect 31212 10852 31236 10854
rect 31292 10852 31316 10854
rect 31372 10852 31378 10854
rect 31070 10843 31378 10852
rect 30932 10736 30984 10742
rect 30932 10678 30984 10684
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30748 10464 30800 10470
rect 30748 10406 30800 10412
rect 30288 10124 30340 10130
rect 30208 10084 30288 10112
rect 30024 9646 30144 9674
rect 30208 9654 30236 10084
rect 30288 10066 30340 10072
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29920 9580 29972 9586
rect 29920 9522 29972 9528
rect 29840 9382 29868 9522
rect 29932 9450 29960 9522
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 29920 9444 29972 9450
rect 29920 9386 29972 9392
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29644 7948 29696 7954
rect 29644 7890 29696 7896
rect 29748 7886 29776 9318
rect 29840 9042 29868 9318
rect 29920 9172 29972 9178
rect 29920 9114 29972 9120
rect 29828 9036 29880 9042
rect 29828 8978 29880 8984
rect 29840 8498 29868 8978
rect 29932 8634 29960 9114
rect 30024 8906 30052 9454
rect 30116 8945 30144 9646
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30102 8936 30158 8945
rect 30012 8900 30064 8906
rect 30102 8871 30158 8880
rect 30012 8842 30064 8848
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 30024 8498 30052 8842
rect 30116 8838 30144 8871
rect 30104 8832 30156 8838
rect 30104 8774 30156 8780
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29564 7546 29592 7686
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29840 7206 29868 7822
rect 30024 7460 30052 8434
rect 30208 8412 30236 9590
rect 30300 9042 30328 9930
rect 30470 9752 30526 9761
rect 30470 9687 30526 9696
rect 30484 9654 30512 9687
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30472 9648 30524 9654
rect 30472 9590 30524 9596
rect 30392 9450 30420 9590
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 30484 9178 30512 9590
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30288 9036 30340 9042
rect 30288 8978 30340 8984
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30392 8498 30420 8774
rect 30472 8560 30524 8566
rect 30472 8502 30524 8508
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30288 8424 30340 8430
rect 30208 8384 30288 8412
rect 30288 8366 30340 8372
rect 30194 7984 30250 7993
rect 30300 7954 30328 8366
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 30194 7919 30250 7928
rect 30288 7948 30340 7954
rect 30104 7472 30156 7478
rect 30024 7432 30104 7460
rect 30104 7414 30156 7420
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 28736 6322 29316 6338
rect 28736 6316 29328 6322
rect 28736 6310 29276 6316
rect 28000 6038 28120 6066
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 28000 5846 28028 6038
rect 28080 5908 28132 5914
rect 28080 5850 28132 5856
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 28000 5642 28028 5782
rect 27988 5636 28040 5642
rect 27988 5578 28040 5584
rect 27896 5296 27948 5302
rect 27896 5238 27948 5244
rect 27436 4752 27488 4758
rect 27436 4694 27488 4700
rect 27448 4185 27476 4694
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27632 4282 27660 4490
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27724 4214 27752 4558
rect 27712 4208 27764 4214
rect 27434 4176 27490 4185
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 27344 4140 27396 4146
rect 27712 4150 27764 4156
rect 27434 4111 27490 4120
rect 27344 4082 27396 4088
rect 27264 3738 27292 4082
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27356 3602 27384 4082
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 27356 3466 27384 3538
rect 27344 3460 27396 3466
rect 27344 3402 27396 3408
rect 27436 3460 27488 3466
rect 27540 3448 27568 4014
rect 27908 3942 27936 5238
rect 27988 4684 28040 4690
rect 28092 4672 28120 5850
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28276 5030 28304 5510
rect 28368 5234 28396 6054
rect 28570 6012 28878 6021
rect 28570 6010 28576 6012
rect 28632 6010 28656 6012
rect 28712 6010 28736 6012
rect 28792 6010 28816 6012
rect 28872 6010 28878 6012
rect 28632 5958 28634 6010
rect 28814 5958 28816 6010
rect 28570 5956 28576 5958
rect 28632 5956 28656 5958
rect 28712 5956 28736 5958
rect 28792 5956 28816 5958
rect 28872 5956 28878 5958
rect 28570 5947 28878 5956
rect 28920 5914 28948 6310
rect 29276 6258 29328 6264
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 28920 5778 28948 5850
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 28448 5568 28500 5574
rect 28920 5556 28948 5714
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 29184 5636 29236 5642
rect 29184 5578 29236 5584
rect 28920 5528 29040 5556
rect 28448 5510 28500 5516
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28264 5024 28316 5030
rect 28264 4966 28316 4972
rect 28040 4644 28120 4672
rect 27988 4626 28040 4632
rect 28000 4078 28028 4626
rect 28276 4282 28304 4966
rect 28368 4622 28396 5170
rect 28460 4729 28488 5510
rect 28570 4924 28878 4933
rect 28570 4922 28576 4924
rect 28632 4922 28656 4924
rect 28712 4922 28736 4924
rect 28792 4922 28816 4924
rect 28872 4922 28878 4924
rect 28632 4870 28634 4922
rect 28814 4870 28816 4922
rect 28570 4868 28576 4870
rect 28632 4868 28656 4870
rect 28712 4868 28736 4870
rect 28792 4868 28816 4870
rect 28872 4868 28878 4870
rect 28570 4859 28878 4868
rect 29012 4842 29040 5528
rect 29104 5370 29132 5578
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29196 5030 29224 5578
rect 29184 5024 29236 5030
rect 29184 4966 29236 4972
rect 29012 4814 29224 4842
rect 28446 4720 28502 4729
rect 28446 4655 28448 4664
rect 28500 4655 28502 4664
rect 28724 4684 28776 4690
rect 28448 4626 28500 4632
rect 28724 4626 28776 4632
rect 28356 4616 28408 4622
rect 28736 4593 28764 4626
rect 28356 4558 28408 4564
rect 28722 4584 28778 4593
rect 28722 4519 28778 4528
rect 29092 4480 29144 4486
rect 29092 4422 29144 4428
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 28724 4208 28776 4214
rect 28776 4168 28948 4196
rect 28724 4150 28776 4156
rect 27988 4072 28040 4078
rect 27988 4014 28040 4020
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27896 3528 27948 3534
rect 28000 3516 28028 4014
rect 28092 3602 28120 4150
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 28184 3602 28212 4082
rect 28644 3942 28672 4082
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28460 3738 28488 3878
rect 28570 3836 28878 3845
rect 28570 3834 28576 3836
rect 28632 3834 28656 3836
rect 28712 3834 28736 3836
rect 28792 3834 28816 3836
rect 28872 3834 28878 3836
rect 28632 3782 28634 3834
rect 28814 3782 28816 3834
rect 28570 3780 28576 3782
rect 28632 3780 28656 3782
rect 28712 3780 28736 3782
rect 28792 3780 28816 3782
rect 28872 3780 28878 3782
rect 28570 3771 28878 3780
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 28540 3664 28592 3670
rect 28920 3618 28948 4168
rect 29104 3670 29132 4422
rect 29196 4282 29224 4814
rect 29288 4622 29316 5714
rect 29472 5148 29500 6190
rect 29564 5370 29592 6598
rect 30116 6390 30144 7414
rect 30104 6384 30156 6390
rect 30104 6326 30156 6332
rect 30208 5817 30236 7919
rect 30288 7890 30340 7896
rect 30392 7834 30420 7958
rect 30484 7857 30512 8502
rect 30300 7806 30420 7834
rect 30470 7848 30526 7857
rect 30300 6934 30328 7806
rect 30576 7834 30604 10406
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30668 10062 30696 10202
rect 30760 10062 30788 10406
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30748 9444 30800 9450
rect 30668 9404 30748 9432
rect 30668 8498 30696 9404
rect 30748 9386 30800 9392
rect 30746 8936 30802 8945
rect 30746 8871 30802 8880
rect 30760 8566 30788 8871
rect 30852 8566 30880 10610
rect 30944 9994 30972 10678
rect 31496 10674 31524 12718
rect 31680 12238 31708 14554
rect 31576 12232 31628 12238
rect 31576 12174 31628 12180
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31496 10470 31524 10610
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 30932 9988 30984 9994
rect 30932 9930 30984 9936
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 30840 8424 30892 8430
rect 30944 8412 30972 9930
rect 31070 9820 31378 9829
rect 31070 9818 31076 9820
rect 31132 9818 31156 9820
rect 31212 9818 31236 9820
rect 31292 9818 31316 9820
rect 31372 9818 31378 9820
rect 31132 9766 31134 9818
rect 31314 9766 31316 9818
rect 31070 9764 31076 9766
rect 31132 9764 31156 9766
rect 31212 9764 31236 9766
rect 31292 9764 31316 9766
rect 31372 9764 31378 9766
rect 31070 9755 31378 9764
rect 31208 9444 31260 9450
rect 31208 9386 31260 9392
rect 31220 9081 31248 9386
rect 31206 9072 31262 9081
rect 31496 9042 31524 10406
rect 31588 9654 31616 12174
rect 31680 11218 31708 12174
rect 31758 11384 31814 11393
rect 31758 11319 31760 11328
rect 31812 11319 31814 11328
rect 31760 11290 31812 11296
rect 31864 11286 31892 15302
rect 31942 15056 31998 15065
rect 31942 14991 31998 15000
rect 32036 15020 32088 15026
rect 31956 13802 31984 14991
rect 32036 14962 32088 14968
rect 31944 13796 31996 13802
rect 31944 13738 31996 13744
rect 31942 12744 31998 12753
rect 31942 12679 31998 12688
rect 31852 11280 31904 11286
rect 31852 11222 31904 11228
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31668 10736 31720 10742
rect 31720 10696 31892 10724
rect 31668 10678 31720 10684
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31206 9007 31262 9016
rect 31300 9036 31352 9042
rect 31484 9036 31536 9042
rect 31352 8996 31432 9024
rect 31300 8978 31352 8984
rect 31404 8786 31432 8996
rect 31484 8978 31536 8984
rect 31484 8832 31536 8838
rect 31404 8758 31448 8786
rect 31484 8774 31536 8780
rect 31070 8732 31378 8741
rect 31070 8730 31076 8732
rect 31132 8730 31156 8732
rect 31212 8730 31236 8732
rect 31292 8730 31316 8732
rect 31372 8730 31378 8732
rect 31132 8678 31134 8730
rect 31314 8678 31316 8730
rect 31070 8676 31076 8678
rect 31132 8676 31156 8678
rect 31212 8676 31236 8678
rect 31292 8676 31316 8678
rect 31372 8676 31378 8678
rect 31070 8667 31378 8676
rect 31420 8650 31448 8758
rect 31404 8622 31448 8650
rect 31404 8498 31432 8622
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 30892 8384 30972 8412
rect 30840 8366 30892 8372
rect 30852 8022 30880 8366
rect 31404 8294 31432 8434
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31312 8266 31432 8294
rect 31220 8090 31248 8230
rect 31208 8084 31260 8090
rect 31208 8026 31260 8032
rect 30840 8016 30892 8022
rect 30840 7958 30892 7964
rect 31312 7954 31340 8266
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 30748 7880 30800 7886
rect 30576 7806 30696 7834
rect 30748 7822 30800 7828
rect 30840 7880 30892 7886
rect 30892 7840 30972 7868
rect 30840 7822 30892 7828
rect 30470 7783 30526 7792
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30392 7546 30420 7686
rect 30380 7540 30432 7546
rect 30380 7482 30432 7488
rect 30288 6928 30340 6934
rect 30288 6870 30340 6876
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30300 6390 30328 6734
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 30194 5808 30250 5817
rect 30194 5743 30250 5752
rect 30300 5710 30328 6326
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 30392 5370 30420 5782
rect 29552 5364 29604 5370
rect 29552 5306 29604 5312
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 29552 5160 29604 5166
rect 29472 5120 29552 5148
rect 29552 5102 29604 5108
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30012 4752 30064 4758
rect 30012 4694 30064 4700
rect 29276 4616 29328 4622
rect 30024 4593 30052 4694
rect 30208 4690 30236 5102
rect 30300 4826 30328 5170
rect 30484 5148 30512 6734
rect 30576 5914 30604 7686
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30668 5658 30696 7806
rect 30760 6798 30788 7822
rect 30838 7304 30894 7313
rect 30838 7239 30840 7248
rect 30892 7239 30894 7248
rect 30840 7210 30892 7216
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30748 6656 30800 6662
rect 30748 6598 30800 6604
rect 30760 6458 30788 6598
rect 30852 6458 30880 6734
rect 30748 6452 30800 6458
rect 30748 6394 30800 6400
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30668 5630 30788 5658
rect 30760 5370 30788 5630
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30564 5160 30616 5166
rect 30484 5120 30564 5148
rect 30564 5102 30616 5108
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30196 4684 30248 4690
rect 30196 4626 30248 4632
rect 29276 4558 29328 4564
rect 30010 4584 30066 4593
rect 29288 4321 29316 4558
rect 30852 4554 30880 6394
rect 30944 5896 30972 7840
rect 31404 7698 31432 7890
rect 31496 7818 31524 8774
rect 31484 7812 31536 7818
rect 31484 7754 31536 7760
rect 31404 7670 31524 7698
rect 31070 7644 31378 7653
rect 31070 7642 31076 7644
rect 31132 7642 31156 7644
rect 31212 7642 31236 7644
rect 31292 7642 31316 7644
rect 31372 7642 31378 7644
rect 31132 7590 31134 7642
rect 31314 7590 31316 7642
rect 31070 7588 31076 7590
rect 31132 7588 31156 7590
rect 31212 7588 31236 7590
rect 31292 7588 31316 7590
rect 31372 7588 31378 7590
rect 31070 7579 31378 7588
rect 31114 7440 31170 7449
rect 31496 7410 31524 7670
rect 31484 7404 31536 7410
rect 31114 7375 31170 7384
rect 31128 7274 31156 7375
rect 31404 7364 31484 7392
rect 31116 7268 31168 7274
rect 31116 7210 31168 7216
rect 31022 6896 31078 6905
rect 31022 6831 31078 6840
rect 31036 6730 31064 6831
rect 31404 6730 31432 7364
rect 31484 7346 31536 7352
rect 31484 6928 31536 6934
rect 31484 6870 31536 6876
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31070 6556 31378 6565
rect 31070 6554 31076 6556
rect 31132 6554 31156 6556
rect 31212 6554 31236 6556
rect 31292 6554 31316 6556
rect 31372 6554 31378 6556
rect 31132 6502 31134 6554
rect 31314 6502 31316 6554
rect 31070 6500 31076 6502
rect 31132 6500 31156 6502
rect 31212 6500 31236 6502
rect 31292 6500 31316 6502
rect 31372 6500 31378 6502
rect 31070 6491 31378 6500
rect 31024 5908 31076 5914
rect 30944 5868 31024 5896
rect 31024 5850 31076 5856
rect 31070 5468 31378 5477
rect 31070 5466 31076 5468
rect 31132 5466 31156 5468
rect 31212 5466 31236 5468
rect 31292 5466 31316 5468
rect 31372 5466 31378 5468
rect 31132 5414 31134 5466
rect 31314 5414 31316 5466
rect 31070 5412 31076 5414
rect 31132 5412 31156 5414
rect 31212 5412 31236 5414
rect 31292 5412 31316 5414
rect 31372 5412 31378 5414
rect 31070 5403 31378 5412
rect 31392 5160 31444 5166
rect 31496 5148 31524 6870
rect 31588 6780 31616 9114
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31680 8566 31708 9046
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 31680 8265 31708 8298
rect 31772 8294 31800 10066
rect 31864 9382 31892 10696
rect 31956 9722 31984 12679
rect 32048 11778 32076 14962
rect 32140 14618 32168 16204
rect 32232 15638 32260 16730
rect 32312 16652 32364 16658
rect 32416 16640 32444 17478
rect 32600 17270 32628 17682
rect 32692 17270 32720 18158
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32680 17264 32732 17270
rect 32680 17206 32732 17212
rect 32784 17202 32812 19110
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32876 18193 32904 18702
rect 32862 18184 32918 18193
rect 32862 18119 32918 18128
rect 32968 17882 32996 19306
rect 33140 19236 33192 19242
rect 33140 19178 33192 19184
rect 33152 18970 33180 19178
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 33244 18358 33272 19314
rect 33428 18952 33456 19366
rect 34060 19304 34112 19310
rect 34060 19246 34112 19252
rect 33570 19068 33878 19077
rect 33570 19066 33576 19068
rect 33632 19066 33656 19068
rect 33712 19066 33736 19068
rect 33792 19066 33816 19068
rect 33872 19066 33878 19068
rect 33632 19014 33634 19066
rect 33814 19014 33816 19066
rect 33570 19012 33576 19014
rect 33632 19012 33656 19014
rect 33712 19012 33736 19014
rect 33792 19012 33816 19014
rect 33872 19012 33878 19014
rect 33570 19003 33878 19012
rect 33428 18924 33548 18952
rect 33520 18834 33548 18924
rect 33416 18828 33468 18834
rect 33416 18770 33468 18776
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33428 18426 33456 18770
rect 33416 18420 33468 18426
rect 33416 18362 33468 18368
rect 33232 18352 33284 18358
rect 33060 18312 33232 18340
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 32876 17338 32904 17818
rect 33060 17542 33088 18312
rect 33232 18294 33284 18300
rect 33232 18080 33284 18086
rect 33520 18068 33548 18770
rect 34072 18630 34100 19246
rect 34256 19242 34284 20334
rect 34334 20295 34390 20304
rect 34244 19236 34296 19242
rect 34244 19178 34296 19184
rect 34242 18728 34298 18737
rect 34152 18692 34204 18698
rect 34242 18663 34298 18672
rect 34152 18634 34204 18640
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 34164 18154 34192 18634
rect 34256 18630 34284 18663
rect 34244 18624 34296 18630
rect 34244 18566 34296 18572
rect 34244 18352 34296 18358
rect 34242 18320 34244 18329
rect 34296 18320 34298 18329
rect 34242 18255 34298 18264
rect 34152 18148 34204 18154
rect 34152 18090 34204 18096
rect 33232 18022 33284 18028
rect 33428 18040 33548 18068
rect 33048 17536 33100 17542
rect 33048 17478 33100 17484
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 32876 17241 32904 17274
rect 32862 17232 32918 17241
rect 32772 17196 32824 17202
rect 32862 17167 32918 17176
rect 32772 17138 32824 17144
rect 32496 17128 32548 17134
rect 32496 17070 32548 17076
rect 32508 16658 32536 17070
rect 32364 16612 32444 16640
rect 32496 16652 32548 16658
rect 32312 16594 32364 16600
rect 32496 16594 32548 16600
rect 32324 16182 32352 16594
rect 32312 16176 32364 16182
rect 32312 16118 32364 16124
rect 32220 15632 32272 15638
rect 32220 15574 32272 15580
rect 32324 15502 32352 16118
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32220 15088 32272 15094
rect 32220 15030 32272 15036
rect 32232 14929 32260 15030
rect 32218 14920 32274 14929
rect 32218 14855 32274 14864
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 32128 14340 32180 14346
rect 32128 14282 32180 14288
rect 32140 11898 32168 14282
rect 32220 13524 32272 13530
rect 32324 13512 32352 15438
rect 32508 14958 32536 16594
rect 32956 16448 33008 16454
rect 32956 16390 33008 16396
rect 33048 16448 33100 16454
rect 33048 16390 33100 16396
rect 32772 16040 32824 16046
rect 32692 16000 32772 16028
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32600 15094 32628 15302
rect 32692 15162 32720 16000
rect 32772 15982 32824 15988
rect 32968 15910 32996 16390
rect 33060 16250 33088 16390
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32956 15904 33008 15910
rect 33152 15858 33180 17274
rect 33244 16998 33272 18022
rect 33232 16992 33284 16998
rect 33232 16934 33284 16940
rect 33324 16720 33376 16726
rect 33324 16662 33376 16668
rect 32956 15846 33008 15852
rect 32864 15632 32916 15638
rect 32864 15574 32916 15580
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32680 15156 32732 15162
rect 32680 15098 32732 15104
rect 32588 15088 32640 15094
rect 32588 15030 32640 15036
rect 32496 14952 32548 14958
rect 32496 14894 32548 14900
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32588 14884 32640 14890
rect 32588 14826 32640 14832
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 32404 14272 32456 14278
rect 32404 14214 32456 14220
rect 32272 13484 32352 13512
rect 32220 13466 32272 13472
rect 32232 12918 32260 13466
rect 32220 12912 32272 12918
rect 32220 12854 32272 12860
rect 32312 12640 32364 12646
rect 32312 12582 32364 12588
rect 32324 12102 32352 12582
rect 32312 12096 32364 12102
rect 32312 12038 32364 12044
rect 32324 11898 32352 12038
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 32220 11824 32272 11830
rect 32048 11750 32168 11778
rect 32220 11766 32272 11772
rect 32036 11144 32088 11150
rect 32036 11086 32088 11092
rect 32048 10062 32076 11086
rect 32140 10470 32168 11750
rect 32232 10996 32260 11766
rect 32324 11150 32352 11834
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32416 11014 32444 14214
rect 32508 14006 32536 14554
rect 32600 14074 32628 14826
rect 32588 14068 32640 14074
rect 32588 14010 32640 14016
rect 32496 14000 32548 14006
rect 32496 13942 32548 13948
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32600 13530 32628 13874
rect 32588 13524 32640 13530
rect 32588 13466 32640 13472
rect 32600 12434 32628 13466
rect 32508 12406 32628 12434
rect 32692 12434 32720 14894
rect 32784 14822 32812 15302
rect 32876 15026 32904 15574
rect 32968 15026 32996 15846
rect 33060 15830 33180 15858
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 33060 14906 33088 15830
rect 33140 15700 33192 15706
rect 33140 15642 33192 15648
rect 33152 15026 33180 15642
rect 33336 15502 33364 16662
rect 33428 16658 33456 18040
rect 33570 17980 33878 17989
rect 33570 17978 33576 17980
rect 33632 17978 33656 17980
rect 33712 17978 33736 17980
rect 33792 17978 33816 17980
rect 33872 17978 33878 17980
rect 33632 17926 33634 17978
rect 33814 17926 33816 17978
rect 33570 17924 33576 17926
rect 33632 17924 33656 17926
rect 33712 17924 33736 17926
rect 33792 17924 33816 17926
rect 33872 17924 33878 17926
rect 33570 17915 33878 17924
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33796 17338 33824 17682
rect 33784 17332 33836 17338
rect 33784 17274 33836 17280
rect 34060 17196 34112 17202
rect 34060 17138 34112 17144
rect 33570 16892 33878 16901
rect 33570 16890 33576 16892
rect 33632 16890 33656 16892
rect 33712 16890 33736 16892
rect 33792 16890 33816 16892
rect 33872 16890 33878 16892
rect 33632 16838 33634 16890
rect 33814 16838 33816 16890
rect 33570 16836 33576 16838
rect 33632 16836 33656 16838
rect 33712 16836 33736 16838
rect 33792 16836 33816 16838
rect 33872 16836 33878 16838
rect 33570 16827 33878 16836
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 34072 16590 34100 17138
rect 34060 16584 34112 16590
rect 33690 16552 33746 16561
rect 34060 16526 34112 16532
rect 33690 16487 33692 16496
rect 33744 16487 33746 16496
rect 33692 16458 33744 16464
rect 34072 16182 34100 16526
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 33416 16040 33468 16046
rect 33416 15982 33468 15988
rect 33428 15706 33456 15982
rect 33570 15804 33878 15813
rect 33570 15802 33576 15804
rect 33632 15802 33656 15804
rect 33712 15802 33736 15804
rect 33792 15802 33816 15804
rect 33872 15802 33878 15804
rect 33632 15750 33634 15802
rect 33814 15750 33816 15802
rect 33570 15748 33576 15750
rect 33632 15748 33656 15750
rect 33712 15748 33736 15750
rect 33792 15748 33816 15750
rect 33872 15748 33878 15750
rect 33570 15739 33878 15748
rect 33416 15700 33468 15706
rect 33416 15642 33468 15648
rect 34072 15502 34100 16118
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33876 15496 33928 15502
rect 33876 15438 33928 15444
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 32968 14878 33088 14906
rect 32772 14816 32824 14822
rect 32772 14758 32824 14764
rect 32968 14550 32996 14878
rect 33048 14816 33100 14822
rect 33048 14758 33100 14764
rect 32956 14544 33008 14550
rect 32876 14504 32956 14532
rect 32876 14074 32904 14504
rect 32956 14486 33008 14492
rect 32956 14408 33008 14414
rect 32956 14350 33008 14356
rect 32864 14068 32916 14074
rect 32784 14028 32864 14056
rect 32784 12646 32812 14028
rect 32864 14010 32916 14016
rect 32968 13841 32996 14350
rect 32954 13832 33010 13841
rect 32954 13767 33010 13776
rect 32772 12640 32824 12646
rect 32772 12582 32824 12588
rect 32864 12640 32916 12646
rect 32864 12582 32916 12588
rect 32692 12406 32812 12434
rect 32508 12238 32536 12406
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 32588 11824 32640 11830
rect 32588 11766 32640 11772
rect 32312 11008 32364 11014
rect 32232 10968 32312 10996
rect 32312 10950 32364 10956
rect 32404 11008 32456 11014
rect 32456 10985 32536 10996
rect 32456 10976 32550 10985
rect 32456 10968 32494 10976
rect 32404 10950 32456 10956
rect 32324 10588 32352 10950
rect 32494 10911 32550 10920
rect 32600 10810 32628 11766
rect 32680 11620 32732 11626
rect 32680 11562 32732 11568
rect 32692 11354 32720 11562
rect 32680 11348 32732 11354
rect 32680 11290 32732 11296
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32496 10600 32548 10606
rect 32324 10560 32444 10588
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32310 10296 32366 10305
rect 32310 10231 32366 10240
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 32034 9616 32090 9625
rect 32034 9551 32036 9560
rect 32088 9551 32090 9560
rect 32036 9522 32088 9528
rect 31852 9376 31904 9382
rect 31852 9318 31904 9324
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32128 9376 32180 9382
rect 32128 9318 32180 9324
rect 32048 9110 32076 9318
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 31852 9036 31904 9042
rect 31852 8978 31904 8984
rect 31864 8566 31892 8978
rect 32140 8838 32168 9318
rect 32220 9104 32272 9110
rect 32220 9046 32272 9052
rect 32128 8832 32180 8838
rect 32128 8774 32180 8780
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31864 8378 31892 8502
rect 32232 8430 32260 9046
rect 32324 8430 32352 10231
rect 32416 10033 32444 10560
rect 32496 10542 32548 10548
rect 32402 10024 32458 10033
rect 32402 9959 32458 9968
rect 32508 9722 32536 10542
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32404 9036 32456 9042
rect 32404 8978 32456 8984
rect 32416 8498 32444 8978
rect 32600 8974 32628 9862
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32508 8634 32536 8774
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32494 8528 32550 8537
rect 32404 8492 32456 8498
rect 32494 8463 32550 8472
rect 32404 8434 32456 8440
rect 32220 8424 32272 8430
rect 32140 8401 32220 8412
rect 32126 8392 32220 8401
rect 31864 8350 32076 8378
rect 31760 8288 31812 8294
rect 31666 8256 31722 8265
rect 31760 8230 31812 8236
rect 31852 8288 31904 8294
rect 31852 8230 31904 8236
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31666 8191 31722 8200
rect 31864 8090 31892 8230
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31852 8084 31904 8090
rect 31852 8026 31904 8032
rect 31680 7546 31708 8026
rect 31760 8016 31812 8022
rect 31956 7970 31984 8230
rect 31812 7964 31984 7970
rect 31760 7958 31984 7964
rect 31772 7942 31984 7958
rect 32048 7954 32076 8350
rect 32182 8384 32220 8392
rect 32220 8366 32272 8372
rect 32312 8424 32364 8430
rect 32312 8366 32364 8372
rect 32126 8327 32182 8336
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31668 7540 31720 7546
rect 31772 7528 31800 7822
rect 32036 7812 32088 7818
rect 32140 7800 32168 8327
rect 32088 7772 32168 7800
rect 32036 7754 32088 7760
rect 31944 7540 31996 7546
rect 31772 7500 31944 7528
rect 31668 7482 31720 7488
rect 31944 7482 31996 7488
rect 31944 6792 31996 6798
rect 31588 6752 31944 6780
rect 31944 6734 31996 6740
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31588 6322 31616 6598
rect 31576 6316 31628 6322
rect 31576 6258 31628 6264
rect 31588 5370 31616 6258
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 31444 5120 31524 5148
rect 31392 5102 31444 5108
rect 31392 5024 31444 5030
rect 31392 4966 31444 4972
rect 31404 4690 31432 4966
rect 31588 4690 31616 5306
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31576 4684 31628 4690
rect 31576 4626 31628 4632
rect 30010 4519 30066 4528
rect 30840 4548 30892 4554
rect 30840 4490 30892 4496
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 30932 4480 30984 4486
rect 30932 4422 30984 4428
rect 31392 4480 31444 4486
rect 31772 4468 31800 5850
rect 32416 5778 32444 8434
rect 32508 6662 32536 8463
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32692 5778 32720 11154
rect 32784 10062 32812 12406
rect 32876 12306 32904 12582
rect 32864 12300 32916 12306
rect 32864 12242 32916 12248
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32876 11529 32904 11630
rect 32862 11520 32918 11529
rect 32862 11455 32918 11464
rect 32968 11218 32996 13767
rect 33060 13394 33088 14758
rect 33244 13977 33272 14962
rect 33336 14958 33364 15438
rect 33888 15162 33916 15438
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 34072 15094 34100 15438
rect 34060 15088 34112 15094
rect 34060 15030 34112 15036
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 34152 14952 34204 14958
rect 34152 14894 34204 14900
rect 33570 14716 33878 14725
rect 33570 14714 33576 14716
rect 33632 14714 33656 14716
rect 33712 14714 33736 14716
rect 33792 14714 33816 14716
rect 33872 14714 33878 14716
rect 33632 14662 33634 14714
rect 33814 14662 33816 14714
rect 33570 14660 33576 14662
rect 33632 14660 33656 14662
rect 33712 14660 33736 14662
rect 33792 14660 33816 14662
rect 33872 14660 33878 14662
rect 33570 14651 33878 14660
rect 33324 14544 33376 14550
rect 33324 14486 33376 14492
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 33336 14074 33364 14486
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 33416 14000 33468 14006
rect 33230 13968 33286 13977
rect 33416 13942 33468 13948
rect 33230 13903 33286 13912
rect 33232 13728 33284 13734
rect 33232 13670 33284 13676
rect 33244 13394 33272 13670
rect 33428 13462 33456 13942
rect 33520 13734 33548 14486
rect 33704 14470 34100 14498
rect 33704 14414 33732 14470
rect 33692 14408 33744 14414
rect 33692 14350 33744 14356
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33796 14074 33824 14350
rect 33968 14272 34020 14278
rect 33968 14214 34020 14220
rect 33784 14068 33836 14074
rect 33784 14010 33836 14016
rect 33508 13728 33560 13734
rect 33508 13670 33560 13676
rect 33570 13628 33878 13637
rect 33570 13626 33576 13628
rect 33632 13626 33656 13628
rect 33712 13626 33736 13628
rect 33792 13626 33816 13628
rect 33872 13626 33878 13628
rect 33632 13574 33634 13626
rect 33814 13574 33816 13626
rect 33570 13572 33576 13574
rect 33632 13572 33656 13574
rect 33712 13572 33736 13574
rect 33792 13572 33816 13574
rect 33872 13572 33878 13574
rect 33570 13563 33878 13572
rect 33416 13456 33468 13462
rect 33416 13398 33468 13404
rect 33876 13456 33928 13462
rect 33876 13398 33928 13404
rect 33048 13388 33100 13394
rect 33048 13330 33100 13336
rect 33232 13388 33284 13394
rect 33232 13330 33284 13336
rect 33324 13388 33376 13394
rect 33324 13330 33376 13336
rect 33048 13184 33100 13190
rect 33048 13126 33100 13132
rect 33060 12646 33088 13126
rect 33232 12912 33284 12918
rect 33230 12880 33232 12889
rect 33284 12880 33286 12889
rect 33336 12850 33364 13330
rect 33888 13258 33916 13398
rect 33980 13326 34008 14214
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 33508 13184 33560 13190
rect 33508 13126 33560 13132
rect 33520 12918 33548 13126
rect 33888 12918 33916 13194
rect 33508 12912 33560 12918
rect 33508 12854 33560 12860
rect 33876 12912 33928 12918
rect 33876 12854 33928 12860
rect 33230 12815 33286 12824
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33138 12744 33194 12753
rect 33138 12679 33194 12688
rect 33048 12640 33100 12646
rect 33048 12582 33100 12588
rect 33152 12102 33180 12679
rect 33336 12442 33364 12786
rect 33416 12640 33468 12646
rect 33416 12582 33468 12588
rect 33324 12436 33376 12442
rect 33244 12396 33324 12424
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 33244 11898 33272 12396
rect 33324 12378 33376 12384
rect 33322 12336 33378 12345
rect 33322 12271 33324 12280
rect 33376 12271 33378 12280
rect 33324 12242 33376 12248
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33336 11898 33364 12038
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 33324 11756 33376 11762
rect 33324 11698 33376 11704
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33140 11552 33192 11558
rect 33140 11494 33192 11500
rect 33232 11552 33284 11558
rect 33232 11494 33284 11500
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 32956 11212 33008 11218
rect 32956 11154 33008 11160
rect 32876 10305 32904 11154
rect 32954 10840 33010 10849
rect 33060 10826 33088 11494
rect 33010 10798 33088 10826
rect 32954 10775 33010 10784
rect 32862 10296 32918 10305
rect 33152 10266 33180 11494
rect 33244 10266 33272 11494
rect 33336 11354 33364 11698
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 33324 11008 33376 11014
rect 33324 10950 33376 10956
rect 33336 10713 33364 10950
rect 33322 10704 33378 10713
rect 33322 10639 33378 10648
rect 32862 10231 32918 10240
rect 33048 10260 33100 10266
rect 33048 10202 33100 10208
rect 33140 10260 33192 10266
rect 33140 10202 33192 10208
rect 33232 10260 33284 10266
rect 33232 10202 33284 10208
rect 32864 10192 32916 10198
rect 32864 10134 32916 10140
rect 32772 10056 32824 10062
rect 32772 9998 32824 10004
rect 32784 9518 32812 9998
rect 32876 9994 32904 10134
rect 32864 9988 32916 9994
rect 32864 9930 32916 9936
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32968 9722 32996 9862
rect 33060 9722 33088 10202
rect 32956 9716 33008 9722
rect 32956 9658 33008 9664
rect 33048 9716 33100 9722
rect 33048 9658 33100 9664
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32784 9178 32812 9454
rect 32864 9376 32916 9382
rect 32864 9318 32916 9324
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 32876 9058 32904 9318
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 32784 9030 32904 9058
rect 32784 6338 32812 9030
rect 33048 8900 33100 8906
rect 33048 8842 33100 8848
rect 33060 8634 33088 8842
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 32864 8424 32916 8430
rect 32864 8366 32916 8372
rect 32876 8090 32904 8366
rect 32864 8084 32916 8090
rect 32864 8026 32916 8032
rect 32956 7948 33008 7954
rect 32956 7890 33008 7896
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 32876 6866 32904 7482
rect 32968 7410 32996 7890
rect 32956 7404 33008 7410
rect 32956 7346 33008 7352
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 32968 6390 32996 7346
rect 32956 6384 33008 6390
rect 32862 6352 32918 6361
rect 32784 6310 32862 6338
rect 32956 6326 33008 6332
rect 32862 6287 32918 6296
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 32680 5636 32732 5642
rect 32680 5578 32732 5584
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 32600 5370 32628 5510
rect 32692 5370 32720 5578
rect 32876 5574 32904 6287
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32864 5568 32916 5574
rect 32864 5510 32916 5516
rect 32588 5364 32640 5370
rect 32588 5306 32640 5312
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 32218 5128 32274 5137
rect 32218 5063 32274 5072
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31444 4440 31800 4468
rect 31392 4422 31444 4428
rect 29274 4312 29330 4321
rect 29184 4276 29236 4282
rect 29274 4247 29330 4256
rect 29644 4276 29696 4282
rect 29184 4218 29236 4224
rect 29644 4218 29696 4224
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 29288 3754 29316 4082
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29196 3726 29316 3754
rect 28540 3606 28592 3612
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 27948 3488 28028 3516
rect 27896 3470 27948 3476
rect 27488 3420 27568 3448
rect 27436 3402 27488 3408
rect 27068 3392 27120 3398
rect 27120 3352 27292 3380
rect 27068 3334 27120 3340
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 26344 2514 26372 2790
rect 25596 2508 25648 2514
rect 26332 2508 26384 2514
rect 25648 2468 25728 2496
rect 25596 2450 25648 2456
rect 25412 2304 25464 2310
rect 25412 2246 25464 2252
rect 25424 1970 25452 2246
rect 25700 2038 25728 2468
rect 26332 2450 26384 2456
rect 26896 2446 26924 3062
rect 27264 2650 27292 3352
rect 27540 3194 27568 3420
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 27252 2644 27304 2650
rect 27252 2586 27304 2592
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 26070 2204 26378 2213
rect 26070 2202 26076 2204
rect 26132 2202 26156 2204
rect 26212 2202 26236 2204
rect 26292 2202 26316 2204
rect 26372 2202 26378 2204
rect 26132 2150 26134 2202
rect 26314 2150 26316 2202
rect 26070 2148 26076 2150
rect 26132 2148 26156 2150
rect 26212 2148 26236 2150
rect 26292 2148 26316 2150
rect 26372 2148 26378 2150
rect 26070 2139 26378 2148
rect 26896 2145 26924 2382
rect 26882 2136 26938 2145
rect 26882 2071 26938 2080
rect 26896 2038 26924 2071
rect 25688 2032 25740 2038
rect 25688 1974 25740 1980
rect 26884 2032 26936 2038
rect 26884 1974 26936 1980
rect 25412 1964 25464 1970
rect 25412 1906 25464 1912
rect 25596 1964 25648 1970
rect 25596 1906 25648 1912
rect 25608 1562 25636 1906
rect 26240 1760 26292 1766
rect 26240 1702 26292 1708
rect 25596 1556 25648 1562
rect 25596 1498 25648 1504
rect 25504 1488 25556 1494
rect 25424 1448 25504 1476
rect 24228 870 24440 898
rect 25228 944 25280 950
rect 25228 886 25280 892
rect 24228 160 24256 870
rect 23386 82 23442 160
rect 23308 54 23442 82
rect 23386 -300 23442 54
rect 24214 -300 24270 160
rect 25042 82 25098 160
rect 25424 82 25452 1448
rect 25504 1430 25556 1436
rect 26148 1420 26200 1426
rect 26148 1362 26200 1368
rect 26160 1204 26188 1362
rect 26252 1358 26280 1702
rect 27172 1358 27200 2518
rect 26240 1352 26292 1358
rect 26240 1294 26292 1300
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 25884 1176 26188 1204
rect 27068 1216 27120 1222
rect 25884 160 25912 1176
rect 27068 1158 27120 1164
rect 26070 1116 26378 1125
rect 26070 1114 26076 1116
rect 26132 1114 26156 1116
rect 26212 1114 26236 1116
rect 26292 1114 26316 1116
rect 26372 1114 26378 1116
rect 26132 1062 26134 1114
rect 26314 1062 26316 1114
rect 26070 1060 26076 1062
rect 26132 1060 26156 1062
rect 26212 1060 26236 1062
rect 26292 1060 26316 1062
rect 26372 1060 26378 1062
rect 26070 1051 26378 1060
rect 25042 54 25452 82
rect 25042 -300 25098 54
rect 25870 -300 25926 160
rect 26698 82 26754 160
rect 27080 82 27108 1158
rect 27264 882 27292 2586
rect 27448 2530 27476 2926
rect 27540 2650 27568 3130
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27448 2502 27568 2530
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27448 2310 27476 2382
rect 27540 2378 27568 2502
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 27632 2106 27660 3334
rect 27724 2553 27752 3402
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 27710 2544 27766 2553
rect 27710 2479 27712 2488
rect 27764 2479 27766 2488
rect 27712 2450 27764 2456
rect 27620 2100 27672 2106
rect 27620 2042 27672 2048
rect 27908 1902 27936 2858
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 28000 1970 28028 2790
rect 28092 2446 28120 3538
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28276 3097 28304 3334
rect 28262 3088 28318 3097
rect 28172 3052 28224 3058
rect 28262 3023 28318 3032
rect 28172 2994 28224 3000
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28078 2136 28134 2145
rect 28078 2071 28080 2080
rect 28132 2071 28134 2080
rect 28080 2042 28132 2048
rect 27988 1964 28040 1970
rect 27988 1906 28040 1912
rect 27896 1896 27948 1902
rect 27896 1838 27948 1844
rect 28184 1766 28212 2994
rect 28264 2984 28316 2990
rect 28368 2961 28396 3470
rect 28264 2926 28316 2932
rect 28354 2952 28410 2961
rect 28080 1760 28132 1766
rect 28080 1702 28132 1708
rect 28172 1760 28224 1766
rect 28172 1702 28224 1708
rect 27540 1562 27660 1578
rect 27540 1556 27672 1562
rect 27540 1550 27620 1556
rect 27252 876 27304 882
rect 27252 818 27304 824
rect 27540 160 27568 1550
rect 27620 1498 27672 1504
rect 28092 1358 28120 1702
rect 28276 1494 28304 2926
rect 28354 2887 28410 2896
rect 28368 2854 28396 2887
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28264 1488 28316 1494
rect 28264 1430 28316 1436
rect 28368 1426 28396 2790
rect 28460 2530 28488 3470
rect 28552 2990 28580 3606
rect 28828 3590 28948 3618
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 28828 3233 28856 3590
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28814 3224 28870 3233
rect 28814 3159 28870 3168
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28570 2748 28878 2757
rect 28570 2746 28576 2748
rect 28632 2746 28656 2748
rect 28712 2746 28736 2748
rect 28792 2746 28816 2748
rect 28872 2746 28878 2748
rect 28632 2694 28634 2746
rect 28814 2694 28816 2746
rect 28570 2692 28576 2694
rect 28632 2692 28656 2694
rect 28712 2692 28736 2694
rect 28792 2692 28816 2694
rect 28872 2692 28878 2694
rect 28570 2683 28878 2692
rect 28460 2502 28672 2530
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28356 1420 28408 1426
rect 28356 1362 28408 1368
rect 28460 1358 28488 2382
rect 28552 1902 28580 2382
rect 28644 1986 28672 2502
rect 28724 2508 28776 2514
rect 28920 2496 28948 3334
rect 29012 2650 29040 3470
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 28776 2468 28948 2496
rect 28724 2450 28776 2456
rect 29104 2310 29132 3470
rect 29196 2854 29224 3726
rect 29274 3496 29330 3505
rect 29380 3466 29408 4014
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29274 3431 29330 3440
rect 29368 3460 29420 3466
rect 29288 3398 29316 3431
rect 29368 3402 29420 3408
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 29092 2304 29144 2310
rect 29092 2246 29144 2252
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 28644 1958 28948 1986
rect 28540 1896 28592 1902
rect 28540 1838 28592 1844
rect 28570 1660 28878 1669
rect 28570 1658 28576 1660
rect 28632 1658 28656 1660
rect 28712 1658 28736 1660
rect 28792 1658 28816 1660
rect 28872 1658 28878 1660
rect 28632 1606 28634 1658
rect 28814 1606 28816 1658
rect 28570 1604 28576 1606
rect 28632 1604 28656 1606
rect 28712 1604 28736 1606
rect 28792 1604 28816 1606
rect 28872 1604 28878 1606
rect 28570 1595 28878 1604
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 28448 1352 28500 1358
rect 28920 1340 28948 1958
rect 29104 1562 29132 2246
rect 29092 1556 29144 1562
rect 29092 1498 29144 1504
rect 28920 1312 29132 1340
rect 28448 1294 28500 1300
rect 29104 1222 29132 1312
rect 29092 1216 29144 1222
rect 29092 1158 29144 1164
rect 28908 672 28960 678
rect 28908 614 28960 620
rect 28920 218 28948 614
rect 28828 190 28948 218
rect 26698 54 27108 82
rect 26698 -300 26754 54
rect 27526 -300 27582 160
rect 28354 82 28410 160
rect 28828 82 28856 190
rect 29196 160 29224 2246
rect 29288 1562 29316 2994
rect 29380 2582 29408 3402
rect 29472 3398 29500 3878
rect 29564 3602 29592 3878
rect 29656 3738 29684 4218
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29552 3460 29604 3466
rect 29604 3420 29684 3448
rect 29552 3402 29604 3408
rect 29460 3392 29512 3398
rect 29460 3334 29512 3340
rect 29472 3074 29500 3334
rect 29472 3058 29592 3074
rect 29472 3052 29604 3058
rect 29472 3046 29552 3052
rect 29552 2994 29604 3000
rect 29656 2938 29684 3420
rect 29748 3194 29776 4082
rect 30012 3936 30064 3942
rect 30012 3878 30064 3884
rect 30024 3738 30052 3878
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 29736 3188 29788 3194
rect 29736 3130 29788 3136
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 29564 2910 29684 2938
rect 30116 2922 30144 2994
rect 30104 2916 30156 2922
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29368 2576 29420 2582
rect 29368 2518 29420 2524
rect 29472 2446 29500 2790
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29564 1970 29592 2910
rect 30104 2858 30156 2864
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29656 1562 29684 2790
rect 30116 2582 30144 2858
rect 30208 2582 30236 4082
rect 30668 4078 30696 4422
rect 30944 4282 30972 4422
rect 31070 4380 31378 4389
rect 31070 4378 31076 4380
rect 31132 4378 31156 4380
rect 31212 4378 31236 4380
rect 31292 4378 31316 4380
rect 31372 4378 31378 4380
rect 31132 4326 31134 4378
rect 31314 4326 31316 4378
rect 31070 4324 31076 4326
rect 31132 4324 31156 4326
rect 31212 4324 31236 4326
rect 31292 4324 31316 4326
rect 31372 4324 31378 4326
rect 31070 4315 31378 4324
rect 30932 4276 30984 4282
rect 30932 4218 30984 4224
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30656 4072 30708 4078
rect 30656 4014 30708 4020
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 30286 3224 30342 3233
rect 30286 3159 30342 3168
rect 30300 3058 30328 3159
rect 30484 3058 30512 3878
rect 30576 3194 30604 3878
rect 30852 3670 30880 4082
rect 30840 3664 30892 3670
rect 30840 3606 30892 3612
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30288 3052 30340 3058
rect 30288 2994 30340 3000
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30392 2961 30420 2994
rect 30378 2952 30434 2961
rect 30378 2887 30434 2896
rect 30392 2774 30420 2887
rect 30300 2746 30420 2774
rect 30104 2576 30156 2582
rect 30104 2518 30156 2524
rect 30196 2576 30248 2582
rect 30196 2518 30248 2524
rect 30300 2446 30328 2746
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30012 2372 30064 2378
rect 30012 2314 30064 2320
rect 30024 2106 30052 2314
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 29736 1964 29788 1970
rect 29736 1906 29788 1912
rect 29276 1556 29328 1562
rect 29276 1498 29328 1504
rect 29644 1556 29696 1562
rect 29644 1498 29696 1504
rect 29276 1420 29328 1426
rect 29276 1362 29328 1368
rect 29288 1290 29316 1362
rect 29748 1290 29776 1906
rect 29920 1896 29972 1902
rect 29920 1838 29972 1844
rect 29932 1562 29960 1838
rect 30024 1766 30052 2042
rect 30576 1834 30604 2450
rect 30668 2446 30696 3538
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 30852 2854 30880 3470
rect 30840 2848 30892 2854
rect 30840 2790 30892 2796
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 30944 2106 30972 4082
rect 31036 3602 31064 4218
rect 31864 4010 31892 4694
rect 32232 4146 32260 5063
rect 32784 5012 32812 5510
rect 32864 5228 32916 5234
rect 32968 5216 32996 6326
rect 33152 5778 33180 9114
rect 33244 9042 33272 9522
rect 33232 9036 33284 9042
rect 33232 8978 33284 8984
rect 33232 8832 33284 8838
rect 33230 8800 33232 8809
rect 33284 8800 33286 8809
rect 33230 8735 33286 8744
rect 33336 8401 33364 9522
rect 33428 9178 33456 12582
rect 33570 12540 33878 12549
rect 33570 12538 33576 12540
rect 33632 12538 33656 12540
rect 33712 12538 33736 12540
rect 33792 12538 33816 12540
rect 33872 12538 33878 12540
rect 33632 12486 33634 12538
rect 33814 12486 33816 12538
rect 33570 12484 33576 12486
rect 33632 12484 33656 12486
rect 33712 12484 33736 12486
rect 33792 12484 33816 12486
rect 33872 12484 33878 12486
rect 33570 12475 33878 12484
rect 34072 12442 34100 14470
rect 34164 12646 34192 14894
rect 34348 14634 34376 20295
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34256 14606 34376 14634
rect 34152 12640 34204 12646
rect 34152 12582 34204 12588
rect 33876 12436 33928 12442
rect 33876 12378 33928 12384
rect 34060 12436 34112 12442
rect 34256 12434 34284 14606
rect 34336 14544 34388 14550
rect 34336 14486 34388 14492
rect 34348 13258 34376 14486
rect 34440 13870 34468 19654
rect 34532 19530 34560 20538
rect 34624 20398 34652 22510
rect 35164 22432 35216 22438
rect 35164 22374 35216 22380
rect 35716 22432 35768 22438
rect 35716 22374 35768 22380
rect 35808 22432 35860 22438
rect 35808 22374 35860 22380
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 36636 22432 36688 22438
rect 36636 22374 36688 22380
rect 34980 21480 35032 21486
rect 34980 21422 35032 21428
rect 34702 20904 34758 20913
rect 34702 20839 34758 20848
rect 34612 20392 34664 20398
rect 34612 20334 34664 20340
rect 34716 20330 34744 20839
rect 34992 20534 35020 21422
rect 35176 20602 35204 22374
rect 35440 22160 35492 22166
rect 35438 22128 35440 22137
rect 35492 22128 35494 22137
rect 35438 22063 35494 22072
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35452 21554 35480 21966
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 35452 20942 35480 21490
rect 35544 21146 35572 21490
rect 35636 21486 35664 21830
rect 35728 21486 35756 22374
rect 35624 21480 35676 21486
rect 35624 21422 35676 21428
rect 35716 21480 35768 21486
rect 35716 21422 35768 21428
rect 35532 21140 35584 21146
rect 35532 21082 35584 21088
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 35164 20596 35216 20602
rect 35164 20538 35216 20544
rect 34980 20528 35032 20534
rect 34980 20470 35032 20476
rect 35728 20398 35756 21422
rect 35072 20392 35124 20398
rect 35072 20334 35124 20340
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 34704 20324 34756 20330
rect 34704 20266 34756 20272
rect 35084 19922 35112 20334
rect 35624 20256 35676 20262
rect 35624 20198 35676 20204
rect 35072 19916 35124 19922
rect 35072 19858 35124 19864
rect 34888 19848 34940 19854
rect 34888 19790 34940 19796
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34532 19502 34652 19530
rect 34624 19446 34652 19502
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34532 18426 34560 19246
rect 34716 18834 34744 19654
rect 34900 19514 34928 19790
rect 35164 19712 35216 19718
rect 35164 19654 35216 19660
rect 34888 19508 34940 19514
rect 34888 19450 34940 19456
rect 35176 18873 35204 19654
rect 35532 19304 35584 19310
rect 35532 19246 35584 19252
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 35162 18864 35218 18873
rect 34704 18828 34756 18834
rect 35162 18799 35218 18808
rect 34704 18770 34756 18776
rect 34612 18624 34664 18630
rect 34612 18566 34664 18572
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34520 18420 34572 18426
rect 34520 18362 34572 18368
rect 34520 18216 34572 18222
rect 34624 18204 34652 18566
rect 34900 18358 34928 18566
rect 34888 18352 34940 18358
rect 34888 18294 34940 18300
rect 34572 18176 34652 18204
rect 34520 18158 34572 18164
rect 34532 17610 34560 18158
rect 34520 17604 34572 17610
rect 34520 17546 34572 17552
rect 34532 17338 34560 17546
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34808 17338 34836 17478
rect 34900 17338 34928 18294
rect 34980 18216 35032 18222
rect 34980 18158 35032 18164
rect 34992 17882 35020 18158
rect 34980 17876 35032 17882
rect 34980 17818 35032 17824
rect 35360 17678 35388 19110
rect 35544 17678 35572 19246
rect 35636 17746 35664 20198
rect 35728 19514 35756 20334
rect 35820 19854 35848 22374
rect 36096 22094 36124 22374
rect 36452 22228 36504 22234
rect 36452 22170 36504 22176
rect 36004 22066 36124 22094
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 35912 20602 35940 21490
rect 36004 20992 36032 22066
rect 36070 21788 36378 21797
rect 36070 21786 36076 21788
rect 36132 21786 36156 21788
rect 36212 21786 36236 21788
rect 36292 21786 36316 21788
rect 36372 21786 36378 21788
rect 36132 21734 36134 21786
rect 36314 21734 36316 21786
rect 36070 21732 36076 21734
rect 36132 21732 36156 21734
rect 36212 21732 36236 21734
rect 36292 21732 36316 21734
rect 36372 21732 36378 21734
rect 36070 21723 36378 21732
rect 36464 21690 36492 22170
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36452 21684 36504 21690
rect 36452 21626 36504 21632
rect 36556 21554 36584 21898
rect 36648 21593 36676 22374
rect 37108 22094 37136 22510
rect 36924 22066 37136 22094
rect 36634 21584 36690 21593
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36544 21548 36596 21554
rect 36634 21519 36690 21528
rect 36544 21490 36596 21496
rect 36176 21004 36228 21010
rect 36004 20964 36176 20992
rect 36176 20946 36228 20952
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 36004 20058 36032 20742
rect 36070 20700 36378 20709
rect 36070 20698 36076 20700
rect 36132 20698 36156 20700
rect 36212 20698 36236 20700
rect 36292 20698 36316 20700
rect 36372 20698 36378 20700
rect 36132 20646 36134 20698
rect 36314 20646 36316 20698
rect 36070 20644 36076 20646
rect 36132 20644 36156 20646
rect 36212 20644 36236 20646
rect 36292 20644 36316 20646
rect 36372 20644 36378 20646
rect 36070 20635 36378 20644
rect 36464 20602 36492 21490
rect 36924 21350 36952 22066
rect 36912 21344 36964 21350
rect 36912 21286 36964 21292
rect 36452 20596 36504 20602
rect 36452 20538 36504 20544
rect 36820 20528 36872 20534
rect 36820 20470 36872 20476
rect 35992 20052 36044 20058
rect 35992 19994 36044 20000
rect 35808 19848 35860 19854
rect 35808 19790 35860 19796
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35716 19508 35768 19514
rect 35716 19450 35768 19456
rect 35820 19310 35848 19654
rect 36070 19612 36378 19621
rect 36070 19610 36076 19612
rect 36132 19610 36156 19612
rect 36212 19610 36236 19612
rect 36292 19610 36316 19612
rect 36372 19610 36378 19612
rect 36132 19558 36134 19610
rect 36314 19558 36316 19610
rect 36070 19556 36076 19558
rect 36132 19556 36156 19558
rect 36212 19556 36236 19558
rect 36292 19556 36316 19558
rect 36372 19556 36378 19558
rect 36070 19547 36378 19556
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35808 19304 35860 19310
rect 35808 19246 35860 19252
rect 35820 18426 35848 19246
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35808 18420 35860 18426
rect 35808 18362 35860 18368
rect 35624 17740 35676 17746
rect 35912 17728 35940 19110
rect 36004 17882 36032 19314
rect 36084 19236 36136 19242
rect 36084 19178 36136 19184
rect 36096 18630 36124 19178
rect 36176 19168 36228 19174
rect 36176 19110 36228 19116
rect 36268 19168 36320 19174
rect 36268 19110 36320 19116
rect 36188 18970 36216 19110
rect 36176 18964 36228 18970
rect 36176 18906 36228 18912
rect 36280 18766 36308 19110
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36832 18630 36860 20470
rect 36924 20466 36952 21286
rect 37292 21146 37320 22578
rect 37556 22568 37608 22574
rect 37556 22510 37608 22516
rect 37372 22500 37424 22506
rect 37372 22442 37424 22448
rect 37384 22166 37412 22442
rect 37372 22160 37424 22166
rect 37372 22102 37424 22108
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 37280 21140 37332 21146
rect 37280 21082 37332 21088
rect 37384 21010 37412 21966
rect 37464 21480 37516 21486
rect 37464 21422 37516 21428
rect 37372 21004 37424 21010
rect 37372 20946 37424 20952
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 36912 20460 36964 20466
rect 36912 20402 36964 20408
rect 37188 20392 37240 20398
rect 37188 20334 37240 20340
rect 37200 19922 37228 20334
rect 37188 19916 37240 19922
rect 37188 19858 37240 19864
rect 36912 19168 36964 19174
rect 36912 19110 36964 19116
rect 37096 19168 37148 19174
rect 37096 19110 37148 19116
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 36452 18624 36504 18630
rect 36452 18566 36504 18572
rect 36820 18624 36872 18630
rect 36820 18566 36872 18572
rect 36070 18524 36378 18533
rect 36070 18522 36076 18524
rect 36132 18522 36156 18524
rect 36212 18522 36236 18524
rect 36292 18522 36316 18524
rect 36372 18522 36378 18524
rect 36132 18470 36134 18522
rect 36314 18470 36316 18522
rect 36070 18468 36076 18470
rect 36132 18468 36156 18470
rect 36212 18468 36236 18470
rect 36292 18468 36316 18470
rect 36372 18468 36378 18470
rect 36070 18459 36378 18468
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35912 17700 36032 17728
rect 35624 17682 35676 17688
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 36004 17610 36032 17700
rect 36176 17672 36228 17678
rect 36464 17660 36492 18566
rect 36924 18222 36952 19110
rect 37004 18828 37056 18834
rect 37004 18770 37056 18776
rect 37016 18698 37044 18770
rect 37004 18692 37056 18698
rect 37004 18634 37056 18640
rect 37108 18358 37136 19110
rect 37096 18352 37148 18358
rect 37096 18294 37148 18300
rect 36912 18216 36964 18222
rect 36912 18158 36964 18164
rect 36924 17882 36952 18158
rect 36912 17876 36964 17882
rect 36912 17818 36964 17824
rect 36228 17632 36492 17660
rect 36176 17614 36228 17620
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34796 17332 34848 17338
rect 34796 17274 34848 17280
rect 34888 17332 34940 17338
rect 34888 17274 34940 17280
rect 34900 17218 34928 17274
rect 34808 17190 34928 17218
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 34428 13728 34480 13734
rect 34428 13670 34480 13676
rect 34336 13252 34388 13258
rect 34336 13194 34388 13200
rect 34060 12378 34112 12384
rect 34164 12406 34284 12434
rect 33888 12238 33916 12378
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33508 12096 33560 12102
rect 33508 12038 33560 12044
rect 33520 11801 33548 12038
rect 33506 11792 33562 11801
rect 33506 11727 33562 11736
rect 33968 11688 34020 11694
rect 33968 11630 34020 11636
rect 33570 11452 33878 11461
rect 33570 11450 33576 11452
rect 33632 11450 33656 11452
rect 33712 11450 33736 11452
rect 33792 11450 33816 11452
rect 33872 11450 33878 11452
rect 33632 11398 33634 11450
rect 33814 11398 33816 11450
rect 33570 11396 33576 11398
rect 33632 11396 33656 11398
rect 33712 11396 33736 11398
rect 33792 11396 33816 11398
rect 33872 11396 33878 11398
rect 33570 11387 33878 11396
rect 33980 11218 34008 11630
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 34072 11218 34100 11494
rect 33968 11212 34020 11218
rect 33968 11154 34020 11160
rect 34060 11212 34112 11218
rect 34060 11154 34112 11160
rect 33876 11008 33928 11014
rect 33876 10950 33928 10956
rect 33966 10976 34022 10985
rect 33888 10742 33916 10950
rect 33966 10911 34022 10920
rect 33876 10736 33928 10742
rect 33876 10678 33928 10684
rect 33570 10364 33878 10373
rect 33570 10362 33576 10364
rect 33632 10362 33656 10364
rect 33712 10362 33736 10364
rect 33792 10362 33816 10364
rect 33872 10362 33878 10364
rect 33632 10310 33634 10362
rect 33814 10310 33816 10362
rect 33570 10308 33576 10310
rect 33632 10308 33656 10310
rect 33712 10308 33736 10310
rect 33792 10308 33816 10310
rect 33872 10308 33878 10310
rect 33570 10299 33878 10308
rect 33506 10160 33562 10169
rect 33506 10095 33562 10104
rect 33600 10124 33652 10130
rect 33520 9994 33548 10095
rect 33600 10066 33652 10072
rect 33612 10033 33640 10066
rect 33598 10024 33654 10033
rect 33508 9988 33560 9994
rect 33598 9959 33654 9968
rect 33508 9930 33560 9936
rect 33612 9489 33640 9959
rect 33980 9654 34008 10911
rect 34164 10826 34192 12406
rect 34440 12374 34468 13670
rect 34532 13530 34560 16934
rect 34808 16522 34836 17190
rect 35912 16794 35940 17546
rect 36924 17542 36952 17818
rect 37200 17746 37228 19858
rect 37292 19854 37320 20538
rect 37372 20392 37424 20398
rect 37476 20380 37504 21422
rect 37424 20352 37504 20380
rect 37372 20334 37424 20340
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37280 19712 37332 19718
rect 37280 19654 37332 19660
rect 37292 19514 37320 19654
rect 37280 19508 37332 19514
rect 37280 19450 37332 19456
rect 37280 19304 37332 19310
rect 37384 19292 37412 20334
rect 37332 19264 37412 19292
rect 37280 19246 37332 19252
rect 37568 18834 37596 22510
rect 37660 20058 37688 22578
rect 37924 22500 37976 22506
rect 37924 22442 37976 22448
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37832 21888 37884 21894
rect 37832 21830 37884 21836
rect 37752 20942 37780 21830
rect 37844 21457 37872 21830
rect 37936 21690 37964 22442
rect 38016 22432 38068 22438
rect 38016 22374 38068 22380
rect 38292 22432 38344 22438
rect 38292 22374 38344 22380
rect 38028 22094 38056 22374
rect 38200 22160 38252 22166
rect 38200 22102 38252 22108
rect 38028 22066 38148 22094
rect 37924 21684 37976 21690
rect 37924 21626 37976 21632
rect 37924 21548 37976 21554
rect 37924 21490 37976 21496
rect 37830 21448 37886 21457
rect 37830 21383 37886 21392
rect 37830 21040 37886 21049
rect 37830 20975 37886 20984
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37752 20602 37780 20878
rect 37844 20874 37872 20975
rect 37936 20942 37964 21490
rect 38016 21412 38068 21418
rect 38016 21354 38068 21360
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37832 20868 37884 20874
rect 37832 20810 37884 20816
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37936 20534 37964 20878
rect 37924 20528 37976 20534
rect 38028 20505 38056 21354
rect 38120 20942 38148 22066
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38108 20528 38160 20534
rect 37924 20470 37976 20476
rect 38014 20496 38070 20505
rect 38108 20470 38160 20476
rect 38014 20431 38070 20440
rect 37648 20052 37700 20058
rect 37648 19994 37700 20000
rect 37924 19712 37976 19718
rect 37924 19654 37976 19660
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37556 18828 37608 18834
rect 37556 18770 37608 18776
rect 37292 18358 37320 18770
rect 37936 18766 37964 19654
rect 38120 19446 38148 20470
rect 38108 19440 38160 19446
rect 38108 19382 38160 19388
rect 38120 19310 38148 19382
rect 38016 19304 38068 19310
rect 38016 19246 38068 19252
rect 38108 19304 38160 19310
rect 38108 19246 38160 19252
rect 37924 18760 37976 18766
rect 37924 18702 37976 18708
rect 38028 18680 38056 19246
rect 38108 18692 38160 18698
rect 38028 18652 38108 18680
rect 38108 18634 38160 18640
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 37292 18086 37320 18294
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 38212 17882 38240 22102
rect 38304 22012 38332 22374
rect 38396 22094 38424 22578
rect 38844 22432 38896 22438
rect 39212 22432 39264 22438
rect 38896 22392 38976 22420
rect 38844 22374 38896 22380
rect 38570 22332 38878 22341
rect 38570 22330 38576 22332
rect 38632 22330 38656 22332
rect 38712 22330 38736 22332
rect 38792 22330 38816 22332
rect 38872 22330 38878 22332
rect 38632 22278 38634 22330
rect 38814 22278 38816 22330
rect 38570 22276 38576 22278
rect 38632 22276 38656 22278
rect 38712 22276 38736 22278
rect 38792 22276 38816 22278
rect 38872 22276 38878 22278
rect 38570 22267 38878 22276
rect 38396 22066 38516 22094
rect 38304 21984 38424 22012
rect 38396 21894 38424 21984
rect 38292 21888 38344 21894
rect 38292 21830 38344 21836
rect 38384 21888 38436 21894
rect 38384 21830 38436 21836
rect 38304 21146 38332 21830
rect 38396 21486 38424 21830
rect 38384 21480 38436 21486
rect 38384 21422 38436 21428
rect 38488 21350 38516 22066
rect 38948 22030 38976 22392
rect 39212 22374 39264 22380
rect 39304 22432 39356 22438
rect 39304 22374 39356 22380
rect 39224 22030 39252 22374
rect 38936 22024 38988 22030
rect 38936 21966 38988 21972
rect 39212 22024 39264 22030
rect 39212 21966 39264 21972
rect 38936 21888 38988 21894
rect 38936 21830 38988 21836
rect 38476 21344 38528 21350
rect 38476 21286 38528 21292
rect 38292 21140 38344 21146
rect 38292 21082 38344 21088
rect 38384 21004 38436 21010
rect 38384 20946 38436 20952
rect 38396 20398 38424 20946
rect 38384 20392 38436 20398
rect 38384 20334 38436 20340
rect 38488 19990 38516 21286
rect 38570 21244 38878 21253
rect 38570 21242 38576 21244
rect 38632 21242 38656 21244
rect 38712 21242 38736 21244
rect 38792 21242 38816 21244
rect 38872 21242 38878 21244
rect 38632 21190 38634 21242
rect 38814 21190 38816 21242
rect 38570 21188 38576 21190
rect 38632 21188 38656 21190
rect 38712 21188 38736 21190
rect 38792 21188 38816 21190
rect 38872 21188 38878 21190
rect 38570 21179 38878 21188
rect 38660 20868 38712 20874
rect 38948 20856 38976 21830
rect 39212 20936 39264 20942
rect 39212 20878 39264 20884
rect 38712 20828 38976 20856
rect 38660 20810 38712 20816
rect 38568 20800 38620 20806
rect 38568 20742 38620 20748
rect 39028 20800 39080 20806
rect 39028 20742 39080 20748
rect 38580 20602 38608 20742
rect 38568 20596 38620 20602
rect 38568 20538 38620 20544
rect 38936 20256 38988 20262
rect 38936 20198 38988 20204
rect 38570 20156 38878 20165
rect 38570 20154 38576 20156
rect 38632 20154 38656 20156
rect 38712 20154 38736 20156
rect 38792 20154 38816 20156
rect 38872 20154 38878 20156
rect 38632 20102 38634 20154
rect 38814 20102 38816 20154
rect 38570 20100 38576 20102
rect 38632 20100 38656 20102
rect 38712 20100 38736 20102
rect 38792 20100 38816 20102
rect 38872 20100 38878 20102
rect 38570 20091 38878 20100
rect 38948 20040 38976 20198
rect 38764 20012 38976 20040
rect 38476 19984 38528 19990
rect 38476 19926 38528 19932
rect 38764 19854 38792 20012
rect 38476 19848 38528 19854
rect 38752 19848 38804 19854
rect 38476 19790 38528 19796
rect 38750 19816 38752 19825
rect 38804 19816 38806 19825
rect 38292 19712 38344 19718
rect 38292 19654 38344 19660
rect 38304 19514 38332 19654
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38488 18970 38516 19790
rect 38750 19751 38806 19760
rect 38934 19272 38990 19281
rect 39040 19258 39068 20742
rect 39224 20398 39252 20878
rect 39212 20392 39264 20398
rect 39212 20334 39264 20340
rect 39224 19786 39252 20334
rect 39212 19780 39264 19786
rect 39212 19722 39264 19728
rect 39224 19310 39252 19722
rect 38990 19230 39068 19258
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 38934 19207 38990 19216
rect 38570 19068 38878 19077
rect 38570 19066 38576 19068
rect 38632 19066 38656 19068
rect 38712 19066 38736 19068
rect 38792 19066 38816 19068
rect 38872 19066 38878 19068
rect 38632 19014 38634 19066
rect 38814 19014 38816 19066
rect 38570 19012 38576 19014
rect 38632 19012 38656 19014
rect 38712 19012 38736 19014
rect 38792 19012 38816 19014
rect 38872 19012 38878 19014
rect 38570 19003 38878 19012
rect 38476 18964 38528 18970
rect 38476 18906 38528 18912
rect 38384 18828 38436 18834
rect 38384 18770 38436 18776
rect 38200 17876 38252 17882
rect 38200 17818 38252 17824
rect 37738 17776 37794 17785
rect 37188 17740 37240 17746
rect 37738 17711 37794 17720
rect 37188 17682 37240 17688
rect 37752 17678 37780 17711
rect 37740 17672 37792 17678
rect 37740 17614 37792 17620
rect 37280 17604 37332 17610
rect 37280 17546 37332 17552
rect 36452 17536 36504 17542
rect 36452 17478 36504 17484
rect 36912 17536 36964 17542
rect 36912 17478 36964 17484
rect 36070 17436 36378 17445
rect 36070 17434 36076 17436
rect 36132 17434 36156 17436
rect 36212 17434 36236 17436
rect 36292 17434 36316 17436
rect 36372 17434 36378 17436
rect 36132 17382 36134 17434
rect 36314 17382 36316 17434
rect 36070 17380 36076 17382
rect 36132 17380 36156 17382
rect 36212 17380 36236 17382
rect 36292 17380 36316 17382
rect 36372 17380 36378 17382
rect 36070 17371 36378 17380
rect 36176 16992 36228 16998
rect 36176 16934 36228 16940
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 35992 16652 36044 16658
rect 35992 16594 36044 16600
rect 35808 16584 35860 16590
rect 35808 16526 35860 16532
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34808 16114 34836 16458
rect 35716 16448 35768 16454
rect 35716 16390 35768 16396
rect 35728 16114 35756 16390
rect 34796 16108 34848 16114
rect 34796 16050 34848 16056
rect 35716 16108 35768 16114
rect 35716 16050 35768 16056
rect 34704 15360 34756 15366
rect 34808 15348 34836 16050
rect 35256 16040 35308 16046
rect 35256 15982 35308 15988
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35072 15904 35124 15910
rect 35072 15846 35124 15852
rect 34756 15320 34836 15348
rect 34704 15302 34756 15308
rect 34612 13728 34664 13734
rect 34612 13670 34664 13676
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34428 12368 34480 12374
rect 34428 12310 34480 12316
rect 34242 12200 34298 12209
rect 34242 12135 34298 12144
rect 34256 12102 34284 12135
rect 34244 12096 34296 12102
rect 34244 12038 34296 12044
rect 34440 11694 34468 12310
rect 34532 11830 34560 13466
rect 34624 12442 34652 13670
rect 34716 13190 34744 15302
rect 35084 15162 35112 15846
rect 35072 15156 35124 15162
rect 35072 15098 35124 15104
rect 35084 15042 35112 15098
rect 35084 15014 35204 15042
rect 35072 14952 35124 14958
rect 35072 14894 35124 14900
rect 34888 14408 34940 14414
rect 34888 14350 34940 14356
rect 34796 13864 34848 13870
rect 34796 13806 34848 13812
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34612 12436 34664 12442
rect 34612 12378 34664 12384
rect 34808 12374 34836 13806
rect 34900 13297 34928 14350
rect 34980 14340 35032 14346
rect 34980 14282 35032 14288
rect 34886 13288 34942 13297
rect 34886 13223 34942 13232
rect 34992 12986 35020 14282
rect 35084 14278 35112 14894
rect 35176 14414 35204 15014
rect 35164 14408 35216 14414
rect 35164 14350 35216 14356
rect 35072 14272 35124 14278
rect 35072 14214 35124 14220
rect 35072 13932 35124 13938
rect 35072 13874 35124 13880
rect 35084 13190 35112 13874
rect 35072 13184 35124 13190
rect 35072 13126 35124 13132
rect 34980 12980 35032 12986
rect 34980 12922 35032 12928
rect 34796 12368 34848 12374
rect 34796 12310 34848 12316
rect 34992 12306 35020 12922
rect 35084 12434 35112 13126
rect 35268 12900 35296 15982
rect 35348 15564 35400 15570
rect 35348 15506 35400 15512
rect 35360 15162 35388 15506
rect 35348 15156 35400 15162
rect 35348 15098 35400 15104
rect 35452 15094 35480 15982
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 35624 14612 35676 14618
rect 35624 14554 35676 14560
rect 35532 14544 35584 14550
rect 35532 14486 35584 14492
rect 35348 12912 35400 12918
rect 35268 12872 35348 12900
rect 35348 12854 35400 12860
rect 35084 12406 35204 12434
rect 34980 12300 35032 12306
rect 34980 12242 35032 12248
rect 35176 12238 35204 12406
rect 35164 12232 35216 12238
rect 35164 12174 35216 12180
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34520 11824 34572 11830
rect 34520 11766 34572 11772
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34428 11212 34480 11218
rect 34428 11154 34480 11160
rect 34336 11076 34388 11082
rect 34336 11018 34388 11024
rect 34164 10798 34284 10826
rect 34060 10260 34112 10266
rect 34060 10202 34112 10208
rect 33968 9648 34020 9654
rect 33968 9590 34020 9596
rect 33598 9480 33654 9489
rect 33598 9415 33654 9424
rect 33968 9376 34020 9382
rect 33968 9318 34020 9324
rect 33570 9276 33878 9285
rect 33570 9274 33576 9276
rect 33632 9274 33656 9276
rect 33712 9274 33736 9276
rect 33792 9274 33816 9276
rect 33872 9274 33878 9276
rect 33632 9222 33634 9274
rect 33814 9222 33816 9274
rect 33570 9220 33576 9222
rect 33632 9220 33656 9222
rect 33712 9220 33736 9222
rect 33792 9220 33816 9222
rect 33872 9220 33878 9222
rect 33570 9211 33878 9220
rect 33980 9178 34008 9318
rect 34072 9217 34100 10202
rect 34058 9208 34114 9217
rect 33416 9172 33468 9178
rect 33416 9114 33468 9120
rect 33968 9172 34020 9178
rect 34058 9143 34114 9152
rect 33968 9114 34020 9120
rect 34072 9058 34100 9143
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 33980 9030 34100 9058
rect 33506 8936 33562 8945
rect 33612 8906 33640 8978
rect 33506 8871 33562 8880
rect 33600 8900 33652 8906
rect 33322 8392 33378 8401
rect 33322 8327 33378 8336
rect 33520 8276 33548 8871
rect 33600 8842 33652 8848
rect 33428 8248 33548 8276
rect 33428 7206 33456 8248
rect 33570 8188 33878 8197
rect 33570 8186 33576 8188
rect 33632 8186 33656 8188
rect 33712 8186 33736 8188
rect 33792 8186 33816 8188
rect 33872 8186 33878 8188
rect 33632 8134 33634 8186
rect 33814 8134 33816 8186
rect 33570 8132 33576 8134
rect 33632 8132 33656 8134
rect 33712 8132 33736 8134
rect 33792 8132 33816 8134
rect 33872 8132 33878 8134
rect 33570 8123 33878 8132
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 33428 6730 33456 7142
rect 33570 7100 33878 7109
rect 33570 7098 33576 7100
rect 33632 7098 33656 7100
rect 33712 7098 33736 7100
rect 33792 7098 33816 7100
rect 33872 7098 33878 7100
rect 33632 7046 33634 7098
rect 33814 7046 33816 7098
rect 33570 7044 33576 7046
rect 33632 7044 33656 7046
rect 33712 7044 33736 7046
rect 33792 7044 33816 7046
rect 33872 7044 33878 7046
rect 33570 7035 33878 7044
rect 33980 7002 34008 9030
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 34060 8560 34112 8566
rect 34060 8502 34112 8508
rect 34072 8022 34100 8502
rect 34060 8016 34112 8022
rect 34060 7958 34112 7964
rect 34060 7880 34112 7886
rect 34060 7822 34112 7828
rect 34072 7546 34100 7822
rect 34164 7546 34192 8570
rect 34256 8276 34284 10798
rect 34348 10266 34376 11018
rect 34440 10810 34468 11154
rect 34532 10810 34560 11630
rect 34428 10804 34480 10810
rect 34428 10746 34480 10752
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34336 10260 34388 10266
rect 34336 10202 34388 10208
rect 34440 9994 34468 10746
rect 34428 9988 34480 9994
rect 34428 9930 34480 9936
rect 34520 9716 34572 9722
rect 34520 9658 34572 9664
rect 34336 9512 34388 9518
rect 34388 9472 34468 9500
rect 34336 9454 34388 9460
rect 34336 9104 34388 9110
rect 34336 9046 34388 9052
rect 34348 8906 34376 9046
rect 34440 9042 34468 9472
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 34336 8900 34388 8906
rect 34336 8842 34388 8848
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34334 8664 34390 8673
rect 34334 8599 34336 8608
rect 34388 8599 34390 8608
rect 34336 8570 34388 8576
rect 34440 8401 34468 8774
rect 34532 8634 34560 9658
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34426 8392 34482 8401
rect 34426 8327 34482 8336
rect 34256 8248 34468 8276
rect 34244 8084 34296 8090
rect 34244 8026 34296 8032
rect 34256 7546 34284 8026
rect 34440 7886 34468 8248
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 34060 7540 34112 7546
rect 34060 7482 34112 7488
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34244 7540 34296 7546
rect 34244 7482 34296 7488
rect 34152 7336 34204 7342
rect 34152 7278 34204 7284
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 33968 6996 34020 7002
rect 33968 6938 34020 6944
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33416 6724 33468 6730
rect 33416 6666 33468 6672
rect 33232 6248 33284 6254
rect 33232 6190 33284 6196
rect 33244 5914 33272 6190
rect 33704 6118 33732 6802
rect 34072 6730 34100 7142
rect 34060 6724 34112 6730
rect 34060 6666 34112 6672
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33968 6656 34020 6662
rect 33968 6598 34020 6604
rect 33796 6361 33824 6598
rect 33782 6352 33838 6361
rect 33782 6287 33838 6296
rect 33416 6112 33468 6118
rect 33416 6054 33468 6060
rect 33692 6112 33744 6118
rect 33692 6054 33744 6060
rect 33232 5908 33284 5914
rect 33232 5850 33284 5856
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33324 5704 33376 5710
rect 33230 5672 33286 5681
rect 33428 5692 33456 6054
rect 33570 6012 33878 6021
rect 33570 6010 33576 6012
rect 33632 6010 33656 6012
rect 33712 6010 33736 6012
rect 33792 6010 33816 6012
rect 33872 6010 33878 6012
rect 33632 5958 33634 6010
rect 33814 5958 33816 6010
rect 33570 5956 33576 5958
rect 33632 5956 33656 5958
rect 33712 5956 33736 5958
rect 33792 5956 33816 5958
rect 33872 5956 33878 5958
rect 33570 5947 33878 5956
rect 33980 5778 34008 6598
rect 34164 6390 34192 7278
rect 34440 7002 34468 7686
rect 34532 7546 34560 8434
rect 34520 7540 34572 7546
rect 34520 7482 34572 7488
rect 34624 7426 34652 11834
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 34716 11665 34744 11698
rect 34702 11656 34758 11665
rect 34702 11591 34758 11600
rect 35072 11552 35124 11558
rect 35072 11494 35124 11500
rect 34980 11076 35032 11082
rect 34980 11018 35032 11024
rect 34888 11008 34940 11014
rect 34888 10950 34940 10956
rect 34794 10840 34850 10849
rect 34794 10775 34850 10784
rect 34702 9616 34758 9625
rect 34808 9602 34836 10775
rect 34900 10606 34928 10950
rect 34992 10742 35020 11018
rect 34980 10736 35032 10742
rect 34980 10678 35032 10684
rect 34888 10600 34940 10606
rect 34888 10542 34940 10548
rect 34900 9994 34928 10542
rect 34888 9988 34940 9994
rect 34888 9930 34940 9936
rect 34900 9722 34928 9930
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 35084 9654 35112 11494
rect 35360 9926 35388 12854
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35452 11218 35480 11834
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35544 10588 35572 14486
rect 35636 13394 35664 14554
rect 35728 14482 35756 16050
rect 35820 16046 35848 16526
rect 35900 16448 35952 16454
rect 35900 16390 35952 16396
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 35808 15360 35860 15366
rect 35808 15302 35860 15308
rect 35820 15162 35848 15302
rect 35808 15156 35860 15162
rect 35808 15098 35860 15104
rect 35820 14482 35848 15098
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 35808 14340 35860 14346
rect 35912 14328 35940 16390
rect 36004 16250 36032 16594
rect 36188 16454 36216 16934
rect 36464 16522 36492 17478
rect 36820 17196 36872 17202
rect 36820 17138 36872 17144
rect 36636 16992 36688 16998
rect 36636 16934 36688 16940
rect 36452 16516 36504 16522
rect 36504 16476 36584 16504
rect 36452 16458 36504 16464
rect 36176 16448 36228 16454
rect 36176 16390 36228 16396
rect 36070 16348 36378 16357
rect 36070 16346 36076 16348
rect 36132 16346 36156 16348
rect 36212 16346 36236 16348
rect 36292 16346 36316 16348
rect 36372 16346 36378 16348
rect 36132 16294 36134 16346
rect 36314 16294 36316 16346
rect 36070 16292 36076 16294
rect 36132 16292 36156 16294
rect 36212 16292 36236 16294
rect 36292 16292 36316 16294
rect 36372 16292 36378 16294
rect 36070 16283 36378 16292
rect 35992 16244 36044 16250
rect 35992 16186 36044 16192
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36070 15260 36378 15269
rect 36070 15258 36076 15260
rect 36132 15258 36156 15260
rect 36212 15258 36236 15260
rect 36292 15258 36316 15260
rect 36372 15258 36378 15260
rect 36132 15206 36134 15258
rect 36314 15206 36316 15258
rect 36070 15204 36076 15206
rect 36132 15204 36156 15206
rect 36212 15204 36236 15206
rect 36292 15204 36316 15206
rect 36372 15204 36378 15206
rect 36070 15195 36378 15204
rect 36464 15162 36492 15370
rect 36452 15156 36504 15162
rect 36452 15098 36504 15104
rect 36556 14482 36584 16476
rect 36648 16182 36676 16934
rect 36832 16794 36860 17138
rect 37292 17066 37320 17546
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 37476 17202 37504 17478
rect 38200 17264 38252 17270
rect 38200 17206 38252 17212
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37280 17060 37332 17066
rect 37280 17002 37332 17008
rect 37188 16992 37240 16998
rect 37188 16934 37240 16940
rect 37200 16794 37228 16934
rect 36820 16788 36872 16794
rect 36820 16730 36872 16736
rect 37188 16788 37240 16794
rect 37188 16730 37240 16736
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 36912 16448 36964 16454
rect 36912 16390 36964 16396
rect 36636 16176 36688 16182
rect 36636 16118 36688 16124
rect 36636 16040 36688 16046
rect 36636 15982 36688 15988
rect 36648 15570 36676 15982
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 36648 14618 36676 15506
rect 36818 14920 36874 14929
rect 36818 14855 36820 14864
rect 36872 14855 36874 14864
rect 36820 14826 36872 14832
rect 36924 14822 36952 16390
rect 37200 15570 37228 16594
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37200 14958 37228 15506
rect 37292 15473 37320 17002
rect 37476 16998 37504 17138
rect 37464 16992 37516 16998
rect 37464 16934 37516 16940
rect 37476 16046 37504 16934
rect 38212 16794 38240 17206
rect 38200 16788 38252 16794
rect 38200 16730 38252 16736
rect 38292 16584 38344 16590
rect 38292 16526 38344 16532
rect 37924 16448 37976 16454
rect 37924 16390 37976 16396
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 37936 16114 37964 16390
rect 37924 16108 37976 16114
rect 37924 16050 37976 16056
rect 37464 16040 37516 16046
rect 37464 15982 37516 15988
rect 37936 15706 37964 16050
rect 38028 15978 38056 16390
rect 38016 15972 38068 15978
rect 38016 15914 38068 15920
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 38212 15502 38240 15846
rect 38304 15706 38332 16526
rect 38292 15700 38344 15706
rect 38292 15642 38344 15648
rect 38200 15496 38252 15502
rect 37278 15464 37334 15473
rect 37830 15464 37886 15473
rect 37278 15399 37334 15408
rect 37556 15428 37608 15434
rect 37886 15422 37964 15450
rect 38200 15438 38252 15444
rect 37830 15399 37886 15408
rect 37556 15370 37608 15376
rect 37568 15094 37596 15370
rect 37648 15360 37700 15366
rect 37648 15302 37700 15308
rect 37660 15162 37688 15302
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37556 15088 37608 15094
rect 37556 15030 37608 15036
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37188 14952 37240 14958
rect 37188 14894 37240 14900
rect 36912 14816 36964 14822
rect 36912 14758 36964 14764
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36544 14476 36596 14482
rect 36544 14418 36596 14424
rect 35992 14408 36044 14414
rect 35992 14350 36044 14356
rect 35860 14300 35940 14328
rect 35808 14282 35860 14288
rect 35716 14272 35768 14278
rect 35716 14214 35768 14220
rect 35728 13870 35756 14214
rect 36004 14074 36032 14350
rect 36452 14272 36504 14278
rect 36452 14214 36504 14220
rect 36070 14172 36378 14181
rect 36070 14170 36076 14172
rect 36132 14170 36156 14172
rect 36212 14170 36236 14172
rect 36292 14170 36316 14172
rect 36372 14170 36378 14172
rect 36132 14118 36134 14170
rect 36314 14118 36316 14170
rect 36070 14116 36076 14118
rect 36132 14116 36156 14118
rect 36212 14116 36236 14118
rect 36292 14116 36316 14118
rect 36372 14116 36378 14118
rect 36070 14107 36378 14116
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 35716 13864 35768 13870
rect 35716 13806 35768 13812
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36372 13530 36400 13806
rect 35900 13524 35952 13530
rect 35820 13484 35900 13512
rect 35624 13388 35676 13394
rect 35624 13330 35676 13336
rect 35636 12850 35664 13330
rect 35820 12986 35848 13484
rect 35900 13466 35952 13472
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 36360 13524 36412 13530
rect 36360 13466 36412 13472
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 35624 12844 35676 12850
rect 35676 12804 35756 12832
rect 35624 12786 35676 12792
rect 35728 12442 35756 12804
rect 36004 12782 36032 13466
rect 36070 13084 36378 13093
rect 36070 13082 36076 13084
rect 36132 13082 36156 13084
rect 36212 13082 36236 13084
rect 36292 13082 36316 13084
rect 36372 13082 36378 13084
rect 36132 13030 36134 13082
rect 36314 13030 36316 13082
rect 36070 13028 36076 13030
rect 36132 13028 36156 13030
rect 36212 13028 36236 13030
rect 36292 13028 36316 13030
rect 36372 13028 36378 13030
rect 36070 13019 36378 13028
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 35716 12436 35768 12442
rect 35716 12378 35768 12384
rect 35728 11898 35756 12378
rect 36464 12306 36492 14214
rect 36556 14074 36584 14418
rect 36924 14074 36952 14758
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 37108 14260 37136 14554
rect 37292 14260 37320 14758
rect 37108 14232 37320 14260
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 36912 14068 36964 14074
rect 36912 14010 36964 14016
rect 37292 13938 37320 14232
rect 37372 14272 37424 14278
rect 37556 14272 37608 14278
rect 37372 14214 37424 14220
rect 37476 14232 37556 14260
rect 36544 13932 36596 13938
rect 36544 13874 36596 13880
rect 37188 13932 37240 13938
rect 37188 13874 37240 13880
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 36556 13394 36584 13874
rect 37096 13864 37148 13870
rect 37096 13806 37148 13812
rect 36544 13388 36596 13394
rect 36544 13330 36596 13336
rect 36556 12986 36584 13330
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 36912 12776 36964 12782
rect 36912 12718 36964 12724
rect 36452 12300 36504 12306
rect 36452 12242 36504 12248
rect 36634 12200 36690 12209
rect 36634 12135 36690 12144
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36070 11996 36378 12005
rect 36070 11994 36076 11996
rect 36132 11994 36156 11996
rect 36212 11994 36236 11996
rect 36292 11994 36316 11996
rect 36372 11994 36378 11996
rect 36132 11942 36134 11994
rect 36314 11942 36316 11994
rect 36070 11940 36076 11942
rect 36132 11940 36156 11942
rect 36212 11940 36236 11942
rect 36292 11940 36316 11942
rect 36372 11940 36378 11942
rect 36070 11931 36378 11940
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35900 11756 35952 11762
rect 35900 11698 35952 11704
rect 35716 11620 35768 11626
rect 35716 11562 35768 11568
rect 35728 11218 35756 11562
rect 35716 11212 35768 11218
rect 35716 11154 35768 11160
rect 35728 10606 35756 11154
rect 35624 10600 35676 10606
rect 35544 10560 35624 10588
rect 35624 10542 35676 10548
rect 35716 10600 35768 10606
rect 35716 10542 35768 10548
rect 35808 10600 35860 10606
rect 35808 10542 35860 10548
rect 35636 9994 35664 10542
rect 35728 10130 35756 10542
rect 35820 10266 35848 10542
rect 35912 10266 35940 11698
rect 36084 11008 36136 11014
rect 36004 10968 36084 10996
rect 36004 10810 36032 10968
rect 36084 10950 36136 10956
rect 36070 10908 36378 10917
rect 36070 10906 36076 10908
rect 36132 10906 36156 10908
rect 36212 10906 36236 10908
rect 36292 10906 36316 10908
rect 36372 10906 36378 10908
rect 36132 10854 36134 10906
rect 36314 10854 36316 10906
rect 36070 10852 36076 10854
rect 36132 10852 36156 10854
rect 36212 10852 36236 10854
rect 36292 10852 36316 10854
rect 36372 10852 36378 10854
rect 36070 10843 36378 10852
rect 36464 10810 36492 12038
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 35992 10804 36044 10810
rect 35992 10746 36044 10752
rect 36452 10804 36504 10810
rect 36452 10746 36504 10752
rect 36004 10690 36032 10746
rect 36004 10662 36124 10690
rect 36556 10674 36584 11630
rect 36648 11150 36676 12135
rect 36924 11558 36952 12718
rect 37108 12442 37136 13806
rect 37200 12442 37228 13874
rect 37280 13728 37332 13734
rect 37280 13670 37332 13676
rect 37292 12986 37320 13670
rect 37384 13530 37412 14214
rect 37372 13524 37424 13530
rect 37372 13466 37424 13472
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37096 12436 37148 12442
rect 37096 12378 37148 12384
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37476 12345 37504 14232
rect 37556 14214 37608 14220
rect 37556 13728 37608 13734
rect 37556 13670 37608 13676
rect 37568 13326 37596 13670
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37648 13252 37700 13258
rect 37648 13194 37700 13200
rect 37660 13138 37688 13194
rect 37568 13110 37688 13138
rect 37462 12336 37518 12345
rect 37462 12271 37518 12280
rect 37568 12238 37596 13110
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 37660 12238 37688 12922
rect 37752 12306 37780 14962
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37844 14006 37872 14214
rect 37832 14000 37884 14006
rect 37832 13942 37884 13948
rect 37936 12594 37964 15422
rect 38108 15360 38160 15366
rect 38108 15302 38160 15308
rect 38120 14414 38148 15302
rect 38200 15088 38252 15094
rect 38200 15030 38252 15036
rect 38016 14408 38068 14414
rect 38016 14350 38068 14356
rect 38108 14408 38160 14414
rect 38108 14350 38160 14356
rect 38028 13530 38056 14350
rect 38212 14006 38240 15030
rect 38200 14000 38252 14006
rect 38200 13942 38252 13948
rect 38016 13524 38068 13530
rect 38016 13466 38068 13472
rect 38212 13394 38240 13942
rect 38200 13388 38252 13394
rect 38200 13330 38252 13336
rect 38212 12918 38240 13330
rect 38200 12912 38252 12918
rect 38200 12854 38252 12860
rect 37936 12566 38148 12594
rect 37740 12300 37792 12306
rect 37740 12242 37792 12248
rect 37556 12232 37608 12238
rect 37476 12192 37556 12220
rect 37096 12164 37148 12170
rect 37096 12106 37148 12112
rect 37108 11898 37136 12106
rect 37280 12096 37332 12102
rect 37280 12038 37332 12044
rect 37292 11898 37320 12038
rect 37476 11914 37504 12192
rect 37556 12174 37608 12180
rect 37648 12232 37700 12238
rect 37648 12174 37700 12180
rect 37476 11898 37688 11914
rect 37096 11892 37148 11898
rect 37096 11834 37148 11840
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 37476 11892 37700 11898
rect 37476 11886 37648 11892
rect 37476 11830 37504 11886
rect 37648 11834 37700 11840
rect 37464 11824 37516 11830
rect 37464 11766 37516 11772
rect 37004 11688 37056 11694
rect 37004 11630 37056 11636
rect 36912 11552 36964 11558
rect 36912 11494 36964 11500
rect 37016 11354 37044 11630
rect 37924 11620 37976 11626
rect 37924 11562 37976 11568
rect 37096 11552 37148 11558
rect 37096 11494 37148 11500
rect 37004 11348 37056 11354
rect 37004 11290 37056 11296
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 37108 11082 37136 11494
rect 37936 11354 37964 11562
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 37096 11076 37148 11082
rect 37096 11018 37148 11024
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37476 10810 37504 10950
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 36818 10704 36874 10713
rect 36096 10470 36124 10662
rect 36268 10668 36320 10674
rect 36268 10610 36320 10616
rect 36544 10668 36596 10674
rect 36818 10639 36874 10648
rect 36544 10610 36596 10616
rect 35992 10464 36044 10470
rect 35992 10406 36044 10412
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 36004 10266 36032 10406
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35900 10260 35952 10266
rect 35900 10202 35952 10208
rect 35992 10260 36044 10266
rect 35992 10202 36044 10208
rect 35716 10124 35768 10130
rect 35716 10066 35768 10072
rect 36280 10062 36308 10610
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 36268 10056 36320 10062
rect 36320 10004 36492 10010
rect 36268 9998 36492 10004
rect 35624 9988 35676 9994
rect 36280 9982 36492 9998
rect 35624 9930 35676 9936
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 36070 9820 36378 9829
rect 36070 9818 36076 9820
rect 36132 9818 36156 9820
rect 36212 9818 36236 9820
rect 36292 9818 36316 9820
rect 36372 9818 36378 9820
rect 36132 9766 36134 9818
rect 36314 9766 36316 9818
rect 36070 9764 36076 9766
rect 36132 9764 36156 9766
rect 36212 9764 36236 9766
rect 36292 9764 36316 9766
rect 36372 9764 36378 9766
rect 36070 9755 36378 9764
rect 36464 9722 36492 9982
rect 36452 9716 36504 9722
rect 36452 9658 36504 9664
rect 35072 9648 35124 9654
rect 34808 9574 34928 9602
rect 35072 9590 35124 9596
rect 34702 9551 34758 9560
rect 34532 7398 34652 7426
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34152 6384 34204 6390
rect 34152 6326 34204 6332
rect 34244 6248 34296 6254
rect 34244 6190 34296 6196
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 33968 5772 34020 5778
rect 33968 5714 34020 5720
rect 34060 5772 34112 5778
rect 34060 5714 34112 5720
rect 33376 5664 33456 5692
rect 33324 5646 33376 5652
rect 33230 5607 33286 5616
rect 32916 5188 33088 5216
rect 32864 5170 32916 5176
rect 32864 5024 32916 5030
rect 32784 4984 32864 5012
rect 32864 4966 32916 4972
rect 32588 4480 32640 4486
rect 32588 4422 32640 4428
rect 32404 4208 32456 4214
rect 32404 4150 32456 4156
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31852 4004 31904 4010
rect 31852 3946 31904 3952
rect 31220 3738 31248 3946
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 31864 3641 31892 3946
rect 32416 3738 32444 4150
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 31850 3632 31906 3641
rect 31024 3596 31076 3602
rect 31850 3567 31906 3576
rect 31024 3538 31076 3544
rect 31956 3534 31984 3674
rect 31944 3528 31996 3534
rect 31298 3496 31354 3505
rect 31354 3466 31432 3482
rect 31944 3470 31996 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 31354 3460 31444 3466
rect 31354 3454 31392 3460
rect 31298 3431 31354 3440
rect 31760 3460 31812 3466
rect 31444 3420 31524 3448
rect 31392 3402 31444 3408
rect 31070 3292 31378 3301
rect 31070 3290 31076 3292
rect 31132 3290 31156 3292
rect 31212 3290 31236 3292
rect 31292 3290 31316 3292
rect 31372 3290 31378 3292
rect 31132 3238 31134 3290
rect 31314 3238 31316 3290
rect 31070 3236 31076 3238
rect 31132 3236 31156 3238
rect 31212 3236 31236 3238
rect 31292 3236 31316 3238
rect 31372 3236 31378 3238
rect 31070 3227 31378 3236
rect 31496 3176 31524 3420
rect 31404 3148 31524 3176
rect 31588 3420 31760 3448
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31206 2680 31262 2689
rect 31206 2615 31262 2624
rect 31220 2514 31248 2615
rect 31312 2582 31340 2926
rect 31300 2576 31352 2582
rect 31300 2518 31352 2524
rect 31208 2508 31260 2514
rect 31208 2450 31260 2456
rect 31404 2417 31432 3148
rect 31588 3074 31616 3420
rect 31760 3402 31812 3408
rect 31496 3058 31616 3074
rect 31484 3052 31616 3058
rect 31536 3046 31616 3052
rect 31484 2994 31536 3000
rect 31484 2916 31536 2922
rect 31484 2858 31536 2864
rect 31390 2408 31446 2417
rect 31390 2343 31392 2352
rect 31444 2343 31446 2352
rect 31392 2314 31444 2320
rect 31496 2310 31524 2858
rect 31588 2836 31616 3046
rect 31668 2848 31720 2854
rect 31588 2808 31668 2836
rect 31484 2304 31536 2310
rect 31484 2246 31536 2252
rect 31070 2204 31378 2213
rect 31070 2202 31076 2204
rect 31132 2202 31156 2204
rect 31212 2202 31236 2204
rect 31292 2202 31316 2204
rect 31372 2202 31378 2204
rect 31132 2150 31134 2202
rect 31314 2150 31316 2202
rect 31070 2148 31076 2150
rect 31132 2148 31156 2150
rect 31212 2148 31236 2150
rect 31292 2148 31316 2150
rect 31372 2148 31378 2150
rect 31070 2139 31378 2148
rect 30932 2100 30984 2106
rect 30932 2042 30984 2048
rect 30564 1828 30616 1834
rect 30564 1770 30616 1776
rect 30012 1760 30064 1766
rect 30012 1702 30064 1708
rect 30472 1760 30524 1766
rect 30472 1702 30524 1708
rect 30840 1760 30892 1766
rect 30840 1702 30892 1708
rect 29920 1556 29972 1562
rect 29920 1498 29972 1504
rect 30012 1556 30064 1562
rect 30012 1498 30064 1504
rect 29276 1284 29328 1290
rect 29276 1226 29328 1232
rect 29736 1284 29788 1290
rect 29736 1226 29788 1232
rect 30024 160 30052 1498
rect 30484 1465 30512 1702
rect 30470 1456 30526 1465
rect 30470 1391 30526 1400
rect 30288 1284 30340 1290
rect 30288 1226 30340 1232
rect 30300 1018 30328 1226
rect 30380 1216 30432 1222
rect 30380 1158 30432 1164
rect 30288 1012 30340 1018
rect 30288 954 30340 960
rect 30392 678 30420 1158
rect 30380 672 30432 678
rect 30380 614 30432 620
rect 30852 160 30880 1702
rect 31496 1358 31524 2246
rect 31588 1834 31616 2808
rect 31668 2790 31720 2796
rect 31956 2689 31984 3470
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 32048 3194 32076 3334
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 31942 2680 31998 2689
rect 31942 2615 31998 2624
rect 32034 2408 32090 2417
rect 31944 2372 31996 2378
rect 32090 2366 32168 2394
rect 32034 2343 32090 2352
rect 31944 2314 31996 2320
rect 31852 2100 31904 2106
rect 31852 2042 31904 2048
rect 31864 1970 31892 2042
rect 31956 2009 31984 2314
rect 31942 2000 31998 2009
rect 31852 1964 31904 1970
rect 31942 1935 31944 1944
rect 31852 1906 31904 1912
rect 31996 1935 31998 1944
rect 31944 1906 31996 1912
rect 31576 1828 31628 1834
rect 31576 1770 31628 1776
rect 31668 1556 31720 1562
rect 31668 1498 31720 1504
rect 31392 1352 31444 1358
rect 31392 1294 31444 1300
rect 31484 1352 31536 1358
rect 31484 1294 31536 1300
rect 31404 1170 31432 1294
rect 31404 1142 31524 1170
rect 31070 1116 31378 1125
rect 31070 1114 31076 1116
rect 31132 1114 31156 1116
rect 31212 1114 31236 1116
rect 31292 1114 31316 1116
rect 31372 1114 31378 1116
rect 31132 1062 31134 1114
rect 31314 1062 31316 1114
rect 31070 1060 31076 1062
rect 31132 1060 31156 1062
rect 31212 1060 31236 1062
rect 31292 1060 31316 1062
rect 31372 1060 31378 1062
rect 31070 1051 31378 1060
rect 31496 882 31524 1142
rect 31484 876 31536 882
rect 31484 818 31536 824
rect 31680 160 31708 1498
rect 32036 1488 32088 1494
rect 32036 1430 32088 1436
rect 32048 1358 32076 1430
rect 32036 1352 32088 1358
rect 32036 1294 32088 1300
rect 32140 1222 32168 2366
rect 32324 2038 32352 3470
rect 32600 2961 32628 4422
rect 32876 3602 32904 4966
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32968 3738 32996 4762
rect 33060 4554 33088 5188
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 32956 3732 33008 3738
rect 32956 3674 33008 3680
rect 33152 3602 33180 4014
rect 33244 3738 33272 5607
rect 33324 5024 33376 5030
rect 33324 4966 33376 4972
rect 33336 4282 33364 4966
rect 33324 4276 33376 4282
rect 33324 4218 33376 4224
rect 33428 4146 33456 5664
rect 33570 4924 33878 4933
rect 33570 4922 33576 4924
rect 33632 4922 33656 4924
rect 33712 4922 33736 4924
rect 33792 4922 33816 4924
rect 33872 4922 33878 4924
rect 33632 4870 33634 4922
rect 33814 4870 33816 4922
rect 33570 4868 33576 4870
rect 33632 4868 33656 4870
rect 33712 4868 33736 4870
rect 33792 4868 33816 4870
rect 33872 4868 33878 4870
rect 33570 4859 33878 4868
rect 33966 4856 34022 4865
rect 33966 4791 34022 4800
rect 33416 4140 33468 4146
rect 33416 4082 33468 4088
rect 33980 4010 34008 4791
rect 34072 4758 34100 5714
rect 34164 5166 34192 6054
rect 34256 5166 34284 6190
rect 34532 5778 34560 7398
rect 34716 7324 34744 9551
rect 34900 9518 34928 9574
rect 34796 9512 34848 9518
rect 34796 9454 34848 9460
rect 34888 9512 34940 9518
rect 34888 9454 34940 9460
rect 35808 9512 35860 9518
rect 35808 9454 35860 9460
rect 34808 8566 34836 9454
rect 34888 9104 34940 9110
rect 34888 9046 34940 9052
rect 34980 9104 35032 9110
rect 34980 9046 35032 9052
rect 35530 9072 35586 9081
rect 34900 8809 34928 9046
rect 34992 8906 35020 9046
rect 35530 9007 35532 9016
rect 35584 9007 35586 9016
rect 35532 8978 35584 8984
rect 35440 8968 35492 8974
rect 35492 8916 35756 8922
rect 35440 8910 35756 8916
rect 34980 8900 35032 8906
rect 35452 8894 35756 8910
rect 35820 8906 35848 9454
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35912 9178 35940 9318
rect 36082 9208 36138 9217
rect 35900 9172 35952 9178
rect 35900 9114 35952 9120
rect 35992 9172 36044 9178
rect 36138 9178 36216 9194
rect 36138 9172 36228 9178
rect 36138 9166 36176 9172
rect 36082 9143 36138 9152
rect 35992 9114 36044 9120
rect 36176 9114 36228 9120
rect 34980 8842 35032 8848
rect 35624 8832 35676 8838
rect 34886 8800 34942 8809
rect 35624 8774 35676 8780
rect 34886 8735 34942 8744
rect 34886 8664 34942 8673
rect 34886 8599 34942 8608
rect 34900 8566 34928 8599
rect 34796 8560 34848 8566
rect 34796 8502 34848 8508
rect 34888 8560 34940 8566
rect 34888 8502 34940 8508
rect 35348 8560 35400 8566
rect 35348 8502 35400 8508
rect 34808 8294 34836 8502
rect 35360 8401 35388 8502
rect 35346 8392 35402 8401
rect 35346 8327 35402 8336
rect 34808 8266 35112 8294
rect 35084 7886 35112 8266
rect 35072 7880 35124 7886
rect 35072 7822 35124 7828
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 34624 7296 34744 7324
rect 34624 6730 34652 7296
rect 34900 7002 34928 7346
rect 34980 7200 35032 7206
rect 34980 7142 35032 7148
rect 34888 6996 34940 7002
rect 34888 6938 34940 6944
rect 34992 6934 35020 7142
rect 34980 6928 35032 6934
rect 34980 6870 35032 6876
rect 34612 6724 34664 6730
rect 34612 6666 34664 6672
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34888 6656 34940 6662
rect 34888 6598 34940 6604
rect 34716 6458 34744 6598
rect 34704 6452 34756 6458
rect 34704 6394 34756 6400
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34624 5914 34652 6190
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34520 5772 34572 5778
rect 34520 5714 34572 5720
rect 34336 5704 34388 5710
rect 34336 5646 34388 5652
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 34348 5370 34376 5646
rect 34336 5364 34388 5370
rect 34336 5306 34388 5312
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 34244 5160 34296 5166
rect 34244 5102 34296 5108
rect 34164 5030 34192 5102
rect 34152 5024 34204 5030
rect 34152 4966 34204 4972
rect 34060 4752 34112 4758
rect 34060 4694 34112 4700
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 34072 4060 34100 4558
rect 34164 4214 34192 4966
rect 34152 4208 34204 4214
rect 34152 4150 34204 4156
rect 34152 4072 34204 4078
rect 34072 4032 34152 4060
rect 34256 4060 34284 5102
rect 34348 4826 34376 5306
rect 34520 5228 34572 5234
rect 34520 5170 34572 5176
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34336 4820 34388 4826
rect 34336 4762 34388 4768
rect 34440 4690 34468 4966
rect 34532 4826 34560 5170
rect 34716 5166 34744 5646
rect 34704 5160 34756 5166
rect 34704 5102 34756 5108
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 34204 4032 34284 4060
rect 34428 4072 34480 4078
rect 34152 4014 34204 4020
rect 34428 4014 34480 4020
rect 33968 4004 34020 4010
rect 33968 3946 34020 3952
rect 33570 3836 33878 3845
rect 33570 3834 33576 3836
rect 33632 3834 33656 3836
rect 33712 3834 33736 3836
rect 33792 3834 33816 3836
rect 33872 3834 33878 3836
rect 33632 3782 33634 3834
rect 33814 3782 33816 3834
rect 33570 3780 33576 3782
rect 33632 3780 33656 3782
rect 33712 3780 33736 3782
rect 33792 3780 33816 3782
rect 33872 3780 33878 3782
rect 33570 3771 33878 3780
rect 33232 3732 33284 3738
rect 33232 3674 33284 3680
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 33140 3596 33192 3602
rect 33140 3538 33192 3544
rect 32692 3194 32720 3538
rect 33416 3528 33468 3534
rect 33244 3488 33416 3516
rect 33140 3460 33192 3466
rect 33140 3402 33192 3408
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32586 2952 32642 2961
rect 32586 2887 32642 2896
rect 32494 2680 32550 2689
rect 32494 2615 32550 2624
rect 32312 2032 32364 2038
rect 32312 1974 32364 1980
rect 32220 1896 32272 1902
rect 32220 1838 32272 1844
rect 32232 1562 32260 1838
rect 32220 1556 32272 1562
rect 32220 1498 32272 1504
rect 32312 1420 32364 1426
rect 32312 1362 32364 1368
rect 32324 1272 32352 1362
rect 32508 1358 32536 2615
rect 32784 2417 32812 3334
rect 33060 3210 33088 3334
rect 32876 3182 33088 3210
rect 32876 2514 32904 3182
rect 32956 3120 33008 3126
rect 32956 3062 33008 3068
rect 32864 2508 32916 2514
rect 32864 2450 32916 2456
rect 32968 2446 32996 3062
rect 33152 2446 33180 3402
rect 33244 2650 33272 3488
rect 33416 3470 33468 3476
rect 33690 3496 33746 3505
rect 33690 3431 33692 3440
rect 33744 3431 33746 3440
rect 33692 3402 33744 3408
rect 33508 3052 33560 3058
rect 33428 3012 33508 3040
rect 33232 2644 33284 2650
rect 33232 2586 33284 2592
rect 32956 2440 33008 2446
rect 32770 2408 32826 2417
rect 32956 2382 33008 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 32770 2343 32826 2352
rect 32968 1902 32996 2382
rect 33232 2304 33284 2310
rect 33232 2246 33284 2252
rect 32956 1896 33008 1902
rect 32956 1838 33008 1844
rect 33244 1358 33272 2246
rect 33324 1760 33376 1766
rect 33324 1702 33376 1708
rect 33336 1494 33364 1702
rect 33324 1488 33376 1494
rect 33324 1430 33376 1436
rect 32496 1352 32548 1358
rect 32496 1294 32548 1300
rect 33048 1352 33100 1358
rect 33048 1294 33100 1300
rect 33232 1352 33284 1358
rect 33232 1294 33284 1300
rect 32404 1284 32456 1290
rect 32324 1244 32404 1272
rect 32404 1226 32456 1232
rect 32864 1284 32916 1290
rect 32864 1226 32916 1232
rect 32128 1216 32180 1222
rect 32128 1158 32180 1164
rect 32876 1018 32904 1226
rect 33060 1222 33088 1294
rect 33428 1222 33456 3012
rect 33508 2994 33560 3000
rect 33796 2922 34008 2938
rect 33784 2916 34008 2922
rect 33836 2910 34008 2916
rect 33784 2858 33836 2864
rect 33570 2748 33878 2757
rect 33570 2746 33576 2748
rect 33632 2746 33656 2748
rect 33712 2746 33736 2748
rect 33792 2746 33816 2748
rect 33872 2746 33878 2748
rect 33632 2694 33634 2746
rect 33814 2694 33816 2746
rect 33570 2692 33576 2694
rect 33632 2692 33656 2694
rect 33712 2692 33736 2694
rect 33792 2692 33816 2694
rect 33872 2692 33878 2694
rect 33570 2683 33878 2692
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33520 2106 33548 2246
rect 33508 2100 33560 2106
rect 33508 2042 33560 2048
rect 33796 2009 33824 2382
rect 33782 2000 33838 2009
rect 33782 1935 33784 1944
rect 33836 1935 33838 1944
rect 33784 1906 33836 1912
rect 33570 1660 33878 1669
rect 33570 1658 33576 1660
rect 33632 1658 33656 1660
rect 33712 1658 33736 1660
rect 33792 1658 33816 1660
rect 33872 1658 33878 1660
rect 33632 1606 33634 1658
rect 33814 1606 33816 1658
rect 33570 1604 33576 1606
rect 33632 1604 33656 1606
rect 33712 1604 33736 1606
rect 33792 1604 33816 1606
rect 33872 1604 33878 1606
rect 33570 1595 33878 1604
rect 33980 1426 34008 2910
rect 34060 2848 34112 2854
rect 34060 2790 34112 2796
rect 34072 2020 34100 2790
rect 34164 2650 34192 4014
rect 34440 3738 34468 4014
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34612 3528 34664 3534
rect 34612 3470 34664 3476
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34440 2774 34468 3334
rect 34624 3194 34652 3470
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 34348 2746 34468 2774
rect 34532 2774 34560 2926
rect 34532 2746 34744 2774
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 34348 2514 34376 2746
rect 34336 2508 34388 2514
rect 34336 2450 34388 2456
rect 34152 2032 34204 2038
rect 34072 1992 34152 2020
rect 34152 1974 34204 1980
rect 34244 1896 34296 1902
rect 34244 1838 34296 1844
rect 33968 1420 34020 1426
rect 33968 1362 34020 1368
rect 34256 1358 34284 1838
rect 34716 1358 34744 2746
rect 34900 1902 34928 6598
rect 35084 6236 35112 7822
rect 35162 7440 35218 7449
rect 35162 7375 35218 7384
rect 35176 7342 35204 7375
rect 35164 7336 35216 7342
rect 35164 7278 35216 7284
rect 35256 6724 35308 6730
rect 35256 6666 35308 6672
rect 35268 6458 35296 6666
rect 35532 6656 35584 6662
rect 35532 6598 35584 6604
rect 35256 6452 35308 6458
rect 35256 6394 35308 6400
rect 35256 6248 35308 6254
rect 35084 6208 35256 6236
rect 35256 6190 35308 6196
rect 35268 5710 35296 6190
rect 35544 5914 35572 6598
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 35256 5704 35308 5710
rect 35256 5646 35308 5652
rect 35348 5024 35400 5030
rect 35348 4966 35400 4972
rect 35360 4758 35388 4966
rect 35348 4752 35400 4758
rect 35348 4694 35400 4700
rect 35348 4480 35400 4486
rect 35400 4440 35480 4468
rect 35348 4422 35400 4428
rect 35256 3120 35308 3126
rect 35256 3062 35308 3068
rect 35268 2825 35296 3062
rect 35254 2816 35310 2825
rect 35176 2774 35254 2802
rect 34888 1896 34940 1902
rect 34888 1838 34940 1844
rect 34980 1556 35032 1562
rect 34980 1498 35032 1504
rect 33876 1352 33928 1358
rect 33874 1320 33876 1329
rect 34244 1352 34296 1358
rect 33928 1320 33930 1329
rect 34244 1294 34296 1300
rect 34704 1352 34756 1358
rect 34704 1294 34756 1300
rect 33874 1255 33930 1264
rect 33048 1216 33100 1222
rect 33048 1158 33100 1164
rect 33416 1216 33468 1222
rect 33416 1158 33468 1164
rect 34336 1216 34388 1222
rect 34336 1158 34388 1164
rect 32864 1012 32916 1018
rect 32864 954 32916 960
rect 34348 950 34376 1158
rect 34336 944 34388 950
rect 34336 886 34388 892
rect 32680 808 32732 814
rect 32508 756 32680 762
rect 32508 750 32732 756
rect 32508 734 32720 750
rect 34428 740 34480 746
rect 32508 160 32536 734
rect 34428 682 34480 688
rect 33508 672 33560 678
rect 33336 620 33508 626
rect 33336 614 33560 620
rect 33336 598 33548 614
rect 33336 160 33364 598
rect 34164 190 34284 218
rect 34164 160 34192 190
rect 28354 54 28856 82
rect 28354 -300 28410 54
rect 29182 -300 29238 160
rect 30010 -300 30066 160
rect 30838 -300 30894 160
rect 31666 -300 31722 160
rect 32494 -300 32550 160
rect 33322 -300 33378 160
rect 34150 -300 34206 160
rect 34256 82 34284 190
rect 34440 82 34468 682
rect 34992 160 35020 1498
rect 35176 1358 35204 2774
rect 35254 2751 35310 2760
rect 35452 2774 35480 4440
rect 35452 2746 35572 2774
rect 35256 2304 35308 2310
rect 35256 2246 35308 2252
rect 35268 1494 35296 2246
rect 35544 2106 35572 2746
rect 35532 2100 35584 2106
rect 35532 2042 35584 2048
rect 35636 1986 35664 8774
rect 35728 8616 35756 8894
rect 35808 8900 35860 8906
rect 35808 8842 35860 8848
rect 35808 8628 35860 8634
rect 35728 8588 35808 8616
rect 36004 8616 36032 9114
rect 36556 8974 36584 10202
rect 36728 9920 36780 9926
rect 36728 9862 36780 9868
rect 36636 9512 36688 9518
rect 36636 9454 36688 9460
rect 36648 8974 36676 9454
rect 36544 8968 36596 8974
rect 36174 8936 36230 8945
rect 36544 8910 36596 8916
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 36174 8871 36176 8880
rect 36228 8871 36230 8880
rect 36176 8842 36228 8848
rect 36544 8832 36596 8838
rect 36544 8774 36596 8780
rect 36070 8732 36378 8741
rect 36070 8730 36076 8732
rect 36132 8730 36156 8732
rect 36212 8730 36236 8732
rect 36292 8730 36316 8732
rect 36372 8730 36378 8732
rect 36132 8678 36134 8730
rect 36314 8678 36316 8730
rect 36070 8676 36076 8678
rect 36132 8676 36156 8678
rect 36212 8676 36236 8678
rect 36292 8676 36316 8678
rect 36372 8676 36378 8678
rect 36070 8667 36378 8676
rect 35860 8588 35940 8616
rect 36004 8588 36124 8616
rect 35808 8570 35860 8576
rect 35716 7744 35768 7750
rect 35716 7686 35768 7692
rect 35808 7744 35860 7750
rect 35808 7686 35860 7692
rect 35728 6769 35756 7686
rect 35714 6760 35770 6769
rect 35714 6695 35770 6704
rect 35728 4554 35756 6695
rect 35820 6186 35848 7686
rect 35912 7528 35940 8588
rect 36096 8430 36124 8588
rect 36176 8560 36228 8566
rect 36556 8537 36584 8774
rect 36176 8502 36228 8508
rect 36542 8528 36598 8537
rect 36084 8424 36136 8430
rect 36188 8401 36216 8502
rect 36648 8498 36676 8910
rect 36542 8463 36598 8472
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 36084 8366 36136 8372
rect 36174 8392 36230 8401
rect 36174 8327 36230 8336
rect 36188 7750 36216 8327
rect 36740 8090 36768 9862
rect 36832 9654 36860 10639
rect 37096 10600 37148 10606
rect 37096 10542 37148 10548
rect 37738 10568 37794 10577
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 36820 9648 36872 9654
rect 36820 9590 36872 9596
rect 36924 8090 36952 9998
rect 37004 9920 37056 9926
rect 37004 9862 37056 9868
rect 37016 9042 37044 9862
rect 37108 9586 37136 10542
rect 37738 10503 37794 10512
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 37292 9654 37320 9862
rect 37280 9648 37332 9654
rect 37280 9590 37332 9596
rect 37464 9648 37516 9654
rect 37464 9590 37516 9596
rect 37096 9580 37148 9586
rect 37096 9522 37148 9528
rect 37188 9376 37240 9382
rect 37188 9318 37240 9324
rect 37004 9036 37056 9042
rect 37004 8978 37056 8984
rect 37096 9036 37148 9042
rect 37096 8978 37148 8984
rect 37108 8294 37136 8978
rect 37096 8288 37148 8294
rect 37096 8230 37148 8236
rect 36728 8084 36780 8090
rect 36728 8026 36780 8032
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 36634 7984 36690 7993
rect 36634 7919 36690 7928
rect 37004 7948 37056 7954
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 36070 7644 36378 7653
rect 36070 7642 36076 7644
rect 36132 7642 36156 7644
rect 36212 7642 36236 7644
rect 36292 7642 36316 7644
rect 36372 7642 36378 7644
rect 36132 7590 36134 7642
rect 36314 7590 36316 7642
rect 36070 7588 36076 7590
rect 36132 7588 36156 7590
rect 36212 7588 36236 7590
rect 36292 7588 36316 7590
rect 36372 7588 36378 7590
rect 36070 7579 36378 7588
rect 35992 7540 36044 7546
rect 35912 7500 35992 7528
rect 35992 7482 36044 7488
rect 35898 7304 35954 7313
rect 35898 7239 35954 7248
rect 36176 7268 36228 7274
rect 35808 6180 35860 6186
rect 35808 6122 35860 6128
rect 35716 4548 35768 4554
rect 35716 4490 35768 4496
rect 35808 4480 35860 4486
rect 35808 4422 35860 4428
rect 35716 3596 35768 3602
rect 35716 3538 35768 3544
rect 35728 2689 35756 3538
rect 35820 3534 35848 4422
rect 35912 4146 35940 7239
rect 36176 7210 36228 7216
rect 35992 6792 36044 6798
rect 35990 6760 35992 6769
rect 36044 6760 36046 6769
rect 36188 6730 36216 7210
rect 35990 6695 36046 6704
rect 36176 6724 36228 6730
rect 36176 6666 36228 6672
rect 36452 6656 36504 6662
rect 36648 6644 36676 7919
rect 37004 7890 37056 7896
rect 36728 7744 36780 7750
rect 36728 7686 36780 7692
rect 36740 6798 36768 7686
rect 37016 7342 37044 7890
rect 37096 7812 37148 7818
rect 37096 7754 37148 7760
rect 37108 7410 37136 7754
rect 37096 7404 37148 7410
rect 37096 7346 37148 7352
rect 37004 7336 37056 7342
rect 37004 7278 37056 7284
rect 37200 7206 37228 9318
rect 37476 8906 37504 9590
rect 37464 8900 37516 8906
rect 37464 8842 37516 8848
rect 37372 8560 37424 8566
rect 37476 8548 37504 8842
rect 37424 8520 37504 8548
rect 37372 8502 37424 8508
rect 37476 8090 37504 8520
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37464 8084 37516 8090
rect 37464 8026 37516 8032
rect 37568 7954 37596 8230
rect 37752 7993 37780 10503
rect 37924 9920 37976 9926
rect 37924 9862 37976 9868
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 37936 8294 37964 9862
rect 38028 9178 38056 9862
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 37924 8288 37976 8294
rect 37924 8230 37976 8236
rect 37738 7984 37794 7993
rect 37556 7948 37608 7954
rect 37556 7890 37608 7896
rect 37648 7948 37700 7954
rect 37738 7919 37794 7928
rect 37648 7890 37700 7896
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37372 7472 37424 7478
rect 37292 7420 37372 7426
rect 37292 7414 37424 7420
rect 37292 7398 37412 7414
rect 37188 7200 37240 7206
rect 37188 7142 37240 7148
rect 37292 6882 37320 7398
rect 37372 7336 37424 7342
rect 37476 7324 37504 7822
rect 37660 7342 37688 7890
rect 37752 7342 37780 7919
rect 37424 7296 37504 7324
rect 37648 7336 37700 7342
rect 37372 7278 37424 7284
rect 37648 7278 37700 7284
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37752 6934 37780 7278
rect 36924 6866 37320 6882
rect 37740 6928 37792 6934
rect 38120 6905 38148 12566
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 38200 12164 38252 12170
rect 38200 12106 38252 12112
rect 38212 11694 38240 12106
rect 38304 11898 38332 12174
rect 38292 11892 38344 11898
rect 38292 11834 38344 11840
rect 38200 11688 38252 11694
rect 38200 11630 38252 11636
rect 38396 10266 38424 18770
rect 38476 18760 38528 18766
rect 38476 18702 38528 18708
rect 38488 18154 38516 18702
rect 38948 18222 38976 19207
rect 39028 19168 39080 19174
rect 39028 19110 39080 19116
rect 39040 18834 39068 19110
rect 39224 18834 39252 19246
rect 39028 18828 39080 18834
rect 39028 18770 39080 18776
rect 39212 18828 39264 18834
rect 39212 18770 39264 18776
rect 39040 18426 39068 18770
rect 39316 18426 39344 22374
rect 39684 21894 39712 22714
rect 40420 22642 40448 23840
rect 41340 23746 41368 23840
rect 41432 23746 41460 23854
rect 41340 23718 41460 23746
rect 40960 23044 41012 23050
rect 40960 22986 41012 22992
rect 40972 22778 41000 22986
rect 41070 22876 41378 22885
rect 41070 22874 41076 22876
rect 41132 22874 41156 22876
rect 41212 22874 41236 22876
rect 41292 22874 41316 22876
rect 41372 22874 41378 22876
rect 41132 22822 41134 22874
rect 41314 22822 41316 22874
rect 41070 22820 41076 22822
rect 41132 22820 41156 22822
rect 41212 22820 41236 22822
rect 41292 22820 41316 22822
rect 41372 22820 41378 22822
rect 41070 22811 41378 22820
rect 40960 22772 41012 22778
rect 40960 22714 41012 22720
rect 41616 22642 41644 23854
rect 42246 23840 42302 24300
rect 43166 23840 43222 24300
rect 44086 23840 44142 24300
rect 45006 23840 45062 24300
rect 42260 22642 42288 23840
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 42812 22778 42840 22918
rect 42800 22772 42852 22778
rect 42800 22714 42852 22720
rect 43180 22642 43208 23840
rect 40408 22636 40460 22642
rect 40408 22578 40460 22584
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 43168 22636 43220 22642
rect 44100 22624 44128 23840
rect 44272 22636 44324 22642
rect 44100 22596 44272 22624
rect 43168 22578 43220 22584
rect 45020 22624 45048 23840
rect 45192 22636 45244 22642
rect 45020 22596 45192 22624
rect 44272 22578 44324 22584
rect 45192 22578 45244 22584
rect 40960 22500 41012 22506
rect 40960 22442 41012 22448
rect 40500 22432 40552 22438
rect 40500 22374 40552 22380
rect 40040 22092 40092 22098
rect 40040 22034 40092 22040
rect 39672 21888 39724 21894
rect 39672 21830 39724 21836
rect 39764 21888 39816 21894
rect 39764 21830 39816 21836
rect 39684 20602 39712 21830
rect 39776 21554 39804 21830
rect 39764 21548 39816 21554
rect 39764 21490 39816 21496
rect 39776 20874 39804 21490
rect 39764 20868 39816 20874
rect 39764 20810 39816 20816
rect 39776 20602 39804 20810
rect 39672 20596 39724 20602
rect 39672 20538 39724 20544
rect 39764 20596 39816 20602
rect 39764 20538 39816 20544
rect 39396 20324 39448 20330
rect 39396 20266 39448 20272
rect 39408 19990 39436 20266
rect 39396 19984 39448 19990
rect 39396 19926 39448 19932
rect 39580 19712 39632 19718
rect 39580 19654 39632 19660
rect 39592 19514 39620 19654
rect 39580 19508 39632 19514
rect 39580 19450 39632 19456
rect 39776 19446 39804 20538
rect 40052 20534 40080 22034
rect 40512 21690 40540 22374
rect 40972 22234 41000 22442
rect 41420 22432 41472 22438
rect 41420 22374 41472 22380
rect 42156 22432 42208 22438
rect 42156 22374 42208 22380
rect 42708 22432 42760 22438
rect 42708 22374 42760 22380
rect 43260 22432 43312 22438
rect 43260 22374 43312 22380
rect 43904 22432 43956 22438
rect 43904 22374 43956 22380
rect 44180 22432 44232 22438
rect 44180 22374 44232 22380
rect 44364 22432 44416 22438
rect 44364 22374 44416 22380
rect 45008 22432 45060 22438
rect 45008 22374 45060 22380
rect 40960 22228 41012 22234
rect 40960 22170 41012 22176
rect 40972 21690 41000 22170
rect 41070 21788 41378 21797
rect 41070 21786 41076 21788
rect 41132 21786 41156 21788
rect 41212 21786 41236 21788
rect 41292 21786 41316 21788
rect 41372 21786 41378 21788
rect 41132 21734 41134 21786
rect 41314 21734 41316 21786
rect 41070 21732 41076 21734
rect 41132 21732 41156 21734
rect 41212 21732 41236 21734
rect 41292 21732 41316 21734
rect 41372 21732 41378 21734
rect 41070 21723 41378 21732
rect 40500 21684 40552 21690
rect 40500 21626 40552 21632
rect 40960 21684 41012 21690
rect 40960 21626 41012 21632
rect 40776 21480 40828 21486
rect 40776 21422 40828 21428
rect 40868 21480 40920 21486
rect 40868 21422 40920 21428
rect 40500 21412 40552 21418
rect 40500 21354 40552 21360
rect 40512 21146 40540 21354
rect 40788 21146 40816 21422
rect 40500 21140 40552 21146
rect 40500 21082 40552 21088
rect 40776 21140 40828 21146
rect 40776 21082 40828 21088
rect 40880 20874 40908 21422
rect 41432 20942 41460 22374
rect 41696 22024 41748 22030
rect 41696 21966 41748 21972
rect 41604 21004 41656 21010
rect 41604 20946 41656 20952
rect 41420 20936 41472 20942
rect 41420 20878 41472 20884
rect 40868 20868 40920 20874
rect 40868 20810 40920 20816
rect 40960 20800 41012 20806
rect 40960 20742 41012 20748
rect 40776 20596 40828 20602
rect 40776 20538 40828 20544
rect 40040 20528 40092 20534
rect 40040 20470 40092 20476
rect 39856 19916 39908 19922
rect 39856 19858 39908 19864
rect 39764 19440 39816 19446
rect 39764 19382 39816 19388
rect 39776 18698 39804 19382
rect 39488 18692 39540 18698
rect 39488 18634 39540 18640
rect 39764 18692 39816 18698
rect 39764 18634 39816 18640
rect 39028 18420 39080 18426
rect 39028 18362 39080 18368
rect 39304 18420 39356 18426
rect 39304 18362 39356 18368
rect 38936 18216 38988 18222
rect 38936 18158 38988 18164
rect 38476 18148 38528 18154
rect 38476 18090 38528 18096
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 39028 18080 39080 18086
rect 39028 18022 39080 18028
rect 38570 17980 38878 17989
rect 38570 17978 38576 17980
rect 38632 17978 38656 17980
rect 38712 17978 38736 17980
rect 38792 17978 38816 17980
rect 38872 17978 38878 17980
rect 38632 17926 38634 17978
rect 38814 17926 38816 17978
rect 38570 17924 38576 17926
rect 38632 17924 38656 17926
rect 38712 17924 38736 17926
rect 38792 17924 38816 17926
rect 38872 17924 38878 17926
rect 38570 17915 38878 17924
rect 38948 17626 38976 18022
rect 39040 17746 39068 18022
rect 39500 17882 39528 18634
rect 39868 18222 39896 19858
rect 40788 19786 40816 20538
rect 40776 19780 40828 19786
rect 40776 19722 40828 19728
rect 39948 19712 40000 19718
rect 39948 19654 40000 19660
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 39960 18970 39988 19654
rect 40880 19514 40908 19654
rect 40868 19508 40920 19514
rect 40868 19450 40920 19456
rect 40972 18970 41000 20742
rect 41070 20700 41378 20709
rect 41070 20698 41076 20700
rect 41132 20698 41156 20700
rect 41212 20698 41236 20700
rect 41292 20698 41316 20700
rect 41372 20698 41378 20700
rect 41132 20646 41134 20698
rect 41314 20646 41316 20698
rect 41070 20644 41076 20646
rect 41132 20644 41156 20646
rect 41212 20644 41236 20646
rect 41292 20644 41316 20646
rect 41372 20644 41378 20646
rect 41070 20635 41378 20644
rect 41420 20460 41472 20466
rect 41420 20402 41472 20408
rect 41432 19922 41460 20402
rect 41420 19916 41472 19922
rect 41420 19858 41472 19864
rect 41070 19612 41378 19621
rect 41070 19610 41076 19612
rect 41132 19610 41156 19612
rect 41212 19610 41236 19612
rect 41292 19610 41316 19612
rect 41372 19610 41378 19612
rect 41132 19558 41134 19610
rect 41314 19558 41316 19610
rect 41070 19556 41076 19558
rect 41132 19556 41156 19558
rect 41212 19556 41236 19558
rect 41292 19556 41316 19558
rect 41372 19556 41378 19558
rect 41070 19547 41378 19556
rect 41432 19242 41460 19858
rect 41512 19372 41564 19378
rect 41512 19314 41564 19320
rect 41420 19236 41472 19242
rect 41420 19178 41472 19184
rect 39948 18964 40000 18970
rect 40960 18964 41012 18970
rect 40000 18924 40080 18952
rect 39948 18906 40000 18912
rect 40052 18426 40080 18924
rect 40960 18906 41012 18912
rect 40960 18828 41012 18834
rect 40960 18770 41012 18776
rect 40040 18420 40092 18426
rect 40040 18362 40092 18368
rect 40972 18358 41000 18770
rect 41432 18766 41460 19178
rect 41524 18970 41552 19314
rect 41616 19310 41644 20946
rect 41708 20262 41736 21966
rect 42168 21894 42196 22374
rect 41972 21888 42024 21894
rect 41972 21830 42024 21836
rect 42156 21888 42208 21894
rect 42156 21830 42208 21836
rect 41984 21690 42012 21830
rect 41972 21684 42024 21690
rect 41972 21626 42024 21632
rect 42168 21350 42196 21830
rect 42156 21344 42208 21350
rect 42156 21286 42208 21292
rect 41878 20904 41934 20913
rect 41878 20839 41934 20848
rect 41892 20806 41920 20839
rect 41880 20800 41932 20806
rect 41880 20742 41932 20748
rect 42340 20800 42392 20806
rect 42340 20742 42392 20748
rect 42352 20602 42380 20742
rect 42340 20596 42392 20602
rect 42340 20538 42392 20544
rect 42064 20528 42116 20534
rect 42064 20470 42116 20476
rect 41788 20392 41840 20398
rect 41788 20334 41840 20340
rect 41696 20256 41748 20262
rect 41696 20198 41748 20204
rect 41696 20052 41748 20058
rect 41696 19994 41748 20000
rect 41708 19514 41736 19994
rect 41800 19514 41828 20334
rect 42076 19854 42104 20470
rect 42340 20392 42392 20398
rect 42340 20334 42392 20340
rect 42064 19848 42116 19854
rect 42064 19790 42116 19796
rect 41696 19508 41748 19514
rect 41696 19450 41748 19456
rect 41788 19508 41840 19514
rect 41788 19450 41840 19456
rect 41604 19304 41656 19310
rect 41604 19246 41656 19252
rect 41616 18970 41644 19246
rect 41512 18964 41564 18970
rect 41512 18906 41564 18912
rect 41604 18964 41656 18970
rect 41604 18906 41656 18912
rect 41616 18850 41644 18906
rect 41616 18822 41920 18850
rect 41420 18760 41472 18766
rect 41420 18702 41472 18708
rect 41512 18760 41564 18766
rect 41512 18702 41564 18708
rect 41070 18524 41378 18533
rect 41070 18522 41076 18524
rect 41132 18522 41156 18524
rect 41212 18522 41236 18524
rect 41292 18522 41316 18524
rect 41372 18522 41378 18524
rect 41132 18470 41134 18522
rect 41314 18470 41316 18522
rect 41070 18468 41076 18470
rect 41132 18468 41156 18470
rect 41212 18468 41236 18470
rect 41292 18468 41316 18470
rect 41372 18468 41378 18470
rect 41070 18459 41378 18468
rect 41524 18426 41552 18702
rect 41696 18624 41748 18630
rect 41696 18566 41748 18572
rect 41512 18420 41564 18426
rect 41512 18362 41564 18368
rect 40960 18352 41012 18358
rect 40960 18294 41012 18300
rect 39856 18216 39908 18222
rect 39856 18158 39908 18164
rect 40316 18216 40368 18222
rect 40316 18158 40368 18164
rect 40328 17882 40356 18158
rect 40592 18080 40644 18086
rect 40592 18022 40644 18028
rect 39488 17876 39540 17882
rect 39488 17818 39540 17824
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 40316 17876 40368 17882
rect 40316 17818 40368 17824
rect 40052 17785 40080 17818
rect 40038 17776 40094 17785
rect 39028 17740 39080 17746
rect 39028 17682 39080 17688
rect 39488 17740 39540 17746
rect 40038 17711 40094 17720
rect 39488 17682 39540 17688
rect 38948 17598 39252 17626
rect 38948 17270 38976 17598
rect 39120 17536 39172 17542
rect 39120 17478 39172 17484
rect 39028 17332 39080 17338
rect 39028 17274 39080 17280
rect 38936 17264 38988 17270
rect 38936 17206 38988 17212
rect 38936 16992 38988 16998
rect 38936 16934 38988 16940
rect 38570 16892 38878 16901
rect 38570 16890 38576 16892
rect 38632 16890 38656 16892
rect 38712 16890 38736 16892
rect 38792 16890 38816 16892
rect 38872 16890 38878 16892
rect 38632 16838 38634 16890
rect 38814 16838 38816 16890
rect 38570 16836 38576 16838
rect 38632 16836 38656 16838
rect 38712 16836 38736 16838
rect 38792 16836 38816 16838
rect 38872 16836 38878 16838
rect 38570 16827 38878 16836
rect 38844 16652 38896 16658
rect 38844 16594 38896 16600
rect 38856 16522 38884 16594
rect 38948 16590 38976 16934
rect 39040 16658 39068 17274
rect 39132 16794 39160 17478
rect 39120 16788 39172 16794
rect 39120 16730 39172 16736
rect 39224 16726 39252 17598
rect 39396 17536 39448 17542
rect 39396 17478 39448 17484
rect 39212 16720 39264 16726
rect 39212 16662 39264 16668
rect 39028 16652 39080 16658
rect 39028 16594 39080 16600
rect 38936 16584 38988 16590
rect 39120 16584 39172 16590
rect 38936 16526 38988 16532
rect 39118 16552 39120 16561
rect 39172 16552 39174 16561
rect 38844 16516 38896 16522
rect 39118 16487 39174 16496
rect 38844 16458 38896 16464
rect 38856 16266 38884 16458
rect 38856 16238 38976 16266
rect 38476 16040 38528 16046
rect 38476 15982 38528 15988
rect 38488 15688 38516 15982
rect 38570 15804 38878 15813
rect 38570 15802 38576 15804
rect 38632 15802 38656 15804
rect 38712 15802 38736 15804
rect 38792 15802 38816 15804
rect 38872 15802 38878 15804
rect 38632 15750 38634 15802
rect 38814 15750 38816 15802
rect 38570 15748 38576 15750
rect 38632 15748 38656 15750
rect 38712 15748 38736 15750
rect 38792 15748 38816 15750
rect 38872 15748 38878 15750
rect 38570 15739 38878 15748
rect 38488 15660 38608 15688
rect 38580 15586 38608 15660
rect 38948 15638 38976 16238
rect 38936 15632 38988 15638
rect 38580 15558 38700 15586
rect 38936 15574 38988 15580
rect 38672 15484 38700 15558
rect 39132 15502 39160 16487
rect 39224 16182 39252 16662
rect 39212 16176 39264 16182
rect 39212 16118 39264 16124
rect 38752 15496 38804 15502
rect 38672 15456 38752 15484
rect 38672 15162 38700 15456
rect 38752 15438 38804 15444
rect 39120 15496 39172 15502
rect 39120 15438 39172 15444
rect 39120 15360 39172 15366
rect 39120 15302 39172 15308
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38672 14822 38700 15098
rect 39028 14952 39080 14958
rect 39028 14894 39080 14900
rect 38660 14816 38712 14822
rect 38488 14776 38660 14804
rect 38488 14414 38516 14776
rect 38660 14758 38712 14764
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 38570 14716 38878 14725
rect 38570 14714 38576 14716
rect 38632 14714 38656 14716
rect 38712 14714 38736 14716
rect 38792 14714 38816 14716
rect 38872 14714 38878 14716
rect 38632 14662 38634 14714
rect 38814 14662 38816 14714
rect 38570 14660 38576 14662
rect 38632 14660 38656 14662
rect 38712 14660 38736 14662
rect 38792 14660 38816 14662
rect 38872 14660 38878 14662
rect 38570 14651 38878 14660
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38844 14408 38896 14414
rect 38844 14350 38896 14356
rect 38476 14068 38528 14074
rect 38476 14010 38528 14016
rect 38488 12288 38516 14010
rect 38856 13802 38884 14350
rect 38844 13796 38896 13802
rect 38844 13738 38896 13744
rect 38570 13628 38878 13637
rect 38570 13626 38576 13628
rect 38632 13626 38656 13628
rect 38712 13626 38736 13628
rect 38792 13626 38816 13628
rect 38872 13626 38878 13628
rect 38632 13574 38634 13626
rect 38814 13574 38816 13626
rect 38570 13572 38576 13574
rect 38632 13572 38656 13574
rect 38712 13572 38736 13574
rect 38792 13572 38816 13574
rect 38872 13572 38878 13574
rect 38570 13563 38878 13572
rect 38844 13184 38896 13190
rect 38844 13126 38896 13132
rect 38856 12730 38884 13126
rect 38948 12986 38976 14758
rect 39040 14482 39068 14894
rect 39028 14476 39080 14482
rect 39028 14418 39080 14424
rect 39040 13462 39068 14418
rect 39132 14278 39160 15302
rect 39408 15094 39436 17478
rect 39500 16522 39528 17682
rect 40052 17626 40080 17711
rect 40604 17678 40632 18022
rect 40592 17672 40644 17678
rect 40052 17610 40172 17626
rect 40592 17614 40644 17620
rect 40052 17604 40184 17610
rect 40052 17598 40132 17604
rect 40184 17564 40356 17592
rect 40132 17546 40184 17552
rect 40040 17536 40092 17542
rect 40040 17478 40092 17484
rect 40052 17270 40080 17478
rect 40040 17264 40092 17270
rect 40040 17206 40092 17212
rect 39580 17196 39632 17202
rect 39580 17138 39632 17144
rect 40132 17196 40184 17202
rect 40132 17138 40184 17144
rect 39592 16998 39620 17138
rect 39764 17060 39816 17066
rect 39764 17002 39816 17008
rect 39580 16992 39632 16998
rect 39580 16934 39632 16940
rect 39488 16516 39540 16522
rect 39488 16458 39540 16464
rect 39500 16046 39528 16458
rect 39488 16040 39540 16046
rect 39488 15982 39540 15988
rect 39776 15910 39804 17002
rect 39856 16992 39908 16998
rect 39856 16934 39908 16940
rect 39868 16266 39896 16934
rect 39948 16788 40000 16794
rect 39948 16730 40000 16736
rect 39960 16522 39988 16730
rect 39948 16516 40000 16522
rect 40000 16476 40080 16504
rect 39948 16458 40000 16464
rect 39868 16238 39988 16266
rect 39764 15904 39816 15910
rect 39764 15846 39816 15852
rect 39960 15552 39988 16238
rect 39868 15524 39988 15552
rect 39868 15366 39896 15524
rect 40052 15434 40080 16476
rect 40144 16250 40172 17138
rect 40132 16244 40184 16250
rect 40132 16186 40184 16192
rect 40040 15428 40092 15434
rect 40040 15370 40092 15376
rect 39856 15360 39908 15366
rect 39856 15302 39908 15308
rect 39396 15088 39448 15094
rect 40052 15076 40080 15370
rect 40224 15088 40276 15094
rect 40052 15048 40224 15076
rect 39396 15030 39448 15036
rect 40224 15030 40276 15036
rect 39212 15020 39264 15026
rect 39212 14962 39264 14968
rect 39672 15020 39724 15026
rect 39672 14962 39724 14968
rect 39224 14822 39252 14962
rect 39212 14816 39264 14822
rect 39212 14758 39264 14764
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39028 13456 39080 13462
rect 39028 13398 39080 13404
rect 39028 13320 39080 13326
rect 39028 13262 39080 13268
rect 38936 12980 38988 12986
rect 38936 12922 38988 12928
rect 38856 12702 38976 12730
rect 38570 12540 38878 12549
rect 38570 12538 38576 12540
rect 38632 12538 38656 12540
rect 38712 12538 38736 12540
rect 38792 12538 38816 12540
rect 38872 12538 38878 12540
rect 38632 12486 38634 12538
rect 38814 12486 38816 12538
rect 38570 12484 38576 12486
rect 38632 12484 38656 12486
rect 38712 12484 38736 12486
rect 38792 12484 38816 12486
rect 38872 12484 38878 12486
rect 38570 12475 38878 12484
rect 38948 12434 38976 12702
rect 39040 12646 39068 13262
rect 39028 12640 39080 12646
rect 39028 12582 39080 12588
rect 38948 12406 39068 12434
rect 38752 12368 38804 12374
rect 38752 12310 38804 12316
rect 38568 12300 38620 12306
rect 38488 12260 38568 12288
rect 38568 12242 38620 12248
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38488 11014 38516 11630
rect 38764 11558 38792 12310
rect 38752 11552 38804 11558
rect 38752 11494 38804 11500
rect 38936 11552 38988 11558
rect 38936 11494 38988 11500
rect 38570 11452 38878 11461
rect 38570 11450 38576 11452
rect 38632 11450 38656 11452
rect 38712 11450 38736 11452
rect 38792 11450 38816 11452
rect 38872 11450 38878 11452
rect 38632 11398 38634 11450
rect 38814 11398 38816 11450
rect 38570 11396 38576 11398
rect 38632 11396 38656 11398
rect 38712 11396 38736 11398
rect 38792 11396 38816 11398
rect 38872 11396 38878 11398
rect 38570 11387 38878 11396
rect 38844 11348 38896 11354
rect 38844 11290 38896 11296
rect 38856 11218 38884 11290
rect 38844 11212 38896 11218
rect 38844 11154 38896 11160
rect 38660 11144 38712 11150
rect 38948 11098 38976 11494
rect 39040 11218 39068 12406
rect 39132 12238 39160 14214
rect 39224 13870 39252 14758
rect 39488 14340 39540 14346
rect 39488 14282 39540 14288
rect 39500 14074 39528 14282
rect 39488 14068 39540 14074
rect 39488 14010 39540 14016
rect 39684 13870 39712 14962
rect 40132 14612 40184 14618
rect 40132 14554 40184 14560
rect 39856 14476 39908 14482
rect 39856 14418 39908 14424
rect 40040 14476 40092 14482
rect 40040 14418 40092 14424
rect 39764 14272 39816 14278
rect 39764 14214 39816 14220
rect 39212 13864 39264 13870
rect 39580 13864 39632 13870
rect 39264 13812 39436 13818
rect 39212 13806 39436 13812
rect 39580 13806 39632 13812
rect 39672 13864 39724 13870
rect 39672 13806 39724 13812
rect 39224 13790 39436 13806
rect 39212 13728 39264 13734
rect 39212 13670 39264 13676
rect 39304 13728 39356 13734
rect 39304 13670 39356 13676
rect 39224 13190 39252 13670
rect 39316 13530 39344 13670
rect 39304 13524 39356 13530
rect 39304 13466 39356 13472
rect 39212 13184 39264 13190
rect 39212 13126 39264 13132
rect 39224 12714 39252 13126
rect 39212 12708 39264 12714
rect 39212 12650 39264 12656
rect 39304 12300 39356 12306
rect 39304 12242 39356 12248
rect 39120 12232 39172 12238
rect 39120 12174 39172 12180
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 39028 11212 39080 11218
rect 39028 11154 39080 11160
rect 38712 11092 38976 11098
rect 38660 11086 38976 11092
rect 38568 11076 38620 11082
rect 38672 11070 38976 11086
rect 39028 11076 39080 11082
rect 38568 11018 38620 11024
rect 39028 11018 39080 11024
rect 38476 11008 38528 11014
rect 38476 10950 38528 10956
rect 38580 10962 38608 11018
rect 38580 10934 38700 10962
rect 38672 10792 38700 10934
rect 38752 10804 38804 10810
rect 38672 10764 38752 10792
rect 38752 10746 38804 10752
rect 38570 10364 38878 10373
rect 38570 10362 38576 10364
rect 38632 10362 38656 10364
rect 38712 10362 38736 10364
rect 38792 10362 38816 10364
rect 38872 10362 38878 10364
rect 38632 10310 38634 10362
rect 38814 10310 38816 10362
rect 38570 10308 38576 10310
rect 38632 10308 38656 10310
rect 38712 10308 38736 10310
rect 38792 10308 38816 10310
rect 38872 10308 38878 10310
rect 38570 10299 38878 10308
rect 38384 10260 38436 10266
rect 38384 10202 38436 10208
rect 39040 10198 39068 11018
rect 39028 10192 39080 10198
rect 39028 10134 39080 10140
rect 39132 10062 39160 12038
rect 39212 11824 39264 11830
rect 39212 11766 39264 11772
rect 39224 10674 39252 11766
rect 39316 11354 39344 12242
rect 39304 11348 39356 11354
rect 39304 11290 39356 11296
rect 39212 10668 39264 10674
rect 39212 10610 39264 10616
rect 39316 10130 39344 11290
rect 39408 10130 39436 13790
rect 39488 13252 39540 13258
rect 39488 13194 39540 13200
rect 39500 12986 39528 13194
rect 39488 12980 39540 12986
rect 39488 12922 39540 12928
rect 39592 12782 39620 13806
rect 39684 12918 39712 13806
rect 39776 13258 39804 14214
rect 39764 13252 39816 13258
rect 39764 13194 39816 13200
rect 39776 12918 39804 13194
rect 39868 12918 39896 14418
rect 39672 12912 39724 12918
rect 39672 12854 39724 12860
rect 39764 12912 39816 12918
rect 39764 12854 39816 12860
rect 39856 12912 39908 12918
rect 39856 12854 39908 12860
rect 40052 12850 40080 14418
rect 40144 12986 40172 14554
rect 40236 14346 40264 15030
rect 40224 14340 40276 14346
rect 40224 14282 40276 14288
rect 40236 14006 40264 14282
rect 40224 14000 40276 14006
rect 40224 13942 40276 13948
rect 40236 13530 40264 13942
rect 40224 13524 40276 13530
rect 40224 13466 40276 13472
rect 40236 13258 40264 13466
rect 40224 13252 40276 13258
rect 40224 13194 40276 13200
rect 40132 12980 40184 12986
rect 40132 12922 40184 12928
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 39580 12776 39632 12782
rect 39580 12718 39632 12724
rect 40328 12434 40356 17564
rect 40972 17320 41000 18294
rect 41708 18290 41736 18566
rect 41696 18284 41748 18290
rect 41696 18226 41748 18232
rect 41708 18170 41736 18226
rect 41432 18142 41736 18170
rect 41432 17898 41460 18142
rect 41512 18080 41564 18086
rect 41512 18022 41564 18028
rect 41340 17870 41460 17898
rect 41340 17746 41368 17870
rect 41328 17740 41380 17746
rect 41328 17682 41380 17688
rect 41420 17604 41472 17610
rect 41420 17546 41472 17552
rect 41070 17436 41378 17445
rect 41070 17434 41076 17436
rect 41132 17434 41156 17436
rect 41212 17434 41236 17436
rect 41292 17434 41316 17436
rect 41372 17434 41378 17436
rect 41132 17382 41134 17434
rect 41314 17382 41316 17434
rect 41070 17380 41076 17382
rect 41132 17380 41156 17382
rect 41212 17380 41236 17382
rect 41292 17380 41316 17382
rect 41372 17380 41378 17382
rect 41070 17371 41378 17380
rect 40972 17292 41092 17320
rect 40960 17196 41012 17202
rect 40960 17138 41012 17144
rect 40592 16992 40644 16998
rect 40592 16934 40644 16940
rect 40604 16794 40632 16934
rect 40972 16794 41000 17138
rect 41064 17134 41092 17292
rect 41052 17128 41104 17134
rect 41052 17070 41104 17076
rect 40592 16788 40644 16794
rect 40592 16730 40644 16736
rect 40960 16788 41012 16794
rect 40960 16730 41012 16736
rect 40960 16584 41012 16590
rect 40958 16552 40960 16561
rect 41012 16552 41014 16561
rect 41432 16538 41460 17546
rect 41524 17338 41552 18022
rect 41512 17332 41564 17338
rect 41512 17274 41564 17280
rect 41604 17196 41656 17202
rect 41604 17138 41656 17144
rect 41512 17128 41564 17134
rect 41512 17070 41564 17076
rect 41340 16522 41460 16538
rect 40958 16487 41014 16496
rect 41328 16516 41460 16522
rect 41380 16510 41460 16516
rect 41328 16458 41380 16464
rect 40776 16448 40828 16454
rect 41524 16402 41552 17070
rect 41616 16454 41644 17138
rect 41892 17134 41920 18822
rect 42076 18222 42104 19790
rect 42156 19712 42208 19718
rect 42156 19654 42208 19660
rect 42168 19514 42196 19654
rect 42156 19508 42208 19514
rect 42156 19450 42208 19456
rect 42168 18834 42196 19450
rect 42352 19310 42380 20334
rect 42616 20256 42668 20262
rect 42616 20198 42668 20204
rect 42628 19922 42656 20198
rect 42616 19916 42668 19922
rect 42616 19858 42668 19864
rect 42720 19446 42748 22374
rect 43168 22092 43220 22098
rect 43168 22034 43220 22040
rect 42800 21888 42852 21894
rect 42800 21830 42852 21836
rect 42812 21690 42840 21830
rect 42800 21684 42852 21690
rect 42800 21626 42852 21632
rect 42812 21146 42840 21626
rect 42800 21140 42852 21146
rect 42800 21082 42852 21088
rect 42812 19786 42840 21082
rect 43180 20874 43208 22034
rect 43168 20868 43220 20874
rect 43168 20810 43220 20816
rect 42800 19780 42852 19786
rect 42800 19722 42852 19728
rect 42708 19440 42760 19446
rect 42708 19382 42760 19388
rect 42340 19304 42392 19310
rect 42340 19246 42392 19252
rect 42812 19242 42840 19722
rect 43180 19310 43208 20810
rect 43168 19304 43220 19310
rect 43088 19264 43168 19292
rect 42800 19236 42852 19242
rect 42800 19178 42852 19184
rect 42156 18828 42208 18834
rect 42156 18770 42208 18776
rect 42248 18624 42300 18630
rect 42248 18566 42300 18572
rect 42708 18624 42760 18630
rect 42708 18566 42760 18572
rect 42064 18216 42116 18222
rect 42064 18158 42116 18164
rect 42260 18086 42288 18566
rect 42720 18426 42748 18566
rect 42708 18420 42760 18426
rect 42708 18362 42760 18368
rect 42812 18358 42840 19178
rect 42984 18692 43036 18698
rect 42984 18634 43036 18640
rect 42996 18426 43024 18634
rect 42984 18420 43036 18426
rect 42984 18362 43036 18368
rect 42800 18352 42852 18358
rect 42800 18294 42852 18300
rect 42812 18222 42840 18294
rect 42800 18216 42852 18222
rect 42800 18158 42852 18164
rect 42248 18080 42300 18086
rect 42248 18022 42300 18028
rect 42260 17882 42288 18022
rect 42248 17876 42300 17882
rect 42248 17818 42300 17824
rect 42432 17604 42484 17610
rect 42432 17546 42484 17552
rect 42444 17270 42472 17546
rect 42812 17338 42840 18158
rect 42996 17746 43024 18362
rect 43088 17746 43116 19264
rect 43168 19246 43220 19252
rect 42984 17740 43036 17746
rect 42984 17682 43036 17688
rect 43076 17740 43128 17746
rect 43076 17682 43128 17688
rect 42800 17332 42852 17338
rect 42800 17274 42852 17280
rect 42432 17264 42484 17270
rect 42432 17206 42484 17212
rect 41880 17128 41932 17134
rect 41880 17070 41932 17076
rect 41788 16992 41840 16998
rect 41788 16934 41840 16940
rect 41800 16574 41828 16934
rect 41708 16546 41828 16574
rect 40776 16390 40828 16396
rect 40684 16244 40736 16250
rect 40684 16186 40736 16192
rect 40500 15904 40552 15910
rect 40500 15846 40552 15852
rect 40512 15706 40540 15846
rect 40696 15706 40724 16186
rect 40788 16114 40816 16390
rect 41432 16374 41552 16402
rect 41604 16448 41656 16454
rect 41604 16390 41656 16396
rect 41070 16348 41378 16357
rect 41070 16346 41076 16348
rect 41132 16346 41156 16348
rect 41212 16346 41236 16348
rect 41292 16346 41316 16348
rect 41372 16346 41378 16348
rect 41132 16294 41134 16346
rect 41314 16294 41316 16346
rect 41070 16292 41076 16294
rect 41132 16292 41156 16294
rect 41212 16292 41236 16294
rect 41292 16292 41316 16294
rect 41372 16292 41378 16294
rect 41070 16283 41378 16292
rect 40776 16108 40828 16114
rect 40776 16050 40828 16056
rect 40500 15700 40552 15706
rect 40500 15642 40552 15648
rect 40684 15700 40736 15706
rect 40684 15642 40736 15648
rect 40788 15638 40816 16050
rect 40776 15632 40828 15638
rect 40776 15574 40828 15580
rect 41432 15570 41460 16374
rect 41616 16266 41644 16390
rect 41524 16238 41644 16266
rect 41524 15994 41552 16238
rect 41604 16108 41656 16114
rect 41708 16096 41736 16546
rect 41656 16068 41736 16096
rect 41604 16050 41656 16056
rect 41788 16040 41840 16046
rect 41524 15966 41736 15994
rect 41788 15982 41840 15988
rect 41420 15564 41472 15570
rect 41420 15506 41472 15512
rect 41708 15502 41736 15966
rect 41696 15496 41748 15502
rect 41696 15438 41748 15444
rect 41052 15360 41104 15366
rect 40972 15320 41052 15348
rect 40972 15162 41000 15320
rect 41052 15302 41104 15308
rect 41512 15360 41564 15366
rect 41512 15302 41564 15308
rect 41604 15360 41656 15366
rect 41604 15302 41656 15308
rect 41070 15260 41378 15269
rect 41070 15258 41076 15260
rect 41132 15258 41156 15260
rect 41212 15258 41236 15260
rect 41292 15258 41316 15260
rect 41372 15258 41378 15260
rect 41132 15206 41134 15258
rect 41314 15206 41316 15258
rect 41070 15204 41076 15206
rect 41132 15204 41156 15206
rect 41212 15204 41236 15206
rect 41292 15204 41316 15206
rect 41372 15204 41378 15206
rect 41070 15195 41378 15204
rect 40960 15156 41012 15162
rect 40960 15098 41012 15104
rect 41236 14884 41288 14890
rect 41236 14826 41288 14832
rect 40776 14816 40828 14822
rect 41144 14816 41196 14822
rect 40828 14776 41144 14804
rect 40776 14758 40828 14764
rect 41144 14758 41196 14764
rect 40960 14476 41012 14482
rect 40960 14418 41012 14424
rect 40868 14272 40920 14278
rect 40868 14214 40920 14220
rect 40880 13818 40908 14214
rect 40972 13938 41000 14418
rect 41248 14278 41276 14826
rect 41524 14822 41552 15302
rect 41616 15094 41644 15302
rect 41604 15088 41656 15094
rect 41604 15030 41656 15036
rect 41800 14958 41828 15982
rect 41788 14952 41840 14958
rect 41788 14894 41840 14900
rect 41420 14816 41472 14822
rect 41420 14758 41472 14764
rect 41512 14816 41564 14822
rect 41512 14758 41564 14764
rect 41432 14550 41460 14758
rect 41420 14544 41472 14550
rect 41420 14486 41472 14492
rect 41236 14272 41288 14278
rect 41236 14214 41288 14220
rect 41070 14172 41378 14181
rect 41070 14170 41076 14172
rect 41132 14170 41156 14172
rect 41212 14170 41236 14172
rect 41292 14170 41316 14172
rect 41372 14170 41378 14172
rect 41132 14118 41134 14170
rect 41314 14118 41316 14170
rect 41070 14116 41076 14118
rect 41132 14116 41156 14118
rect 41212 14116 41236 14118
rect 41292 14116 41316 14118
rect 41372 14116 41378 14118
rect 41070 14107 41378 14116
rect 40960 13932 41012 13938
rect 40960 13874 41012 13880
rect 40880 13790 41000 13818
rect 40972 13462 41000 13790
rect 41432 13546 41460 14486
rect 41524 14278 41552 14758
rect 41892 14482 41920 17070
rect 42248 15632 42300 15638
rect 42248 15574 42300 15580
rect 42064 15564 42116 15570
rect 42064 15506 42116 15512
rect 41880 14476 41932 14482
rect 41708 14436 41880 14464
rect 41512 14272 41564 14278
rect 41512 14214 41564 14220
rect 41340 13530 41460 13546
rect 41328 13524 41460 13530
rect 41380 13518 41460 13524
rect 41328 13466 41380 13472
rect 40960 13456 41012 13462
rect 40960 13398 41012 13404
rect 40776 13388 40828 13394
rect 40776 13330 40828 13336
rect 40500 12640 40552 12646
rect 40500 12582 40552 12588
rect 40236 12406 40356 12434
rect 39948 12096 40000 12102
rect 39948 12038 40000 12044
rect 39764 11688 39816 11694
rect 39764 11630 39816 11636
rect 39672 11008 39724 11014
rect 39672 10950 39724 10956
rect 39684 10606 39712 10950
rect 39776 10810 39804 11630
rect 39960 11354 39988 12038
rect 39948 11348 40000 11354
rect 39948 11290 40000 11296
rect 39948 11076 40000 11082
rect 39948 11018 40000 11024
rect 39764 10804 39816 10810
rect 39764 10746 39816 10752
rect 39960 10742 39988 11018
rect 39948 10736 40000 10742
rect 39948 10678 40000 10684
rect 39672 10600 39724 10606
rect 39672 10542 39724 10548
rect 39948 10600 40000 10606
rect 39948 10542 40000 10548
rect 39304 10124 39356 10130
rect 39304 10066 39356 10072
rect 39396 10124 39448 10130
rect 39396 10066 39448 10072
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 39120 10056 39172 10062
rect 39120 9998 39172 10004
rect 38672 9722 38700 9998
rect 39684 9926 39712 10542
rect 39960 10266 39988 10542
rect 39948 10260 40000 10266
rect 39948 10202 40000 10208
rect 39672 9920 39724 9926
rect 39672 9862 39724 9868
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 38476 9444 38528 9450
rect 38476 9386 38528 9392
rect 38292 8968 38344 8974
rect 38292 8910 38344 8916
rect 38200 8424 38252 8430
rect 38200 8366 38252 8372
rect 38212 7750 38240 8366
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38304 7546 38332 8910
rect 38384 8288 38436 8294
rect 38384 8230 38436 8236
rect 38396 7886 38424 8230
rect 38488 8090 38516 9386
rect 38570 9276 38878 9285
rect 38570 9274 38576 9276
rect 38632 9274 38656 9276
rect 38712 9274 38736 9276
rect 38792 9274 38816 9276
rect 38872 9274 38878 9276
rect 38632 9222 38634 9274
rect 38814 9222 38816 9274
rect 38570 9220 38576 9222
rect 38632 9220 38656 9222
rect 38712 9220 38736 9222
rect 38792 9220 38816 9222
rect 38872 9220 38878 9222
rect 38570 9211 38878 9220
rect 39684 8974 39712 9862
rect 40132 9512 40184 9518
rect 40132 9454 40184 9460
rect 39764 9376 39816 9382
rect 39764 9318 39816 9324
rect 39776 9178 39804 9318
rect 39764 9172 39816 9178
rect 39764 9114 39816 9120
rect 39672 8968 39724 8974
rect 39672 8910 39724 8916
rect 39764 8968 39816 8974
rect 39764 8910 39816 8916
rect 38844 8832 38896 8838
rect 38844 8774 38896 8780
rect 38752 8628 38804 8634
rect 38752 8570 38804 8576
rect 38764 8537 38792 8570
rect 38750 8528 38806 8537
rect 38750 8463 38806 8472
rect 38856 8294 38884 8774
rect 38844 8288 38896 8294
rect 38844 8230 38896 8236
rect 38570 8188 38878 8197
rect 38570 8186 38576 8188
rect 38632 8186 38656 8188
rect 38712 8186 38736 8188
rect 38792 8186 38816 8188
rect 38872 8186 38878 8188
rect 38632 8134 38634 8186
rect 38814 8134 38816 8186
rect 38570 8132 38576 8134
rect 38632 8132 38656 8134
rect 38712 8132 38736 8134
rect 38792 8132 38816 8134
rect 38872 8132 38878 8134
rect 38570 8123 38878 8132
rect 38476 8084 38528 8090
rect 38476 8026 38528 8032
rect 39684 7886 39712 8910
rect 39776 8362 39804 8910
rect 40040 8560 40092 8566
rect 40038 8528 40040 8537
rect 40092 8528 40094 8537
rect 40038 8463 40094 8472
rect 40144 8430 40172 9454
rect 40236 8566 40264 12406
rect 40512 12102 40540 12582
rect 40500 12096 40552 12102
rect 40500 12038 40552 12044
rect 40788 11898 40816 13330
rect 40972 12782 41000 13398
rect 41070 13084 41378 13093
rect 41070 13082 41076 13084
rect 41132 13082 41156 13084
rect 41212 13082 41236 13084
rect 41292 13082 41316 13084
rect 41372 13082 41378 13084
rect 41132 13030 41134 13082
rect 41314 13030 41316 13082
rect 41070 13028 41076 13030
rect 41132 13028 41156 13030
rect 41212 13028 41236 13030
rect 41292 13028 41316 13030
rect 41372 13028 41378 13030
rect 41070 13019 41378 13028
rect 40960 12776 41012 12782
rect 40960 12718 41012 12724
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 40776 11892 40828 11898
rect 40776 11834 40828 11840
rect 40408 11688 40460 11694
rect 40408 11630 40460 11636
rect 40420 11098 40448 11630
rect 40972 11558 41000 12038
rect 41070 11996 41378 12005
rect 41070 11994 41076 11996
rect 41132 11994 41156 11996
rect 41212 11994 41236 11996
rect 41292 11994 41316 11996
rect 41372 11994 41378 11996
rect 41132 11942 41134 11994
rect 41314 11942 41316 11994
rect 41070 11940 41076 11942
rect 41132 11940 41156 11942
rect 41212 11940 41236 11942
rect 41292 11940 41316 11942
rect 41372 11940 41378 11942
rect 41070 11931 41378 11940
rect 41432 11762 41460 12174
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 40960 11552 41012 11558
rect 40960 11494 41012 11500
rect 40328 11070 40448 11098
rect 40776 11076 40828 11082
rect 40328 11014 40356 11070
rect 40776 11018 40828 11024
rect 40316 11008 40368 11014
rect 40316 10950 40368 10956
rect 40328 10062 40356 10950
rect 40316 10056 40368 10062
rect 40316 9998 40368 10004
rect 40408 10056 40460 10062
rect 40408 9998 40460 10004
rect 40420 9926 40448 9998
rect 40788 9994 40816 11018
rect 40776 9988 40828 9994
rect 40776 9930 40828 9936
rect 40972 9926 41000 11494
rect 41070 10908 41378 10917
rect 41070 10906 41076 10908
rect 41132 10906 41156 10908
rect 41212 10906 41236 10908
rect 41292 10906 41316 10908
rect 41372 10906 41378 10908
rect 41132 10854 41134 10906
rect 41314 10854 41316 10906
rect 41070 10852 41076 10854
rect 41132 10852 41156 10854
rect 41212 10852 41236 10854
rect 41292 10852 41316 10854
rect 41372 10852 41378 10854
rect 41070 10843 41378 10852
rect 41432 10810 41460 11698
rect 41524 11150 41552 14214
rect 41604 12300 41656 12306
rect 41604 12242 41656 12248
rect 41616 11898 41644 12242
rect 41604 11892 41656 11898
rect 41604 11834 41656 11840
rect 41604 11688 41656 11694
rect 41604 11630 41656 11636
rect 41616 11218 41644 11630
rect 41604 11212 41656 11218
rect 41604 11154 41656 11160
rect 41512 11144 41564 11150
rect 41512 11086 41564 11092
rect 41420 10804 41472 10810
rect 41420 10746 41472 10752
rect 40408 9920 40460 9926
rect 40408 9862 40460 9868
rect 40960 9920 41012 9926
rect 40960 9862 41012 9868
rect 40420 9722 40448 9862
rect 41070 9820 41378 9829
rect 41070 9818 41076 9820
rect 41132 9818 41156 9820
rect 41212 9818 41236 9820
rect 41292 9818 41316 9820
rect 41372 9818 41378 9820
rect 41132 9766 41134 9818
rect 41314 9766 41316 9818
rect 41070 9764 41076 9766
rect 41132 9764 41156 9766
rect 41212 9764 41236 9766
rect 41292 9764 41316 9766
rect 41372 9764 41378 9766
rect 41070 9755 41378 9764
rect 40408 9716 40460 9722
rect 40408 9658 40460 9664
rect 41512 9648 41564 9654
rect 41512 9590 41564 9596
rect 40868 9580 40920 9586
rect 40868 9522 40920 9528
rect 40592 9036 40644 9042
rect 40592 8978 40644 8984
rect 40224 8560 40276 8566
rect 40224 8502 40276 8508
rect 40604 8498 40632 8978
rect 40592 8492 40644 8498
rect 40592 8434 40644 8440
rect 40776 8492 40828 8498
rect 40776 8434 40828 8440
rect 40132 8424 40184 8430
rect 40132 8366 40184 8372
rect 39764 8356 39816 8362
rect 39764 8298 39816 8304
rect 38384 7880 38436 7886
rect 38384 7822 38436 7828
rect 39580 7880 39632 7886
rect 39580 7822 39632 7828
rect 39672 7880 39724 7886
rect 39672 7822 39724 7828
rect 39212 7812 39264 7818
rect 39212 7754 39264 7760
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 39120 7404 39172 7410
rect 39120 7346 39172 7352
rect 38200 7200 38252 7206
rect 38200 7142 38252 7148
rect 37740 6870 37792 6876
rect 38106 6896 38162 6905
rect 36912 6860 37320 6866
rect 36964 6854 37320 6860
rect 37924 6860 37976 6866
rect 36912 6802 36964 6808
rect 36728 6792 36780 6798
rect 36726 6760 36728 6769
rect 36780 6760 36782 6769
rect 36726 6695 36782 6704
rect 36820 6656 36872 6662
rect 36648 6616 36768 6644
rect 36452 6598 36504 6604
rect 36070 6556 36378 6565
rect 36070 6554 36076 6556
rect 36132 6554 36156 6556
rect 36212 6554 36236 6556
rect 36292 6554 36316 6556
rect 36372 6554 36378 6556
rect 36132 6502 36134 6554
rect 36314 6502 36316 6554
rect 36070 6500 36076 6502
rect 36132 6500 36156 6502
rect 36212 6500 36236 6502
rect 36292 6500 36316 6502
rect 36372 6500 36378 6502
rect 36070 6491 36378 6500
rect 36464 6458 36492 6598
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 36004 6186 36032 6258
rect 35992 6180 36044 6186
rect 35992 6122 36044 6128
rect 36004 4758 36032 6122
rect 36176 6112 36228 6118
rect 36176 6054 36228 6060
rect 36188 5778 36216 6054
rect 36176 5772 36228 5778
rect 36176 5714 36228 5720
rect 36636 5704 36688 5710
rect 36636 5646 36688 5652
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36070 5468 36378 5477
rect 36070 5466 36076 5468
rect 36132 5466 36156 5468
rect 36212 5466 36236 5468
rect 36292 5466 36316 5468
rect 36372 5466 36378 5468
rect 36132 5414 36134 5466
rect 36314 5414 36316 5466
rect 36070 5412 36076 5414
rect 36132 5412 36156 5414
rect 36212 5412 36236 5414
rect 36292 5412 36316 5414
rect 36372 5412 36378 5414
rect 36070 5403 36378 5412
rect 36360 5364 36412 5370
rect 36360 5306 36412 5312
rect 36084 5228 36136 5234
rect 36084 5170 36136 5176
rect 35992 4752 36044 4758
rect 35992 4694 36044 4700
rect 36096 4622 36124 5170
rect 36372 4690 36400 5306
rect 36464 5030 36492 5510
rect 36648 5234 36676 5646
rect 36636 5228 36688 5234
rect 36636 5170 36688 5176
rect 36740 5166 36768 6616
rect 36820 6598 36872 6604
rect 36832 5914 36860 6598
rect 36912 6452 36964 6458
rect 36912 6394 36964 6400
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36832 5778 36860 5850
rect 36820 5772 36872 5778
rect 36820 5714 36872 5720
rect 36924 5710 36952 6394
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 37016 6225 37044 6258
rect 37096 6248 37148 6254
rect 37002 6216 37058 6225
rect 37096 6190 37148 6196
rect 37002 6151 37058 6160
rect 37108 5914 37136 6190
rect 37096 5908 37148 5914
rect 37096 5850 37148 5856
rect 37200 5794 37228 6854
rect 38106 6831 38162 6840
rect 37924 6802 37976 6808
rect 37280 6656 37332 6662
rect 37280 6598 37332 6604
rect 37292 6390 37320 6598
rect 37280 6384 37332 6390
rect 37280 6326 37332 6332
rect 37280 5908 37332 5914
rect 37280 5850 37332 5856
rect 37016 5766 37228 5794
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 36820 5636 36872 5642
rect 36820 5578 36872 5584
rect 36832 5370 36860 5578
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 36728 5160 36780 5166
rect 36728 5102 36780 5108
rect 36452 5024 36504 5030
rect 36452 4966 36504 4972
rect 36452 4752 36504 4758
rect 36452 4694 36504 4700
rect 36360 4684 36412 4690
rect 36360 4626 36412 4632
rect 36084 4616 36136 4622
rect 36004 4576 36084 4604
rect 36004 4214 36032 4576
rect 36084 4558 36136 4564
rect 36070 4380 36378 4389
rect 36070 4378 36076 4380
rect 36132 4378 36156 4380
rect 36212 4378 36236 4380
rect 36292 4378 36316 4380
rect 36372 4378 36378 4380
rect 36132 4326 36134 4378
rect 36314 4326 36316 4378
rect 36070 4324 36076 4326
rect 36132 4324 36156 4326
rect 36212 4324 36236 4326
rect 36292 4324 36316 4326
rect 36372 4324 36378 4326
rect 36070 4315 36378 4324
rect 35992 4208 36044 4214
rect 35992 4150 36044 4156
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 36464 4078 36492 4694
rect 37016 4690 37044 5766
rect 37188 5704 37240 5710
rect 37188 5646 37240 5652
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 37108 5234 37136 5510
rect 37096 5228 37148 5234
rect 37096 5170 37148 5176
rect 36544 4684 36596 4690
rect 36544 4626 36596 4632
rect 37004 4684 37056 4690
rect 37004 4626 37056 4632
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35912 3738 35940 3878
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 36556 3602 36584 4626
rect 36912 4616 36964 4622
rect 36912 4558 36964 4564
rect 36818 4040 36874 4049
rect 36818 3975 36820 3984
rect 36872 3975 36874 3984
rect 36820 3946 36872 3952
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35820 3194 35848 3470
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 35912 2990 35940 3470
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 3194 36032 3334
rect 36070 3292 36378 3301
rect 36070 3290 36076 3292
rect 36132 3290 36156 3292
rect 36212 3290 36236 3292
rect 36292 3290 36316 3292
rect 36372 3290 36378 3292
rect 36132 3238 36134 3290
rect 36314 3238 36316 3290
rect 36070 3236 36076 3238
rect 36132 3236 36156 3238
rect 36212 3236 36236 3238
rect 36292 3236 36316 3238
rect 36372 3236 36378 3238
rect 36070 3227 36378 3236
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 36360 2984 36412 2990
rect 36412 2944 36492 2972
rect 36360 2926 36412 2932
rect 35808 2848 35860 2854
rect 35992 2848 36044 2854
rect 35808 2790 35860 2796
rect 35898 2816 35954 2825
rect 35714 2680 35770 2689
rect 35714 2615 35770 2624
rect 35728 2310 35756 2615
rect 35820 2514 35848 2790
rect 35992 2790 36044 2796
rect 35898 2751 35954 2760
rect 35912 2650 35940 2751
rect 35900 2644 35952 2650
rect 35900 2586 35952 2592
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 36004 2394 36032 2790
rect 35820 2366 36032 2394
rect 36464 2378 36492 2944
rect 36452 2372 36504 2378
rect 35716 2304 35768 2310
rect 35716 2246 35768 2252
rect 35636 1958 35756 1986
rect 35624 1896 35676 1902
rect 35624 1838 35676 1844
rect 35256 1488 35308 1494
rect 35256 1430 35308 1436
rect 35636 1426 35664 1838
rect 35624 1420 35676 1426
rect 35624 1362 35676 1368
rect 35728 1358 35756 1958
rect 35164 1352 35216 1358
rect 35164 1294 35216 1300
rect 35716 1352 35768 1358
rect 35716 1294 35768 1300
rect 35624 1216 35676 1222
rect 35624 1158 35676 1164
rect 35636 1018 35664 1158
rect 35624 1012 35676 1018
rect 35624 954 35676 960
rect 35820 160 35848 2366
rect 36452 2314 36504 2320
rect 35900 2304 35952 2310
rect 35900 2246 35952 2252
rect 35912 2106 35940 2246
rect 36070 2204 36378 2213
rect 36070 2202 36076 2204
rect 36132 2202 36156 2204
rect 36212 2202 36236 2204
rect 36292 2202 36316 2204
rect 36372 2202 36378 2204
rect 36132 2150 36134 2202
rect 36314 2150 36316 2202
rect 36070 2148 36076 2150
rect 36132 2148 36156 2150
rect 36212 2148 36236 2150
rect 36292 2148 36316 2150
rect 36372 2148 36378 2150
rect 36070 2139 36378 2148
rect 35900 2100 35952 2106
rect 35900 2042 35952 2048
rect 36464 1970 36492 2314
rect 36452 1964 36504 1970
rect 36452 1906 36504 1912
rect 36464 1494 36492 1906
rect 36556 1902 36584 3538
rect 36728 3392 36780 3398
rect 36728 3334 36780 3340
rect 36820 3392 36872 3398
rect 36820 3334 36872 3340
rect 36740 3097 36768 3334
rect 36832 3194 36860 3334
rect 36820 3188 36872 3194
rect 36820 3130 36872 3136
rect 36726 3088 36782 3097
rect 36726 3023 36782 3032
rect 36924 2514 36952 4558
rect 37016 3534 37044 4626
rect 37200 4622 37228 5646
rect 37292 5574 37320 5850
rect 37936 5778 37964 6802
rect 38016 6724 38068 6730
rect 38120 6712 38148 6831
rect 38068 6684 38148 6712
rect 38016 6666 38068 6672
rect 38106 6352 38162 6361
rect 38106 6287 38162 6296
rect 38120 5914 38148 6287
rect 38108 5908 38160 5914
rect 38108 5850 38160 5856
rect 37924 5772 37976 5778
rect 37924 5714 37976 5720
rect 37280 5568 37332 5574
rect 37280 5510 37332 5516
rect 37292 5234 37320 5510
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 37292 4214 37320 5170
rect 37936 4758 37964 5714
rect 38212 5710 38240 7142
rect 38570 7100 38878 7109
rect 38570 7098 38576 7100
rect 38632 7098 38656 7100
rect 38712 7098 38736 7100
rect 38792 7098 38816 7100
rect 38872 7098 38878 7100
rect 38632 7046 38634 7098
rect 38814 7046 38816 7098
rect 38570 7044 38576 7046
rect 38632 7044 38656 7046
rect 38712 7044 38736 7046
rect 38792 7044 38816 7046
rect 38872 7044 38878 7046
rect 38570 7035 38878 7044
rect 39132 6798 39160 7346
rect 39224 6866 39252 7754
rect 39592 7546 39620 7822
rect 40604 7818 40632 8434
rect 40684 8424 40736 8430
rect 40684 8366 40736 8372
rect 40592 7812 40644 7818
rect 40592 7754 40644 7760
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 40500 7472 40552 7478
rect 40500 7414 40552 7420
rect 39580 7336 39632 7342
rect 39580 7278 39632 7284
rect 39212 6860 39264 6866
rect 39212 6802 39264 6808
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 38844 6656 38896 6662
rect 38844 6598 38896 6604
rect 38856 6458 38884 6598
rect 39132 6458 39160 6734
rect 38844 6452 38896 6458
rect 39120 6452 39172 6458
rect 38896 6412 38976 6440
rect 38844 6394 38896 6400
rect 38476 6316 38528 6322
rect 38476 6258 38528 6264
rect 38660 6316 38712 6322
rect 38660 6258 38712 6264
rect 38488 5914 38516 6258
rect 38672 6186 38700 6258
rect 38660 6180 38712 6186
rect 38660 6122 38712 6128
rect 38570 6012 38878 6021
rect 38570 6010 38576 6012
rect 38632 6010 38656 6012
rect 38712 6010 38736 6012
rect 38792 6010 38816 6012
rect 38872 6010 38878 6012
rect 38632 5958 38634 6010
rect 38814 5958 38816 6010
rect 38570 5956 38576 5958
rect 38632 5956 38656 5958
rect 38712 5956 38736 5958
rect 38792 5956 38816 5958
rect 38872 5956 38878 5958
rect 38570 5947 38878 5956
rect 38476 5908 38528 5914
rect 38476 5850 38528 5856
rect 38200 5704 38252 5710
rect 38200 5646 38252 5652
rect 38948 5574 38976 6412
rect 39120 6394 39172 6400
rect 39224 6390 39252 6802
rect 39212 6384 39264 6390
rect 39212 6326 39264 6332
rect 39224 6202 39252 6326
rect 39132 6174 39252 6202
rect 39028 5908 39080 5914
rect 39028 5850 39080 5856
rect 38476 5568 38528 5574
rect 38476 5510 38528 5516
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 38028 4826 38056 5102
rect 38382 4856 38438 4865
rect 38016 4820 38068 4826
rect 38382 4791 38384 4800
rect 38016 4762 38068 4768
rect 38436 4791 38438 4800
rect 38384 4762 38436 4768
rect 37924 4752 37976 4758
rect 37924 4694 37976 4700
rect 37738 4584 37794 4593
rect 37738 4519 37740 4528
rect 37792 4519 37794 4528
rect 37740 4490 37792 4496
rect 37280 4208 37332 4214
rect 37280 4150 37332 4156
rect 38292 4208 38344 4214
rect 38292 4150 38344 4156
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37004 3528 37056 3534
rect 37004 3470 37056 3476
rect 37188 3460 37240 3466
rect 37188 3402 37240 3408
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 36544 1896 36596 1902
rect 36544 1838 36596 1844
rect 36452 1488 36504 1494
rect 36082 1456 36138 1465
rect 36452 1430 36504 1436
rect 36082 1391 36138 1400
rect 36096 1358 36124 1391
rect 36084 1352 36136 1358
rect 36176 1352 36228 1358
rect 36084 1294 36136 1300
rect 36174 1320 36176 1329
rect 36360 1352 36412 1358
rect 36228 1320 36230 1329
rect 36820 1352 36872 1358
rect 36412 1312 36492 1340
rect 36360 1294 36412 1300
rect 36174 1255 36230 1264
rect 35992 1216 36044 1222
rect 35898 1184 35954 1193
rect 35954 1164 35992 1170
rect 35954 1158 36044 1164
rect 35954 1142 36032 1158
rect 35898 1119 35954 1128
rect 36070 1116 36378 1125
rect 36070 1114 36076 1116
rect 36132 1114 36156 1116
rect 36212 1114 36236 1116
rect 36292 1114 36316 1116
rect 36372 1114 36378 1116
rect 36132 1062 36134 1114
rect 36314 1062 36316 1114
rect 36070 1060 36076 1062
rect 36132 1060 36156 1062
rect 36212 1060 36236 1062
rect 36292 1060 36316 1062
rect 36372 1060 36378 1062
rect 36070 1051 36378 1060
rect 36464 814 36492 1312
rect 36820 1294 36872 1300
rect 36452 808 36504 814
rect 36452 750 36504 756
rect 36832 678 36860 1294
rect 36820 672 36872 678
rect 36820 614 36872 620
rect 36648 190 36768 218
rect 36648 160 36676 190
rect 34256 54 34468 82
rect 34978 -300 35034 160
rect 35806 -300 35862 160
rect 36634 -300 36690 160
rect 36740 82 36768 190
rect 37016 82 37044 3130
rect 37200 2666 37228 3402
rect 37280 3392 37332 3398
rect 37280 3334 37332 3340
rect 37292 2990 37320 3334
rect 37476 3126 37504 4082
rect 37924 3936 37976 3942
rect 37924 3878 37976 3884
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 37936 3641 37964 3878
rect 37922 3632 37978 3641
rect 38212 3602 38240 3878
rect 37922 3567 37978 3576
rect 38200 3596 38252 3602
rect 38200 3538 38252 3544
rect 37648 3392 37700 3398
rect 37648 3334 37700 3340
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38108 3392 38160 3398
rect 38108 3334 38160 3340
rect 37464 3120 37516 3126
rect 37464 3062 37516 3068
rect 37280 2984 37332 2990
rect 37280 2926 37332 2932
rect 37200 2650 37320 2666
rect 37200 2644 37332 2650
rect 37200 2638 37280 2644
rect 37280 2586 37332 2592
rect 37476 2378 37504 3062
rect 37660 2961 37688 3334
rect 38028 3233 38056 3334
rect 38014 3224 38070 3233
rect 38014 3159 38070 3168
rect 37646 2952 37702 2961
rect 37646 2887 37702 2896
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37660 2378 37688 2586
rect 38120 2514 38148 3334
rect 38304 3058 38332 4150
rect 38384 4072 38436 4078
rect 38384 4014 38436 4020
rect 38396 3738 38424 4014
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 38292 2848 38344 2854
rect 38344 2808 38424 2836
rect 38292 2790 38344 2796
rect 38290 2680 38346 2689
rect 38290 2615 38346 2624
rect 38304 2514 38332 2615
rect 38108 2508 38160 2514
rect 38108 2450 38160 2456
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 37464 2372 37516 2378
rect 37464 2314 37516 2320
rect 37648 2372 37700 2378
rect 37648 2314 37700 2320
rect 37476 2038 37504 2314
rect 37832 2304 37884 2310
rect 37832 2246 37884 2252
rect 37464 2032 37516 2038
rect 37464 1974 37516 1980
rect 37096 1352 37148 1358
rect 37096 1294 37148 1300
rect 37108 746 37136 1294
rect 37844 1290 37872 2246
rect 38120 1834 38148 2450
rect 38396 2446 38424 2808
rect 38384 2440 38436 2446
rect 38384 2382 38436 2388
rect 38200 1964 38252 1970
rect 38200 1906 38252 1912
rect 38108 1828 38160 1834
rect 38108 1770 38160 1776
rect 38212 1562 38240 1906
rect 38200 1556 38252 1562
rect 38200 1498 38252 1504
rect 37832 1284 37884 1290
rect 37832 1226 37884 1232
rect 38292 1012 38344 1018
rect 38292 954 38344 960
rect 37096 740 37148 746
rect 37096 682 37148 688
rect 37832 740 37884 746
rect 37832 682 37884 688
rect 36740 54 37044 82
rect 37462 82 37518 160
rect 37844 82 37872 682
rect 38304 160 38332 954
rect 38488 882 38516 5510
rect 39040 5234 39068 5850
rect 39132 5642 39160 6174
rect 39592 6118 39620 7278
rect 39856 7200 39908 7206
rect 39856 7142 39908 7148
rect 39868 7002 39896 7142
rect 40512 7002 40540 7414
rect 40696 7342 40724 8366
rect 40788 7750 40816 8434
rect 40880 7993 40908 9522
rect 41524 8974 41552 9590
rect 41708 9518 41736 14436
rect 41880 14418 41932 14424
rect 41972 13184 42024 13190
rect 41972 13126 42024 13132
rect 41984 12646 42012 13126
rect 41972 12640 42024 12646
rect 41972 12582 42024 12588
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 41800 10606 41828 12038
rect 41972 11280 42024 11286
rect 41972 11222 42024 11228
rect 41880 11008 41932 11014
rect 41880 10950 41932 10956
rect 41788 10600 41840 10606
rect 41788 10542 41840 10548
rect 41788 10464 41840 10470
rect 41788 10406 41840 10412
rect 41800 10266 41828 10406
rect 41892 10266 41920 10950
rect 41984 10674 42012 11222
rect 42076 11218 42104 15506
rect 42260 14074 42288 15574
rect 42248 14068 42300 14074
rect 42248 14010 42300 14016
rect 42260 12374 42288 14010
rect 42444 12986 42472 17206
rect 42800 16992 42852 16998
rect 42800 16934 42852 16940
rect 42812 16574 42840 16934
rect 43088 16794 43116 17682
rect 43272 17678 43300 22374
rect 43570 22332 43878 22341
rect 43570 22330 43576 22332
rect 43632 22330 43656 22332
rect 43712 22330 43736 22332
rect 43792 22330 43816 22332
rect 43872 22330 43878 22332
rect 43632 22278 43634 22330
rect 43814 22278 43816 22330
rect 43570 22276 43576 22278
rect 43632 22276 43656 22278
rect 43712 22276 43736 22278
rect 43792 22276 43816 22278
rect 43872 22276 43878 22278
rect 43570 22267 43878 22276
rect 43916 22030 43944 22374
rect 43904 22024 43956 22030
rect 43904 21966 43956 21972
rect 43916 21622 43944 21966
rect 44192 21690 44220 22374
rect 44180 21684 44232 21690
rect 44180 21626 44232 21632
rect 43904 21616 43956 21622
rect 43904 21558 43956 21564
rect 44272 21344 44324 21350
rect 44272 21286 44324 21292
rect 43570 21244 43878 21253
rect 43570 21242 43576 21244
rect 43632 21242 43656 21244
rect 43712 21242 43736 21244
rect 43792 21242 43816 21244
rect 43872 21242 43878 21244
rect 43632 21190 43634 21242
rect 43814 21190 43816 21242
rect 43570 21188 43576 21190
rect 43632 21188 43656 21190
rect 43712 21188 43736 21190
rect 43792 21188 43816 21190
rect 43872 21188 43878 21190
rect 43570 21179 43878 21188
rect 44180 20868 44232 20874
rect 44180 20810 44232 20816
rect 43444 20800 43496 20806
rect 43444 20742 43496 20748
rect 43456 20534 43484 20742
rect 43444 20528 43496 20534
rect 43444 20470 43496 20476
rect 43456 19446 43484 20470
rect 43810 20360 43866 20369
rect 43810 20295 43812 20304
rect 43864 20295 43866 20304
rect 43812 20266 43864 20272
rect 44192 20262 44220 20810
rect 44284 20806 44312 21286
rect 44272 20800 44324 20806
rect 44272 20742 44324 20748
rect 44180 20256 44232 20262
rect 44180 20198 44232 20204
rect 44272 20256 44324 20262
rect 44272 20198 44324 20204
rect 43570 20156 43878 20165
rect 43570 20154 43576 20156
rect 43632 20154 43656 20156
rect 43712 20154 43736 20156
rect 43792 20154 43816 20156
rect 43872 20154 43878 20156
rect 43632 20102 43634 20154
rect 43814 20102 43816 20154
rect 43570 20100 43576 20102
rect 43632 20100 43656 20102
rect 43712 20100 43736 20102
rect 43792 20100 43816 20102
rect 43872 20100 43878 20102
rect 43570 20091 43878 20100
rect 44192 20058 44220 20198
rect 44180 20052 44232 20058
rect 44180 19994 44232 20000
rect 43996 19712 44048 19718
rect 43996 19654 44048 19660
rect 44008 19514 44036 19654
rect 43996 19508 44048 19514
rect 43996 19450 44048 19456
rect 43444 19440 43496 19446
rect 43444 19382 43496 19388
rect 43570 19068 43878 19077
rect 43570 19066 43576 19068
rect 43632 19066 43656 19068
rect 43712 19066 43736 19068
rect 43792 19066 43816 19068
rect 43872 19066 43878 19068
rect 43632 19014 43634 19066
rect 43814 19014 43816 19066
rect 43570 19012 43576 19014
rect 43632 19012 43656 19014
rect 43712 19012 43736 19014
rect 43792 19012 43816 19014
rect 43872 19012 43878 19014
rect 43570 19003 43878 19012
rect 43720 18624 43772 18630
rect 43720 18566 43772 18572
rect 43812 18624 43864 18630
rect 43812 18566 43864 18572
rect 43732 18426 43760 18566
rect 43720 18420 43772 18426
rect 43720 18362 43772 18368
rect 43732 18068 43760 18362
rect 43824 18222 43852 18566
rect 43812 18216 43864 18222
rect 43812 18158 43864 18164
rect 43732 18040 43944 18068
rect 43570 17980 43878 17989
rect 43570 17978 43576 17980
rect 43632 17978 43656 17980
rect 43712 17978 43736 17980
rect 43792 17978 43816 17980
rect 43872 17978 43878 17980
rect 43632 17926 43634 17978
rect 43814 17926 43816 17978
rect 43570 17924 43576 17926
rect 43632 17924 43656 17926
rect 43712 17924 43736 17926
rect 43792 17924 43816 17926
rect 43872 17924 43878 17926
rect 43570 17915 43878 17924
rect 43260 17672 43312 17678
rect 43260 17614 43312 17620
rect 43916 17542 43944 18040
rect 43536 17536 43588 17542
rect 43536 17478 43588 17484
rect 43904 17536 43956 17542
rect 43904 17478 43956 17484
rect 43168 17332 43220 17338
rect 43168 17274 43220 17280
rect 43076 16788 43128 16794
rect 43076 16730 43128 16736
rect 42812 16546 43116 16574
rect 42708 16516 42760 16522
rect 42708 16458 42760 16464
rect 42720 15570 42748 16458
rect 42892 16448 42944 16454
rect 42892 16390 42944 16396
rect 42904 16250 42932 16390
rect 42892 16244 42944 16250
rect 42892 16186 42944 16192
rect 42708 15564 42760 15570
rect 42708 15506 42760 15512
rect 42616 15360 42668 15366
rect 42616 15302 42668 15308
rect 42628 14822 42656 15302
rect 42616 14816 42668 14822
rect 42616 14758 42668 14764
rect 42628 14414 42656 14758
rect 42616 14408 42668 14414
rect 42616 14350 42668 14356
rect 42432 12980 42484 12986
rect 42432 12922 42484 12928
rect 42248 12368 42300 12374
rect 42248 12310 42300 12316
rect 42340 11892 42392 11898
rect 42340 11834 42392 11840
rect 42064 11212 42116 11218
rect 42064 11154 42116 11160
rect 41972 10668 42024 10674
rect 41972 10610 42024 10616
rect 41788 10260 41840 10266
rect 41788 10202 41840 10208
rect 41880 10260 41932 10266
rect 41880 10202 41932 10208
rect 41892 10146 41920 10202
rect 41800 10118 41920 10146
rect 41800 9722 41828 10118
rect 41788 9716 41840 9722
rect 41788 9658 41840 9664
rect 41696 9512 41748 9518
rect 41696 9454 41748 9460
rect 41972 9512 42024 9518
rect 41972 9454 42024 9460
rect 41984 9081 42012 9454
rect 42076 9450 42104 11154
rect 42352 10810 42380 11834
rect 42444 11694 42472 12922
rect 42616 12640 42668 12646
rect 42616 12582 42668 12588
rect 42628 12102 42656 12582
rect 42616 12096 42668 12102
rect 42616 12038 42668 12044
rect 42720 11778 42748 15506
rect 42800 15496 42852 15502
rect 42800 15438 42852 15444
rect 42812 14618 42840 15438
rect 43088 15366 43116 16546
rect 43180 16114 43208 17274
rect 43352 17196 43404 17202
rect 43352 17138 43404 17144
rect 43364 16658 43392 17138
rect 43548 16998 43576 17478
rect 43904 17332 43956 17338
rect 43904 17274 43956 17280
rect 43536 16992 43588 16998
rect 43536 16934 43588 16940
rect 43570 16892 43878 16901
rect 43570 16890 43576 16892
rect 43632 16890 43656 16892
rect 43712 16890 43736 16892
rect 43792 16890 43816 16892
rect 43872 16890 43878 16892
rect 43632 16838 43634 16890
rect 43814 16838 43816 16890
rect 43570 16836 43576 16838
rect 43632 16836 43656 16838
rect 43712 16836 43736 16838
rect 43792 16836 43816 16838
rect 43872 16836 43878 16838
rect 43570 16827 43878 16836
rect 43916 16794 43944 17274
rect 43904 16788 43956 16794
rect 43904 16730 43956 16736
rect 43352 16652 43404 16658
rect 43352 16594 43404 16600
rect 44180 16652 44232 16658
rect 44180 16594 44232 16600
rect 43364 16250 43392 16594
rect 43352 16244 43404 16250
rect 43352 16186 43404 16192
rect 43168 16108 43220 16114
rect 43168 16050 43220 16056
rect 43904 15904 43956 15910
rect 43904 15846 43956 15852
rect 43570 15804 43878 15813
rect 43570 15802 43576 15804
rect 43632 15802 43656 15804
rect 43712 15802 43736 15804
rect 43792 15802 43816 15804
rect 43872 15802 43878 15804
rect 43632 15750 43634 15802
rect 43814 15750 43816 15802
rect 43570 15748 43576 15750
rect 43632 15748 43656 15750
rect 43712 15748 43736 15750
rect 43792 15748 43816 15750
rect 43872 15748 43878 15750
rect 43570 15739 43878 15748
rect 43444 15496 43496 15502
rect 43444 15438 43496 15444
rect 42984 15360 43036 15366
rect 42984 15302 43036 15308
rect 43076 15360 43128 15366
rect 43076 15302 43128 15308
rect 42996 15162 43024 15302
rect 42984 15156 43036 15162
rect 42984 15098 43036 15104
rect 42800 14612 42852 14618
rect 42800 14554 42852 14560
rect 43088 14278 43116 15302
rect 43456 14278 43484 15438
rect 43916 15366 43944 15846
rect 43904 15360 43956 15366
rect 43904 15302 43956 15308
rect 43916 14822 43944 15302
rect 43904 14816 43956 14822
rect 43904 14758 43956 14764
rect 43570 14716 43878 14725
rect 43570 14714 43576 14716
rect 43632 14714 43656 14716
rect 43712 14714 43736 14716
rect 43792 14714 43816 14716
rect 43872 14714 43878 14716
rect 43632 14662 43634 14714
rect 43814 14662 43816 14714
rect 43570 14660 43576 14662
rect 43632 14660 43656 14662
rect 43712 14660 43736 14662
rect 43792 14660 43816 14662
rect 43872 14660 43878 14662
rect 43570 14651 43878 14660
rect 42800 14272 42852 14278
rect 42800 14214 42852 14220
rect 43076 14272 43128 14278
rect 43076 14214 43128 14220
rect 43444 14272 43496 14278
rect 43444 14214 43496 14220
rect 42812 13870 42840 14214
rect 42800 13864 42852 13870
rect 42800 13806 42852 13812
rect 42628 11750 42748 11778
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 42340 10804 42392 10810
rect 42340 10746 42392 10752
rect 42524 10600 42576 10606
rect 42524 10542 42576 10548
rect 42536 9994 42564 10542
rect 42524 9988 42576 9994
rect 42524 9930 42576 9936
rect 42536 9625 42564 9930
rect 42522 9616 42578 9625
rect 42522 9551 42578 9560
rect 42064 9444 42116 9450
rect 42064 9386 42116 9392
rect 41970 9072 42026 9081
rect 41970 9007 42026 9016
rect 41512 8968 41564 8974
rect 41512 8910 41564 8916
rect 42536 8906 42564 9551
rect 42628 9518 42656 11750
rect 42708 11688 42760 11694
rect 42708 11630 42760 11636
rect 42720 11286 42748 11630
rect 42812 11354 42840 13806
rect 43088 13734 43116 14214
rect 43352 13796 43404 13802
rect 43352 13738 43404 13744
rect 43076 13728 43128 13734
rect 43076 13670 43128 13676
rect 43088 13462 43116 13670
rect 43076 13456 43128 13462
rect 43076 13398 43128 13404
rect 43364 13190 43392 13738
rect 43352 13184 43404 13190
rect 43352 13126 43404 13132
rect 42892 12776 42944 12782
rect 42892 12718 42944 12724
rect 42904 12434 42932 12718
rect 43456 12442 43484 14214
rect 43916 13802 43944 14758
rect 44192 14346 44220 16594
rect 44284 14618 44312 20198
rect 44376 16590 44404 22374
rect 44548 21684 44600 21690
rect 44548 21626 44600 21632
rect 44560 21146 44588 21626
rect 44916 21344 44968 21350
rect 44916 21286 44968 21292
rect 44548 21140 44600 21146
rect 44548 21082 44600 21088
rect 44732 20800 44784 20806
rect 44732 20742 44784 20748
rect 44744 19310 44772 20742
rect 44928 20058 44956 21286
rect 44916 20052 44968 20058
rect 44916 19994 44968 20000
rect 44732 19304 44784 19310
rect 44732 19246 44784 19252
rect 44824 18624 44876 18630
rect 44824 18566 44876 18572
rect 44836 18426 44864 18566
rect 44824 18420 44876 18426
rect 44824 18362 44876 18368
rect 44928 17882 44956 19994
rect 44916 17876 44968 17882
rect 44916 17818 44968 17824
rect 44916 17536 44968 17542
rect 44916 17478 44968 17484
rect 44928 17202 44956 17478
rect 44916 17196 44968 17202
rect 44916 17138 44968 17144
rect 44640 16992 44692 16998
rect 44640 16934 44692 16940
rect 44652 16794 44680 16934
rect 44640 16788 44692 16794
rect 44640 16730 44692 16736
rect 44364 16584 44416 16590
rect 44364 16526 44416 16532
rect 44364 15904 44416 15910
rect 44364 15846 44416 15852
rect 44376 15366 44404 15846
rect 45020 15502 45048 22374
rect 45192 20868 45244 20874
rect 45192 20810 45244 20816
rect 45204 20777 45232 20810
rect 45190 20768 45246 20777
rect 45190 20703 45246 20712
rect 45008 15496 45060 15502
rect 45008 15438 45060 15444
rect 44364 15360 44416 15366
rect 44364 15302 44416 15308
rect 44376 14822 44404 15302
rect 45192 15020 45244 15026
rect 45192 14962 45244 14968
rect 44364 14816 44416 14822
rect 44364 14758 44416 14764
rect 45008 14816 45060 14822
rect 45204 14793 45232 14962
rect 45008 14758 45060 14764
rect 45190 14784 45246 14793
rect 44272 14612 44324 14618
rect 44272 14554 44324 14560
rect 44180 14340 44232 14346
rect 44180 14282 44232 14288
rect 43904 13796 43956 13802
rect 43904 13738 43956 13744
rect 43570 13628 43878 13637
rect 43570 13626 43576 13628
rect 43632 13626 43656 13628
rect 43712 13626 43736 13628
rect 43792 13626 43816 13628
rect 43872 13626 43878 13628
rect 43632 13574 43634 13626
rect 43814 13574 43816 13626
rect 43570 13572 43576 13574
rect 43632 13572 43656 13574
rect 43712 13572 43736 13574
rect 43792 13572 43816 13574
rect 43872 13572 43878 13574
rect 43570 13563 43878 13572
rect 43570 12540 43878 12549
rect 43570 12538 43576 12540
rect 43632 12538 43656 12540
rect 43712 12538 43736 12540
rect 43792 12538 43816 12540
rect 43872 12538 43878 12540
rect 43632 12486 43634 12538
rect 43814 12486 43816 12538
rect 43570 12484 43576 12486
rect 43632 12484 43656 12486
rect 43712 12484 43736 12486
rect 43792 12484 43816 12486
rect 43872 12484 43878 12486
rect 43570 12475 43878 12484
rect 43444 12436 43496 12442
rect 42904 12406 43116 12434
rect 43088 12170 43116 12406
rect 43444 12378 43496 12384
rect 43076 12164 43128 12170
rect 43076 12106 43128 12112
rect 43088 11762 43116 12106
rect 43076 11756 43128 11762
rect 43076 11698 43128 11704
rect 42800 11348 42852 11354
rect 42800 11290 42852 11296
rect 42708 11280 42760 11286
rect 42708 11222 42760 11228
rect 42812 11082 42840 11290
rect 43456 11150 43484 12378
rect 43570 11452 43878 11461
rect 43570 11450 43576 11452
rect 43632 11450 43656 11452
rect 43712 11450 43736 11452
rect 43792 11450 43816 11452
rect 43872 11450 43878 11452
rect 43632 11398 43634 11450
rect 43814 11398 43816 11450
rect 43570 11396 43576 11398
rect 43632 11396 43656 11398
rect 43712 11396 43736 11398
rect 43792 11396 43816 11398
rect 43872 11396 43878 11398
rect 43570 11387 43878 11396
rect 43444 11144 43496 11150
rect 43444 11086 43496 11092
rect 42800 11076 42852 11082
rect 42800 11018 42852 11024
rect 42984 11008 43036 11014
rect 42984 10950 43036 10956
rect 42996 10742 43024 10950
rect 44284 10810 44312 14554
rect 44376 14278 44404 14758
rect 44364 14272 44416 14278
rect 44364 14214 44416 14220
rect 44732 14272 44784 14278
rect 44732 14214 44784 14220
rect 44376 13734 44404 14214
rect 44744 13802 44772 14214
rect 44732 13796 44784 13802
rect 44732 13738 44784 13744
rect 44364 13728 44416 13734
rect 44364 13670 44416 13676
rect 44548 13728 44600 13734
rect 44548 13670 44600 13676
rect 44560 13190 44588 13670
rect 44548 13184 44600 13190
rect 44548 13126 44600 13132
rect 44364 12640 44416 12646
rect 44364 12582 44416 12588
rect 44376 12102 44404 12582
rect 44560 12374 44588 13126
rect 44548 12368 44600 12374
rect 44548 12310 44600 12316
rect 44364 12096 44416 12102
rect 44364 12038 44416 12044
rect 44560 11354 44588 12310
rect 44640 12096 44692 12102
rect 44640 12038 44692 12044
rect 44548 11348 44600 11354
rect 44548 11290 44600 11296
rect 44548 11008 44600 11014
rect 44548 10950 44600 10956
rect 44560 10810 44588 10950
rect 43260 10804 43312 10810
rect 43260 10746 43312 10752
rect 44272 10804 44324 10810
rect 44272 10746 44324 10752
rect 44548 10804 44600 10810
rect 44548 10746 44600 10752
rect 42984 10736 43036 10742
rect 42984 10678 43036 10684
rect 42984 10260 43036 10266
rect 42984 10202 43036 10208
rect 42996 9722 43024 10202
rect 43272 10198 43300 10746
rect 43570 10364 43878 10373
rect 43570 10362 43576 10364
rect 43632 10362 43656 10364
rect 43712 10362 43736 10364
rect 43792 10362 43816 10364
rect 43872 10362 43878 10364
rect 43632 10310 43634 10362
rect 43814 10310 43816 10362
rect 43570 10308 43576 10310
rect 43632 10308 43656 10310
rect 43712 10308 43736 10310
rect 43792 10308 43816 10310
rect 43872 10308 43878 10310
rect 43570 10299 43878 10308
rect 44560 10266 44588 10746
rect 44548 10260 44600 10266
rect 44548 10202 44600 10208
rect 43260 10192 43312 10198
rect 44652 10146 44680 12038
rect 44732 11824 44784 11830
rect 44732 11766 44784 11772
rect 44744 11014 44772 11766
rect 45020 11762 45048 14758
rect 45190 14719 45246 14728
rect 45008 11756 45060 11762
rect 45008 11698 45060 11704
rect 44824 11688 44876 11694
rect 44824 11630 44876 11636
rect 44836 11257 44864 11630
rect 44822 11248 44878 11257
rect 44822 11183 44878 11192
rect 44732 11008 44784 11014
rect 44732 10950 44784 10956
rect 44744 10470 44772 10950
rect 44732 10464 44784 10470
rect 44732 10406 44784 10412
rect 44824 10464 44876 10470
rect 44824 10406 44876 10412
rect 43260 10134 43312 10140
rect 43272 9722 43300 10134
rect 44560 10118 44680 10146
rect 42984 9716 43036 9722
rect 42984 9658 43036 9664
rect 43260 9716 43312 9722
rect 43260 9658 43312 9664
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 42616 9512 42668 9518
rect 42616 9454 42668 9460
rect 42524 8900 42576 8906
rect 42524 8842 42576 8848
rect 40960 8832 41012 8838
rect 40960 8774 41012 8780
rect 41880 8832 41932 8838
rect 41880 8774 41932 8780
rect 40972 8634 41000 8774
rect 41070 8732 41378 8741
rect 41070 8730 41076 8732
rect 41132 8730 41156 8732
rect 41212 8730 41236 8732
rect 41292 8730 41316 8732
rect 41372 8730 41378 8732
rect 41132 8678 41134 8730
rect 41314 8678 41316 8730
rect 41070 8676 41076 8678
rect 41132 8676 41156 8678
rect 41212 8676 41236 8678
rect 41292 8676 41316 8678
rect 41372 8676 41378 8678
rect 41070 8667 41378 8676
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 41420 8492 41472 8498
rect 41420 8434 41472 8440
rect 41432 8090 41460 8434
rect 41420 8084 41472 8090
rect 41420 8026 41472 8032
rect 40866 7984 40922 7993
rect 40922 7942 41368 7970
rect 40866 7919 40922 7928
rect 41340 7750 41368 7942
rect 41892 7886 41920 8774
rect 42536 8566 42564 8842
rect 42524 8560 42576 8566
rect 42524 8502 42576 8508
rect 42064 7948 42116 7954
rect 42064 7890 42116 7896
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 40776 7744 40828 7750
rect 40776 7686 40828 7692
rect 41328 7744 41380 7750
rect 41328 7686 41380 7692
rect 40788 7546 40816 7686
rect 41070 7644 41378 7653
rect 41070 7642 41076 7644
rect 41132 7642 41156 7644
rect 41212 7642 41236 7644
rect 41292 7642 41316 7644
rect 41372 7642 41378 7644
rect 41132 7590 41134 7642
rect 41314 7590 41316 7642
rect 41070 7588 41076 7590
rect 41132 7588 41156 7590
rect 41212 7588 41236 7590
rect 41292 7588 41316 7590
rect 41372 7588 41378 7590
rect 41070 7579 41378 7588
rect 40776 7540 40828 7546
rect 40776 7482 40828 7488
rect 41420 7404 41472 7410
rect 41420 7346 41472 7352
rect 41512 7404 41564 7410
rect 41512 7346 41564 7352
rect 40684 7336 40736 7342
rect 40684 7278 40736 7284
rect 41432 7206 41460 7346
rect 40960 7200 41012 7206
rect 40960 7142 41012 7148
rect 41328 7200 41380 7206
rect 41328 7142 41380 7148
rect 41420 7200 41472 7206
rect 41420 7142 41472 7148
rect 39856 6996 39908 7002
rect 39856 6938 39908 6944
rect 40500 6996 40552 7002
rect 40500 6938 40552 6944
rect 40316 6656 40368 6662
rect 40316 6598 40368 6604
rect 40328 6322 40356 6598
rect 40512 6390 40540 6938
rect 40684 6860 40736 6866
rect 40684 6802 40736 6808
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40316 6316 40368 6322
rect 40316 6258 40368 6264
rect 40592 6316 40644 6322
rect 40592 6258 40644 6264
rect 39304 6112 39356 6118
rect 39304 6054 39356 6060
rect 39580 6112 39632 6118
rect 39580 6054 39632 6060
rect 39120 5636 39172 5642
rect 39120 5578 39172 5584
rect 39028 5228 39080 5234
rect 39028 5170 39080 5176
rect 39316 5166 39344 6054
rect 39488 5636 39540 5642
rect 39488 5578 39540 5584
rect 39396 5228 39448 5234
rect 39396 5170 39448 5176
rect 39304 5160 39356 5166
rect 39304 5102 39356 5108
rect 39212 5024 39264 5030
rect 39212 4966 39264 4972
rect 38570 4924 38878 4933
rect 38570 4922 38576 4924
rect 38632 4922 38656 4924
rect 38712 4922 38736 4924
rect 38792 4922 38816 4924
rect 38872 4922 38878 4924
rect 38632 4870 38634 4922
rect 38814 4870 38816 4922
rect 38570 4868 38576 4870
rect 38632 4868 38656 4870
rect 38712 4868 38736 4870
rect 38792 4868 38816 4870
rect 38872 4868 38878 4870
rect 38570 4859 38878 4868
rect 39224 4690 39252 4966
rect 39212 4684 39264 4690
rect 39212 4626 39264 4632
rect 39408 4146 39436 5170
rect 39500 4826 39528 5578
rect 39592 5166 39620 6054
rect 39856 5772 39908 5778
rect 39856 5714 39908 5720
rect 39580 5160 39632 5166
rect 39580 5102 39632 5108
rect 39592 4842 39620 5102
rect 39488 4820 39540 4826
rect 39592 4814 39804 4842
rect 39488 4762 39540 4768
rect 39396 4140 39448 4146
rect 39396 4082 39448 4088
rect 38570 3836 38878 3845
rect 38570 3834 38576 3836
rect 38632 3834 38656 3836
rect 38712 3834 38736 3836
rect 38792 3834 38816 3836
rect 38872 3834 38878 3836
rect 38632 3782 38634 3834
rect 38814 3782 38816 3834
rect 38570 3780 38576 3782
rect 38632 3780 38656 3782
rect 38712 3780 38736 3782
rect 38792 3780 38816 3782
rect 38872 3780 38878 3782
rect 38570 3771 38878 3780
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 38764 3126 38792 3402
rect 39408 3126 39436 4082
rect 39776 4078 39804 4814
rect 39868 4758 39896 5714
rect 40224 5636 40276 5642
rect 40328 5624 40356 6258
rect 40276 5596 40356 5624
rect 40224 5578 40276 5584
rect 40604 5370 40632 6258
rect 40696 6254 40724 6802
rect 40868 6792 40920 6798
rect 40868 6734 40920 6740
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 40774 6216 40830 6225
rect 40774 6151 40776 6160
rect 40828 6151 40830 6160
rect 40776 6122 40828 6128
rect 40880 5710 40908 6734
rect 40972 5846 41000 7142
rect 41340 7002 41368 7142
rect 41328 6996 41380 7002
rect 41328 6938 41380 6944
rect 41070 6556 41378 6565
rect 41070 6554 41076 6556
rect 41132 6554 41156 6556
rect 41212 6554 41236 6556
rect 41292 6554 41316 6556
rect 41372 6554 41378 6556
rect 41132 6502 41134 6554
rect 41314 6502 41316 6554
rect 41070 6500 41076 6502
rect 41132 6500 41156 6502
rect 41212 6500 41236 6502
rect 41292 6500 41316 6502
rect 41372 6500 41378 6502
rect 41070 6491 41378 6500
rect 41524 6458 41552 7346
rect 42076 7342 42104 7890
rect 42064 7336 42116 7342
rect 42064 7278 42116 7284
rect 41880 7200 41932 7206
rect 41880 7142 41932 7148
rect 41892 6866 41920 7142
rect 41880 6860 41932 6866
rect 41880 6802 41932 6808
rect 41512 6452 41564 6458
rect 41512 6394 41564 6400
rect 42076 6254 42104 7278
rect 42536 6866 42564 8502
rect 42720 7954 42748 9522
rect 43272 9178 43300 9658
rect 44560 9382 44588 10118
rect 44744 9625 44772 10406
rect 44836 10198 44864 10406
rect 44824 10192 44876 10198
rect 44824 10134 44876 10140
rect 44730 9616 44786 9625
rect 44640 9580 44692 9586
rect 44730 9551 44786 9560
rect 44640 9522 44692 9528
rect 44548 9376 44600 9382
rect 44548 9318 44600 9324
rect 43570 9276 43878 9285
rect 43570 9274 43576 9276
rect 43632 9274 43656 9276
rect 43712 9274 43736 9276
rect 43792 9274 43816 9276
rect 43872 9274 43878 9276
rect 43632 9222 43634 9274
rect 43814 9222 43816 9274
rect 43570 9220 43576 9222
rect 43632 9220 43656 9222
rect 43712 9220 43736 9222
rect 43792 9220 43816 9222
rect 43872 9220 43878 9222
rect 43570 9211 43878 9220
rect 43260 9172 43312 9178
rect 43260 9114 43312 9120
rect 42800 8288 42852 8294
rect 42800 8230 42852 8236
rect 42812 7954 42840 8230
rect 43272 8090 43300 9114
rect 44560 8838 44588 9318
rect 44548 8832 44600 8838
rect 44652 8809 44680 9522
rect 44744 9450 44772 9551
rect 44732 9444 44784 9450
rect 44732 9386 44784 9392
rect 44916 8832 44968 8838
rect 44548 8774 44600 8780
rect 44638 8800 44694 8809
rect 44560 8650 44588 8774
rect 44916 8774 44968 8780
rect 44638 8735 44694 8744
rect 44560 8622 44680 8650
rect 43444 8424 43496 8430
rect 43444 8366 43496 8372
rect 43260 8084 43312 8090
rect 43260 8026 43312 8032
rect 42708 7948 42760 7954
rect 42708 7890 42760 7896
rect 42800 7948 42852 7954
rect 42800 7890 42852 7896
rect 42720 6905 42748 7890
rect 42890 7848 42946 7857
rect 42890 7783 42946 7792
rect 42706 6896 42762 6905
rect 42524 6860 42576 6866
rect 42706 6831 42762 6840
rect 42800 6860 42852 6866
rect 42524 6802 42576 6808
rect 42064 6248 42116 6254
rect 42064 6190 42116 6196
rect 40960 5840 41012 5846
rect 40960 5782 41012 5788
rect 42536 5778 42564 6802
rect 42720 6254 42748 6831
rect 42800 6802 42852 6808
rect 42812 6458 42840 6802
rect 42904 6798 42932 7783
rect 43272 7546 43300 8026
rect 43456 7750 43484 8366
rect 44548 8288 44600 8294
rect 44548 8230 44600 8236
rect 43570 8188 43878 8197
rect 43570 8186 43576 8188
rect 43632 8186 43656 8188
rect 43712 8186 43736 8188
rect 43792 8186 43816 8188
rect 43872 8186 43878 8188
rect 43632 8134 43634 8186
rect 43814 8134 43816 8186
rect 43570 8132 43576 8134
rect 43632 8132 43656 8134
rect 43712 8132 43736 8134
rect 43792 8132 43816 8134
rect 43872 8132 43878 8134
rect 43570 8123 43878 8132
rect 44560 7750 44588 8230
rect 43444 7744 43496 7750
rect 43444 7686 43496 7692
rect 44180 7744 44232 7750
rect 44180 7686 44232 7692
rect 44548 7744 44600 7750
rect 44548 7686 44600 7692
rect 43260 7540 43312 7546
rect 43312 7500 43392 7528
rect 43260 7482 43312 7488
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 42892 6792 42944 6798
rect 42892 6734 42944 6740
rect 43088 6458 43116 7346
rect 43260 6656 43312 6662
rect 43260 6598 43312 6604
rect 42800 6452 42852 6458
rect 42800 6394 42852 6400
rect 43076 6452 43128 6458
rect 43076 6394 43128 6400
rect 42708 6248 42760 6254
rect 42708 6190 42760 6196
rect 42984 6112 43036 6118
rect 42984 6054 43036 6060
rect 42524 5772 42576 5778
rect 42524 5714 42576 5720
rect 40868 5704 40920 5710
rect 40920 5664 41000 5692
rect 40868 5646 40920 5652
rect 40868 5568 40920 5574
rect 40868 5510 40920 5516
rect 40040 5364 40092 5370
rect 40040 5306 40092 5312
rect 40592 5364 40644 5370
rect 40592 5306 40644 5312
rect 39948 5228 40000 5234
rect 39948 5170 40000 5176
rect 39856 4752 39908 4758
rect 39856 4694 39908 4700
rect 39960 4622 39988 5170
rect 40052 4690 40080 5306
rect 40132 5296 40184 5302
rect 40132 5238 40184 5244
rect 40040 4684 40092 4690
rect 40040 4626 40092 4632
rect 39948 4616 40000 4622
rect 39948 4558 40000 4564
rect 39960 4282 39988 4558
rect 40040 4480 40092 4486
rect 40040 4422 40092 4428
rect 39948 4276 40000 4282
rect 39948 4218 40000 4224
rect 39764 4072 39816 4078
rect 39764 4014 39816 4020
rect 38752 3120 38804 3126
rect 38752 3062 38804 3068
rect 39028 3120 39080 3126
rect 39028 3062 39080 3068
rect 39396 3120 39448 3126
rect 39448 3080 39528 3108
rect 39396 3062 39448 3068
rect 38752 2984 38804 2990
rect 38804 2944 38976 2972
rect 38752 2926 38804 2932
rect 38570 2748 38878 2757
rect 38570 2746 38576 2748
rect 38632 2746 38656 2748
rect 38712 2746 38736 2748
rect 38792 2746 38816 2748
rect 38872 2746 38878 2748
rect 38632 2694 38634 2746
rect 38814 2694 38816 2746
rect 38570 2692 38576 2694
rect 38632 2692 38656 2694
rect 38712 2692 38736 2694
rect 38792 2692 38816 2694
rect 38872 2692 38878 2694
rect 38570 2683 38878 2692
rect 38948 2650 38976 2944
rect 38936 2644 38988 2650
rect 38936 2586 38988 2592
rect 39040 2106 39068 3062
rect 39396 2848 39448 2854
rect 39396 2790 39448 2796
rect 39408 2446 39436 2790
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39500 2106 39528 3080
rect 39580 2576 39632 2582
rect 39580 2518 39632 2524
rect 39028 2100 39080 2106
rect 39028 2042 39080 2048
rect 39488 2100 39540 2106
rect 39488 2042 39540 2048
rect 38844 1760 38896 1766
rect 38896 1720 38976 1748
rect 38844 1702 38896 1708
rect 38570 1660 38878 1669
rect 38570 1658 38576 1660
rect 38632 1658 38656 1660
rect 38712 1658 38736 1660
rect 38792 1658 38816 1660
rect 38872 1658 38878 1660
rect 38632 1606 38634 1658
rect 38814 1606 38816 1658
rect 38570 1604 38576 1606
rect 38632 1604 38656 1606
rect 38712 1604 38736 1606
rect 38792 1604 38816 1606
rect 38872 1604 38878 1606
rect 38570 1595 38878 1604
rect 38948 1562 38976 1720
rect 38936 1556 38988 1562
rect 38936 1498 38988 1504
rect 39500 1358 39528 2042
rect 39592 1358 39620 2518
rect 39776 2514 39804 4014
rect 39948 3936 40000 3942
rect 39948 3878 40000 3884
rect 39960 3738 39988 3878
rect 39948 3732 40000 3738
rect 39948 3674 40000 3680
rect 40052 3602 40080 4422
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 40144 3058 40172 5238
rect 40880 5166 40908 5510
rect 40972 5370 41000 5664
rect 41070 5468 41378 5477
rect 41070 5466 41076 5468
rect 41132 5466 41156 5468
rect 41212 5466 41236 5468
rect 41292 5466 41316 5468
rect 41372 5466 41378 5468
rect 41132 5414 41134 5466
rect 41314 5414 41316 5466
rect 41070 5412 41076 5414
rect 41132 5412 41156 5414
rect 41212 5412 41236 5414
rect 41292 5412 41316 5414
rect 41372 5412 41378 5414
rect 41070 5403 41378 5412
rect 40960 5364 41012 5370
rect 40960 5306 41012 5312
rect 41788 5364 41840 5370
rect 41788 5306 41840 5312
rect 40868 5160 40920 5166
rect 40868 5102 40920 5108
rect 40960 5160 41012 5166
rect 40960 5102 41012 5108
rect 40592 4820 40644 4826
rect 40592 4762 40644 4768
rect 40408 4752 40460 4758
rect 40408 4694 40460 4700
rect 40224 4140 40276 4146
rect 40224 4082 40276 4088
rect 40316 4140 40368 4146
rect 40316 4082 40368 4088
rect 40236 3602 40264 4082
rect 40224 3596 40276 3602
rect 40224 3538 40276 3544
rect 40328 3194 40356 4082
rect 40316 3188 40368 3194
rect 40316 3130 40368 3136
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 40328 2514 40356 3130
rect 40420 2650 40448 4694
rect 40500 4480 40552 4486
rect 40500 4422 40552 4428
rect 40512 4282 40540 4422
rect 40500 4276 40552 4282
rect 40500 4218 40552 4224
rect 40604 3670 40632 4762
rect 40880 4554 40908 5102
rect 40868 4548 40920 4554
rect 40868 4490 40920 4496
rect 40972 4434 41000 5102
rect 41800 4826 41828 5306
rect 42064 5228 42116 5234
rect 42064 5170 42116 5176
rect 41972 5024 42024 5030
rect 41972 4966 42024 4972
rect 41788 4820 41840 4826
rect 41840 4780 41920 4808
rect 41788 4762 41840 4768
rect 41512 4548 41564 4554
rect 41512 4490 41564 4496
rect 40880 4406 41000 4434
rect 40880 3942 40908 4406
rect 41070 4380 41378 4389
rect 41070 4378 41076 4380
rect 41132 4378 41156 4380
rect 41212 4378 41236 4380
rect 41292 4378 41316 4380
rect 41372 4378 41378 4380
rect 41132 4326 41134 4378
rect 41314 4326 41316 4378
rect 41070 4324 41076 4326
rect 41132 4324 41156 4326
rect 41212 4324 41236 4326
rect 41292 4324 41316 4326
rect 41372 4324 41378 4326
rect 41070 4315 41378 4324
rect 40960 4276 41012 4282
rect 40960 4218 41012 4224
rect 40868 3936 40920 3942
rect 40868 3878 40920 3884
rect 40592 3664 40644 3670
rect 40592 3606 40644 3612
rect 40592 3120 40644 3126
rect 40592 3062 40644 3068
rect 40682 3088 40738 3097
rect 40500 2984 40552 2990
rect 40500 2926 40552 2932
rect 40408 2644 40460 2650
rect 40408 2586 40460 2592
rect 39764 2508 39816 2514
rect 39764 2450 39816 2456
rect 40316 2508 40368 2514
rect 40316 2450 40368 2456
rect 39764 2372 39816 2378
rect 39764 2314 39816 2320
rect 40132 2372 40184 2378
rect 40132 2314 40184 2320
rect 39776 1358 39804 2314
rect 40040 2100 40092 2106
rect 40040 2042 40092 2048
rect 40052 1408 40080 2042
rect 39868 1380 40080 1408
rect 39488 1352 39540 1358
rect 39488 1294 39540 1300
rect 39580 1352 39632 1358
rect 39580 1294 39632 1300
rect 39672 1352 39724 1358
rect 39672 1294 39724 1300
rect 39764 1352 39816 1358
rect 39764 1294 39816 1300
rect 39028 1216 39080 1222
rect 39684 1204 39712 1294
rect 39868 1204 39896 1380
rect 39948 1284 40000 1290
rect 39948 1226 40000 1232
rect 39684 1176 39896 1204
rect 39028 1158 39080 1164
rect 39040 950 39068 1158
rect 39028 944 39080 950
rect 39028 886 39080 892
rect 38476 876 38528 882
rect 38476 818 38528 824
rect 39396 808 39448 814
rect 39396 750 39448 756
rect 39132 190 39252 218
rect 39132 160 39160 190
rect 37462 54 37872 82
rect 37462 -300 37518 54
rect 38290 -300 38346 160
rect 39118 -300 39174 160
rect 39224 82 39252 190
rect 39408 82 39436 750
rect 39960 160 39988 1226
rect 40144 950 40172 2314
rect 40316 2304 40368 2310
rect 40316 2246 40368 2252
rect 40224 1760 40276 1766
rect 40224 1702 40276 1708
rect 40236 1562 40264 1702
rect 40224 1556 40276 1562
rect 40224 1498 40276 1504
rect 40328 1358 40356 2246
rect 40512 2106 40540 2926
rect 40500 2100 40552 2106
rect 40500 2042 40552 2048
rect 40408 2032 40460 2038
rect 40408 1974 40460 1980
rect 40316 1352 40368 1358
rect 40316 1294 40368 1300
rect 40420 1222 40448 1974
rect 40604 1970 40632 3062
rect 40682 3023 40738 3032
rect 40696 2106 40724 3023
rect 40880 2990 40908 3878
rect 40972 3738 41000 4218
rect 41524 4185 41552 4490
rect 41892 4282 41920 4780
rect 41984 4729 42012 4966
rect 41970 4720 42026 4729
rect 41970 4655 42026 4664
rect 41984 4282 42012 4655
rect 41880 4276 41932 4282
rect 41880 4218 41932 4224
rect 41972 4276 42024 4282
rect 41972 4218 42024 4224
rect 41788 4208 41840 4214
rect 41510 4176 41566 4185
rect 41788 4150 41840 4156
rect 41510 4111 41566 4120
rect 40960 3732 41012 3738
rect 40960 3674 41012 3680
rect 41070 3292 41378 3301
rect 41070 3290 41076 3292
rect 41132 3290 41156 3292
rect 41212 3290 41236 3292
rect 41292 3290 41316 3292
rect 41372 3290 41378 3292
rect 41132 3238 41134 3290
rect 41314 3238 41316 3290
rect 41070 3236 41076 3238
rect 41132 3236 41156 3238
rect 41212 3236 41236 3238
rect 41292 3236 41316 3238
rect 41372 3236 41378 3238
rect 41070 3227 41378 3236
rect 41420 3052 41472 3058
rect 41420 2994 41472 3000
rect 40868 2984 40920 2990
rect 40868 2926 40920 2932
rect 40880 2514 40908 2926
rect 40868 2508 40920 2514
rect 40868 2450 40920 2456
rect 40866 2408 40922 2417
rect 40866 2343 40922 2352
rect 40880 2310 40908 2343
rect 40868 2304 40920 2310
rect 40868 2246 40920 2252
rect 40960 2304 41012 2310
rect 40960 2246 41012 2252
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 40592 1964 40644 1970
rect 40592 1906 40644 1912
rect 40972 1562 41000 2246
rect 41070 2204 41378 2213
rect 41070 2202 41076 2204
rect 41132 2202 41156 2204
rect 41212 2202 41236 2204
rect 41292 2202 41316 2204
rect 41372 2202 41378 2204
rect 41132 2150 41134 2202
rect 41314 2150 41316 2202
rect 41070 2148 41076 2150
rect 41132 2148 41156 2150
rect 41212 2148 41236 2150
rect 41292 2148 41316 2150
rect 41372 2148 41378 2150
rect 41070 2139 41378 2148
rect 40960 1556 41012 1562
rect 40960 1498 41012 1504
rect 40776 1352 40828 1358
rect 40498 1320 40554 1329
rect 40554 1278 40724 1306
rect 40776 1294 40828 1300
rect 40868 1352 40920 1358
rect 41328 1352 41380 1358
rect 40868 1294 40920 1300
rect 40972 1312 41328 1340
rect 40498 1255 40554 1264
rect 40696 1222 40724 1278
rect 40408 1216 40460 1222
rect 40408 1158 40460 1164
rect 40684 1216 40736 1222
rect 40684 1158 40736 1164
rect 40132 944 40184 950
rect 40132 886 40184 892
rect 40788 746 40816 1294
rect 40880 1018 40908 1294
rect 40868 1012 40920 1018
rect 40868 954 40920 960
rect 40972 814 41000 1312
rect 41328 1294 41380 1300
rect 41432 1222 41460 2994
rect 41510 2544 41566 2553
rect 41510 2479 41566 2488
rect 41524 2038 41552 2479
rect 41512 2032 41564 2038
rect 41512 1974 41564 1980
rect 41696 1284 41748 1290
rect 41616 1244 41696 1272
rect 41420 1216 41472 1222
rect 41420 1158 41472 1164
rect 41070 1116 41378 1125
rect 41070 1114 41076 1116
rect 41132 1114 41156 1116
rect 41212 1114 41236 1116
rect 41292 1114 41316 1116
rect 41372 1114 41378 1116
rect 41132 1062 41134 1114
rect 41314 1062 41316 1114
rect 41070 1060 41076 1062
rect 41132 1060 41156 1062
rect 41212 1060 41236 1062
rect 41292 1060 41316 1062
rect 41372 1060 41378 1062
rect 41070 1051 41378 1060
rect 40960 808 41012 814
rect 40960 750 41012 756
rect 40776 740 40828 746
rect 40776 682 40828 688
rect 40960 672 41012 678
rect 40960 614 41012 620
rect 40972 354 41000 614
rect 40788 326 41000 354
rect 40788 160 40816 326
rect 41616 160 41644 1244
rect 41696 1226 41748 1232
rect 41800 1222 41828 4150
rect 41892 3738 41920 4218
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41892 3194 41920 3674
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41892 2650 41920 3130
rect 41880 2644 41932 2650
rect 41880 2586 41932 2592
rect 41972 1352 42024 1358
rect 41972 1294 42024 1300
rect 41788 1216 41840 1222
rect 41788 1158 41840 1164
rect 41984 678 42012 1294
rect 42076 1222 42104 5170
rect 42248 4820 42300 4826
rect 42248 4762 42300 4768
rect 42260 3670 42288 4762
rect 42536 4690 42564 5714
rect 42892 5296 42944 5302
rect 42892 5238 42944 5244
rect 42904 4826 42932 5238
rect 42996 4826 43024 6054
rect 43088 5914 43116 6394
rect 43076 5908 43128 5914
rect 43076 5850 43128 5856
rect 43076 5568 43128 5574
rect 43076 5510 43128 5516
rect 43088 5370 43116 5510
rect 43076 5364 43128 5370
rect 43076 5306 43128 5312
rect 42892 4820 42944 4826
rect 42892 4762 42944 4768
rect 42984 4820 43036 4826
rect 42984 4762 43036 4768
rect 42524 4684 42576 4690
rect 42524 4626 42576 4632
rect 42536 3670 42564 4626
rect 42996 4282 43024 4762
rect 42984 4276 43036 4282
rect 42984 4218 43036 4224
rect 42248 3664 42300 3670
rect 42248 3606 42300 3612
rect 42524 3664 42576 3670
rect 42524 3606 42576 3612
rect 42260 3126 42288 3606
rect 42248 3120 42300 3126
rect 42248 3062 42300 3068
rect 42260 2582 42288 3062
rect 42432 2644 42484 2650
rect 42432 2586 42484 2592
rect 42248 2576 42300 2582
rect 42248 2518 42300 2524
rect 42260 2106 42288 2518
rect 42248 2100 42300 2106
rect 42248 2042 42300 2048
rect 42444 2038 42472 2586
rect 42984 2100 43036 2106
rect 42984 2042 43036 2048
rect 42432 2032 42484 2038
rect 42432 1974 42484 1980
rect 42996 1562 43024 2042
rect 42984 1556 43036 1562
rect 42984 1498 43036 1504
rect 43272 1358 43300 6598
rect 43364 6458 43392 7500
rect 43456 7206 43484 7686
rect 44192 7478 44220 7686
rect 44560 7546 44588 7686
rect 44548 7540 44600 7546
rect 44548 7482 44600 7488
rect 44180 7472 44232 7478
rect 44178 7440 44180 7449
rect 44232 7440 44234 7449
rect 44178 7375 44234 7384
rect 44548 7268 44600 7274
rect 44548 7210 44600 7216
rect 43444 7200 43496 7206
rect 43444 7142 43496 7148
rect 43456 7002 43484 7142
rect 43570 7100 43878 7109
rect 43570 7098 43576 7100
rect 43632 7098 43656 7100
rect 43712 7098 43736 7100
rect 43792 7098 43816 7100
rect 43872 7098 43878 7100
rect 43632 7046 43634 7098
rect 43814 7046 43816 7098
rect 43570 7044 43576 7046
rect 43632 7044 43656 7046
rect 43712 7044 43736 7046
rect 43792 7044 43816 7046
rect 43872 7044 43878 7046
rect 43570 7035 43878 7044
rect 43444 6996 43496 7002
rect 43444 6938 43496 6944
rect 44180 6860 44232 6866
rect 44180 6802 44232 6808
rect 43352 6452 43404 6458
rect 43352 6394 43404 6400
rect 43364 5914 43392 6394
rect 44192 6254 44220 6802
rect 44364 6316 44416 6322
rect 44364 6258 44416 6264
rect 44180 6248 44232 6254
rect 44180 6190 44232 6196
rect 43996 6112 44048 6118
rect 43996 6054 44048 6060
rect 43570 6012 43878 6021
rect 43570 6010 43576 6012
rect 43632 6010 43656 6012
rect 43712 6010 43736 6012
rect 43792 6010 43816 6012
rect 43872 6010 43878 6012
rect 43632 5958 43634 6010
rect 43814 5958 43816 6010
rect 43570 5956 43576 5958
rect 43632 5956 43656 5958
rect 43712 5956 43736 5958
rect 43792 5956 43816 5958
rect 43872 5956 43878 5958
rect 43570 5947 43878 5956
rect 43352 5908 43404 5914
rect 43352 5850 43404 5856
rect 43364 5302 43392 5850
rect 44008 5370 44036 6054
rect 43996 5364 44048 5370
rect 43996 5306 44048 5312
rect 43352 5296 43404 5302
rect 43352 5238 43404 5244
rect 43570 4924 43878 4933
rect 43570 4922 43576 4924
rect 43632 4922 43656 4924
rect 43712 4922 43736 4924
rect 43792 4922 43816 4924
rect 43872 4922 43878 4924
rect 43632 4870 43634 4922
rect 43814 4870 43816 4922
rect 43570 4868 43576 4870
rect 43632 4868 43656 4870
rect 43712 4868 43736 4870
rect 43792 4868 43816 4870
rect 43872 4868 43878 4870
rect 43570 4859 43878 4868
rect 44008 4758 44036 5306
rect 44192 5030 44220 6190
rect 44088 5024 44140 5030
rect 44088 4966 44140 4972
rect 44180 5024 44232 5030
rect 44180 4966 44232 4972
rect 44100 4826 44128 4966
rect 44088 4820 44140 4826
rect 44088 4762 44140 4768
rect 43996 4752 44048 4758
rect 43996 4694 44048 4700
rect 43444 4684 43496 4690
rect 43444 4626 43496 4632
rect 43456 4282 43484 4626
rect 44008 4282 44036 4694
rect 43444 4276 43496 4282
rect 43444 4218 43496 4224
rect 43996 4276 44048 4282
rect 43996 4218 44048 4224
rect 43570 3836 43878 3845
rect 43570 3834 43576 3836
rect 43632 3834 43656 3836
rect 43712 3834 43736 3836
rect 43792 3834 43816 3836
rect 43872 3834 43878 3836
rect 43632 3782 43634 3834
rect 43814 3782 43816 3834
rect 43570 3780 43576 3782
rect 43632 3780 43656 3782
rect 43712 3780 43736 3782
rect 43792 3780 43816 3782
rect 43872 3780 43878 3782
rect 43570 3771 43878 3780
rect 43352 3664 43404 3670
rect 43352 3606 43404 3612
rect 43364 2650 43392 3606
rect 43570 2748 43878 2757
rect 43570 2746 43576 2748
rect 43632 2746 43656 2748
rect 43712 2746 43736 2748
rect 43792 2746 43816 2748
rect 43872 2746 43878 2748
rect 43632 2694 43634 2746
rect 43814 2694 43816 2746
rect 43570 2692 43576 2694
rect 43632 2692 43656 2694
rect 43712 2692 43736 2694
rect 43792 2692 43816 2694
rect 43872 2692 43878 2694
rect 43570 2683 43878 2692
rect 44192 2650 44220 4966
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 43812 2508 43864 2514
rect 43812 2450 43864 2456
rect 43824 2106 43852 2450
rect 43812 2100 43864 2106
rect 43864 2060 43944 2088
rect 43812 2042 43864 2048
rect 43570 1660 43878 1669
rect 43570 1658 43576 1660
rect 43632 1658 43656 1660
rect 43712 1658 43736 1660
rect 43792 1658 43816 1660
rect 43872 1658 43878 1660
rect 43632 1606 43634 1658
rect 43814 1606 43816 1658
rect 43570 1604 43576 1606
rect 43632 1604 43656 1606
rect 43712 1604 43736 1606
rect 43792 1604 43816 1606
rect 43872 1604 43878 1606
rect 43570 1595 43878 1604
rect 43916 1562 43944 2060
rect 43904 1556 43956 1562
rect 43904 1498 43956 1504
rect 44376 1358 44404 6258
rect 44560 5370 44588 7210
rect 44548 5364 44600 5370
rect 44548 5306 44600 5312
rect 44560 3738 44588 5306
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 44652 3618 44680 8622
rect 44928 8430 44956 8774
rect 44916 8424 44968 8430
rect 44916 8366 44968 8372
rect 45008 7812 45060 7818
rect 45008 7754 45060 7760
rect 44916 7744 44968 7750
rect 44916 7686 44968 7692
rect 44732 7472 44784 7478
rect 44732 7414 44784 7420
rect 44744 6458 44772 7414
rect 44928 7002 44956 7686
rect 44916 6996 44968 7002
rect 44916 6938 44968 6944
rect 44732 6452 44784 6458
rect 44732 6394 44784 6400
rect 44916 5908 44968 5914
rect 44916 5850 44968 5856
rect 44732 4276 44784 4282
rect 44732 4218 44784 4224
rect 44744 3670 44772 4218
rect 44928 3738 44956 5850
rect 44824 3732 44876 3738
rect 44824 3674 44876 3680
rect 44916 3732 44968 3738
rect 44916 3674 44968 3680
rect 44560 3590 44680 3618
rect 44732 3664 44784 3670
rect 44732 3606 44784 3612
rect 44560 2106 44588 3590
rect 44744 3194 44772 3606
rect 44732 3188 44784 3194
rect 44732 3130 44784 3136
rect 44640 3052 44692 3058
rect 44640 2994 44692 3000
rect 44652 2825 44680 2994
rect 44638 2816 44694 2825
rect 44638 2751 44694 2760
rect 44744 2650 44772 3130
rect 44732 2644 44784 2650
rect 44732 2586 44784 2592
rect 44744 2106 44772 2586
rect 44548 2100 44600 2106
rect 44548 2042 44600 2048
rect 44732 2100 44784 2106
rect 44732 2042 44784 2048
rect 44836 1358 44864 3674
rect 45020 1358 45048 7754
rect 42708 1352 42760 1358
rect 42708 1294 42760 1300
rect 43260 1352 43312 1358
rect 43260 1294 43312 1300
rect 43536 1352 43588 1358
rect 43536 1294 43588 1300
rect 44364 1352 44416 1358
rect 44364 1294 44416 1300
rect 44548 1352 44600 1358
rect 44548 1294 44600 1300
rect 44824 1352 44876 1358
rect 44824 1294 44876 1300
rect 45008 1352 45060 1358
rect 45008 1294 45060 1300
rect 45192 1352 45244 1358
rect 45192 1294 45244 1300
rect 42064 1216 42116 1222
rect 42064 1158 42116 1164
rect 42524 1216 42576 1222
rect 42524 1158 42576 1164
rect 42536 882 42564 1158
rect 42524 876 42576 882
rect 42524 818 42576 824
rect 41972 672 42024 678
rect 41972 614 42024 620
rect 39224 54 39436 82
rect 39946 -300 40002 160
rect 40774 -300 40830 160
rect 41602 -300 41658 160
rect 42430 82 42486 160
rect 42720 82 42748 1294
rect 42430 54 42748 82
rect 43258 82 43314 160
rect 43548 82 43576 1294
rect 43258 54 43576 82
rect 44086 82 44142 160
rect 44560 82 44588 1294
rect 44086 54 44588 82
rect 44914 82 44970 160
rect 45204 82 45232 1294
rect 44914 54 45232 82
rect 42430 -300 42486 54
rect 43258 -300 43314 54
rect 44086 -300 44142 54
rect 44914 -300 44970 54
<< via2 >>
rect 3576 22330 3632 22332
rect 3656 22330 3712 22332
rect 3736 22330 3792 22332
rect 3816 22330 3872 22332
rect 3576 22278 3622 22330
rect 3622 22278 3632 22330
rect 3656 22278 3686 22330
rect 3686 22278 3698 22330
rect 3698 22278 3712 22330
rect 3736 22278 3750 22330
rect 3750 22278 3762 22330
rect 3762 22278 3792 22330
rect 3816 22278 3826 22330
rect 3826 22278 3872 22330
rect 3576 22276 3632 22278
rect 3656 22276 3712 22278
rect 3736 22276 3792 22278
rect 3816 22276 3872 22278
rect 6076 22874 6132 22876
rect 6156 22874 6212 22876
rect 6236 22874 6292 22876
rect 6316 22874 6372 22876
rect 6076 22822 6122 22874
rect 6122 22822 6132 22874
rect 6156 22822 6186 22874
rect 6186 22822 6198 22874
rect 6198 22822 6212 22874
rect 6236 22822 6250 22874
rect 6250 22822 6262 22874
rect 6262 22822 6292 22874
rect 6316 22822 6326 22874
rect 6326 22822 6372 22874
rect 6076 22820 6132 22822
rect 6156 22820 6212 22822
rect 6236 22820 6292 22822
rect 6316 22820 6372 22822
rect 11076 22874 11132 22876
rect 11156 22874 11212 22876
rect 11236 22874 11292 22876
rect 11316 22874 11372 22876
rect 11076 22822 11122 22874
rect 11122 22822 11132 22874
rect 11156 22822 11186 22874
rect 11186 22822 11198 22874
rect 11198 22822 11212 22874
rect 11236 22822 11250 22874
rect 11250 22822 11262 22874
rect 11262 22822 11292 22874
rect 11316 22822 11326 22874
rect 11326 22822 11372 22874
rect 11076 22820 11132 22822
rect 11156 22820 11212 22822
rect 11236 22820 11292 22822
rect 11316 22820 11372 22822
rect 5078 22072 5134 22128
rect 4434 21972 4436 21992
rect 4436 21972 4488 21992
rect 4488 21972 4490 21992
rect 938 20712 994 20768
rect 938 14728 994 14784
rect 938 8780 940 8800
rect 940 8780 992 8800
rect 992 8780 994 8800
rect 938 8744 994 8780
rect 4434 21936 4490 21972
rect 3576 21242 3632 21244
rect 3656 21242 3712 21244
rect 3736 21242 3792 21244
rect 3816 21242 3872 21244
rect 3576 21190 3622 21242
rect 3622 21190 3632 21242
rect 3656 21190 3686 21242
rect 3686 21190 3698 21242
rect 3698 21190 3712 21242
rect 3736 21190 3750 21242
rect 3750 21190 3762 21242
rect 3762 21190 3792 21242
rect 3816 21190 3826 21242
rect 3826 21190 3872 21242
rect 3576 21188 3632 21190
rect 3656 21188 3712 21190
rect 3736 21188 3792 21190
rect 3816 21188 3872 21190
rect 3576 20154 3632 20156
rect 3656 20154 3712 20156
rect 3736 20154 3792 20156
rect 3816 20154 3872 20156
rect 3576 20102 3622 20154
rect 3622 20102 3632 20154
rect 3656 20102 3686 20154
rect 3686 20102 3698 20154
rect 3698 20102 3712 20154
rect 3736 20102 3750 20154
rect 3750 20102 3762 20154
rect 3762 20102 3792 20154
rect 3816 20102 3826 20154
rect 3826 20102 3872 20154
rect 3576 20100 3632 20102
rect 3656 20100 3712 20102
rect 3736 20100 3792 20102
rect 3816 20100 3872 20102
rect 3576 19066 3632 19068
rect 3656 19066 3712 19068
rect 3736 19066 3792 19068
rect 3816 19066 3872 19068
rect 3576 19014 3622 19066
rect 3622 19014 3632 19066
rect 3656 19014 3686 19066
rect 3686 19014 3698 19066
rect 3698 19014 3712 19066
rect 3736 19014 3750 19066
rect 3750 19014 3762 19066
rect 3762 19014 3792 19066
rect 3816 19014 3826 19066
rect 3826 19014 3872 19066
rect 3576 19012 3632 19014
rect 3656 19012 3712 19014
rect 3736 19012 3792 19014
rect 3816 19012 3872 19014
rect 3576 17978 3632 17980
rect 3656 17978 3712 17980
rect 3736 17978 3792 17980
rect 3816 17978 3872 17980
rect 3576 17926 3622 17978
rect 3622 17926 3632 17978
rect 3656 17926 3686 17978
rect 3686 17926 3698 17978
rect 3698 17926 3712 17978
rect 3736 17926 3750 17978
rect 3750 17926 3762 17978
rect 3762 17926 3792 17978
rect 3816 17926 3826 17978
rect 3826 17926 3872 17978
rect 3576 17924 3632 17926
rect 3656 17924 3712 17926
rect 3736 17924 3792 17926
rect 3816 17924 3872 17926
rect 3576 16890 3632 16892
rect 3656 16890 3712 16892
rect 3736 16890 3792 16892
rect 3816 16890 3872 16892
rect 3576 16838 3622 16890
rect 3622 16838 3632 16890
rect 3656 16838 3686 16890
rect 3686 16838 3698 16890
rect 3698 16838 3712 16890
rect 3736 16838 3750 16890
rect 3750 16838 3762 16890
rect 3762 16838 3792 16890
rect 3816 16838 3826 16890
rect 3826 16838 3872 16890
rect 3576 16836 3632 16838
rect 3656 16836 3712 16838
rect 3736 16836 3792 16838
rect 3816 16836 3872 16838
rect 3576 15802 3632 15804
rect 3656 15802 3712 15804
rect 3736 15802 3792 15804
rect 3816 15802 3872 15804
rect 3576 15750 3622 15802
rect 3622 15750 3632 15802
rect 3656 15750 3686 15802
rect 3686 15750 3698 15802
rect 3698 15750 3712 15802
rect 3736 15750 3750 15802
rect 3750 15750 3762 15802
rect 3762 15750 3792 15802
rect 3816 15750 3826 15802
rect 3826 15750 3872 15802
rect 3576 15748 3632 15750
rect 3656 15748 3712 15750
rect 3736 15748 3792 15750
rect 3816 15748 3872 15750
rect 3576 14714 3632 14716
rect 3656 14714 3712 14716
rect 3736 14714 3792 14716
rect 3816 14714 3872 14716
rect 3576 14662 3622 14714
rect 3622 14662 3632 14714
rect 3656 14662 3686 14714
rect 3686 14662 3698 14714
rect 3698 14662 3712 14714
rect 3736 14662 3750 14714
rect 3750 14662 3762 14714
rect 3762 14662 3792 14714
rect 3816 14662 3826 14714
rect 3826 14662 3872 14714
rect 3576 14660 3632 14662
rect 3656 14660 3712 14662
rect 3736 14660 3792 14662
rect 3816 14660 3872 14662
rect 3576 13626 3632 13628
rect 3656 13626 3712 13628
rect 3736 13626 3792 13628
rect 3816 13626 3872 13628
rect 3576 13574 3622 13626
rect 3622 13574 3632 13626
rect 3656 13574 3686 13626
rect 3686 13574 3698 13626
rect 3698 13574 3712 13626
rect 3736 13574 3750 13626
rect 3750 13574 3762 13626
rect 3762 13574 3792 13626
rect 3816 13574 3826 13626
rect 3826 13574 3872 13626
rect 3576 13572 3632 13574
rect 3656 13572 3712 13574
rect 3736 13572 3792 13574
rect 3816 13572 3872 13574
rect 3576 12538 3632 12540
rect 3656 12538 3712 12540
rect 3736 12538 3792 12540
rect 3816 12538 3872 12540
rect 3576 12486 3622 12538
rect 3622 12486 3632 12538
rect 3656 12486 3686 12538
rect 3686 12486 3698 12538
rect 3698 12486 3712 12538
rect 3736 12486 3750 12538
rect 3750 12486 3762 12538
rect 3762 12486 3792 12538
rect 3816 12486 3826 12538
rect 3826 12486 3872 12538
rect 3576 12484 3632 12486
rect 3656 12484 3712 12486
rect 3736 12484 3792 12486
rect 3816 12484 3872 12486
rect 8576 22330 8632 22332
rect 8656 22330 8712 22332
rect 8736 22330 8792 22332
rect 8816 22330 8872 22332
rect 8576 22278 8622 22330
rect 8622 22278 8632 22330
rect 8656 22278 8686 22330
rect 8686 22278 8698 22330
rect 8698 22278 8712 22330
rect 8736 22278 8750 22330
rect 8750 22278 8762 22330
rect 8762 22278 8792 22330
rect 8816 22278 8826 22330
rect 8826 22278 8872 22330
rect 8576 22276 8632 22278
rect 8656 22276 8712 22278
rect 8736 22276 8792 22278
rect 8816 22276 8872 22278
rect 5354 21936 5410 21992
rect 6076 21786 6132 21788
rect 6156 21786 6212 21788
rect 6236 21786 6292 21788
rect 6316 21786 6372 21788
rect 6076 21734 6122 21786
rect 6122 21734 6132 21786
rect 6156 21734 6186 21786
rect 6186 21734 6198 21786
rect 6198 21734 6212 21786
rect 6236 21734 6250 21786
rect 6250 21734 6262 21786
rect 6262 21734 6292 21786
rect 6316 21734 6326 21786
rect 6326 21734 6372 21786
rect 6076 21732 6132 21734
rect 6156 21732 6212 21734
rect 6236 21732 6292 21734
rect 6316 21732 6372 21734
rect 6458 21528 6514 21584
rect 5446 19896 5502 19952
rect 6076 20698 6132 20700
rect 6156 20698 6212 20700
rect 6236 20698 6292 20700
rect 6316 20698 6372 20700
rect 6076 20646 6122 20698
rect 6122 20646 6132 20698
rect 6156 20646 6186 20698
rect 6186 20646 6198 20698
rect 6198 20646 6212 20698
rect 6236 20646 6250 20698
rect 6250 20646 6262 20698
rect 6262 20646 6292 20698
rect 6316 20646 6326 20698
rect 6326 20646 6372 20698
rect 6076 20644 6132 20646
rect 6156 20644 6212 20646
rect 6236 20644 6292 20646
rect 6316 20644 6372 20646
rect 6076 19610 6132 19612
rect 6156 19610 6212 19612
rect 6236 19610 6292 19612
rect 6316 19610 6372 19612
rect 6076 19558 6122 19610
rect 6122 19558 6132 19610
rect 6156 19558 6186 19610
rect 6186 19558 6198 19610
rect 6198 19558 6212 19610
rect 6236 19558 6250 19610
rect 6250 19558 6262 19610
rect 6262 19558 6292 19610
rect 6316 19558 6326 19610
rect 6326 19558 6372 19610
rect 6076 19556 6132 19558
rect 6156 19556 6212 19558
rect 6236 19556 6292 19558
rect 6316 19556 6372 19558
rect 6076 18522 6132 18524
rect 6156 18522 6212 18524
rect 6236 18522 6292 18524
rect 6316 18522 6372 18524
rect 6076 18470 6122 18522
rect 6122 18470 6132 18522
rect 6156 18470 6186 18522
rect 6186 18470 6198 18522
rect 6198 18470 6212 18522
rect 6236 18470 6250 18522
rect 6250 18470 6262 18522
rect 6262 18470 6292 18522
rect 6316 18470 6326 18522
rect 6326 18470 6372 18522
rect 6076 18468 6132 18470
rect 6156 18468 6212 18470
rect 6236 18468 6292 18470
rect 6316 18468 6372 18470
rect 6076 17434 6132 17436
rect 6156 17434 6212 17436
rect 6236 17434 6292 17436
rect 6316 17434 6372 17436
rect 6076 17382 6122 17434
rect 6122 17382 6132 17434
rect 6156 17382 6186 17434
rect 6186 17382 6198 17434
rect 6198 17382 6212 17434
rect 6236 17382 6250 17434
rect 6250 17382 6262 17434
rect 6262 17382 6292 17434
rect 6316 17382 6326 17434
rect 6326 17382 6372 17434
rect 6076 17380 6132 17382
rect 6156 17380 6212 17382
rect 6236 17380 6292 17382
rect 6316 17380 6372 17382
rect 6076 16346 6132 16348
rect 6156 16346 6212 16348
rect 6236 16346 6292 16348
rect 6316 16346 6372 16348
rect 6076 16294 6122 16346
rect 6122 16294 6132 16346
rect 6156 16294 6186 16346
rect 6186 16294 6198 16346
rect 6198 16294 6212 16346
rect 6236 16294 6250 16346
rect 6250 16294 6262 16346
rect 6262 16294 6292 16346
rect 6316 16294 6326 16346
rect 6326 16294 6372 16346
rect 6076 16292 6132 16294
rect 6156 16292 6212 16294
rect 6236 16292 6292 16294
rect 6316 16292 6372 16294
rect 6076 15258 6132 15260
rect 6156 15258 6212 15260
rect 6236 15258 6292 15260
rect 6316 15258 6372 15260
rect 6076 15206 6122 15258
rect 6122 15206 6132 15258
rect 6156 15206 6186 15258
rect 6186 15206 6198 15258
rect 6198 15206 6212 15258
rect 6236 15206 6250 15258
rect 6250 15206 6262 15258
rect 6262 15206 6292 15258
rect 6316 15206 6326 15258
rect 6326 15206 6372 15258
rect 6076 15204 6132 15206
rect 6156 15204 6212 15206
rect 6236 15204 6292 15206
rect 6316 15204 6372 15206
rect 6076 14170 6132 14172
rect 6156 14170 6212 14172
rect 6236 14170 6292 14172
rect 6316 14170 6372 14172
rect 6076 14118 6122 14170
rect 6122 14118 6132 14170
rect 6156 14118 6186 14170
rect 6186 14118 6198 14170
rect 6198 14118 6212 14170
rect 6236 14118 6250 14170
rect 6250 14118 6262 14170
rect 6262 14118 6292 14170
rect 6316 14118 6326 14170
rect 6326 14118 6372 14170
rect 6076 14116 6132 14118
rect 6156 14116 6212 14118
rect 6236 14116 6292 14118
rect 6316 14116 6372 14118
rect 6076 13082 6132 13084
rect 6156 13082 6212 13084
rect 6236 13082 6292 13084
rect 6316 13082 6372 13084
rect 6076 13030 6122 13082
rect 6122 13030 6132 13082
rect 6156 13030 6186 13082
rect 6186 13030 6198 13082
rect 6198 13030 6212 13082
rect 6236 13030 6250 13082
rect 6250 13030 6262 13082
rect 6262 13030 6292 13082
rect 6316 13030 6326 13082
rect 6326 13030 6372 13082
rect 6076 13028 6132 13030
rect 6156 13028 6212 13030
rect 6236 13028 6292 13030
rect 6316 13028 6372 13030
rect 3576 11450 3632 11452
rect 3656 11450 3712 11452
rect 3736 11450 3792 11452
rect 3816 11450 3872 11452
rect 3576 11398 3622 11450
rect 3622 11398 3632 11450
rect 3656 11398 3686 11450
rect 3686 11398 3698 11450
rect 3698 11398 3712 11450
rect 3736 11398 3750 11450
rect 3750 11398 3762 11450
rect 3762 11398 3792 11450
rect 3816 11398 3826 11450
rect 3826 11398 3872 11450
rect 3576 11396 3632 11398
rect 3656 11396 3712 11398
rect 3736 11396 3792 11398
rect 3816 11396 3872 11398
rect 3576 10362 3632 10364
rect 3656 10362 3712 10364
rect 3736 10362 3792 10364
rect 3816 10362 3872 10364
rect 3576 10310 3622 10362
rect 3622 10310 3632 10362
rect 3656 10310 3686 10362
rect 3686 10310 3698 10362
rect 3698 10310 3712 10362
rect 3736 10310 3750 10362
rect 3750 10310 3762 10362
rect 3762 10310 3792 10362
rect 3816 10310 3826 10362
rect 3826 10310 3872 10362
rect 3576 10308 3632 10310
rect 3656 10308 3712 10310
rect 3736 10308 3792 10310
rect 3816 10308 3872 10310
rect 3576 9274 3632 9276
rect 3656 9274 3712 9276
rect 3736 9274 3792 9276
rect 3816 9274 3872 9276
rect 3576 9222 3622 9274
rect 3622 9222 3632 9274
rect 3656 9222 3686 9274
rect 3686 9222 3698 9274
rect 3698 9222 3712 9274
rect 3736 9222 3750 9274
rect 3750 9222 3762 9274
rect 3762 9222 3792 9274
rect 3816 9222 3826 9274
rect 3826 9222 3872 9274
rect 3576 9220 3632 9222
rect 3656 9220 3712 9222
rect 3736 9220 3792 9222
rect 3816 9220 3872 9222
rect 3576 8186 3632 8188
rect 3656 8186 3712 8188
rect 3736 8186 3792 8188
rect 3816 8186 3872 8188
rect 3576 8134 3622 8186
rect 3622 8134 3632 8186
rect 3656 8134 3686 8186
rect 3686 8134 3698 8186
rect 3698 8134 3712 8186
rect 3736 8134 3750 8186
rect 3750 8134 3762 8186
rect 3762 8134 3792 8186
rect 3816 8134 3826 8186
rect 3826 8134 3872 8186
rect 3576 8132 3632 8134
rect 3656 8132 3712 8134
rect 3736 8132 3792 8134
rect 3816 8132 3872 8134
rect 3576 7098 3632 7100
rect 3656 7098 3712 7100
rect 3736 7098 3792 7100
rect 3816 7098 3872 7100
rect 3576 7046 3622 7098
rect 3622 7046 3632 7098
rect 3656 7046 3686 7098
rect 3686 7046 3698 7098
rect 3698 7046 3712 7098
rect 3736 7046 3750 7098
rect 3750 7046 3762 7098
rect 3762 7046 3792 7098
rect 3816 7046 3826 7098
rect 3826 7046 3872 7098
rect 3576 7044 3632 7046
rect 3656 7044 3712 7046
rect 3736 7044 3792 7046
rect 3816 7044 3872 7046
rect 3576 6010 3632 6012
rect 3656 6010 3712 6012
rect 3736 6010 3792 6012
rect 3816 6010 3872 6012
rect 3576 5958 3622 6010
rect 3622 5958 3632 6010
rect 3656 5958 3686 6010
rect 3686 5958 3698 6010
rect 3698 5958 3712 6010
rect 3736 5958 3750 6010
rect 3750 5958 3762 6010
rect 3762 5958 3792 6010
rect 3816 5958 3826 6010
rect 3826 5958 3872 6010
rect 3576 5956 3632 5958
rect 3656 5956 3712 5958
rect 3736 5956 3792 5958
rect 3816 5956 3872 5958
rect 754 2760 810 2816
rect 3422 5616 3478 5672
rect 3576 4922 3632 4924
rect 3656 4922 3712 4924
rect 3736 4922 3792 4924
rect 3816 4922 3872 4924
rect 3576 4870 3622 4922
rect 3622 4870 3632 4922
rect 3656 4870 3686 4922
rect 3686 4870 3698 4922
rect 3698 4870 3712 4922
rect 3736 4870 3750 4922
rect 3750 4870 3762 4922
rect 3762 4870 3792 4922
rect 3816 4870 3826 4922
rect 3826 4870 3872 4922
rect 3576 4868 3632 4870
rect 3656 4868 3712 4870
rect 3736 4868 3792 4870
rect 3816 4868 3872 4870
rect 3514 4564 3516 4584
rect 3516 4564 3568 4584
rect 3568 4564 3570 4584
rect 3514 4528 3570 4564
rect 3576 3834 3632 3836
rect 3656 3834 3712 3836
rect 3736 3834 3792 3836
rect 3816 3834 3872 3836
rect 3576 3782 3622 3834
rect 3622 3782 3632 3834
rect 3656 3782 3686 3834
rect 3686 3782 3698 3834
rect 3698 3782 3712 3834
rect 3736 3782 3750 3834
rect 3750 3782 3762 3834
rect 3762 3782 3792 3834
rect 3816 3782 3826 3834
rect 3826 3782 3872 3834
rect 3576 3780 3632 3782
rect 3656 3780 3712 3782
rect 3736 3780 3792 3782
rect 3816 3780 3872 3782
rect 4986 11872 5042 11928
rect 5170 11772 5172 11792
rect 5172 11772 5224 11792
rect 5224 11772 5226 11792
rect 5170 11736 5226 11772
rect 5538 11872 5594 11928
rect 6076 11994 6132 11996
rect 6156 11994 6212 11996
rect 6236 11994 6292 11996
rect 6316 11994 6372 11996
rect 6076 11942 6122 11994
rect 6122 11942 6132 11994
rect 6156 11942 6186 11994
rect 6186 11942 6198 11994
rect 6198 11942 6212 11994
rect 6236 11942 6250 11994
rect 6250 11942 6262 11994
rect 6262 11942 6292 11994
rect 6316 11942 6326 11994
rect 6326 11942 6372 11994
rect 6076 11940 6132 11942
rect 6156 11940 6212 11942
rect 6236 11940 6292 11942
rect 6316 11940 6372 11942
rect 5722 11772 5724 11792
rect 5724 11772 5776 11792
rect 5776 11772 5778 11792
rect 5722 11736 5778 11772
rect 6076 10906 6132 10908
rect 6156 10906 6212 10908
rect 6236 10906 6292 10908
rect 6316 10906 6372 10908
rect 6076 10854 6122 10906
rect 6122 10854 6132 10906
rect 6156 10854 6186 10906
rect 6186 10854 6198 10906
rect 6198 10854 6212 10906
rect 6236 10854 6250 10906
rect 6250 10854 6262 10906
rect 6262 10854 6292 10906
rect 6316 10854 6326 10906
rect 6326 10854 6372 10906
rect 6076 10852 6132 10854
rect 6156 10852 6212 10854
rect 6236 10852 6292 10854
rect 6316 10852 6372 10854
rect 6076 9818 6132 9820
rect 6156 9818 6212 9820
rect 6236 9818 6292 9820
rect 6316 9818 6372 9820
rect 6076 9766 6122 9818
rect 6122 9766 6132 9818
rect 6156 9766 6186 9818
rect 6186 9766 6198 9818
rect 6198 9766 6212 9818
rect 6236 9766 6250 9818
rect 6250 9766 6262 9818
rect 6262 9766 6292 9818
rect 6316 9766 6326 9818
rect 6326 9766 6372 9818
rect 6076 9764 6132 9766
rect 6156 9764 6212 9766
rect 6236 9764 6292 9766
rect 6316 9764 6372 9766
rect 6076 8730 6132 8732
rect 6156 8730 6212 8732
rect 6236 8730 6292 8732
rect 6316 8730 6372 8732
rect 6076 8678 6122 8730
rect 6122 8678 6132 8730
rect 6156 8678 6186 8730
rect 6186 8678 6198 8730
rect 6198 8678 6212 8730
rect 6236 8678 6250 8730
rect 6250 8678 6262 8730
rect 6262 8678 6292 8730
rect 6316 8678 6326 8730
rect 6326 8678 6372 8730
rect 6076 8676 6132 8678
rect 6156 8676 6212 8678
rect 6236 8676 6292 8678
rect 6316 8676 6372 8678
rect 6076 7642 6132 7644
rect 6156 7642 6212 7644
rect 6236 7642 6292 7644
rect 6316 7642 6372 7644
rect 6076 7590 6122 7642
rect 6122 7590 6132 7642
rect 6156 7590 6186 7642
rect 6186 7590 6198 7642
rect 6198 7590 6212 7642
rect 6236 7590 6250 7642
rect 6250 7590 6262 7642
rect 6262 7590 6292 7642
rect 6316 7590 6326 7642
rect 6326 7590 6372 7642
rect 6076 7588 6132 7590
rect 6156 7588 6212 7590
rect 6236 7588 6292 7590
rect 6316 7588 6372 7590
rect 6076 6554 6132 6556
rect 6156 6554 6212 6556
rect 6236 6554 6292 6556
rect 6316 6554 6372 6556
rect 6076 6502 6122 6554
rect 6122 6502 6132 6554
rect 6156 6502 6186 6554
rect 6186 6502 6198 6554
rect 6198 6502 6212 6554
rect 6236 6502 6250 6554
rect 6250 6502 6262 6554
rect 6262 6502 6292 6554
rect 6316 6502 6326 6554
rect 6326 6502 6372 6554
rect 6076 6500 6132 6502
rect 6156 6500 6212 6502
rect 6236 6500 6292 6502
rect 6316 6500 6372 6502
rect 3576 2746 3632 2748
rect 3656 2746 3712 2748
rect 3736 2746 3792 2748
rect 3816 2746 3872 2748
rect 3576 2694 3622 2746
rect 3622 2694 3632 2746
rect 3656 2694 3686 2746
rect 3686 2694 3698 2746
rect 3698 2694 3712 2746
rect 3736 2694 3750 2746
rect 3750 2694 3762 2746
rect 3762 2694 3792 2746
rect 3816 2694 3826 2746
rect 3826 2694 3872 2746
rect 3576 2692 3632 2694
rect 3656 2692 3712 2694
rect 3736 2692 3792 2694
rect 3816 2692 3872 2694
rect 5446 4664 5502 4720
rect 6076 5466 6132 5468
rect 6156 5466 6212 5468
rect 6236 5466 6292 5468
rect 6316 5466 6372 5468
rect 6076 5414 6122 5466
rect 6122 5414 6132 5466
rect 6156 5414 6186 5466
rect 6186 5414 6198 5466
rect 6198 5414 6212 5466
rect 6236 5414 6250 5466
rect 6250 5414 6262 5466
rect 6262 5414 6292 5466
rect 6316 5414 6326 5466
rect 6326 5414 6372 5466
rect 6076 5412 6132 5414
rect 6156 5412 6212 5414
rect 6236 5412 6292 5414
rect 6316 5412 6372 5414
rect 6734 19252 6736 19272
rect 6736 19252 6788 19272
rect 6788 19252 6790 19272
rect 6734 19216 6790 19252
rect 8576 21242 8632 21244
rect 8656 21242 8712 21244
rect 8736 21242 8792 21244
rect 8816 21242 8872 21244
rect 8576 21190 8622 21242
rect 8622 21190 8632 21242
rect 8656 21190 8686 21242
rect 8686 21190 8698 21242
rect 8698 21190 8712 21242
rect 8736 21190 8750 21242
rect 8750 21190 8762 21242
rect 8762 21190 8792 21242
rect 8816 21190 8826 21242
rect 8826 21190 8872 21242
rect 8576 21188 8632 21190
rect 8656 21188 8712 21190
rect 8736 21188 8792 21190
rect 8816 21188 8872 21190
rect 8942 20712 8998 20768
rect 8576 20154 8632 20156
rect 8656 20154 8712 20156
rect 8736 20154 8792 20156
rect 8816 20154 8872 20156
rect 8576 20102 8622 20154
rect 8622 20102 8632 20154
rect 8656 20102 8686 20154
rect 8686 20102 8698 20154
rect 8698 20102 8712 20154
rect 8736 20102 8750 20154
rect 8750 20102 8762 20154
rect 8762 20102 8792 20154
rect 8816 20102 8826 20154
rect 8826 20102 8872 20154
rect 8576 20100 8632 20102
rect 8656 20100 8712 20102
rect 8736 20100 8792 20102
rect 8816 20100 8872 20102
rect 8576 19066 8632 19068
rect 8656 19066 8712 19068
rect 8736 19066 8792 19068
rect 8816 19066 8872 19068
rect 8576 19014 8622 19066
rect 8622 19014 8632 19066
rect 8656 19014 8686 19066
rect 8686 19014 8698 19066
rect 8698 19014 8712 19066
rect 8736 19014 8750 19066
rect 8750 19014 8762 19066
rect 8762 19014 8792 19066
rect 8816 19014 8826 19066
rect 8826 19014 8872 19066
rect 8576 19012 8632 19014
rect 8656 19012 8712 19014
rect 8736 19012 8792 19014
rect 8816 19012 8872 19014
rect 8576 17978 8632 17980
rect 8656 17978 8712 17980
rect 8736 17978 8792 17980
rect 8816 17978 8872 17980
rect 8576 17926 8622 17978
rect 8622 17926 8632 17978
rect 8656 17926 8686 17978
rect 8686 17926 8698 17978
rect 8698 17926 8712 17978
rect 8736 17926 8750 17978
rect 8750 17926 8762 17978
rect 8762 17926 8792 17978
rect 8816 17926 8826 17978
rect 8826 17926 8872 17978
rect 8576 17924 8632 17926
rect 8656 17924 8712 17926
rect 8736 17924 8792 17926
rect 8816 17924 8872 17926
rect 8206 17040 8262 17096
rect 8576 16890 8632 16892
rect 8656 16890 8712 16892
rect 8736 16890 8792 16892
rect 8816 16890 8872 16892
rect 8576 16838 8622 16890
rect 8622 16838 8632 16890
rect 8656 16838 8686 16890
rect 8686 16838 8698 16890
rect 8698 16838 8712 16890
rect 8736 16838 8750 16890
rect 8750 16838 8762 16890
rect 8762 16838 8792 16890
rect 8816 16838 8826 16890
rect 8826 16838 8872 16890
rect 8576 16836 8632 16838
rect 8656 16836 8712 16838
rect 8736 16836 8792 16838
rect 8816 16836 8872 16838
rect 8576 15802 8632 15804
rect 8656 15802 8712 15804
rect 8736 15802 8792 15804
rect 8816 15802 8872 15804
rect 8576 15750 8622 15802
rect 8622 15750 8632 15802
rect 8656 15750 8686 15802
rect 8686 15750 8698 15802
rect 8698 15750 8712 15802
rect 8736 15750 8750 15802
rect 8750 15750 8762 15802
rect 8762 15750 8792 15802
rect 8816 15750 8826 15802
rect 8826 15750 8872 15802
rect 8576 15748 8632 15750
rect 8656 15748 8712 15750
rect 8736 15748 8792 15750
rect 8816 15748 8872 15750
rect 8576 14714 8632 14716
rect 8656 14714 8712 14716
rect 8736 14714 8792 14716
rect 8816 14714 8872 14716
rect 8576 14662 8622 14714
rect 8622 14662 8632 14714
rect 8656 14662 8686 14714
rect 8686 14662 8698 14714
rect 8698 14662 8712 14714
rect 8736 14662 8750 14714
rect 8750 14662 8762 14714
rect 8762 14662 8792 14714
rect 8816 14662 8826 14714
rect 8826 14662 8872 14714
rect 8576 14660 8632 14662
rect 8656 14660 8712 14662
rect 8736 14660 8792 14662
rect 8816 14660 8872 14662
rect 8576 13626 8632 13628
rect 8656 13626 8712 13628
rect 8736 13626 8792 13628
rect 8816 13626 8872 13628
rect 8576 13574 8622 13626
rect 8622 13574 8632 13626
rect 8656 13574 8686 13626
rect 8686 13574 8698 13626
rect 8698 13574 8712 13626
rect 8736 13574 8750 13626
rect 8750 13574 8762 13626
rect 8762 13574 8792 13626
rect 8816 13574 8826 13626
rect 8826 13574 8872 13626
rect 8576 13572 8632 13574
rect 8656 13572 8712 13574
rect 8736 13572 8792 13574
rect 8816 13572 8872 13574
rect 9402 12824 9458 12880
rect 8576 12538 8632 12540
rect 8656 12538 8712 12540
rect 8736 12538 8792 12540
rect 8816 12538 8872 12540
rect 8576 12486 8622 12538
rect 8622 12486 8632 12538
rect 8656 12486 8686 12538
rect 8686 12486 8698 12538
rect 8698 12486 8712 12538
rect 8736 12486 8750 12538
rect 8750 12486 8762 12538
rect 8762 12486 8792 12538
rect 8816 12486 8826 12538
rect 8826 12486 8872 12538
rect 8576 12484 8632 12486
rect 8656 12484 8712 12486
rect 8736 12484 8792 12486
rect 8816 12484 8872 12486
rect 8576 11450 8632 11452
rect 8656 11450 8712 11452
rect 8736 11450 8792 11452
rect 8816 11450 8872 11452
rect 8576 11398 8622 11450
rect 8622 11398 8632 11450
rect 8656 11398 8686 11450
rect 8686 11398 8698 11450
rect 8698 11398 8712 11450
rect 8736 11398 8750 11450
rect 8750 11398 8762 11450
rect 8762 11398 8792 11450
rect 8816 11398 8826 11450
rect 8826 11398 8872 11450
rect 8576 11396 8632 11398
rect 8656 11396 8712 11398
rect 8736 11396 8792 11398
rect 8816 11396 8872 11398
rect 8576 10362 8632 10364
rect 8656 10362 8712 10364
rect 8736 10362 8792 10364
rect 8816 10362 8872 10364
rect 8576 10310 8622 10362
rect 8622 10310 8632 10362
rect 8656 10310 8686 10362
rect 8686 10310 8698 10362
rect 8698 10310 8712 10362
rect 8736 10310 8750 10362
rect 8750 10310 8762 10362
rect 8762 10310 8792 10362
rect 8816 10310 8826 10362
rect 8826 10310 8872 10362
rect 8576 10308 8632 10310
rect 8656 10308 8712 10310
rect 8736 10308 8792 10310
rect 8816 10308 8872 10310
rect 6076 4378 6132 4380
rect 6156 4378 6212 4380
rect 6236 4378 6292 4380
rect 6316 4378 6372 4380
rect 6076 4326 6122 4378
rect 6122 4326 6132 4378
rect 6156 4326 6186 4378
rect 6186 4326 6198 4378
rect 6198 4326 6212 4378
rect 6236 4326 6250 4378
rect 6250 4326 6262 4378
rect 6262 4326 6292 4378
rect 6316 4326 6326 4378
rect 6326 4326 6372 4378
rect 6076 4324 6132 4326
rect 6156 4324 6212 4326
rect 6236 4324 6292 4326
rect 6316 4324 6372 4326
rect 6076 3290 6132 3292
rect 6156 3290 6212 3292
rect 6236 3290 6292 3292
rect 6316 3290 6372 3292
rect 6076 3238 6122 3290
rect 6122 3238 6132 3290
rect 6156 3238 6186 3290
rect 6186 3238 6198 3290
rect 6198 3238 6212 3290
rect 6236 3238 6250 3290
rect 6250 3238 6262 3290
rect 6262 3238 6292 3290
rect 6316 3238 6326 3290
rect 6326 3238 6372 3290
rect 6076 3236 6132 3238
rect 6156 3236 6212 3238
rect 6236 3236 6292 3238
rect 6316 3236 6372 3238
rect 3576 1658 3632 1660
rect 3656 1658 3712 1660
rect 3736 1658 3792 1660
rect 3816 1658 3872 1660
rect 3576 1606 3622 1658
rect 3622 1606 3632 1658
rect 3656 1606 3686 1658
rect 3686 1606 3698 1658
rect 3698 1606 3712 1658
rect 3736 1606 3750 1658
rect 3750 1606 3762 1658
rect 3762 1606 3792 1658
rect 3816 1606 3826 1658
rect 3826 1606 3872 1658
rect 3576 1604 3632 1606
rect 3656 1604 3712 1606
rect 3736 1604 3792 1606
rect 3816 1604 3872 1606
rect 6076 2202 6132 2204
rect 6156 2202 6212 2204
rect 6236 2202 6292 2204
rect 6316 2202 6372 2204
rect 6076 2150 6122 2202
rect 6122 2150 6132 2202
rect 6156 2150 6186 2202
rect 6186 2150 6198 2202
rect 6198 2150 6212 2202
rect 6236 2150 6250 2202
rect 6250 2150 6262 2202
rect 6262 2150 6292 2202
rect 6316 2150 6326 2202
rect 6326 2150 6372 2202
rect 6076 2148 6132 2150
rect 6156 2148 6212 2150
rect 6236 2148 6292 2150
rect 6316 2148 6372 2150
rect 8576 9274 8632 9276
rect 8656 9274 8712 9276
rect 8736 9274 8792 9276
rect 8816 9274 8872 9276
rect 8576 9222 8622 9274
rect 8622 9222 8632 9274
rect 8656 9222 8686 9274
rect 8686 9222 8698 9274
rect 8698 9222 8712 9274
rect 8736 9222 8750 9274
rect 8750 9222 8762 9274
rect 8762 9222 8792 9274
rect 8816 9222 8826 9274
rect 8826 9222 8872 9274
rect 8576 9220 8632 9222
rect 8656 9220 8712 9222
rect 8736 9220 8792 9222
rect 8816 9220 8872 9222
rect 8576 8186 8632 8188
rect 8656 8186 8712 8188
rect 8736 8186 8792 8188
rect 8816 8186 8872 8188
rect 8576 8134 8622 8186
rect 8622 8134 8632 8186
rect 8656 8134 8686 8186
rect 8686 8134 8698 8186
rect 8698 8134 8712 8186
rect 8736 8134 8750 8186
rect 8750 8134 8762 8186
rect 8762 8134 8792 8186
rect 8816 8134 8826 8186
rect 8826 8134 8872 8186
rect 8576 8132 8632 8134
rect 8656 8132 8712 8134
rect 8736 8132 8792 8134
rect 8816 8132 8872 8134
rect 8576 7098 8632 7100
rect 8656 7098 8712 7100
rect 8736 7098 8792 7100
rect 8816 7098 8872 7100
rect 8576 7046 8622 7098
rect 8622 7046 8632 7098
rect 8656 7046 8686 7098
rect 8686 7046 8698 7098
rect 8698 7046 8712 7098
rect 8736 7046 8750 7098
rect 8750 7046 8762 7098
rect 8762 7046 8792 7098
rect 8816 7046 8826 7098
rect 8826 7046 8872 7098
rect 8576 7044 8632 7046
rect 8656 7044 8712 7046
rect 8736 7044 8792 7046
rect 8816 7044 8872 7046
rect 9218 6840 9274 6896
rect 11076 21786 11132 21788
rect 11156 21786 11212 21788
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11076 21734 11122 21786
rect 11122 21734 11132 21786
rect 11156 21734 11186 21786
rect 11186 21734 11198 21786
rect 11198 21734 11212 21786
rect 11236 21734 11250 21786
rect 11250 21734 11262 21786
rect 11262 21734 11292 21786
rect 11316 21734 11326 21786
rect 11326 21734 11372 21786
rect 11076 21732 11132 21734
rect 11156 21732 11212 21734
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11076 20698 11132 20700
rect 11156 20698 11212 20700
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11076 20646 11122 20698
rect 11122 20646 11132 20698
rect 11156 20646 11186 20698
rect 11186 20646 11198 20698
rect 11198 20646 11212 20698
rect 11236 20646 11250 20698
rect 11250 20646 11262 20698
rect 11262 20646 11292 20698
rect 11316 20646 11326 20698
rect 11326 20646 11372 20698
rect 11076 20644 11132 20646
rect 11156 20644 11212 20646
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11702 21392 11758 21448
rect 12806 22516 12808 22536
rect 12808 22516 12860 22536
rect 12860 22516 12862 22536
rect 12806 22480 12862 22516
rect 13576 22330 13632 22332
rect 13656 22330 13712 22332
rect 13736 22330 13792 22332
rect 13816 22330 13872 22332
rect 13576 22278 13622 22330
rect 13622 22278 13632 22330
rect 13656 22278 13686 22330
rect 13686 22278 13698 22330
rect 13698 22278 13712 22330
rect 13736 22278 13750 22330
rect 13750 22278 13762 22330
rect 13762 22278 13792 22330
rect 13816 22278 13826 22330
rect 13826 22278 13872 22330
rect 13576 22276 13632 22278
rect 13656 22276 13712 22278
rect 13736 22276 13792 22278
rect 13816 22276 13872 22278
rect 16076 22874 16132 22876
rect 16156 22874 16212 22876
rect 16236 22874 16292 22876
rect 16316 22874 16372 22876
rect 16076 22822 16122 22874
rect 16122 22822 16132 22874
rect 16156 22822 16186 22874
rect 16186 22822 16198 22874
rect 16198 22822 16212 22874
rect 16236 22822 16250 22874
rect 16250 22822 16262 22874
rect 16262 22822 16292 22874
rect 16316 22822 16326 22874
rect 16326 22822 16372 22874
rect 16076 22820 16132 22822
rect 16156 22820 16212 22822
rect 16236 22820 16292 22822
rect 16316 22820 16372 22822
rect 11610 20304 11666 20360
rect 11076 19610 11132 19612
rect 11156 19610 11212 19612
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11076 19558 11122 19610
rect 11122 19558 11132 19610
rect 11156 19558 11186 19610
rect 11186 19558 11198 19610
rect 11198 19558 11212 19610
rect 11236 19558 11250 19610
rect 11250 19558 11262 19610
rect 11262 19558 11292 19610
rect 11316 19558 11326 19610
rect 11326 19558 11372 19610
rect 11076 19556 11132 19558
rect 11156 19556 11212 19558
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 12622 20984 12678 21040
rect 12070 19760 12126 19816
rect 11076 18522 11132 18524
rect 11156 18522 11212 18524
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11076 18470 11122 18522
rect 11122 18470 11132 18522
rect 11156 18470 11186 18522
rect 11186 18470 11198 18522
rect 11198 18470 11212 18522
rect 11236 18470 11250 18522
rect 11250 18470 11262 18522
rect 11262 18470 11292 18522
rect 11316 18470 11326 18522
rect 11326 18470 11372 18522
rect 11076 18468 11132 18470
rect 11156 18468 11212 18470
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11076 17434 11132 17436
rect 11156 17434 11212 17436
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11076 17382 11122 17434
rect 11122 17382 11132 17434
rect 11156 17382 11186 17434
rect 11186 17382 11198 17434
rect 11198 17382 11212 17434
rect 11236 17382 11250 17434
rect 11250 17382 11262 17434
rect 11262 17382 11292 17434
rect 11316 17382 11326 17434
rect 11326 17382 11372 17434
rect 11076 17380 11132 17382
rect 11156 17380 11212 17382
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11076 16346 11132 16348
rect 11156 16346 11212 16348
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11076 16294 11122 16346
rect 11122 16294 11132 16346
rect 11156 16294 11186 16346
rect 11186 16294 11198 16346
rect 11198 16294 11212 16346
rect 11236 16294 11250 16346
rect 11250 16294 11262 16346
rect 11262 16294 11292 16346
rect 11316 16294 11326 16346
rect 11326 16294 11372 16346
rect 11076 16292 11132 16294
rect 11156 16292 11212 16294
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11076 15258 11132 15260
rect 11156 15258 11212 15260
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11076 15206 11122 15258
rect 11122 15206 11132 15258
rect 11156 15206 11186 15258
rect 11186 15206 11198 15258
rect 11198 15206 11212 15258
rect 11236 15206 11250 15258
rect 11250 15206 11262 15258
rect 11262 15206 11292 15258
rect 11316 15206 11326 15258
rect 11326 15206 11372 15258
rect 11076 15204 11132 15206
rect 11156 15204 11212 15206
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 13082 17176 13138 17232
rect 11076 14170 11132 14172
rect 11156 14170 11212 14172
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11076 14118 11122 14170
rect 11122 14118 11132 14170
rect 11156 14118 11186 14170
rect 11186 14118 11198 14170
rect 11198 14118 11212 14170
rect 11236 14118 11250 14170
rect 11250 14118 11262 14170
rect 11262 14118 11292 14170
rect 11316 14118 11326 14170
rect 11326 14118 11372 14170
rect 11076 14116 11132 14118
rect 11156 14116 11212 14118
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11076 13082 11132 13084
rect 11156 13082 11212 13084
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11076 13030 11122 13082
rect 11122 13030 11132 13082
rect 11156 13030 11186 13082
rect 11186 13030 11198 13082
rect 11198 13030 11212 13082
rect 11236 13030 11250 13082
rect 11250 13030 11262 13082
rect 11262 13030 11292 13082
rect 11316 13030 11326 13082
rect 11326 13030 11372 13082
rect 11076 13028 11132 13030
rect 11156 13028 11212 13030
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 8576 6010 8632 6012
rect 8656 6010 8712 6012
rect 8736 6010 8792 6012
rect 8816 6010 8872 6012
rect 8576 5958 8622 6010
rect 8622 5958 8632 6010
rect 8656 5958 8686 6010
rect 8686 5958 8698 6010
rect 8698 5958 8712 6010
rect 8736 5958 8750 6010
rect 8750 5958 8762 6010
rect 8762 5958 8792 6010
rect 8816 5958 8826 6010
rect 8826 5958 8872 6010
rect 8576 5956 8632 5958
rect 8656 5956 8712 5958
rect 8736 5956 8792 5958
rect 8816 5956 8872 5958
rect 8576 4922 8632 4924
rect 8656 4922 8712 4924
rect 8736 4922 8792 4924
rect 8816 4922 8872 4924
rect 8576 4870 8622 4922
rect 8622 4870 8632 4922
rect 8656 4870 8686 4922
rect 8686 4870 8698 4922
rect 8698 4870 8712 4922
rect 8736 4870 8750 4922
rect 8750 4870 8762 4922
rect 8762 4870 8792 4922
rect 8816 4870 8826 4922
rect 8826 4870 8872 4922
rect 8576 4868 8632 4870
rect 8656 4868 8712 4870
rect 8736 4868 8792 4870
rect 8816 4868 8872 4870
rect 6076 1114 6132 1116
rect 6156 1114 6212 1116
rect 6236 1114 6292 1116
rect 6316 1114 6372 1116
rect 6076 1062 6122 1114
rect 6122 1062 6132 1114
rect 6156 1062 6186 1114
rect 6186 1062 6198 1114
rect 6198 1062 6212 1114
rect 6236 1062 6250 1114
rect 6250 1062 6262 1114
rect 6262 1062 6292 1114
rect 6316 1062 6326 1114
rect 6326 1062 6372 1114
rect 6076 1060 6132 1062
rect 6156 1060 6212 1062
rect 6236 1060 6292 1062
rect 6316 1060 6372 1062
rect 8298 2916 8354 2952
rect 8298 2896 8300 2916
rect 8300 2896 8352 2916
rect 8352 2896 8354 2916
rect 8576 3834 8632 3836
rect 8656 3834 8712 3836
rect 8736 3834 8792 3836
rect 8816 3834 8872 3836
rect 8576 3782 8622 3834
rect 8622 3782 8632 3834
rect 8656 3782 8686 3834
rect 8686 3782 8698 3834
rect 8698 3782 8712 3834
rect 8736 3782 8750 3834
rect 8750 3782 8762 3834
rect 8762 3782 8792 3834
rect 8816 3782 8826 3834
rect 8826 3782 8872 3834
rect 8576 3780 8632 3782
rect 8656 3780 8712 3782
rect 8736 3780 8792 3782
rect 8816 3780 8872 3782
rect 8576 2746 8632 2748
rect 8656 2746 8712 2748
rect 8736 2746 8792 2748
rect 8816 2746 8872 2748
rect 8576 2694 8622 2746
rect 8622 2694 8632 2746
rect 8656 2694 8686 2746
rect 8686 2694 8698 2746
rect 8698 2694 8712 2746
rect 8736 2694 8750 2746
rect 8750 2694 8762 2746
rect 8762 2694 8792 2746
rect 8816 2694 8826 2746
rect 8826 2694 8872 2746
rect 8576 2692 8632 2694
rect 8656 2692 8712 2694
rect 8736 2692 8792 2694
rect 8816 2692 8872 2694
rect 10414 3576 10470 3632
rect 11076 11994 11132 11996
rect 11156 11994 11212 11996
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11076 11942 11122 11994
rect 11122 11942 11132 11994
rect 11156 11942 11186 11994
rect 11186 11942 11198 11994
rect 11198 11942 11212 11994
rect 11236 11942 11250 11994
rect 11250 11942 11262 11994
rect 11262 11942 11292 11994
rect 11316 11942 11326 11994
rect 11326 11942 11372 11994
rect 11076 11940 11132 11942
rect 11156 11940 11212 11942
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 12714 12844 12770 12880
rect 12714 12824 12716 12844
rect 12716 12824 12768 12844
rect 12768 12824 12770 12844
rect 11076 10906 11132 10908
rect 11156 10906 11212 10908
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11076 10854 11122 10906
rect 11122 10854 11132 10906
rect 11156 10854 11186 10906
rect 11186 10854 11198 10906
rect 11198 10854 11212 10906
rect 11236 10854 11250 10906
rect 11250 10854 11262 10906
rect 11262 10854 11292 10906
rect 11316 10854 11326 10906
rect 11326 10854 11372 10906
rect 11076 10852 11132 10854
rect 11156 10852 11212 10854
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11076 9818 11132 9820
rect 11156 9818 11212 9820
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11076 9766 11122 9818
rect 11122 9766 11132 9818
rect 11156 9766 11186 9818
rect 11186 9766 11198 9818
rect 11198 9766 11212 9818
rect 11236 9766 11250 9818
rect 11250 9766 11262 9818
rect 11262 9766 11292 9818
rect 11316 9766 11326 9818
rect 11326 9766 11372 9818
rect 11076 9764 11132 9766
rect 11156 9764 11212 9766
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 13266 10512 13322 10568
rect 13576 21242 13632 21244
rect 13656 21242 13712 21244
rect 13736 21242 13792 21244
rect 13816 21242 13872 21244
rect 13576 21190 13622 21242
rect 13622 21190 13632 21242
rect 13656 21190 13686 21242
rect 13686 21190 13698 21242
rect 13698 21190 13712 21242
rect 13736 21190 13750 21242
rect 13750 21190 13762 21242
rect 13762 21190 13792 21242
rect 13816 21190 13826 21242
rect 13826 21190 13872 21242
rect 13576 21188 13632 21190
rect 13656 21188 13712 21190
rect 13736 21188 13792 21190
rect 13816 21188 13872 21190
rect 14002 21140 14058 21176
rect 14002 21120 14004 21140
rect 14004 21120 14056 21140
rect 14056 21120 14058 21140
rect 13576 20154 13632 20156
rect 13656 20154 13712 20156
rect 13736 20154 13792 20156
rect 13816 20154 13872 20156
rect 13576 20102 13622 20154
rect 13622 20102 13632 20154
rect 13656 20102 13686 20154
rect 13686 20102 13698 20154
rect 13698 20102 13712 20154
rect 13736 20102 13750 20154
rect 13750 20102 13762 20154
rect 13762 20102 13792 20154
rect 13816 20102 13826 20154
rect 13826 20102 13872 20154
rect 13576 20100 13632 20102
rect 13656 20100 13712 20102
rect 13736 20100 13792 20102
rect 13816 20100 13872 20102
rect 13576 19066 13632 19068
rect 13656 19066 13712 19068
rect 13736 19066 13792 19068
rect 13816 19066 13872 19068
rect 13576 19014 13622 19066
rect 13622 19014 13632 19066
rect 13656 19014 13686 19066
rect 13686 19014 13698 19066
rect 13698 19014 13712 19066
rect 13736 19014 13750 19066
rect 13750 19014 13762 19066
rect 13762 19014 13792 19066
rect 13816 19014 13826 19066
rect 13826 19014 13872 19066
rect 13576 19012 13632 19014
rect 13656 19012 13712 19014
rect 13736 19012 13792 19014
rect 13816 19012 13872 19014
rect 14002 18808 14058 18864
rect 13576 17978 13632 17980
rect 13656 17978 13712 17980
rect 13736 17978 13792 17980
rect 13816 17978 13872 17980
rect 13576 17926 13622 17978
rect 13622 17926 13632 17978
rect 13656 17926 13686 17978
rect 13686 17926 13698 17978
rect 13698 17926 13712 17978
rect 13736 17926 13750 17978
rect 13750 17926 13762 17978
rect 13762 17926 13792 17978
rect 13816 17926 13826 17978
rect 13826 17926 13872 17978
rect 13576 17924 13632 17926
rect 13656 17924 13712 17926
rect 13736 17924 13792 17926
rect 13816 17924 13872 17926
rect 13576 16890 13632 16892
rect 13656 16890 13712 16892
rect 13736 16890 13792 16892
rect 13816 16890 13872 16892
rect 13576 16838 13622 16890
rect 13622 16838 13632 16890
rect 13656 16838 13686 16890
rect 13686 16838 13698 16890
rect 13698 16838 13712 16890
rect 13736 16838 13750 16890
rect 13750 16838 13762 16890
rect 13762 16838 13792 16890
rect 13816 16838 13826 16890
rect 13826 16838 13872 16890
rect 13576 16836 13632 16838
rect 13656 16836 13712 16838
rect 13736 16836 13792 16838
rect 13816 16836 13872 16838
rect 13576 15802 13632 15804
rect 13656 15802 13712 15804
rect 13736 15802 13792 15804
rect 13816 15802 13872 15804
rect 13576 15750 13622 15802
rect 13622 15750 13632 15802
rect 13656 15750 13686 15802
rect 13686 15750 13698 15802
rect 13698 15750 13712 15802
rect 13736 15750 13750 15802
rect 13750 15750 13762 15802
rect 13762 15750 13792 15802
rect 13816 15750 13826 15802
rect 13826 15750 13872 15802
rect 13576 15748 13632 15750
rect 13656 15748 13712 15750
rect 13736 15748 13792 15750
rect 13816 15748 13872 15750
rect 14278 21256 14334 21312
rect 14278 20440 14334 20496
rect 14462 20476 14464 20496
rect 14464 20476 14516 20496
rect 14516 20476 14518 20496
rect 14462 20440 14518 20476
rect 14186 20032 14242 20088
rect 13576 14714 13632 14716
rect 13656 14714 13712 14716
rect 13736 14714 13792 14716
rect 13816 14714 13872 14716
rect 13576 14662 13622 14714
rect 13622 14662 13632 14714
rect 13656 14662 13686 14714
rect 13686 14662 13698 14714
rect 13698 14662 13712 14714
rect 13736 14662 13750 14714
rect 13750 14662 13762 14714
rect 13762 14662 13792 14714
rect 13816 14662 13826 14714
rect 13826 14662 13872 14714
rect 13576 14660 13632 14662
rect 13656 14660 13712 14662
rect 13736 14660 13792 14662
rect 13816 14660 13872 14662
rect 13634 13776 13690 13832
rect 13576 13626 13632 13628
rect 13656 13626 13712 13628
rect 13736 13626 13792 13628
rect 13816 13626 13872 13628
rect 13576 13574 13622 13626
rect 13622 13574 13632 13626
rect 13656 13574 13686 13626
rect 13686 13574 13698 13626
rect 13698 13574 13712 13626
rect 13736 13574 13750 13626
rect 13750 13574 13762 13626
rect 13762 13574 13792 13626
rect 13816 13574 13826 13626
rect 13826 13574 13872 13626
rect 13576 13572 13632 13574
rect 13656 13572 13712 13574
rect 13736 13572 13792 13574
rect 13816 13572 13872 13574
rect 13576 12538 13632 12540
rect 13656 12538 13712 12540
rect 13736 12538 13792 12540
rect 13816 12538 13872 12540
rect 13576 12486 13622 12538
rect 13622 12486 13632 12538
rect 13656 12486 13686 12538
rect 13686 12486 13698 12538
rect 13698 12486 13712 12538
rect 13736 12486 13750 12538
rect 13750 12486 13762 12538
rect 13762 12486 13792 12538
rect 13816 12486 13826 12538
rect 13826 12486 13872 12538
rect 13576 12484 13632 12486
rect 13656 12484 13712 12486
rect 13736 12484 13792 12486
rect 13816 12484 13872 12486
rect 14278 13776 14334 13832
rect 13576 11450 13632 11452
rect 13656 11450 13712 11452
rect 13736 11450 13792 11452
rect 13816 11450 13872 11452
rect 13576 11398 13622 11450
rect 13622 11398 13632 11450
rect 13656 11398 13686 11450
rect 13686 11398 13698 11450
rect 13698 11398 13712 11450
rect 13736 11398 13750 11450
rect 13750 11398 13762 11450
rect 13762 11398 13792 11450
rect 13816 11398 13826 11450
rect 13826 11398 13872 11450
rect 13576 11396 13632 11398
rect 13656 11396 13712 11398
rect 13736 11396 13792 11398
rect 13816 11396 13872 11398
rect 13726 10920 13782 10976
rect 13576 10362 13632 10364
rect 13656 10362 13712 10364
rect 13736 10362 13792 10364
rect 13816 10362 13872 10364
rect 13576 10310 13622 10362
rect 13622 10310 13632 10362
rect 13656 10310 13686 10362
rect 13686 10310 13698 10362
rect 13698 10310 13712 10362
rect 13736 10310 13750 10362
rect 13750 10310 13762 10362
rect 13762 10310 13792 10362
rect 13816 10310 13826 10362
rect 13826 10310 13872 10362
rect 13576 10308 13632 10310
rect 13656 10308 13712 10310
rect 13736 10308 13792 10310
rect 13816 10308 13872 10310
rect 11242 9152 11298 9208
rect 11076 8730 11132 8732
rect 11156 8730 11212 8732
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11076 8678 11122 8730
rect 11122 8678 11132 8730
rect 11156 8678 11186 8730
rect 11186 8678 11198 8730
rect 11198 8678 11212 8730
rect 11236 8678 11250 8730
rect 11250 8678 11262 8730
rect 11262 8678 11292 8730
rect 11316 8678 11326 8730
rect 11326 8678 11372 8730
rect 11076 8676 11132 8678
rect 11156 8676 11212 8678
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11978 8880 12034 8936
rect 11076 7642 11132 7644
rect 11156 7642 11212 7644
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11076 7590 11122 7642
rect 11122 7590 11132 7642
rect 11156 7590 11186 7642
rect 11186 7590 11198 7642
rect 11198 7590 11212 7642
rect 11236 7590 11250 7642
rect 11250 7590 11262 7642
rect 11262 7590 11292 7642
rect 11316 7590 11326 7642
rect 11326 7590 11372 7642
rect 11076 7588 11132 7590
rect 11156 7588 11212 7590
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 13266 9152 13322 9208
rect 13082 9016 13138 9072
rect 17130 22516 17132 22536
rect 17132 22516 17184 22536
rect 17184 22516 17186 22536
rect 17130 22480 17186 22516
rect 21076 22874 21132 22876
rect 21156 22874 21212 22876
rect 21236 22874 21292 22876
rect 21316 22874 21372 22876
rect 21076 22822 21122 22874
rect 21122 22822 21132 22874
rect 21156 22822 21186 22874
rect 21186 22822 21198 22874
rect 21198 22822 21212 22874
rect 21236 22822 21250 22874
rect 21250 22822 21262 22874
rect 21262 22822 21292 22874
rect 21316 22822 21326 22874
rect 21326 22822 21372 22874
rect 21076 22820 21132 22822
rect 21156 22820 21212 22822
rect 21236 22820 21292 22822
rect 21316 22820 21372 22822
rect 17958 22480 18014 22536
rect 18576 22330 18632 22332
rect 18656 22330 18712 22332
rect 18736 22330 18792 22332
rect 18816 22330 18872 22332
rect 18576 22278 18622 22330
rect 18622 22278 18632 22330
rect 18656 22278 18686 22330
rect 18686 22278 18698 22330
rect 18698 22278 18712 22330
rect 18736 22278 18750 22330
rect 18750 22278 18762 22330
rect 18762 22278 18792 22330
rect 18816 22278 18826 22330
rect 18826 22278 18872 22330
rect 18576 22276 18632 22278
rect 18656 22276 18712 22278
rect 18736 22276 18792 22278
rect 18816 22276 18872 22278
rect 16076 21786 16132 21788
rect 16156 21786 16212 21788
rect 16236 21786 16292 21788
rect 16316 21786 16372 21788
rect 16076 21734 16122 21786
rect 16122 21734 16132 21786
rect 16156 21734 16186 21786
rect 16186 21734 16198 21786
rect 16198 21734 16212 21786
rect 16236 21734 16250 21786
rect 16250 21734 16262 21786
rect 16262 21734 16292 21786
rect 16316 21734 16326 21786
rect 16326 21734 16372 21786
rect 16076 21732 16132 21734
rect 16156 21732 16212 21734
rect 16236 21732 16292 21734
rect 16316 21732 16372 21734
rect 15290 20848 15346 20904
rect 14922 20168 14978 20224
rect 15750 20440 15806 20496
rect 16302 20848 16358 20904
rect 16486 20884 16488 20904
rect 16488 20884 16540 20904
rect 16540 20884 16542 20904
rect 16486 20848 16542 20884
rect 16076 20698 16132 20700
rect 16156 20698 16212 20700
rect 16236 20698 16292 20700
rect 16316 20698 16372 20700
rect 16076 20646 16122 20698
rect 16122 20646 16132 20698
rect 16156 20646 16186 20698
rect 16186 20646 16198 20698
rect 16198 20646 16212 20698
rect 16236 20646 16250 20698
rect 16250 20646 16262 20698
rect 16262 20646 16292 20698
rect 16316 20646 16326 20698
rect 16326 20646 16372 20698
rect 16076 20644 16132 20646
rect 16156 20644 16212 20646
rect 16236 20644 16292 20646
rect 16316 20644 16372 20646
rect 16578 20440 16634 20496
rect 15290 18128 15346 18184
rect 16076 19610 16132 19612
rect 16156 19610 16212 19612
rect 16236 19610 16292 19612
rect 16316 19610 16372 19612
rect 16076 19558 16122 19610
rect 16122 19558 16132 19610
rect 16156 19558 16186 19610
rect 16186 19558 16198 19610
rect 16198 19558 16212 19610
rect 16236 19558 16250 19610
rect 16250 19558 16262 19610
rect 16262 19558 16292 19610
rect 16316 19558 16326 19610
rect 16326 19558 16372 19610
rect 16076 19556 16132 19558
rect 16156 19556 16212 19558
rect 16236 19556 16292 19558
rect 16316 19556 16372 19558
rect 16076 18522 16132 18524
rect 16156 18522 16212 18524
rect 16236 18522 16292 18524
rect 16316 18522 16372 18524
rect 16076 18470 16122 18522
rect 16122 18470 16132 18522
rect 16156 18470 16186 18522
rect 16186 18470 16198 18522
rect 16198 18470 16212 18522
rect 16236 18470 16250 18522
rect 16250 18470 16262 18522
rect 16262 18470 16292 18522
rect 16316 18470 16326 18522
rect 16326 18470 16372 18522
rect 16076 18468 16132 18470
rect 16156 18468 16212 18470
rect 16236 18468 16292 18470
rect 16316 18468 16372 18470
rect 16946 20460 17002 20496
rect 16946 20440 16948 20460
rect 16948 20440 17000 20460
rect 17000 20440 17002 20460
rect 16670 20032 16726 20088
rect 17314 21392 17370 21448
rect 17130 20712 17186 20768
rect 17498 21256 17554 21312
rect 17406 20868 17462 20904
rect 17406 20848 17408 20868
rect 17408 20848 17460 20868
rect 17460 20848 17462 20868
rect 18326 21956 18382 21992
rect 18326 21936 18328 21956
rect 18328 21936 18380 21956
rect 18380 21936 18382 21956
rect 17866 20984 17922 21040
rect 17498 20712 17554 20768
rect 17038 20168 17094 20224
rect 16486 18284 16542 18320
rect 16486 18264 16488 18284
rect 16488 18264 16540 18284
rect 16540 18264 16542 18284
rect 16578 17992 16634 18048
rect 16394 17856 16450 17912
rect 16394 17720 16450 17776
rect 16076 17434 16132 17436
rect 16156 17434 16212 17436
rect 16236 17434 16292 17436
rect 16316 17434 16372 17436
rect 16076 17382 16122 17434
rect 16122 17382 16132 17434
rect 16156 17382 16186 17434
rect 16186 17382 16198 17434
rect 16198 17382 16212 17434
rect 16236 17382 16250 17434
rect 16250 17382 16262 17434
rect 16262 17382 16292 17434
rect 16316 17382 16326 17434
rect 16326 17382 16372 17434
rect 16076 17380 16132 17382
rect 16156 17380 16212 17382
rect 16236 17380 16292 17382
rect 16316 17380 16372 17382
rect 14738 15408 14794 15464
rect 15198 15408 15254 15464
rect 13576 9274 13632 9276
rect 13656 9274 13712 9276
rect 13736 9274 13792 9276
rect 13816 9274 13872 9276
rect 13576 9222 13622 9274
rect 13622 9222 13632 9274
rect 13656 9222 13686 9274
rect 13686 9222 13698 9274
rect 13698 9222 13712 9274
rect 13736 9222 13750 9274
rect 13750 9222 13762 9274
rect 13762 9222 13792 9274
rect 13816 9222 13826 9274
rect 13826 9222 13872 9274
rect 13576 9220 13632 9222
rect 13656 9220 13712 9222
rect 13736 9220 13792 9222
rect 13816 9220 13872 9222
rect 13542 9016 13598 9072
rect 13818 8880 13874 8936
rect 13576 8186 13632 8188
rect 13656 8186 13712 8188
rect 13736 8186 13792 8188
rect 13816 8186 13872 8188
rect 13576 8134 13622 8186
rect 13622 8134 13632 8186
rect 13656 8134 13686 8186
rect 13686 8134 13698 8186
rect 13698 8134 13712 8186
rect 13736 8134 13750 8186
rect 13750 8134 13762 8186
rect 13762 8134 13792 8186
rect 13816 8134 13826 8186
rect 13826 8134 13872 8186
rect 13576 8132 13632 8134
rect 13656 8132 13712 8134
rect 13736 8132 13792 8134
rect 13816 8132 13872 8134
rect 15106 10920 15162 10976
rect 16076 16346 16132 16348
rect 16156 16346 16212 16348
rect 16236 16346 16292 16348
rect 16316 16346 16372 16348
rect 16076 16294 16122 16346
rect 16122 16294 16132 16346
rect 16156 16294 16186 16346
rect 16186 16294 16198 16346
rect 16198 16294 16212 16346
rect 16236 16294 16250 16346
rect 16250 16294 16262 16346
rect 16262 16294 16292 16346
rect 16316 16294 16326 16346
rect 16326 16294 16372 16346
rect 16076 16292 16132 16294
rect 16156 16292 16212 16294
rect 16236 16292 16292 16294
rect 16316 16292 16372 16294
rect 16210 16088 16266 16144
rect 16076 15258 16132 15260
rect 16156 15258 16212 15260
rect 16236 15258 16292 15260
rect 16316 15258 16372 15260
rect 16076 15206 16122 15258
rect 16122 15206 16132 15258
rect 16156 15206 16186 15258
rect 16186 15206 16198 15258
rect 16198 15206 16212 15258
rect 16236 15206 16250 15258
rect 16250 15206 16262 15258
rect 16262 15206 16292 15258
rect 16316 15206 16326 15258
rect 16326 15206 16372 15258
rect 16076 15204 16132 15206
rect 16156 15204 16212 15206
rect 16236 15204 16292 15206
rect 16316 15204 16372 15206
rect 16302 15000 16358 15056
rect 17222 19896 17278 19952
rect 17590 19916 17646 19952
rect 17590 19896 17592 19916
rect 17592 19896 17644 19916
rect 17644 19896 17646 19916
rect 17222 19352 17278 19408
rect 17038 18264 17094 18320
rect 17130 18128 17186 18184
rect 17314 18028 17316 18048
rect 17316 18028 17368 18048
rect 17368 18028 17370 18048
rect 17314 17992 17370 18028
rect 16076 14170 16132 14172
rect 16156 14170 16212 14172
rect 16236 14170 16292 14172
rect 16316 14170 16372 14172
rect 16076 14118 16122 14170
rect 16122 14118 16132 14170
rect 16156 14118 16186 14170
rect 16186 14118 16198 14170
rect 16198 14118 16212 14170
rect 16236 14118 16250 14170
rect 16250 14118 16262 14170
rect 16262 14118 16292 14170
rect 16316 14118 16326 14170
rect 16326 14118 16372 14170
rect 16076 14116 16132 14118
rect 16156 14116 16212 14118
rect 16236 14116 16292 14118
rect 16316 14116 16372 14118
rect 17498 18128 17554 18184
rect 18142 21392 18198 21448
rect 18576 21242 18632 21244
rect 18656 21242 18712 21244
rect 18736 21242 18792 21244
rect 18816 21242 18872 21244
rect 18576 21190 18622 21242
rect 18622 21190 18632 21242
rect 18656 21190 18686 21242
rect 18686 21190 18698 21242
rect 18698 21190 18712 21242
rect 18736 21190 18750 21242
rect 18750 21190 18762 21242
rect 18762 21190 18792 21242
rect 18816 21190 18826 21242
rect 18826 21190 18872 21242
rect 18576 21188 18632 21190
rect 18656 21188 18712 21190
rect 18736 21188 18792 21190
rect 18816 21188 18872 21190
rect 18234 21120 18290 21176
rect 18970 21120 19026 21176
rect 19062 20984 19118 21040
rect 18050 20848 18106 20904
rect 18234 20848 18290 20904
rect 18576 20154 18632 20156
rect 18656 20154 18712 20156
rect 18736 20154 18792 20156
rect 18816 20154 18872 20156
rect 18576 20102 18622 20154
rect 18622 20102 18632 20154
rect 18656 20102 18686 20154
rect 18686 20102 18698 20154
rect 18698 20102 18712 20154
rect 18736 20102 18750 20154
rect 18750 20102 18762 20154
rect 18762 20102 18792 20154
rect 18816 20102 18826 20154
rect 18826 20102 18872 20154
rect 18576 20100 18632 20102
rect 18656 20100 18712 20102
rect 18736 20100 18792 20102
rect 18816 20100 18872 20102
rect 18326 19624 18382 19680
rect 17774 18128 17830 18184
rect 17958 18672 18014 18728
rect 17958 18284 18014 18320
rect 17958 18264 17960 18284
rect 17960 18264 18012 18284
rect 18012 18264 18014 18284
rect 17958 17876 18014 17912
rect 17958 17856 17960 17876
rect 17960 17856 18012 17876
rect 18012 17856 18014 17876
rect 19798 21936 19854 21992
rect 19522 21664 19578 21720
rect 19062 19624 19118 19680
rect 19522 21020 19524 21040
rect 19524 21020 19576 21040
rect 19576 21020 19578 21040
rect 19522 20984 19578 21020
rect 19430 19896 19486 19952
rect 18576 19066 18632 19068
rect 18656 19066 18712 19068
rect 18736 19066 18792 19068
rect 18816 19066 18872 19068
rect 18576 19014 18622 19066
rect 18622 19014 18632 19066
rect 18656 19014 18686 19066
rect 18686 19014 18698 19066
rect 18698 19014 18712 19066
rect 18736 19014 18750 19066
rect 18750 19014 18762 19066
rect 18762 19014 18792 19066
rect 18816 19014 18826 19066
rect 18826 19014 18872 19066
rect 18576 19012 18632 19014
rect 18656 19012 18712 19014
rect 18736 19012 18792 19014
rect 18816 19012 18872 19014
rect 18576 17978 18632 17980
rect 18656 17978 18712 17980
rect 18736 17978 18792 17980
rect 18816 17978 18872 17980
rect 18576 17926 18622 17978
rect 18622 17926 18632 17978
rect 18656 17926 18686 17978
rect 18686 17926 18698 17978
rect 18698 17926 18712 17978
rect 18736 17926 18750 17978
rect 18750 17926 18762 17978
rect 18762 17926 18792 17978
rect 18816 17926 18826 17978
rect 18826 17926 18872 17978
rect 18576 17924 18632 17926
rect 18656 17924 18712 17926
rect 18736 17924 18792 17926
rect 18816 17924 18872 17926
rect 18234 17720 18290 17776
rect 16026 13232 16082 13288
rect 16076 13082 16132 13084
rect 16156 13082 16212 13084
rect 16236 13082 16292 13084
rect 16316 13082 16372 13084
rect 16076 13030 16122 13082
rect 16122 13030 16132 13082
rect 16156 13030 16186 13082
rect 16186 13030 16198 13082
rect 16198 13030 16212 13082
rect 16236 13030 16250 13082
rect 16250 13030 16262 13082
rect 16262 13030 16292 13082
rect 16316 13030 16326 13082
rect 16326 13030 16372 13082
rect 16076 13028 16132 13030
rect 16156 13028 16212 13030
rect 16236 13028 16292 13030
rect 16316 13028 16372 13030
rect 16076 11994 16132 11996
rect 16156 11994 16212 11996
rect 16236 11994 16292 11996
rect 16316 11994 16372 11996
rect 16076 11942 16122 11994
rect 16122 11942 16132 11994
rect 16156 11942 16186 11994
rect 16186 11942 16198 11994
rect 16198 11942 16212 11994
rect 16236 11942 16250 11994
rect 16250 11942 16262 11994
rect 16262 11942 16292 11994
rect 16316 11942 16326 11994
rect 16326 11942 16372 11994
rect 16076 11940 16132 11942
rect 16156 11940 16212 11942
rect 16236 11940 16292 11942
rect 16316 11940 16372 11942
rect 16076 10906 16132 10908
rect 16156 10906 16212 10908
rect 16236 10906 16292 10908
rect 16316 10906 16372 10908
rect 16076 10854 16122 10906
rect 16122 10854 16132 10906
rect 16156 10854 16186 10906
rect 16186 10854 16198 10906
rect 16198 10854 16212 10906
rect 16236 10854 16250 10906
rect 16250 10854 16262 10906
rect 16262 10854 16292 10906
rect 16316 10854 16326 10906
rect 16326 10854 16372 10906
rect 16076 10852 16132 10854
rect 16156 10852 16212 10854
rect 16236 10852 16292 10854
rect 16316 10852 16372 10854
rect 17406 12316 17408 12336
rect 17408 12316 17460 12336
rect 17460 12316 17462 12336
rect 17406 12280 17462 12316
rect 18576 16890 18632 16892
rect 18656 16890 18712 16892
rect 18736 16890 18792 16892
rect 18816 16890 18872 16892
rect 18576 16838 18622 16890
rect 18622 16838 18632 16890
rect 18656 16838 18686 16890
rect 18686 16838 18698 16890
rect 18698 16838 18712 16890
rect 18736 16838 18750 16890
rect 18750 16838 18762 16890
rect 18762 16838 18792 16890
rect 18816 16838 18826 16890
rect 18826 16838 18872 16890
rect 18576 16836 18632 16838
rect 18656 16836 18712 16838
rect 18736 16836 18792 16838
rect 18816 16836 18872 16838
rect 19062 18672 19118 18728
rect 19430 18672 19486 18728
rect 18970 16496 19026 16552
rect 18234 16088 18290 16144
rect 18576 15802 18632 15804
rect 18656 15802 18712 15804
rect 18736 15802 18792 15804
rect 18816 15802 18872 15804
rect 18576 15750 18622 15802
rect 18622 15750 18632 15802
rect 18656 15750 18686 15802
rect 18686 15750 18698 15802
rect 18698 15750 18712 15802
rect 18736 15750 18750 15802
rect 18750 15750 18762 15802
rect 18762 15750 18792 15802
rect 18816 15750 18826 15802
rect 18826 15750 18872 15802
rect 18576 15748 18632 15750
rect 18656 15748 18712 15750
rect 18736 15748 18792 15750
rect 18816 15748 18872 15750
rect 18576 14714 18632 14716
rect 18656 14714 18712 14716
rect 18736 14714 18792 14716
rect 18816 14714 18872 14716
rect 18576 14662 18622 14714
rect 18622 14662 18632 14714
rect 18656 14662 18686 14714
rect 18686 14662 18698 14714
rect 18698 14662 18712 14714
rect 18736 14662 18750 14714
rect 18750 14662 18762 14714
rect 18762 14662 18792 14714
rect 18816 14662 18826 14714
rect 18826 14662 18872 14714
rect 18576 14660 18632 14662
rect 18656 14660 18712 14662
rect 18736 14660 18792 14662
rect 18816 14660 18872 14662
rect 18970 14456 19026 14512
rect 20258 21800 20314 21856
rect 19798 20712 19854 20768
rect 20258 21392 20314 21448
rect 20074 20440 20130 20496
rect 19706 19624 19762 19680
rect 20074 19896 20130 19952
rect 20258 18944 20314 19000
rect 21076 21786 21132 21788
rect 21156 21786 21212 21788
rect 21236 21786 21292 21788
rect 21316 21786 21372 21788
rect 21076 21734 21122 21786
rect 21122 21734 21132 21786
rect 21156 21734 21186 21786
rect 21186 21734 21198 21786
rect 21198 21734 21212 21786
rect 21236 21734 21250 21786
rect 21250 21734 21262 21786
rect 21262 21734 21292 21786
rect 21316 21734 21326 21786
rect 21326 21734 21372 21786
rect 21076 21732 21132 21734
rect 21156 21732 21212 21734
rect 21236 21732 21292 21734
rect 21316 21732 21372 21734
rect 21178 21120 21234 21176
rect 21076 20698 21132 20700
rect 21156 20698 21212 20700
rect 21236 20698 21292 20700
rect 21316 20698 21372 20700
rect 21076 20646 21122 20698
rect 21122 20646 21132 20698
rect 21156 20646 21186 20698
rect 21186 20646 21198 20698
rect 21198 20646 21212 20698
rect 21236 20646 21250 20698
rect 21250 20646 21262 20698
rect 21262 20646 21292 20698
rect 21316 20646 21326 20698
rect 21326 20646 21372 20698
rect 21076 20644 21132 20646
rect 21156 20644 21212 20646
rect 21236 20644 21292 20646
rect 21316 20644 21372 20646
rect 21638 21120 21694 21176
rect 20534 19624 20590 19680
rect 19338 16904 19394 16960
rect 19798 17584 19854 17640
rect 19706 17312 19762 17368
rect 16076 9818 16132 9820
rect 16156 9818 16212 9820
rect 16236 9818 16292 9820
rect 16316 9818 16372 9820
rect 16076 9766 16122 9818
rect 16122 9766 16132 9818
rect 16156 9766 16186 9818
rect 16186 9766 16198 9818
rect 16198 9766 16212 9818
rect 16236 9766 16250 9818
rect 16250 9766 16262 9818
rect 16262 9766 16292 9818
rect 16316 9766 16326 9818
rect 16326 9766 16372 9818
rect 16076 9764 16132 9766
rect 16156 9764 16212 9766
rect 16236 9764 16292 9766
rect 16316 9764 16372 9766
rect 17682 12144 17738 12200
rect 15842 8880 15898 8936
rect 11076 6554 11132 6556
rect 11156 6554 11212 6556
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11076 6502 11122 6554
rect 11122 6502 11132 6554
rect 11156 6502 11186 6554
rect 11186 6502 11198 6554
rect 11198 6502 11212 6554
rect 11236 6502 11250 6554
rect 11250 6502 11262 6554
rect 11262 6502 11292 6554
rect 11316 6502 11326 6554
rect 11326 6502 11372 6554
rect 11076 6500 11132 6502
rect 11156 6500 11212 6502
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11076 5466 11132 5468
rect 11156 5466 11212 5468
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11076 5414 11122 5466
rect 11122 5414 11132 5466
rect 11156 5414 11186 5466
rect 11186 5414 11198 5466
rect 11198 5414 11212 5466
rect 11236 5414 11250 5466
rect 11250 5414 11262 5466
rect 11262 5414 11292 5466
rect 11316 5414 11326 5466
rect 11326 5414 11372 5466
rect 11076 5412 11132 5414
rect 11156 5412 11212 5414
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11076 4378 11132 4380
rect 11156 4378 11212 4380
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11076 4326 11122 4378
rect 11122 4326 11132 4378
rect 11156 4326 11186 4378
rect 11186 4326 11198 4378
rect 11198 4326 11212 4378
rect 11236 4326 11250 4378
rect 11250 4326 11262 4378
rect 11262 4326 11292 4378
rect 11316 4326 11326 4378
rect 11326 4326 11372 4378
rect 11076 4324 11132 4326
rect 11156 4324 11212 4326
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 8576 1658 8632 1660
rect 8656 1658 8712 1660
rect 8736 1658 8792 1660
rect 8816 1658 8872 1660
rect 8576 1606 8622 1658
rect 8622 1606 8632 1658
rect 8656 1606 8686 1658
rect 8686 1606 8698 1658
rect 8698 1606 8712 1658
rect 8736 1606 8750 1658
rect 8750 1606 8762 1658
rect 8762 1606 8792 1658
rect 8816 1606 8826 1658
rect 8826 1606 8872 1658
rect 8576 1604 8632 1606
rect 8656 1604 8712 1606
rect 8736 1604 8792 1606
rect 8816 1604 8872 1606
rect 11076 3290 11132 3292
rect 11156 3290 11212 3292
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11076 3238 11122 3290
rect 11122 3238 11132 3290
rect 11156 3238 11186 3290
rect 11186 3238 11198 3290
rect 11198 3238 11212 3290
rect 11236 3238 11250 3290
rect 11250 3238 11262 3290
rect 11262 3238 11292 3290
rect 11316 3238 11326 3290
rect 11326 3238 11372 3290
rect 11076 3236 11132 3238
rect 11156 3236 11212 3238
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11334 3052 11390 3088
rect 11334 3032 11336 3052
rect 11336 3032 11388 3052
rect 11388 3032 11390 3052
rect 11076 2202 11132 2204
rect 11156 2202 11212 2204
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11076 2150 11122 2202
rect 11122 2150 11132 2202
rect 11156 2150 11186 2202
rect 11186 2150 11198 2202
rect 11198 2150 11212 2202
rect 11236 2150 11250 2202
rect 11250 2150 11262 2202
rect 11262 2150 11292 2202
rect 11316 2150 11326 2202
rect 11326 2150 11372 2202
rect 11076 2148 11132 2150
rect 11156 2148 11212 2150
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 13576 7098 13632 7100
rect 13656 7098 13712 7100
rect 13736 7098 13792 7100
rect 13816 7098 13872 7100
rect 13576 7046 13622 7098
rect 13622 7046 13632 7098
rect 13656 7046 13686 7098
rect 13686 7046 13698 7098
rect 13698 7046 13712 7098
rect 13736 7046 13750 7098
rect 13750 7046 13762 7098
rect 13762 7046 13792 7098
rect 13816 7046 13826 7098
rect 13826 7046 13872 7098
rect 13576 7044 13632 7046
rect 13656 7044 13712 7046
rect 13736 7044 13792 7046
rect 13816 7044 13872 7046
rect 16076 8730 16132 8732
rect 16156 8730 16212 8732
rect 16236 8730 16292 8732
rect 16316 8730 16372 8732
rect 16076 8678 16122 8730
rect 16122 8678 16132 8730
rect 16156 8678 16186 8730
rect 16186 8678 16198 8730
rect 16198 8678 16212 8730
rect 16236 8678 16250 8730
rect 16250 8678 16262 8730
rect 16262 8678 16292 8730
rect 16316 8678 16326 8730
rect 16326 8678 16372 8730
rect 16076 8676 16132 8678
rect 16156 8676 16212 8678
rect 16236 8676 16292 8678
rect 16316 8676 16372 8678
rect 18576 13626 18632 13628
rect 18656 13626 18712 13628
rect 18736 13626 18792 13628
rect 18816 13626 18872 13628
rect 18576 13574 18622 13626
rect 18622 13574 18632 13626
rect 18656 13574 18686 13626
rect 18686 13574 18698 13626
rect 18698 13574 18712 13626
rect 18736 13574 18750 13626
rect 18750 13574 18762 13626
rect 18762 13574 18792 13626
rect 18816 13574 18826 13626
rect 18826 13574 18872 13626
rect 18576 13572 18632 13574
rect 18656 13572 18712 13574
rect 18736 13572 18792 13574
rect 18816 13572 18872 13574
rect 18576 12538 18632 12540
rect 18656 12538 18712 12540
rect 18736 12538 18792 12540
rect 18816 12538 18872 12540
rect 18576 12486 18622 12538
rect 18622 12486 18632 12538
rect 18656 12486 18686 12538
rect 18686 12486 18698 12538
rect 18698 12486 18712 12538
rect 18736 12486 18750 12538
rect 18750 12486 18762 12538
rect 18762 12486 18792 12538
rect 18816 12486 18826 12538
rect 18826 12486 18872 12538
rect 18576 12484 18632 12486
rect 18656 12484 18712 12486
rect 18736 12484 18792 12486
rect 18816 12484 18872 12486
rect 20994 19916 21050 19952
rect 20994 19896 20996 19916
rect 20996 19896 21048 19916
rect 21048 19896 21050 19916
rect 21076 19610 21132 19612
rect 21156 19610 21212 19612
rect 21236 19610 21292 19612
rect 21316 19610 21372 19612
rect 21076 19558 21122 19610
rect 21122 19558 21132 19610
rect 21156 19558 21186 19610
rect 21186 19558 21198 19610
rect 21198 19558 21212 19610
rect 21236 19558 21250 19610
rect 21250 19558 21262 19610
rect 21262 19558 21292 19610
rect 21316 19558 21326 19610
rect 21326 19558 21372 19610
rect 21076 19556 21132 19558
rect 21156 19556 21212 19558
rect 21236 19556 21292 19558
rect 21316 19556 21372 19558
rect 21178 18944 21234 19000
rect 21076 18522 21132 18524
rect 21156 18522 21212 18524
rect 21236 18522 21292 18524
rect 21316 18522 21372 18524
rect 21076 18470 21122 18522
rect 21122 18470 21132 18522
rect 21156 18470 21186 18522
rect 21186 18470 21198 18522
rect 21198 18470 21212 18522
rect 21236 18470 21250 18522
rect 21250 18470 21262 18522
rect 21262 18470 21292 18522
rect 21316 18470 21326 18522
rect 21326 18470 21372 18522
rect 21076 18468 21132 18470
rect 21156 18468 21212 18470
rect 21236 18468 21292 18470
rect 21316 18468 21372 18470
rect 20442 17332 20498 17368
rect 20442 17312 20444 17332
rect 20444 17312 20496 17332
rect 20496 17312 20498 17332
rect 19890 16904 19946 16960
rect 21076 17434 21132 17436
rect 21156 17434 21212 17436
rect 21236 17434 21292 17436
rect 21316 17434 21372 17436
rect 21076 17382 21122 17434
rect 21122 17382 21132 17434
rect 21156 17382 21186 17434
rect 21186 17382 21198 17434
rect 21198 17382 21212 17434
rect 21236 17382 21250 17434
rect 21250 17382 21262 17434
rect 21262 17382 21292 17434
rect 21316 17382 21326 17434
rect 21326 17382 21372 17434
rect 21076 17380 21132 17382
rect 21156 17380 21212 17382
rect 21236 17380 21292 17382
rect 21316 17380 21372 17382
rect 20902 17060 20958 17096
rect 20902 17040 20904 17060
rect 20904 17040 20956 17060
rect 20956 17040 20958 17060
rect 20534 16904 20590 16960
rect 19798 13232 19854 13288
rect 18694 12044 18696 12064
rect 18696 12044 18748 12064
rect 18748 12044 18750 12064
rect 18694 12008 18750 12044
rect 18576 11450 18632 11452
rect 18656 11450 18712 11452
rect 18736 11450 18792 11452
rect 18816 11450 18872 11452
rect 18576 11398 18622 11450
rect 18622 11398 18632 11450
rect 18656 11398 18686 11450
rect 18686 11398 18698 11450
rect 18698 11398 18712 11450
rect 18736 11398 18750 11450
rect 18750 11398 18762 11450
rect 18762 11398 18792 11450
rect 18816 11398 18826 11450
rect 18826 11398 18872 11450
rect 18576 11396 18632 11398
rect 18656 11396 18712 11398
rect 18736 11396 18792 11398
rect 18816 11396 18872 11398
rect 19154 12164 19210 12200
rect 19154 12144 19156 12164
rect 19156 12144 19208 12164
rect 19208 12144 19210 12164
rect 19430 11736 19486 11792
rect 20166 13368 20222 13424
rect 20166 12844 20222 12880
rect 20166 12824 20168 12844
rect 20168 12824 20220 12844
rect 20220 12824 20222 12844
rect 20166 12416 20222 12472
rect 19982 11620 20038 11656
rect 19982 11600 19984 11620
rect 19984 11600 20036 11620
rect 20036 11600 20038 11620
rect 21076 16346 21132 16348
rect 21156 16346 21212 16348
rect 21236 16346 21292 16348
rect 21316 16346 21372 16348
rect 21076 16294 21122 16346
rect 21122 16294 21132 16346
rect 21156 16294 21186 16346
rect 21186 16294 21198 16346
rect 21198 16294 21212 16346
rect 21236 16294 21250 16346
rect 21250 16294 21262 16346
rect 21262 16294 21292 16346
rect 21316 16294 21326 16346
rect 21326 16294 21372 16346
rect 21076 16292 21132 16294
rect 21156 16292 21212 16294
rect 21236 16292 21292 16294
rect 21316 16292 21372 16294
rect 21076 15258 21132 15260
rect 21156 15258 21212 15260
rect 21236 15258 21292 15260
rect 21316 15258 21372 15260
rect 21076 15206 21122 15258
rect 21122 15206 21132 15258
rect 21156 15206 21186 15258
rect 21186 15206 21198 15258
rect 21198 15206 21212 15258
rect 21236 15206 21250 15258
rect 21250 15206 21262 15258
rect 21262 15206 21292 15258
rect 21316 15206 21326 15258
rect 21326 15206 21372 15258
rect 21076 15204 21132 15206
rect 21156 15204 21212 15206
rect 21236 15204 21292 15206
rect 21316 15204 21372 15206
rect 20442 12280 20498 12336
rect 21730 16632 21786 16688
rect 21076 14170 21132 14172
rect 21156 14170 21212 14172
rect 21236 14170 21292 14172
rect 21316 14170 21372 14172
rect 21076 14118 21122 14170
rect 21122 14118 21132 14170
rect 21156 14118 21186 14170
rect 21186 14118 21198 14170
rect 21198 14118 21212 14170
rect 21236 14118 21250 14170
rect 21250 14118 21262 14170
rect 21262 14118 21292 14170
rect 21316 14118 21326 14170
rect 21326 14118 21372 14170
rect 21076 14116 21132 14118
rect 21156 14116 21212 14118
rect 21236 14116 21292 14118
rect 21316 14116 21372 14118
rect 20810 13368 20866 13424
rect 21546 13912 21602 13968
rect 21076 13082 21132 13084
rect 21156 13082 21212 13084
rect 21236 13082 21292 13084
rect 21316 13082 21372 13084
rect 21076 13030 21122 13082
rect 21122 13030 21132 13082
rect 21156 13030 21186 13082
rect 21186 13030 21198 13082
rect 21198 13030 21212 13082
rect 21236 13030 21250 13082
rect 21250 13030 21262 13082
rect 21262 13030 21292 13082
rect 21316 13030 21326 13082
rect 21326 13030 21372 13082
rect 21076 13028 21132 13030
rect 21156 13028 21212 13030
rect 21236 13028 21292 13030
rect 21316 13028 21372 13030
rect 20626 12044 20628 12064
rect 20628 12044 20680 12064
rect 20680 12044 20682 12064
rect 20626 12008 20682 12044
rect 19062 11192 19118 11248
rect 18576 10362 18632 10364
rect 18656 10362 18712 10364
rect 18736 10362 18792 10364
rect 18816 10362 18872 10364
rect 18576 10310 18622 10362
rect 18622 10310 18632 10362
rect 18656 10310 18686 10362
rect 18686 10310 18698 10362
rect 18698 10310 18712 10362
rect 18736 10310 18750 10362
rect 18750 10310 18762 10362
rect 18762 10310 18792 10362
rect 18816 10310 18826 10362
rect 18826 10310 18872 10362
rect 18576 10308 18632 10310
rect 18656 10308 18712 10310
rect 18736 10308 18792 10310
rect 18816 10308 18872 10310
rect 16076 7642 16132 7644
rect 16156 7642 16212 7644
rect 16236 7642 16292 7644
rect 16316 7642 16372 7644
rect 16076 7590 16122 7642
rect 16122 7590 16132 7642
rect 16156 7590 16186 7642
rect 16186 7590 16198 7642
rect 16198 7590 16212 7642
rect 16236 7590 16250 7642
rect 16250 7590 16262 7642
rect 16262 7590 16292 7642
rect 16316 7590 16326 7642
rect 16326 7590 16372 7642
rect 16076 7588 16132 7590
rect 16156 7588 16212 7590
rect 16236 7588 16292 7590
rect 16316 7588 16372 7590
rect 13358 6296 13414 6352
rect 13634 6180 13690 6216
rect 13634 6160 13636 6180
rect 13636 6160 13688 6180
rect 13688 6160 13690 6180
rect 13576 6010 13632 6012
rect 13656 6010 13712 6012
rect 13736 6010 13792 6012
rect 13816 6010 13872 6012
rect 13576 5958 13622 6010
rect 13622 5958 13632 6010
rect 13656 5958 13686 6010
rect 13686 5958 13698 6010
rect 13698 5958 13712 6010
rect 13736 5958 13750 6010
rect 13750 5958 13762 6010
rect 13762 5958 13792 6010
rect 13816 5958 13826 6010
rect 13826 5958 13872 6010
rect 13576 5956 13632 5958
rect 13656 5956 13712 5958
rect 13736 5956 13792 5958
rect 13816 5956 13872 5958
rect 13726 5228 13782 5264
rect 13726 5208 13728 5228
rect 13728 5208 13780 5228
rect 13780 5208 13782 5228
rect 14002 5092 14058 5128
rect 14002 5072 14004 5092
rect 14004 5072 14056 5092
rect 14056 5072 14058 5092
rect 13576 4922 13632 4924
rect 13656 4922 13712 4924
rect 13736 4922 13792 4924
rect 13816 4922 13872 4924
rect 13576 4870 13622 4922
rect 13622 4870 13632 4922
rect 13656 4870 13686 4922
rect 13686 4870 13698 4922
rect 13698 4870 13712 4922
rect 13736 4870 13750 4922
rect 13750 4870 13762 4922
rect 13762 4870 13792 4922
rect 13816 4870 13826 4922
rect 13826 4870 13872 4922
rect 13576 4868 13632 4870
rect 13656 4868 13712 4870
rect 13736 4868 13792 4870
rect 13816 4868 13872 4870
rect 14462 5888 14518 5944
rect 14278 5752 14334 5808
rect 13576 3834 13632 3836
rect 13656 3834 13712 3836
rect 13736 3834 13792 3836
rect 13816 3834 13872 3836
rect 13576 3782 13622 3834
rect 13622 3782 13632 3834
rect 13656 3782 13686 3834
rect 13686 3782 13698 3834
rect 13698 3782 13712 3834
rect 13736 3782 13750 3834
rect 13750 3782 13762 3834
rect 13762 3782 13792 3834
rect 13816 3782 13826 3834
rect 13826 3782 13872 3834
rect 13576 3780 13632 3782
rect 13656 3780 13712 3782
rect 13736 3780 13792 3782
rect 13816 3780 13872 3782
rect 14462 5636 14518 5672
rect 14462 5616 14464 5636
rect 14464 5616 14516 5636
rect 14516 5616 14518 5636
rect 14830 4120 14886 4176
rect 16076 6554 16132 6556
rect 16156 6554 16212 6556
rect 16236 6554 16292 6556
rect 16316 6554 16372 6556
rect 16076 6502 16122 6554
rect 16122 6502 16132 6554
rect 16156 6502 16186 6554
rect 16186 6502 16198 6554
rect 16198 6502 16212 6554
rect 16236 6502 16250 6554
rect 16250 6502 16262 6554
rect 16262 6502 16292 6554
rect 16316 6502 16326 6554
rect 16326 6502 16372 6554
rect 16076 6500 16132 6502
rect 16156 6500 16212 6502
rect 16236 6500 16292 6502
rect 16316 6500 16372 6502
rect 18576 9274 18632 9276
rect 18656 9274 18712 9276
rect 18736 9274 18792 9276
rect 18816 9274 18872 9276
rect 18576 9222 18622 9274
rect 18622 9222 18632 9274
rect 18656 9222 18686 9274
rect 18686 9222 18698 9274
rect 18698 9222 18712 9274
rect 18736 9222 18750 9274
rect 18750 9222 18762 9274
rect 18762 9222 18792 9274
rect 18816 9222 18826 9274
rect 18826 9222 18872 9274
rect 18576 9220 18632 9222
rect 18656 9220 18712 9222
rect 18736 9220 18792 9222
rect 18816 9220 18872 9222
rect 18576 8186 18632 8188
rect 18656 8186 18712 8188
rect 18736 8186 18792 8188
rect 18816 8186 18872 8188
rect 18576 8134 18622 8186
rect 18622 8134 18632 8186
rect 18656 8134 18686 8186
rect 18686 8134 18698 8186
rect 18698 8134 18712 8186
rect 18736 8134 18750 8186
rect 18750 8134 18762 8186
rect 18762 8134 18792 8186
rect 18816 8134 18826 8186
rect 18826 8134 18872 8186
rect 18576 8132 18632 8134
rect 18656 8132 18712 8134
rect 18736 8132 18792 8134
rect 18816 8132 18872 8134
rect 18576 7098 18632 7100
rect 18656 7098 18712 7100
rect 18736 7098 18792 7100
rect 18816 7098 18872 7100
rect 18576 7046 18622 7098
rect 18622 7046 18632 7098
rect 18656 7046 18686 7098
rect 18686 7046 18698 7098
rect 18698 7046 18712 7098
rect 18736 7046 18750 7098
rect 18750 7046 18762 7098
rect 18762 7046 18792 7098
rect 18816 7046 18826 7098
rect 18826 7046 18872 7098
rect 18576 7044 18632 7046
rect 18656 7044 18712 7046
rect 18736 7044 18792 7046
rect 18816 7044 18872 7046
rect 16118 6024 16174 6080
rect 16854 6024 16910 6080
rect 16076 5466 16132 5468
rect 16156 5466 16212 5468
rect 16236 5466 16292 5468
rect 16316 5466 16372 5468
rect 16076 5414 16122 5466
rect 16122 5414 16132 5466
rect 16156 5414 16186 5466
rect 16186 5414 16198 5466
rect 16198 5414 16212 5466
rect 16236 5414 16250 5466
rect 16250 5414 16262 5466
rect 16262 5414 16292 5466
rect 16316 5414 16326 5466
rect 16326 5414 16372 5466
rect 16076 5412 16132 5414
rect 16156 5412 16212 5414
rect 16236 5412 16292 5414
rect 16316 5412 16372 5414
rect 13576 2746 13632 2748
rect 13656 2746 13712 2748
rect 13736 2746 13792 2748
rect 13816 2746 13872 2748
rect 13576 2694 13622 2746
rect 13622 2694 13632 2746
rect 13656 2694 13686 2746
rect 13686 2694 13698 2746
rect 13698 2694 13712 2746
rect 13736 2694 13750 2746
rect 13750 2694 13762 2746
rect 13762 2694 13792 2746
rect 13816 2694 13826 2746
rect 13826 2694 13872 2746
rect 13576 2692 13632 2694
rect 13656 2692 13712 2694
rect 13736 2692 13792 2694
rect 13816 2692 13872 2694
rect 17774 5908 17830 5944
rect 17774 5888 17776 5908
rect 17776 5888 17828 5908
rect 17828 5888 17830 5908
rect 16486 4664 16542 4720
rect 16394 4528 16450 4584
rect 16076 4378 16132 4380
rect 16156 4378 16212 4380
rect 16236 4378 16292 4380
rect 16316 4378 16372 4380
rect 16076 4326 16122 4378
rect 16122 4326 16132 4378
rect 16156 4326 16186 4378
rect 16186 4326 16198 4378
rect 16198 4326 16212 4378
rect 16236 4326 16250 4378
rect 16250 4326 16262 4378
rect 16262 4326 16292 4378
rect 16316 4326 16326 4378
rect 16326 4326 16372 4378
rect 16076 4324 16132 4326
rect 16156 4324 16212 4326
rect 16236 4324 16292 4326
rect 16316 4324 16372 4326
rect 17222 5480 17278 5536
rect 16076 3290 16132 3292
rect 16156 3290 16212 3292
rect 16236 3290 16292 3292
rect 16316 3290 16372 3292
rect 16076 3238 16122 3290
rect 16122 3238 16132 3290
rect 16156 3238 16186 3290
rect 16186 3238 16198 3290
rect 16198 3238 16212 3290
rect 16236 3238 16250 3290
rect 16250 3238 16262 3290
rect 16262 3238 16292 3290
rect 16316 3238 16326 3290
rect 16326 3238 16372 3290
rect 16076 3236 16132 3238
rect 16156 3236 16212 3238
rect 16236 3236 16292 3238
rect 16316 3236 16372 3238
rect 16394 2896 16450 2952
rect 13576 1658 13632 1660
rect 13656 1658 13712 1660
rect 13736 1658 13792 1660
rect 13816 1658 13872 1660
rect 13576 1606 13622 1658
rect 13622 1606 13632 1658
rect 13656 1606 13686 1658
rect 13686 1606 13698 1658
rect 13698 1606 13712 1658
rect 13736 1606 13750 1658
rect 13750 1606 13762 1658
rect 13762 1606 13792 1658
rect 13816 1606 13826 1658
rect 13826 1606 13872 1658
rect 13576 1604 13632 1606
rect 13656 1604 13712 1606
rect 13736 1604 13792 1606
rect 13816 1604 13872 1606
rect 11076 1114 11132 1116
rect 11156 1114 11212 1116
rect 11236 1114 11292 1116
rect 11316 1114 11372 1116
rect 11076 1062 11122 1114
rect 11122 1062 11132 1114
rect 11156 1062 11186 1114
rect 11186 1062 11198 1114
rect 11198 1062 11212 1114
rect 11236 1062 11250 1114
rect 11250 1062 11262 1114
rect 11262 1062 11292 1114
rect 11316 1062 11326 1114
rect 11326 1062 11372 1114
rect 11076 1060 11132 1062
rect 11156 1060 11212 1062
rect 11236 1060 11292 1062
rect 11316 1060 11372 1062
rect 16076 2202 16132 2204
rect 16156 2202 16212 2204
rect 16236 2202 16292 2204
rect 16316 2202 16372 2204
rect 16076 2150 16122 2202
rect 16122 2150 16132 2202
rect 16156 2150 16186 2202
rect 16186 2150 16198 2202
rect 16198 2150 16212 2202
rect 16236 2150 16250 2202
rect 16250 2150 16262 2202
rect 16262 2150 16292 2202
rect 16316 2150 16326 2202
rect 16326 2150 16372 2202
rect 16076 2148 16132 2150
rect 16156 2148 16212 2150
rect 16236 2148 16292 2150
rect 16316 2148 16372 2150
rect 18576 6010 18632 6012
rect 18656 6010 18712 6012
rect 18736 6010 18792 6012
rect 18816 6010 18872 6012
rect 18576 5958 18622 6010
rect 18622 5958 18632 6010
rect 18656 5958 18686 6010
rect 18686 5958 18698 6010
rect 18698 5958 18712 6010
rect 18736 5958 18750 6010
rect 18750 5958 18762 6010
rect 18762 5958 18792 6010
rect 18816 5958 18826 6010
rect 18826 5958 18872 6010
rect 18576 5956 18632 5958
rect 18656 5956 18712 5958
rect 18736 5956 18792 5958
rect 18816 5956 18872 5958
rect 19062 6024 19118 6080
rect 18576 4922 18632 4924
rect 18656 4922 18712 4924
rect 18736 4922 18792 4924
rect 18816 4922 18872 4924
rect 18576 4870 18622 4922
rect 18622 4870 18632 4922
rect 18656 4870 18686 4922
rect 18686 4870 18698 4922
rect 18698 4870 18712 4922
rect 18736 4870 18750 4922
rect 18750 4870 18762 4922
rect 18762 4870 18792 4922
rect 18816 4870 18826 4922
rect 18826 4870 18872 4922
rect 18576 4868 18632 4870
rect 18656 4868 18712 4870
rect 18736 4868 18792 4870
rect 18816 4868 18872 4870
rect 18576 3834 18632 3836
rect 18656 3834 18712 3836
rect 18736 3834 18792 3836
rect 18816 3834 18872 3836
rect 18576 3782 18622 3834
rect 18622 3782 18632 3834
rect 18656 3782 18686 3834
rect 18686 3782 18698 3834
rect 18698 3782 18712 3834
rect 18736 3782 18750 3834
rect 18750 3782 18762 3834
rect 18762 3782 18792 3834
rect 18816 3782 18826 3834
rect 18826 3782 18872 3834
rect 18576 3780 18632 3782
rect 18656 3780 18712 3782
rect 18736 3780 18792 3782
rect 18816 3780 18872 3782
rect 19154 4020 19156 4040
rect 19156 4020 19208 4040
rect 19208 4020 19210 4040
rect 19154 3984 19210 4020
rect 18576 2746 18632 2748
rect 18656 2746 18712 2748
rect 18736 2746 18792 2748
rect 18816 2746 18872 2748
rect 18576 2694 18622 2746
rect 18622 2694 18632 2746
rect 18656 2694 18686 2746
rect 18686 2694 18698 2746
rect 18698 2694 18712 2746
rect 18736 2694 18750 2746
rect 18750 2694 18762 2746
rect 18762 2694 18792 2746
rect 18816 2694 18826 2746
rect 18826 2694 18872 2746
rect 18576 2692 18632 2694
rect 18656 2692 18712 2694
rect 18736 2692 18792 2694
rect 18816 2692 18872 2694
rect 16076 1114 16132 1116
rect 16156 1114 16212 1116
rect 16236 1114 16292 1116
rect 16316 1114 16372 1116
rect 16076 1062 16122 1114
rect 16122 1062 16132 1114
rect 16156 1062 16186 1114
rect 16186 1062 16198 1114
rect 16198 1062 16212 1114
rect 16236 1062 16250 1114
rect 16250 1062 16262 1114
rect 16262 1062 16292 1114
rect 16316 1062 16326 1114
rect 16326 1062 16372 1114
rect 16076 1060 16132 1062
rect 16156 1060 16212 1062
rect 16236 1060 16292 1062
rect 16316 1060 16372 1062
rect 21076 11994 21132 11996
rect 21156 11994 21212 11996
rect 21236 11994 21292 11996
rect 21316 11994 21372 11996
rect 21076 11942 21122 11994
rect 21122 11942 21132 11994
rect 21156 11942 21186 11994
rect 21186 11942 21198 11994
rect 21198 11942 21212 11994
rect 21236 11942 21250 11994
rect 21250 11942 21262 11994
rect 21262 11942 21292 11994
rect 21316 11942 21326 11994
rect 21326 11942 21372 11994
rect 21076 11940 21132 11942
rect 21156 11940 21212 11942
rect 21236 11940 21292 11942
rect 21316 11940 21372 11942
rect 21076 10906 21132 10908
rect 21156 10906 21212 10908
rect 21236 10906 21292 10908
rect 21316 10906 21372 10908
rect 21076 10854 21122 10906
rect 21122 10854 21132 10906
rect 21156 10854 21186 10906
rect 21186 10854 21198 10906
rect 21198 10854 21212 10906
rect 21236 10854 21250 10906
rect 21250 10854 21262 10906
rect 21262 10854 21292 10906
rect 21316 10854 21326 10906
rect 21326 10854 21372 10906
rect 21076 10852 21132 10854
rect 21156 10852 21212 10854
rect 21236 10852 21292 10854
rect 21316 10852 21372 10854
rect 21076 9818 21132 9820
rect 21156 9818 21212 9820
rect 21236 9818 21292 9820
rect 21316 9818 21372 9820
rect 21076 9766 21122 9818
rect 21122 9766 21132 9818
rect 21156 9766 21186 9818
rect 21186 9766 21198 9818
rect 21198 9766 21212 9818
rect 21236 9766 21250 9818
rect 21250 9766 21262 9818
rect 21262 9766 21292 9818
rect 21316 9766 21326 9818
rect 21326 9766 21372 9818
rect 21076 9764 21132 9766
rect 21156 9764 21212 9766
rect 21236 9764 21292 9766
rect 21316 9764 21372 9766
rect 22098 20440 22154 20496
rect 22374 20712 22430 20768
rect 23576 22330 23632 22332
rect 23656 22330 23712 22332
rect 23736 22330 23792 22332
rect 23816 22330 23872 22332
rect 23576 22278 23622 22330
rect 23622 22278 23632 22330
rect 23656 22278 23686 22330
rect 23686 22278 23698 22330
rect 23698 22278 23712 22330
rect 23736 22278 23750 22330
rect 23750 22278 23762 22330
rect 23762 22278 23792 22330
rect 23816 22278 23826 22330
rect 23826 22278 23872 22330
rect 23576 22276 23632 22278
rect 23656 22276 23712 22278
rect 23736 22276 23792 22278
rect 23816 22276 23872 22278
rect 23294 21528 23350 21584
rect 23018 21392 23074 21448
rect 23018 20848 23074 20904
rect 23386 21392 23442 21448
rect 23662 21528 23718 21584
rect 23576 21242 23632 21244
rect 23656 21242 23712 21244
rect 23736 21242 23792 21244
rect 23816 21242 23872 21244
rect 23576 21190 23622 21242
rect 23622 21190 23632 21242
rect 23656 21190 23686 21242
rect 23686 21190 23698 21242
rect 23698 21190 23712 21242
rect 23736 21190 23750 21242
rect 23750 21190 23762 21242
rect 23762 21190 23792 21242
rect 23816 21190 23826 21242
rect 23826 21190 23872 21242
rect 23576 21188 23632 21190
rect 23656 21188 23712 21190
rect 23736 21188 23792 21190
rect 23816 21188 23872 21190
rect 23294 20712 23350 20768
rect 26076 22874 26132 22876
rect 26156 22874 26212 22876
rect 26236 22874 26292 22876
rect 26316 22874 26372 22876
rect 26076 22822 26122 22874
rect 26122 22822 26132 22874
rect 26156 22822 26186 22874
rect 26186 22822 26198 22874
rect 26198 22822 26212 22874
rect 26236 22822 26250 22874
rect 26250 22822 26262 22874
rect 26262 22822 26292 22874
rect 26316 22822 26326 22874
rect 26326 22822 26372 22874
rect 26076 22820 26132 22822
rect 26156 22820 26212 22822
rect 26236 22820 26292 22822
rect 26316 22820 26372 22822
rect 25594 22072 25650 22128
rect 24858 20712 24914 20768
rect 25686 21664 25742 21720
rect 25686 21120 25742 21176
rect 26076 21786 26132 21788
rect 26156 21786 26212 21788
rect 26236 21786 26292 21788
rect 26316 21786 26372 21788
rect 26076 21734 26122 21786
rect 26122 21734 26132 21786
rect 26156 21734 26186 21786
rect 26186 21734 26198 21786
rect 26198 21734 26212 21786
rect 26236 21734 26250 21786
rect 26250 21734 26262 21786
rect 26262 21734 26292 21786
rect 26316 21734 26326 21786
rect 26326 21734 26372 21786
rect 26076 21732 26132 21734
rect 26156 21732 26212 21734
rect 26236 21732 26292 21734
rect 26316 21732 26372 21734
rect 23576 20154 23632 20156
rect 23656 20154 23712 20156
rect 23736 20154 23792 20156
rect 23816 20154 23872 20156
rect 23576 20102 23622 20154
rect 23622 20102 23632 20154
rect 23656 20102 23686 20154
rect 23686 20102 23698 20154
rect 23698 20102 23712 20154
rect 23736 20102 23750 20154
rect 23750 20102 23762 20154
rect 23762 20102 23792 20154
rect 23816 20102 23826 20154
rect 23826 20102 23872 20154
rect 23576 20100 23632 20102
rect 23656 20100 23712 20102
rect 23736 20100 23792 20102
rect 23816 20100 23872 20102
rect 23202 18400 23258 18456
rect 23576 19066 23632 19068
rect 23656 19066 23712 19068
rect 23736 19066 23792 19068
rect 23816 19066 23872 19068
rect 23576 19014 23622 19066
rect 23622 19014 23632 19066
rect 23656 19014 23686 19066
rect 23686 19014 23698 19066
rect 23698 19014 23712 19066
rect 23736 19014 23750 19066
rect 23750 19014 23762 19066
rect 23762 19014 23792 19066
rect 23816 19014 23826 19066
rect 23826 19014 23872 19066
rect 23576 19012 23632 19014
rect 23656 19012 23712 19014
rect 23736 19012 23792 19014
rect 23816 19012 23872 19014
rect 23938 18400 23994 18456
rect 23576 17978 23632 17980
rect 23656 17978 23712 17980
rect 23736 17978 23792 17980
rect 23816 17978 23872 17980
rect 23576 17926 23622 17978
rect 23622 17926 23632 17978
rect 23656 17926 23686 17978
rect 23686 17926 23698 17978
rect 23698 17926 23712 17978
rect 23736 17926 23750 17978
rect 23750 17926 23762 17978
rect 23762 17926 23792 17978
rect 23816 17926 23826 17978
rect 23826 17926 23872 17978
rect 23576 17924 23632 17926
rect 23656 17924 23712 17926
rect 23736 17924 23792 17926
rect 23816 17924 23872 17926
rect 22558 15952 22614 16008
rect 21914 13388 21970 13424
rect 21914 13368 21916 13388
rect 21916 13368 21968 13388
rect 21968 13368 21970 13388
rect 22282 12960 22338 13016
rect 23576 16890 23632 16892
rect 23656 16890 23712 16892
rect 23736 16890 23792 16892
rect 23816 16890 23872 16892
rect 23576 16838 23622 16890
rect 23622 16838 23632 16890
rect 23656 16838 23686 16890
rect 23686 16838 23698 16890
rect 23698 16838 23712 16890
rect 23736 16838 23750 16890
rect 23750 16838 23762 16890
rect 23762 16838 23792 16890
rect 23816 16838 23826 16890
rect 23826 16838 23872 16890
rect 23576 16836 23632 16838
rect 23656 16836 23712 16838
rect 23736 16836 23792 16838
rect 23816 16836 23872 16838
rect 23754 16496 23810 16552
rect 23576 15802 23632 15804
rect 23656 15802 23712 15804
rect 23736 15802 23792 15804
rect 23816 15802 23872 15804
rect 23576 15750 23622 15802
rect 23622 15750 23632 15802
rect 23656 15750 23686 15802
rect 23686 15750 23698 15802
rect 23698 15750 23712 15802
rect 23736 15750 23750 15802
rect 23750 15750 23762 15802
rect 23762 15750 23792 15802
rect 23816 15750 23826 15802
rect 23826 15750 23872 15802
rect 23576 15748 23632 15750
rect 23656 15748 23712 15750
rect 23736 15748 23792 15750
rect 23816 15748 23872 15750
rect 26698 21392 26754 21448
rect 24858 19896 24914 19952
rect 23386 14456 23442 14512
rect 23938 15544 23994 15600
rect 24214 15000 24270 15056
rect 23576 14714 23632 14716
rect 23656 14714 23712 14716
rect 23736 14714 23792 14716
rect 23816 14714 23872 14716
rect 23576 14662 23622 14714
rect 23622 14662 23632 14714
rect 23656 14662 23686 14714
rect 23686 14662 23698 14714
rect 23698 14662 23712 14714
rect 23736 14662 23750 14714
rect 23750 14662 23762 14714
rect 23762 14662 23792 14714
rect 23816 14662 23826 14714
rect 23826 14662 23872 14714
rect 23576 14660 23632 14662
rect 23656 14660 23712 14662
rect 23736 14660 23792 14662
rect 23816 14660 23872 14662
rect 23294 12960 23350 13016
rect 23576 13626 23632 13628
rect 23656 13626 23712 13628
rect 23736 13626 23792 13628
rect 23816 13626 23872 13628
rect 23576 13574 23622 13626
rect 23622 13574 23632 13626
rect 23656 13574 23686 13626
rect 23686 13574 23698 13626
rect 23698 13574 23712 13626
rect 23736 13574 23750 13626
rect 23750 13574 23762 13626
rect 23762 13574 23792 13626
rect 23816 13574 23826 13626
rect 23826 13574 23872 13626
rect 23576 13572 23632 13574
rect 23656 13572 23712 13574
rect 23736 13572 23792 13574
rect 23816 13572 23872 13574
rect 23846 13268 23848 13288
rect 23848 13268 23900 13288
rect 23900 13268 23902 13288
rect 23846 13232 23902 13268
rect 23846 12824 23902 12880
rect 23576 12538 23632 12540
rect 23656 12538 23712 12540
rect 23736 12538 23792 12540
rect 23816 12538 23872 12540
rect 23576 12486 23622 12538
rect 23622 12486 23632 12538
rect 23656 12486 23686 12538
rect 23686 12486 23698 12538
rect 23698 12486 23712 12538
rect 23736 12486 23750 12538
rect 23750 12486 23762 12538
rect 23762 12486 23792 12538
rect 23816 12486 23826 12538
rect 23826 12486 23872 12538
rect 23576 12484 23632 12486
rect 23656 12484 23712 12486
rect 23736 12484 23792 12486
rect 23816 12484 23872 12486
rect 24582 14612 24638 14648
rect 24582 14592 24584 14612
rect 24584 14592 24636 14612
rect 24636 14592 24638 14612
rect 24858 18284 24914 18320
rect 24858 18264 24860 18284
rect 24860 18264 24912 18284
rect 24912 18264 24914 18284
rect 24582 13096 24638 13152
rect 23576 11450 23632 11452
rect 23656 11450 23712 11452
rect 23736 11450 23792 11452
rect 23816 11450 23872 11452
rect 23576 11398 23622 11450
rect 23622 11398 23632 11450
rect 23656 11398 23686 11450
rect 23686 11398 23698 11450
rect 23698 11398 23712 11450
rect 23736 11398 23750 11450
rect 23750 11398 23762 11450
rect 23762 11398 23792 11450
rect 23816 11398 23826 11450
rect 23826 11398 23872 11450
rect 23576 11396 23632 11398
rect 23656 11396 23712 11398
rect 23736 11396 23792 11398
rect 23816 11396 23872 11398
rect 21178 9444 21234 9480
rect 21178 9424 21180 9444
rect 21180 9424 21232 9444
rect 21232 9424 21234 9444
rect 21076 8730 21132 8732
rect 21156 8730 21212 8732
rect 21236 8730 21292 8732
rect 21316 8730 21372 8732
rect 21076 8678 21122 8730
rect 21122 8678 21132 8730
rect 21156 8678 21186 8730
rect 21186 8678 21198 8730
rect 21198 8678 21212 8730
rect 21236 8678 21250 8730
rect 21250 8678 21262 8730
rect 21262 8678 21292 8730
rect 21316 8678 21326 8730
rect 21326 8678 21372 8730
rect 21076 8676 21132 8678
rect 21156 8676 21212 8678
rect 21236 8676 21292 8678
rect 21316 8676 21372 8678
rect 19798 6840 19854 6896
rect 19614 4800 19670 4856
rect 19890 5480 19946 5536
rect 19890 4664 19946 4720
rect 19430 3168 19486 3224
rect 19246 2352 19302 2408
rect 18576 1658 18632 1660
rect 18656 1658 18712 1660
rect 18736 1658 18792 1660
rect 18816 1658 18872 1660
rect 18576 1606 18622 1658
rect 18622 1606 18632 1658
rect 18656 1606 18686 1658
rect 18686 1606 18698 1658
rect 18698 1606 18712 1658
rect 18736 1606 18750 1658
rect 18750 1606 18762 1658
rect 18762 1606 18792 1658
rect 18816 1606 18826 1658
rect 18826 1606 18872 1658
rect 18576 1604 18632 1606
rect 18656 1604 18712 1606
rect 18736 1604 18792 1606
rect 18816 1604 18872 1606
rect 22006 9016 22062 9072
rect 21546 8336 21602 8392
rect 21076 7642 21132 7644
rect 21156 7642 21212 7644
rect 21236 7642 21292 7644
rect 21316 7642 21372 7644
rect 21076 7590 21122 7642
rect 21122 7590 21132 7642
rect 21156 7590 21186 7642
rect 21186 7590 21198 7642
rect 21198 7590 21212 7642
rect 21236 7590 21250 7642
rect 21250 7590 21262 7642
rect 21262 7590 21292 7642
rect 21316 7590 21326 7642
rect 21326 7590 21372 7642
rect 21076 7588 21132 7590
rect 21156 7588 21212 7590
rect 21236 7588 21292 7590
rect 21316 7588 21372 7590
rect 20902 6432 20958 6488
rect 21076 6554 21132 6556
rect 21156 6554 21212 6556
rect 21236 6554 21292 6556
rect 21316 6554 21372 6556
rect 21076 6502 21122 6554
rect 21122 6502 21132 6554
rect 21156 6502 21186 6554
rect 21186 6502 21198 6554
rect 21198 6502 21212 6554
rect 21236 6502 21250 6554
rect 21250 6502 21262 6554
rect 21262 6502 21292 6554
rect 21316 6502 21326 6554
rect 21326 6502 21372 6554
rect 21076 6500 21132 6502
rect 21156 6500 21212 6502
rect 21236 6500 21292 6502
rect 21316 6500 21372 6502
rect 20810 5344 20866 5400
rect 21076 5466 21132 5468
rect 21156 5466 21212 5468
rect 21236 5466 21292 5468
rect 21316 5466 21372 5468
rect 21076 5414 21122 5466
rect 21122 5414 21132 5466
rect 21156 5414 21186 5466
rect 21186 5414 21198 5466
rect 21198 5414 21212 5466
rect 21236 5414 21250 5466
rect 21250 5414 21262 5466
rect 21262 5414 21292 5466
rect 21316 5414 21326 5466
rect 21326 5414 21372 5466
rect 21076 5412 21132 5414
rect 21156 5412 21212 5414
rect 21236 5412 21292 5414
rect 21316 5412 21372 5414
rect 21454 4528 21510 4584
rect 21076 4378 21132 4380
rect 21156 4378 21212 4380
rect 21236 4378 21292 4380
rect 21316 4378 21372 4380
rect 21076 4326 21122 4378
rect 21122 4326 21132 4378
rect 21156 4326 21186 4378
rect 21186 4326 21198 4378
rect 21198 4326 21212 4378
rect 21236 4326 21250 4378
rect 21250 4326 21262 4378
rect 21262 4326 21292 4378
rect 21316 4326 21326 4378
rect 21326 4326 21372 4378
rect 21076 4324 21132 4326
rect 21156 4324 21212 4326
rect 21236 4324 21292 4326
rect 21316 4324 21372 4326
rect 20350 3984 20406 4040
rect 22834 9832 22890 9888
rect 23576 10362 23632 10364
rect 23656 10362 23712 10364
rect 23736 10362 23792 10364
rect 23816 10362 23872 10364
rect 23576 10310 23622 10362
rect 23622 10310 23632 10362
rect 23656 10310 23686 10362
rect 23686 10310 23698 10362
rect 23698 10310 23712 10362
rect 23736 10310 23750 10362
rect 23750 10310 23762 10362
rect 23762 10310 23792 10362
rect 23816 10310 23826 10362
rect 23826 10310 23872 10362
rect 23576 10308 23632 10310
rect 23656 10308 23712 10310
rect 23736 10308 23792 10310
rect 23816 10308 23872 10310
rect 24858 12416 24914 12472
rect 25318 19352 25374 19408
rect 25686 18420 25742 18456
rect 25686 18400 25688 18420
rect 25688 18400 25740 18420
rect 25740 18400 25742 18420
rect 25502 13368 25558 13424
rect 25502 13232 25558 13288
rect 25870 19896 25926 19952
rect 26076 20698 26132 20700
rect 26156 20698 26212 20700
rect 26236 20698 26292 20700
rect 26316 20698 26372 20700
rect 26076 20646 26122 20698
rect 26122 20646 26132 20698
rect 26156 20646 26186 20698
rect 26186 20646 26198 20698
rect 26198 20646 26212 20698
rect 26236 20646 26250 20698
rect 26250 20646 26262 20698
rect 26262 20646 26292 20698
rect 26316 20646 26326 20698
rect 26326 20646 26372 20698
rect 26076 20644 26132 20646
rect 26156 20644 26212 20646
rect 26236 20644 26292 20646
rect 26316 20644 26372 20646
rect 26146 19760 26202 19816
rect 26076 19610 26132 19612
rect 26156 19610 26212 19612
rect 26236 19610 26292 19612
rect 26316 19610 26372 19612
rect 26076 19558 26122 19610
rect 26122 19558 26132 19610
rect 26156 19558 26186 19610
rect 26186 19558 26198 19610
rect 26198 19558 26212 19610
rect 26236 19558 26250 19610
rect 26250 19558 26262 19610
rect 26262 19558 26292 19610
rect 26316 19558 26326 19610
rect 26326 19558 26372 19610
rect 26076 19556 26132 19558
rect 26156 19556 26212 19558
rect 26236 19556 26292 19558
rect 26316 19556 26372 19558
rect 26076 18522 26132 18524
rect 26156 18522 26212 18524
rect 26236 18522 26292 18524
rect 26316 18522 26372 18524
rect 26076 18470 26122 18522
rect 26122 18470 26132 18522
rect 26156 18470 26186 18522
rect 26186 18470 26198 18522
rect 26198 18470 26212 18522
rect 26236 18470 26250 18522
rect 26250 18470 26262 18522
rect 26262 18470 26292 18522
rect 26316 18470 26326 18522
rect 26326 18470 26372 18522
rect 26076 18468 26132 18470
rect 26156 18468 26212 18470
rect 26236 18468 26292 18470
rect 26316 18468 26372 18470
rect 25962 18264 26018 18320
rect 24858 12144 24914 12200
rect 23386 9832 23442 9888
rect 22374 8744 22430 8800
rect 22558 7284 22560 7304
rect 22560 7284 22612 7304
rect 22612 7284 22614 7304
rect 22558 7248 22614 7284
rect 22466 6568 22522 6624
rect 23478 9444 23534 9480
rect 23478 9424 23480 9444
rect 23480 9424 23532 9444
rect 23532 9424 23534 9444
rect 23576 9274 23632 9276
rect 23656 9274 23712 9276
rect 23736 9274 23792 9276
rect 23816 9274 23872 9276
rect 23576 9222 23622 9274
rect 23622 9222 23632 9274
rect 23656 9222 23686 9274
rect 23686 9222 23698 9274
rect 23698 9222 23712 9274
rect 23736 9222 23750 9274
rect 23750 9222 23762 9274
rect 23762 9222 23792 9274
rect 23816 9222 23826 9274
rect 23826 9222 23872 9274
rect 23576 9220 23632 9222
rect 23656 9220 23712 9222
rect 23736 9220 23792 9222
rect 23816 9220 23872 9222
rect 23386 8780 23388 8800
rect 23388 8780 23440 8800
rect 23440 8780 23442 8800
rect 23386 8744 23442 8780
rect 22466 5888 22522 5944
rect 22006 5344 22062 5400
rect 21730 3984 21786 4040
rect 21730 3732 21786 3768
rect 22466 4936 22522 4992
rect 23018 6976 23074 7032
rect 23018 6840 23074 6896
rect 23576 8186 23632 8188
rect 23656 8186 23712 8188
rect 23736 8186 23792 8188
rect 23816 8186 23872 8188
rect 23576 8134 23622 8186
rect 23622 8134 23632 8186
rect 23656 8134 23686 8186
rect 23686 8134 23698 8186
rect 23698 8134 23712 8186
rect 23736 8134 23750 8186
rect 23750 8134 23762 8186
rect 23762 8134 23792 8186
rect 23816 8134 23826 8186
rect 23826 8134 23872 8186
rect 23576 8132 23632 8134
rect 23656 8132 23712 8134
rect 23736 8132 23792 8134
rect 23816 8132 23872 8134
rect 24122 7248 24178 7304
rect 23576 7098 23632 7100
rect 23656 7098 23712 7100
rect 23736 7098 23792 7100
rect 23816 7098 23872 7100
rect 23576 7046 23622 7098
rect 23622 7046 23632 7098
rect 23656 7046 23686 7098
rect 23686 7046 23698 7098
rect 23698 7046 23712 7098
rect 23736 7046 23750 7098
rect 23750 7046 23762 7098
rect 23762 7046 23792 7098
rect 23816 7046 23826 7098
rect 23826 7046 23872 7098
rect 23576 7044 23632 7046
rect 23656 7044 23712 7046
rect 23736 7044 23792 7046
rect 23816 7044 23872 7046
rect 24306 6840 24362 6896
rect 24122 6568 24178 6624
rect 23110 6296 23166 6352
rect 23576 6010 23632 6012
rect 23656 6010 23712 6012
rect 23736 6010 23792 6012
rect 23816 6010 23872 6012
rect 23576 5958 23622 6010
rect 23622 5958 23632 6010
rect 23656 5958 23686 6010
rect 23686 5958 23698 6010
rect 23698 5958 23712 6010
rect 23736 5958 23750 6010
rect 23750 5958 23762 6010
rect 23762 5958 23792 6010
rect 23816 5958 23826 6010
rect 23826 5958 23872 6010
rect 23576 5956 23632 5958
rect 23656 5956 23712 5958
rect 23736 5956 23792 5958
rect 23816 5956 23872 5958
rect 23386 5888 23442 5944
rect 23202 5480 23258 5536
rect 22742 4800 22798 4856
rect 23294 5228 23350 5264
rect 23294 5208 23296 5228
rect 23296 5208 23348 5228
rect 23348 5208 23350 5228
rect 22926 4664 22982 4720
rect 22282 4392 22338 4448
rect 21730 3712 21732 3732
rect 21732 3712 21784 3732
rect 21784 3712 21786 3732
rect 21076 3290 21132 3292
rect 21156 3290 21212 3292
rect 21236 3290 21292 3292
rect 21316 3290 21372 3292
rect 21076 3238 21122 3290
rect 21122 3238 21132 3290
rect 21156 3238 21186 3290
rect 21186 3238 21198 3290
rect 21198 3238 21212 3290
rect 21236 3238 21250 3290
rect 21250 3238 21262 3290
rect 21262 3238 21292 3290
rect 21316 3238 21326 3290
rect 21326 3238 21372 3290
rect 21076 3236 21132 3238
rect 21156 3236 21212 3238
rect 21236 3236 21292 3238
rect 21316 3236 21372 3238
rect 21178 3032 21234 3088
rect 21076 2202 21132 2204
rect 21156 2202 21212 2204
rect 21236 2202 21292 2204
rect 21316 2202 21372 2204
rect 21076 2150 21122 2202
rect 21122 2150 21132 2202
rect 21156 2150 21186 2202
rect 21186 2150 21198 2202
rect 21198 2150 21212 2202
rect 21236 2150 21250 2202
rect 21250 2150 21262 2202
rect 21262 2150 21292 2202
rect 21316 2150 21326 2202
rect 21326 2150 21372 2202
rect 21076 2148 21132 2150
rect 21156 2148 21212 2150
rect 21236 2148 21292 2150
rect 21316 2148 21372 2150
rect 21546 1964 21602 2000
rect 21546 1944 21548 1964
rect 21548 1944 21600 1964
rect 21600 1944 21602 1964
rect 21076 1114 21132 1116
rect 21156 1114 21212 1116
rect 21236 1114 21292 1116
rect 21316 1114 21372 1116
rect 21076 1062 21122 1114
rect 21122 1062 21132 1114
rect 21156 1062 21186 1114
rect 21186 1062 21198 1114
rect 21198 1062 21212 1114
rect 21236 1062 21250 1114
rect 21250 1062 21262 1114
rect 21262 1062 21292 1114
rect 21316 1062 21326 1114
rect 21326 1062 21372 1114
rect 21076 1060 21132 1062
rect 21156 1060 21212 1062
rect 21236 1060 21292 1062
rect 21316 1060 21372 1062
rect 23294 4528 23350 4584
rect 23576 4922 23632 4924
rect 23656 4922 23712 4924
rect 23736 4922 23792 4924
rect 23816 4922 23872 4924
rect 23576 4870 23622 4922
rect 23622 4870 23632 4922
rect 23656 4870 23686 4922
rect 23686 4870 23698 4922
rect 23698 4870 23712 4922
rect 23736 4870 23750 4922
rect 23750 4870 23762 4922
rect 23762 4870 23792 4922
rect 23816 4870 23826 4922
rect 23826 4870 23872 4922
rect 23576 4868 23632 4870
rect 23656 4868 23712 4870
rect 23736 4868 23792 4870
rect 23816 4868 23872 4870
rect 23846 4140 23902 4176
rect 23846 4120 23848 4140
rect 23848 4120 23900 4140
rect 23900 4120 23902 4140
rect 23576 3834 23632 3836
rect 23656 3834 23712 3836
rect 23736 3834 23792 3836
rect 23816 3834 23872 3836
rect 23576 3782 23622 3834
rect 23622 3782 23632 3834
rect 23656 3782 23686 3834
rect 23686 3782 23698 3834
rect 23698 3782 23712 3834
rect 23736 3782 23750 3834
rect 23750 3782 23762 3834
rect 23762 3782 23792 3834
rect 23816 3782 23826 3834
rect 23826 3782 23872 3834
rect 23576 3780 23632 3782
rect 23656 3780 23712 3782
rect 23736 3780 23792 3782
rect 23816 3780 23872 3782
rect 23386 3732 23442 3768
rect 23386 3712 23388 3732
rect 23388 3712 23440 3732
rect 23440 3712 23442 3732
rect 23386 3576 23442 3632
rect 24214 6024 24270 6080
rect 24122 5072 24178 5128
rect 24122 4428 24124 4448
rect 24124 4428 24176 4448
rect 24176 4428 24178 4448
rect 24122 4392 24178 4428
rect 23576 2746 23632 2748
rect 23656 2746 23712 2748
rect 23736 2746 23792 2748
rect 23816 2746 23872 2748
rect 23576 2694 23622 2746
rect 23622 2694 23632 2746
rect 23656 2694 23686 2746
rect 23686 2694 23698 2746
rect 23698 2694 23712 2746
rect 23736 2694 23750 2746
rect 23750 2694 23762 2746
rect 23762 2694 23792 2746
rect 23816 2694 23826 2746
rect 23826 2694 23872 2746
rect 23576 2692 23632 2694
rect 23656 2692 23712 2694
rect 23736 2692 23792 2694
rect 23816 2692 23872 2694
rect 25318 13096 25374 13152
rect 25410 12860 25412 12880
rect 25412 12860 25464 12880
rect 25464 12860 25466 12880
rect 25226 12724 25228 12744
rect 25228 12724 25280 12744
rect 25280 12724 25282 12744
rect 25226 12688 25282 12724
rect 25410 12824 25466 12860
rect 25318 11736 25374 11792
rect 25042 9016 25098 9072
rect 24766 6840 24822 6896
rect 24306 5652 24308 5672
rect 24308 5652 24360 5672
rect 24360 5652 24362 5672
rect 24306 5616 24362 5652
rect 24490 5616 24546 5672
rect 24582 5480 24638 5536
rect 24490 5072 24546 5128
rect 24306 3576 24362 3632
rect 23576 1658 23632 1660
rect 23656 1658 23712 1660
rect 23736 1658 23792 1660
rect 23816 1658 23872 1660
rect 23576 1606 23622 1658
rect 23622 1606 23632 1658
rect 23656 1606 23686 1658
rect 23686 1606 23698 1658
rect 23698 1606 23712 1658
rect 23736 1606 23750 1658
rect 23750 1606 23762 1658
rect 23762 1606 23792 1658
rect 23816 1606 23826 1658
rect 23826 1606 23872 1658
rect 23576 1604 23632 1606
rect 23656 1604 23712 1606
rect 23736 1604 23792 1606
rect 23816 1604 23872 1606
rect 24582 4936 24638 4992
rect 25042 6840 25098 6896
rect 25594 8336 25650 8392
rect 25502 7792 25558 7848
rect 25134 6296 25190 6352
rect 25042 5888 25098 5944
rect 25778 7248 25834 7304
rect 25594 6704 25650 6760
rect 25410 6432 25466 6488
rect 25134 5752 25190 5808
rect 25042 5344 25098 5400
rect 25134 5208 25190 5264
rect 25042 4528 25098 4584
rect 25226 3984 25282 4040
rect 25134 3032 25190 3088
rect 25594 6160 25650 6216
rect 25594 5752 25650 5808
rect 26076 17434 26132 17436
rect 26156 17434 26212 17436
rect 26236 17434 26292 17436
rect 26316 17434 26372 17436
rect 26076 17382 26122 17434
rect 26122 17382 26132 17434
rect 26156 17382 26186 17434
rect 26186 17382 26198 17434
rect 26198 17382 26212 17434
rect 26236 17382 26250 17434
rect 26250 17382 26262 17434
rect 26262 17382 26292 17434
rect 26316 17382 26326 17434
rect 26326 17382 26372 17434
rect 26076 17380 26132 17382
rect 26156 17380 26212 17382
rect 26236 17380 26292 17382
rect 26316 17380 26372 17382
rect 26076 16346 26132 16348
rect 26156 16346 26212 16348
rect 26236 16346 26292 16348
rect 26316 16346 26372 16348
rect 26076 16294 26122 16346
rect 26122 16294 26132 16346
rect 26156 16294 26186 16346
rect 26186 16294 26198 16346
rect 26198 16294 26212 16346
rect 26236 16294 26250 16346
rect 26250 16294 26262 16346
rect 26262 16294 26292 16346
rect 26316 16294 26326 16346
rect 26326 16294 26372 16346
rect 26076 16292 26132 16294
rect 26156 16292 26212 16294
rect 26236 16292 26292 16294
rect 26316 16292 26372 16294
rect 27158 21004 27214 21040
rect 27158 20984 27160 21004
rect 27160 20984 27212 21004
rect 27212 20984 27214 21004
rect 26882 18808 26938 18864
rect 26882 16496 26938 16552
rect 26514 15972 26570 16008
rect 26514 15952 26516 15972
rect 26516 15952 26568 15972
rect 26568 15952 26570 15972
rect 26076 15258 26132 15260
rect 26156 15258 26212 15260
rect 26236 15258 26292 15260
rect 26316 15258 26372 15260
rect 26076 15206 26122 15258
rect 26122 15206 26132 15258
rect 26156 15206 26186 15258
rect 26186 15206 26198 15258
rect 26198 15206 26212 15258
rect 26236 15206 26250 15258
rect 26250 15206 26262 15258
rect 26262 15206 26292 15258
rect 26316 15206 26326 15258
rect 26326 15206 26372 15258
rect 26076 15204 26132 15206
rect 26156 15204 26212 15206
rect 26236 15204 26292 15206
rect 26316 15204 26372 15206
rect 26238 14592 26294 14648
rect 26076 14170 26132 14172
rect 26156 14170 26212 14172
rect 26236 14170 26292 14172
rect 26316 14170 26372 14172
rect 26076 14118 26122 14170
rect 26122 14118 26132 14170
rect 26156 14118 26186 14170
rect 26186 14118 26198 14170
rect 26198 14118 26212 14170
rect 26236 14118 26250 14170
rect 26250 14118 26262 14170
rect 26262 14118 26292 14170
rect 26316 14118 26326 14170
rect 26326 14118 26372 14170
rect 26076 14116 26132 14118
rect 26156 14116 26212 14118
rect 26236 14116 26292 14118
rect 26316 14116 26372 14118
rect 27066 14320 27122 14376
rect 26076 13082 26132 13084
rect 26156 13082 26212 13084
rect 26236 13082 26292 13084
rect 26316 13082 26372 13084
rect 26076 13030 26122 13082
rect 26122 13030 26132 13082
rect 26156 13030 26186 13082
rect 26186 13030 26198 13082
rect 26198 13030 26212 13082
rect 26236 13030 26250 13082
rect 26250 13030 26262 13082
rect 26262 13030 26292 13082
rect 26316 13030 26326 13082
rect 26326 13030 26372 13082
rect 26076 13028 26132 13030
rect 26156 13028 26212 13030
rect 26236 13028 26292 13030
rect 26316 13028 26372 13030
rect 26054 12824 26110 12880
rect 27158 13524 27214 13560
rect 27158 13504 27160 13524
rect 27160 13504 27212 13524
rect 27212 13504 27214 13524
rect 26422 12280 26478 12336
rect 26076 11994 26132 11996
rect 26156 11994 26212 11996
rect 26236 11994 26292 11996
rect 26316 11994 26372 11996
rect 26076 11942 26122 11994
rect 26122 11942 26132 11994
rect 26156 11942 26186 11994
rect 26186 11942 26198 11994
rect 26198 11942 26212 11994
rect 26236 11942 26250 11994
rect 26250 11942 26262 11994
rect 26262 11942 26292 11994
rect 26316 11942 26326 11994
rect 26326 11942 26372 11994
rect 26076 11940 26132 11942
rect 26156 11940 26212 11942
rect 26236 11940 26292 11942
rect 26316 11940 26372 11942
rect 26076 10906 26132 10908
rect 26156 10906 26212 10908
rect 26236 10906 26292 10908
rect 26316 10906 26372 10908
rect 26076 10854 26122 10906
rect 26122 10854 26132 10906
rect 26156 10854 26186 10906
rect 26186 10854 26198 10906
rect 26198 10854 26212 10906
rect 26236 10854 26250 10906
rect 26250 10854 26262 10906
rect 26262 10854 26292 10906
rect 26316 10854 26326 10906
rect 26326 10854 26372 10906
rect 26076 10852 26132 10854
rect 26156 10852 26212 10854
rect 26236 10852 26292 10854
rect 26316 10852 26372 10854
rect 26076 9818 26132 9820
rect 26156 9818 26212 9820
rect 26236 9818 26292 9820
rect 26316 9818 26372 9820
rect 26076 9766 26122 9818
rect 26122 9766 26132 9818
rect 26156 9766 26186 9818
rect 26186 9766 26198 9818
rect 26198 9766 26212 9818
rect 26236 9766 26250 9818
rect 26250 9766 26262 9818
rect 26262 9766 26292 9818
rect 26316 9766 26326 9818
rect 26326 9766 26372 9818
rect 26076 9764 26132 9766
rect 26156 9764 26212 9766
rect 26236 9764 26292 9766
rect 26316 9764 26372 9766
rect 26514 8900 26570 8936
rect 26514 8880 26516 8900
rect 26516 8880 26568 8900
rect 26568 8880 26570 8900
rect 26076 8730 26132 8732
rect 26156 8730 26212 8732
rect 26236 8730 26292 8732
rect 26316 8730 26372 8732
rect 26076 8678 26122 8730
rect 26122 8678 26132 8730
rect 26156 8678 26186 8730
rect 26186 8678 26198 8730
rect 26198 8678 26212 8730
rect 26236 8678 26250 8730
rect 26250 8678 26262 8730
rect 26262 8678 26292 8730
rect 26316 8678 26326 8730
rect 26326 8678 26372 8730
rect 26076 8676 26132 8678
rect 26156 8676 26212 8678
rect 26236 8676 26292 8678
rect 26316 8676 26372 8678
rect 26974 12708 27030 12744
rect 26974 12688 26976 12708
rect 26976 12688 27028 12708
rect 27028 12688 27030 12708
rect 26882 11192 26938 11248
rect 26790 7928 26846 7984
rect 26514 7792 26570 7848
rect 26076 7642 26132 7644
rect 26156 7642 26212 7644
rect 26236 7642 26292 7644
rect 26316 7642 26372 7644
rect 26076 7590 26122 7642
rect 26122 7590 26132 7642
rect 26156 7590 26186 7642
rect 26186 7590 26198 7642
rect 26198 7590 26212 7642
rect 26236 7590 26250 7642
rect 26250 7590 26262 7642
rect 26262 7590 26292 7642
rect 26316 7590 26326 7642
rect 26326 7590 26372 7642
rect 26076 7588 26132 7590
rect 26156 7588 26212 7590
rect 26236 7588 26292 7590
rect 26316 7588 26372 7590
rect 26146 6840 26202 6896
rect 26076 6554 26132 6556
rect 26156 6554 26212 6556
rect 26236 6554 26292 6556
rect 26316 6554 26372 6556
rect 26076 6502 26122 6554
rect 26122 6502 26132 6554
rect 26156 6502 26186 6554
rect 26186 6502 26198 6554
rect 26198 6502 26212 6554
rect 26236 6502 26250 6554
rect 26250 6502 26262 6554
rect 26262 6502 26292 6554
rect 26316 6502 26326 6554
rect 26326 6502 26372 6554
rect 26076 6500 26132 6502
rect 26156 6500 26212 6502
rect 26236 6500 26292 6502
rect 26316 6500 26372 6502
rect 26076 5466 26132 5468
rect 26156 5466 26212 5468
rect 26236 5466 26292 5468
rect 26316 5466 26372 5468
rect 26076 5414 26122 5466
rect 26122 5414 26132 5466
rect 26156 5414 26186 5466
rect 26186 5414 26198 5466
rect 26198 5414 26212 5466
rect 26236 5414 26250 5466
rect 26250 5414 26262 5466
rect 26262 5414 26292 5466
rect 26316 5414 26326 5466
rect 26326 5414 26372 5466
rect 26076 5412 26132 5414
rect 26156 5412 26212 5414
rect 26236 5412 26292 5414
rect 26316 5412 26372 5414
rect 26054 4800 26110 4856
rect 26076 4378 26132 4380
rect 26156 4378 26212 4380
rect 26236 4378 26292 4380
rect 26316 4378 26372 4380
rect 26076 4326 26122 4378
rect 26122 4326 26132 4378
rect 26156 4326 26186 4378
rect 26186 4326 26198 4378
rect 26198 4326 26212 4378
rect 26236 4326 26250 4378
rect 26250 4326 26262 4378
rect 26262 4326 26292 4378
rect 26316 4326 26326 4378
rect 26326 4326 26372 4378
rect 26076 4324 26132 4326
rect 26156 4324 26212 4326
rect 26236 4324 26292 4326
rect 26316 4324 26372 4326
rect 28576 22330 28632 22332
rect 28656 22330 28712 22332
rect 28736 22330 28792 22332
rect 28816 22330 28872 22332
rect 28576 22278 28622 22330
rect 28622 22278 28632 22330
rect 28656 22278 28686 22330
rect 28686 22278 28698 22330
rect 28698 22278 28712 22330
rect 28736 22278 28750 22330
rect 28750 22278 28762 22330
rect 28762 22278 28792 22330
rect 28816 22278 28826 22330
rect 28826 22278 28872 22330
rect 28576 22276 28632 22278
rect 28656 22276 28712 22278
rect 28736 22276 28792 22278
rect 28816 22276 28872 22278
rect 27618 21936 27674 21992
rect 27710 21664 27766 21720
rect 28354 21956 28410 21992
rect 28354 21936 28356 21956
rect 28356 21936 28408 21956
rect 28408 21936 28410 21956
rect 27710 20440 27766 20496
rect 27342 15544 27398 15600
rect 28576 21242 28632 21244
rect 28656 21242 28712 21244
rect 28736 21242 28792 21244
rect 28816 21242 28872 21244
rect 28576 21190 28622 21242
rect 28622 21190 28632 21242
rect 28656 21190 28686 21242
rect 28686 21190 28698 21242
rect 28698 21190 28712 21242
rect 28736 21190 28750 21242
rect 28750 21190 28762 21242
rect 28762 21190 28792 21242
rect 28816 21190 28826 21242
rect 28826 21190 28872 21242
rect 28576 21188 28632 21190
rect 28656 21188 28712 21190
rect 28736 21188 28792 21190
rect 28816 21188 28872 21190
rect 28354 19896 28410 19952
rect 28078 19488 28134 19544
rect 28262 19352 28318 19408
rect 27894 16632 27950 16688
rect 27434 14456 27490 14512
rect 27618 12980 27674 13016
rect 27618 12960 27620 12980
rect 27620 12960 27672 12980
rect 27672 12960 27674 12980
rect 27894 15272 27950 15328
rect 27158 6840 27214 6896
rect 27434 7384 27490 7440
rect 26974 5208 27030 5264
rect 28576 20154 28632 20156
rect 28656 20154 28712 20156
rect 28736 20154 28792 20156
rect 28816 20154 28872 20156
rect 28576 20102 28622 20154
rect 28622 20102 28632 20154
rect 28656 20102 28686 20154
rect 28686 20102 28698 20154
rect 28698 20102 28712 20154
rect 28736 20102 28750 20154
rect 28750 20102 28762 20154
rect 28762 20102 28792 20154
rect 28816 20102 28826 20154
rect 28826 20102 28872 20154
rect 28576 20100 28632 20102
rect 28656 20100 28712 20102
rect 28736 20100 28792 20102
rect 28816 20100 28872 20102
rect 28630 19896 28686 19952
rect 31076 22874 31132 22876
rect 31156 22874 31212 22876
rect 31236 22874 31292 22876
rect 31316 22874 31372 22876
rect 31076 22822 31122 22874
rect 31122 22822 31132 22874
rect 31156 22822 31186 22874
rect 31186 22822 31198 22874
rect 31198 22822 31212 22874
rect 31236 22822 31250 22874
rect 31250 22822 31262 22874
rect 31262 22822 31292 22874
rect 31316 22822 31326 22874
rect 31326 22822 31372 22874
rect 31076 22820 31132 22822
rect 31156 22820 31212 22822
rect 31236 22820 31292 22822
rect 31316 22820 31372 22822
rect 30010 21528 30066 21584
rect 29090 20712 29146 20768
rect 28630 19488 28686 19544
rect 28576 19066 28632 19068
rect 28656 19066 28712 19068
rect 28736 19066 28792 19068
rect 28816 19066 28872 19068
rect 28576 19014 28622 19066
rect 28622 19014 28632 19066
rect 28656 19014 28686 19066
rect 28686 19014 28698 19066
rect 28698 19014 28712 19066
rect 28736 19014 28750 19066
rect 28750 19014 28762 19066
rect 28762 19014 28792 19066
rect 28816 19014 28826 19066
rect 28826 19014 28872 19066
rect 28576 19012 28632 19014
rect 28656 19012 28712 19014
rect 28736 19012 28792 19014
rect 28816 19012 28872 19014
rect 30378 21120 30434 21176
rect 29918 20848 29974 20904
rect 29182 20440 29238 20496
rect 29642 19488 29698 19544
rect 29090 18264 29146 18320
rect 28576 17978 28632 17980
rect 28656 17978 28712 17980
rect 28736 17978 28792 17980
rect 28816 17978 28872 17980
rect 28576 17926 28622 17978
rect 28622 17926 28632 17978
rect 28656 17926 28686 17978
rect 28686 17926 28698 17978
rect 28698 17926 28712 17978
rect 28736 17926 28750 17978
rect 28750 17926 28762 17978
rect 28762 17926 28792 17978
rect 28816 17926 28826 17978
rect 28826 17926 28872 17978
rect 28576 17924 28632 17926
rect 28656 17924 28712 17926
rect 28736 17924 28792 17926
rect 28816 17924 28872 17926
rect 28576 16890 28632 16892
rect 28656 16890 28712 16892
rect 28736 16890 28792 16892
rect 28816 16890 28872 16892
rect 28576 16838 28622 16890
rect 28622 16838 28632 16890
rect 28656 16838 28686 16890
rect 28686 16838 28698 16890
rect 28698 16838 28712 16890
rect 28736 16838 28750 16890
rect 28750 16838 28762 16890
rect 28762 16838 28792 16890
rect 28816 16838 28826 16890
rect 28826 16838 28872 16890
rect 28576 16836 28632 16838
rect 28656 16836 28712 16838
rect 28736 16836 28792 16838
rect 28816 16836 28872 16838
rect 28576 15802 28632 15804
rect 28656 15802 28712 15804
rect 28736 15802 28792 15804
rect 28816 15802 28872 15804
rect 28576 15750 28622 15802
rect 28622 15750 28632 15802
rect 28656 15750 28686 15802
rect 28686 15750 28698 15802
rect 28698 15750 28712 15802
rect 28736 15750 28750 15802
rect 28750 15750 28762 15802
rect 28762 15750 28792 15802
rect 28816 15750 28826 15802
rect 28826 15750 28872 15802
rect 28576 15748 28632 15750
rect 28656 15748 28712 15750
rect 28736 15748 28792 15750
rect 28816 15748 28872 15750
rect 29826 18808 29882 18864
rect 29090 15988 29092 16008
rect 29092 15988 29144 16008
rect 29144 15988 29146 16008
rect 29090 15952 29146 15988
rect 28078 14320 28134 14376
rect 28354 14068 28410 14104
rect 28576 14714 28632 14716
rect 28656 14714 28712 14716
rect 28736 14714 28792 14716
rect 28816 14714 28872 14716
rect 28576 14662 28622 14714
rect 28622 14662 28632 14714
rect 28656 14662 28686 14714
rect 28686 14662 28698 14714
rect 28698 14662 28712 14714
rect 28736 14662 28750 14714
rect 28750 14662 28762 14714
rect 28762 14662 28792 14714
rect 28816 14662 28826 14714
rect 28826 14662 28872 14714
rect 28576 14660 28632 14662
rect 28656 14660 28712 14662
rect 28736 14660 28792 14662
rect 28816 14660 28872 14662
rect 29090 15272 29146 15328
rect 28354 14048 28356 14068
rect 28356 14048 28408 14068
rect 28408 14048 28410 14068
rect 28576 13626 28632 13628
rect 28656 13626 28712 13628
rect 28736 13626 28792 13628
rect 28816 13626 28872 13628
rect 28576 13574 28622 13626
rect 28622 13574 28632 13626
rect 28656 13574 28686 13626
rect 28686 13574 28698 13626
rect 28698 13574 28712 13626
rect 28736 13574 28750 13626
rect 28750 13574 28762 13626
rect 28762 13574 28792 13626
rect 28816 13574 28826 13626
rect 28826 13574 28872 13626
rect 28576 13572 28632 13574
rect 28656 13572 28712 13574
rect 28736 13572 28792 13574
rect 28816 13572 28872 13574
rect 28262 12960 28318 13016
rect 28354 12824 28410 12880
rect 29090 13776 29146 13832
rect 28576 12538 28632 12540
rect 28656 12538 28712 12540
rect 28736 12538 28792 12540
rect 28816 12538 28872 12540
rect 28576 12486 28622 12538
rect 28622 12486 28632 12538
rect 28656 12486 28686 12538
rect 28686 12486 28698 12538
rect 28698 12486 28712 12538
rect 28736 12486 28750 12538
rect 28750 12486 28762 12538
rect 28762 12486 28792 12538
rect 28816 12486 28826 12538
rect 28826 12486 28872 12538
rect 28576 12484 28632 12486
rect 28656 12484 28712 12486
rect 28736 12484 28792 12486
rect 28816 12484 28872 12486
rect 28576 11450 28632 11452
rect 28656 11450 28712 11452
rect 28736 11450 28792 11452
rect 28816 11450 28872 11452
rect 28576 11398 28622 11450
rect 28622 11398 28632 11450
rect 28656 11398 28686 11450
rect 28686 11398 28698 11450
rect 28698 11398 28712 11450
rect 28736 11398 28750 11450
rect 28750 11398 28762 11450
rect 28762 11398 28792 11450
rect 28816 11398 28826 11450
rect 28826 11398 28872 11450
rect 28576 11396 28632 11398
rect 28656 11396 28712 11398
rect 28736 11396 28792 11398
rect 28816 11396 28872 11398
rect 29366 14864 29422 14920
rect 29274 13368 29330 13424
rect 29182 12144 29238 12200
rect 29918 17584 29974 17640
rect 30746 21548 30802 21584
rect 30746 21528 30748 21548
rect 30748 21528 30800 21548
rect 30800 21528 30802 21548
rect 30378 20032 30434 20088
rect 30470 19352 30526 19408
rect 30746 20576 30802 20632
rect 31076 21786 31132 21788
rect 31156 21786 31212 21788
rect 31236 21786 31292 21788
rect 31316 21786 31372 21788
rect 31076 21734 31122 21786
rect 31122 21734 31132 21786
rect 31156 21734 31186 21786
rect 31186 21734 31198 21786
rect 31198 21734 31212 21786
rect 31236 21734 31250 21786
rect 31250 21734 31262 21786
rect 31262 21734 31292 21786
rect 31316 21734 31326 21786
rect 31326 21734 31372 21786
rect 31076 21732 31132 21734
rect 31156 21732 31212 21734
rect 31236 21732 31292 21734
rect 31316 21732 31372 21734
rect 31114 21392 31170 21448
rect 31076 20698 31132 20700
rect 31156 20698 31212 20700
rect 31236 20698 31292 20700
rect 31316 20698 31372 20700
rect 31076 20646 31122 20698
rect 31122 20646 31132 20698
rect 31156 20646 31186 20698
rect 31186 20646 31198 20698
rect 31198 20646 31212 20698
rect 31236 20646 31250 20698
rect 31250 20646 31262 20698
rect 31262 20646 31292 20698
rect 31316 20646 31326 20698
rect 31326 20646 31372 20698
rect 31076 20644 31132 20646
rect 31156 20644 31212 20646
rect 31236 20644 31292 20646
rect 31316 20644 31372 20646
rect 32402 22072 32458 22128
rect 32954 22072 33010 22128
rect 30746 20168 30802 20224
rect 31022 20032 31078 20088
rect 30470 17448 30526 17504
rect 31076 19610 31132 19612
rect 31156 19610 31212 19612
rect 31236 19610 31292 19612
rect 31316 19610 31372 19612
rect 31076 19558 31122 19610
rect 31122 19558 31132 19610
rect 31156 19558 31186 19610
rect 31186 19558 31198 19610
rect 31198 19558 31212 19610
rect 31236 19558 31250 19610
rect 31250 19558 31262 19610
rect 31262 19558 31292 19610
rect 31316 19558 31326 19610
rect 31326 19558 31372 19610
rect 31076 19556 31132 19558
rect 31156 19556 31212 19558
rect 31236 19556 31292 19558
rect 31316 19556 31372 19558
rect 30930 19488 30986 19544
rect 30746 18944 30802 19000
rect 31666 20168 31722 20224
rect 32126 20984 32182 21040
rect 32034 20440 32090 20496
rect 31076 18522 31132 18524
rect 31156 18522 31212 18524
rect 31236 18522 31292 18524
rect 31316 18522 31372 18524
rect 31076 18470 31122 18522
rect 31122 18470 31132 18522
rect 31156 18470 31186 18522
rect 31186 18470 31198 18522
rect 31198 18470 31212 18522
rect 31236 18470 31250 18522
rect 31250 18470 31262 18522
rect 31262 18470 31292 18522
rect 31316 18470 31326 18522
rect 31326 18470 31372 18522
rect 31076 18468 31132 18470
rect 31156 18468 31212 18470
rect 31236 18468 31292 18470
rect 31316 18468 31372 18470
rect 31574 18944 31630 19000
rect 31206 18128 31262 18184
rect 32310 20324 32366 20360
rect 32310 20304 32312 20324
rect 32312 20304 32364 20324
rect 32364 20304 32366 20324
rect 31574 17584 31630 17640
rect 31076 17434 31132 17436
rect 31156 17434 31212 17436
rect 31236 17434 31292 17436
rect 31316 17434 31372 17436
rect 31076 17382 31122 17434
rect 31122 17382 31132 17434
rect 31156 17382 31186 17434
rect 31186 17382 31198 17434
rect 31198 17382 31212 17434
rect 31236 17382 31250 17434
rect 31250 17382 31262 17434
rect 31262 17382 31292 17434
rect 31316 17382 31326 17434
rect 31326 17382 31372 17434
rect 31076 17380 31132 17382
rect 31156 17380 31212 17382
rect 31236 17380 31292 17382
rect 31316 17380 31372 17382
rect 29734 14320 29790 14376
rect 31758 17196 31814 17232
rect 32586 20984 32642 21040
rect 36076 22874 36132 22876
rect 36156 22874 36212 22876
rect 36236 22874 36292 22876
rect 36316 22874 36372 22876
rect 36076 22822 36122 22874
rect 36122 22822 36132 22874
rect 36156 22822 36186 22874
rect 36186 22822 36198 22874
rect 36198 22822 36212 22874
rect 36236 22822 36250 22874
rect 36250 22822 36262 22874
rect 36262 22822 36292 22874
rect 36316 22822 36326 22874
rect 36326 22822 36372 22874
rect 36076 22820 36132 22822
rect 36156 22820 36212 22822
rect 36236 22820 36292 22822
rect 36316 22820 36372 22822
rect 33576 22330 33632 22332
rect 33656 22330 33712 22332
rect 33736 22330 33792 22332
rect 33816 22330 33872 22332
rect 33576 22278 33622 22330
rect 33622 22278 33632 22330
rect 33656 22278 33686 22330
rect 33686 22278 33698 22330
rect 33698 22278 33712 22330
rect 33736 22278 33750 22330
rect 33750 22278 33762 22330
rect 33762 22278 33792 22330
rect 33816 22278 33826 22330
rect 33826 22278 33872 22330
rect 33576 22276 33632 22278
rect 33656 22276 33712 22278
rect 33736 22276 33792 22278
rect 33816 22276 33872 22278
rect 33414 21936 33470 21992
rect 33230 20984 33286 21040
rect 33576 21242 33632 21244
rect 33656 21242 33712 21244
rect 33736 21242 33792 21244
rect 33816 21242 33872 21244
rect 33576 21190 33622 21242
rect 33622 21190 33632 21242
rect 33656 21190 33686 21242
rect 33686 21190 33698 21242
rect 33698 21190 33712 21242
rect 33736 21190 33750 21242
rect 33750 21190 33762 21242
rect 33762 21190 33792 21242
rect 33816 21190 33826 21242
rect 33826 21190 33872 21242
rect 33576 21188 33632 21190
rect 33656 21188 33712 21190
rect 33736 21188 33792 21190
rect 33816 21188 33872 21190
rect 32954 20712 33010 20768
rect 32770 20576 32826 20632
rect 32494 19760 32550 19816
rect 32954 20476 32956 20496
rect 32956 20476 33008 20496
rect 33008 20476 33010 20496
rect 32954 20440 33010 20476
rect 33230 20304 33286 20360
rect 33322 20032 33378 20088
rect 33576 20154 33632 20156
rect 33656 20154 33712 20156
rect 33736 20154 33792 20156
rect 33816 20154 33872 20156
rect 33576 20102 33622 20154
rect 33622 20102 33632 20154
rect 33656 20102 33686 20154
rect 33686 20102 33698 20154
rect 33698 20102 33712 20154
rect 33736 20102 33750 20154
rect 33750 20102 33762 20154
rect 33762 20102 33792 20154
rect 33816 20102 33826 20154
rect 33826 20102 33872 20154
rect 33576 20100 33632 20102
rect 33656 20100 33712 20102
rect 33736 20100 33792 20102
rect 33816 20100 33872 20102
rect 34150 19780 34206 19816
rect 34150 19760 34152 19780
rect 34152 19760 34204 19780
rect 34204 19760 34206 19780
rect 31758 17176 31760 17196
rect 31760 17176 31812 17196
rect 31812 17176 31814 17196
rect 31076 16346 31132 16348
rect 31156 16346 31212 16348
rect 31236 16346 31292 16348
rect 31316 16346 31372 16348
rect 31076 16294 31122 16346
rect 31122 16294 31132 16346
rect 31156 16294 31186 16346
rect 31186 16294 31198 16346
rect 31198 16294 31212 16346
rect 31236 16294 31250 16346
rect 31250 16294 31262 16346
rect 31262 16294 31292 16346
rect 31316 16294 31326 16346
rect 31326 16294 31372 16346
rect 31076 16292 31132 16294
rect 31156 16292 31212 16294
rect 31236 16292 31292 16294
rect 31316 16292 31372 16294
rect 31076 15258 31132 15260
rect 31156 15258 31212 15260
rect 31236 15258 31292 15260
rect 31316 15258 31372 15260
rect 31076 15206 31122 15258
rect 31122 15206 31132 15258
rect 31156 15206 31186 15258
rect 31186 15206 31198 15258
rect 31198 15206 31212 15258
rect 31236 15206 31250 15258
rect 31250 15206 31262 15258
rect 31262 15206 31292 15258
rect 31316 15206 31326 15258
rect 31326 15206 31372 15258
rect 31076 15204 31132 15206
rect 31156 15204 31212 15206
rect 31236 15204 31292 15206
rect 31316 15204 31372 15206
rect 30102 13232 30158 13288
rect 29918 12824 29974 12880
rect 29458 11328 29514 11384
rect 29366 10920 29422 10976
rect 28576 10362 28632 10364
rect 28656 10362 28712 10364
rect 28736 10362 28792 10364
rect 28816 10362 28872 10364
rect 28576 10310 28622 10362
rect 28622 10310 28632 10362
rect 28656 10310 28686 10362
rect 28686 10310 28698 10362
rect 28698 10310 28712 10362
rect 28736 10310 28750 10362
rect 28750 10310 28762 10362
rect 28762 10310 28792 10362
rect 28816 10310 28826 10362
rect 28826 10310 28872 10362
rect 28576 10308 28632 10310
rect 28656 10308 28712 10310
rect 28736 10308 28792 10310
rect 28816 10308 28872 10310
rect 28170 9560 28226 9616
rect 27986 8336 28042 8392
rect 28576 9274 28632 9276
rect 28656 9274 28712 9276
rect 28736 9274 28792 9276
rect 28816 9274 28872 9276
rect 28576 9222 28622 9274
rect 28622 9222 28632 9274
rect 28656 9222 28686 9274
rect 28686 9222 28698 9274
rect 28698 9222 28712 9274
rect 28736 9222 28750 9274
rect 28750 9222 28762 9274
rect 28762 9222 28792 9274
rect 28816 9222 28826 9274
rect 28826 9222 28872 9274
rect 28576 9220 28632 9222
rect 28656 9220 28712 9222
rect 28736 9220 28792 9222
rect 28816 9220 28872 9222
rect 28722 8472 28778 8528
rect 28538 8372 28540 8392
rect 28540 8372 28592 8392
rect 28592 8372 28594 8392
rect 27158 4800 27214 4856
rect 26076 3290 26132 3292
rect 26156 3290 26212 3292
rect 26236 3290 26292 3292
rect 26316 3290 26372 3292
rect 26076 3238 26122 3290
rect 26122 3238 26132 3290
rect 26156 3238 26186 3290
rect 26186 3238 26198 3290
rect 26198 3238 26212 3290
rect 26236 3238 26250 3290
rect 26250 3238 26262 3290
rect 26262 3238 26292 3290
rect 26316 3238 26326 3290
rect 26326 3238 26372 3290
rect 26076 3236 26132 3238
rect 26156 3236 26212 3238
rect 26236 3236 26292 3238
rect 26316 3236 26372 3238
rect 28538 8336 28594 8372
rect 28576 8186 28632 8188
rect 28656 8186 28712 8188
rect 28736 8186 28792 8188
rect 28816 8186 28872 8188
rect 28576 8134 28622 8186
rect 28622 8134 28632 8186
rect 28656 8134 28686 8186
rect 28686 8134 28698 8186
rect 28698 8134 28712 8186
rect 28736 8134 28750 8186
rect 28750 8134 28762 8186
rect 28762 8134 28792 8186
rect 28816 8134 28826 8186
rect 28826 8134 28872 8186
rect 28576 8132 28632 8134
rect 28656 8132 28712 8134
rect 28736 8132 28792 8134
rect 28816 8132 28872 8134
rect 28446 7928 28502 7984
rect 29366 10104 29422 10160
rect 29826 11500 29828 11520
rect 29828 11500 29880 11520
rect 29880 11500 29882 11520
rect 29826 11464 29882 11500
rect 29182 8336 29238 8392
rect 28576 7098 28632 7100
rect 28656 7098 28712 7100
rect 28736 7098 28792 7100
rect 28816 7098 28872 7100
rect 28576 7046 28622 7098
rect 28622 7046 28632 7098
rect 28656 7046 28686 7098
rect 28686 7046 28698 7098
rect 28698 7046 28712 7098
rect 28736 7046 28750 7098
rect 28750 7046 28762 7098
rect 28762 7046 28792 7098
rect 28816 7046 28826 7098
rect 28826 7046 28872 7098
rect 28576 7044 28632 7046
rect 28656 7044 28712 7046
rect 28736 7044 28792 7046
rect 28816 7044 28872 7046
rect 29550 9016 29606 9072
rect 31758 14884 31814 14920
rect 31758 14864 31760 14884
rect 31760 14864 31812 14884
rect 31812 14864 31814 14884
rect 31114 14320 31170 14376
rect 31076 14170 31132 14172
rect 31156 14170 31212 14172
rect 31236 14170 31292 14172
rect 31316 14170 31372 14172
rect 31076 14118 31122 14170
rect 31122 14118 31132 14170
rect 31156 14118 31186 14170
rect 31186 14118 31198 14170
rect 31198 14118 31212 14170
rect 31236 14118 31250 14170
rect 31250 14118 31262 14170
rect 31262 14118 31292 14170
rect 31316 14118 31326 14170
rect 31326 14118 31372 14170
rect 31076 14116 31132 14118
rect 31156 14116 31212 14118
rect 31236 14116 31292 14118
rect 31316 14116 31372 14118
rect 31076 13082 31132 13084
rect 31156 13082 31212 13084
rect 31236 13082 31292 13084
rect 31316 13082 31372 13084
rect 31076 13030 31122 13082
rect 31122 13030 31132 13082
rect 31156 13030 31186 13082
rect 31186 13030 31198 13082
rect 31198 13030 31212 13082
rect 31236 13030 31250 13082
rect 31250 13030 31262 13082
rect 31262 13030 31292 13082
rect 31316 13030 31326 13082
rect 31326 13030 31372 13082
rect 31076 13028 31132 13030
rect 31156 13028 31212 13030
rect 31236 13028 31292 13030
rect 31316 13028 31372 13030
rect 31076 11994 31132 11996
rect 31156 11994 31212 11996
rect 31236 11994 31292 11996
rect 31316 11994 31372 11996
rect 31076 11942 31122 11994
rect 31122 11942 31132 11994
rect 31156 11942 31186 11994
rect 31186 11942 31198 11994
rect 31198 11942 31212 11994
rect 31236 11942 31250 11994
rect 31250 11942 31262 11994
rect 31262 11942 31292 11994
rect 31316 11942 31326 11994
rect 31326 11942 31372 11994
rect 31076 11940 31132 11942
rect 31156 11940 31212 11942
rect 31236 11940 31292 11942
rect 31316 11940 31372 11942
rect 30838 11056 30894 11112
rect 31076 10906 31132 10908
rect 31156 10906 31212 10908
rect 31236 10906 31292 10908
rect 31316 10906 31372 10908
rect 31076 10854 31122 10906
rect 31122 10854 31132 10906
rect 31156 10854 31186 10906
rect 31186 10854 31198 10906
rect 31198 10854 31212 10906
rect 31236 10854 31250 10906
rect 31250 10854 31262 10906
rect 31262 10854 31292 10906
rect 31316 10854 31326 10906
rect 31326 10854 31372 10906
rect 31076 10852 31132 10854
rect 31156 10852 31212 10854
rect 31236 10852 31292 10854
rect 31316 10852 31372 10854
rect 30102 8880 30158 8936
rect 30470 9696 30526 9752
rect 30194 7928 30250 7984
rect 27434 4120 27490 4176
rect 28576 6010 28632 6012
rect 28656 6010 28712 6012
rect 28736 6010 28792 6012
rect 28816 6010 28872 6012
rect 28576 5958 28622 6010
rect 28622 5958 28632 6010
rect 28656 5958 28686 6010
rect 28686 5958 28698 6010
rect 28698 5958 28712 6010
rect 28736 5958 28750 6010
rect 28750 5958 28762 6010
rect 28762 5958 28792 6010
rect 28816 5958 28826 6010
rect 28826 5958 28872 6010
rect 28576 5956 28632 5958
rect 28656 5956 28712 5958
rect 28736 5956 28792 5958
rect 28816 5956 28872 5958
rect 28576 4922 28632 4924
rect 28656 4922 28712 4924
rect 28736 4922 28792 4924
rect 28816 4922 28872 4924
rect 28576 4870 28622 4922
rect 28622 4870 28632 4922
rect 28656 4870 28686 4922
rect 28686 4870 28698 4922
rect 28698 4870 28712 4922
rect 28736 4870 28750 4922
rect 28750 4870 28762 4922
rect 28762 4870 28792 4922
rect 28816 4870 28826 4922
rect 28826 4870 28872 4922
rect 28576 4868 28632 4870
rect 28656 4868 28712 4870
rect 28736 4868 28792 4870
rect 28816 4868 28872 4870
rect 28446 4684 28502 4720
rect 28446 4664 28448 4684
rect 28448 4664 28500 4684
rect 28500 4664 28502 4684
rect 28722 4528 28778 4584
rect 28576 3834 28632 3836
rect 28656 3834 28712 3836
rect 28736 3834 28792 3836
rect 28816 3834 28872 3836
rect 28576 3782 28622 3834
rect 28622 3782 28632 3834
rect 28656 3782 28686 3834
rect 28686 3782 28698 3834
rect 28698 3782 28712 3834
rect 28736 3782 28750 3834
rect 28750 3782 28762 3834
rect 28762 3782 28792 3834
rect 28816 3782 28826 3834
rect 28826 3782 28872 3834
rect 28576 3780 28632 3782
rect 28656 3780 28712 3782
rect 28736 3780 28792 3782
rect 28816 3780 28872 3782
rect 30470 7792 30526 7848
rect 30746 8880 30802 8936
rect 31076 9818 31132 9820
rect 31156 9818 31212 9820
rect 31236 9818 31292 9820
rect 31316 9818 31372 9820
rect 31076 9766 31122 9818
rect 31122 9766 31132 9818
rect 31156 9766 31186 9818
rect 31186 9766 31198 9818
rect 31198 9766 31212 9818
rect 31236 9766 31250 9818
rect 31250 9766 31262 9818
rect 31262 9766 31292 9818
rect 31316 9766 31326 9818
rect 31326 9766 31372 9818
rect 31076 9764 31132 9766
rect 31156 9764 31212 9766
rect 31236 9764 31292 9766
rect 31316 9764 31372 9766
rect 31206 9016 31262 9072
rect 31758 11348 31814 11384
rect 31758 11328 31760 11348
rect 31760 11328 31812 11348
rect 31812 11328 31814 11348
rect 31942 15000 31998 15056
rect 31942 12688 31998 12744
rect 31076 8730 31132 8732
rect 31156 8730 31212 8732
rect 31236 8730 31292 8732
rect 31316 8730 31372 8732
rect 31076 8678 31122 8730
rect 31122 8678 31132 8730
rect 31156 8678 31186 8730
rect 31186 8678 31198 8730
rect 31198 8678 31212 8730
rect 31236 8678 31250 8730
rect 31250 8678 31262 8730
rect 31262 8678 31292 8730
rect 31316 8678 31326 8730
rect 31326 8678 31372 8730
rect 31076 8676 31132 8678
rect 31156 8676 31212 8678
rect 31236 8676 31292 8678
rect 31316 8676 31372 8678
rect 30194 5752 30250 5808
rect 30838 7268 30894 7304
rect 30838 7248 30840 7268
rect 30840 7248 30892 7268
rect 30892 7248 30894 7268
rect 30010 4528 30066 4584
rect 31076 7642 31132 7644
rect 31156 7642 31212 7644
rect 31236 7642 31292 7644
rect 31316 7642 31372 7644
rect 31076 7590 31122 7642
rect 31122 7590 31132 7642
rect 31156 7590 31186 7642
rect 31186 7590 31198 7642
rect 31198 7590 31212 7642
rect 31236 7590 31250 7642
rect 31250 7590 31262 7642
rect 31262 7590 31292 7642
rect 31316 7590 31326 7642
rect 31326 7590 31372 7642
rect 31076 7588 31132 7590
rect 31156 7588 31212 7590
rect 31236 7588 31292 7590
rect 31316 7588 31372 7590
rect 31114 7384 31170 7440
rect 31022 6840 31078 6896
rect 31076 6554 31132 6556
rect 31156 6554 31212 6556
rect 31236 6554 31292 6556
rect 31316 6554 31372 6556
rect 31076 6502 31122 6554
rect 31122 6502 31132 6554
rect 31156 6502 31186 6554
rect 31186 6502 31198 6554
rect 31198 6502 31212 6554
rect 31236 6502 31250 6554
rect 31250 6502 31262 6554
rect 31262 6502 31292 6554
rect 31316 6502 31326 6554
rect 31326 6502 31372 6554
rect 31076 6500 31132 6502
rect 31156 6500 31212 6502
rect 31236 6500 31292 6502
rect 31316 6500 31372 6502
rect 31076 5466 31132 5468
rect 31156 5466 31212 5468
rect 31236 5466 31292 5468
rect 31316 5466 31372 5468
rect 31076 5414 31122 5466
rect 31122 5414 31132 5466
rect 31156 5414 31186 5466
rect 31186 5414 31198 5466
rect 31198 5414 31212 5466
rect 31236 5414 31250 5466
rect 31250 5414 31262 5466
rect 31262 5414 31292 5466
rect 31316 5414 31326 5466
rect 31326 5414 31372 5466
rect 31076 5412 31132 5414
rect 31156 5412 31212 5414
rect 31236 5412 31292 5414
rect 31316 5412 31372 5414
rect 32862 18128 32918 18184
rect 33576 19066 33632 19068
rect 33656 19066 33712 19068
rect 33736 19066 33792 19068
rect 33816 19066 33872 19068
rect 33576 19014 33622 19066
rect 33622 19014 33632 19066
rect 33656 19014 33686 19066
rect 33686 19014 33698 19066
rect 33698 19014 33712 19066
rect 33736 19014 33750 19066
rect 33750 19014 33762 19066
rect 33762 19014 33792 19066
rect 33816 19014 33826 19066
rect 33826 19014 33872 19066
rect 33576 19012 33632 19014
rect 33656 19012 33712 19014
rect 33736 19012 33792 19014
rect 33816 19012 33872 19014
rect 34334 20304 34390 20360
rect 34242 18672 34298 18728
rect 34242 18300 34244 18320
rect 34244 18300 34296 18320
rect 34296 18300 34298 18320
rect 34242 18264 34298 18300
rect 32862 17176 32918 17232
rect 32218 14864 32274 14920
rect 33576 17978 33632 17980
rect 33656 17978 33712 17980
rect 33736 17978 33792 17980
rect 33816 17978 33872 17980
rect 33576 17926 33622 17978
rect 33622 17926 33632 17978
rect 33656 17926 33686 17978
rect 33686 17926 33698 17978
rect 33698 17926 33712 17978
rect 33736 17926 33750 17978
rect 33750 17926 33762 17978
rect 33762 17926 33792 17978
rect 33816 17926 33826 17978
rect 33826 17926 33872 17978
rect 33576 17924 33632 17926
rect 33656 17924 33712 17926
rect 33736 17924 33792 17926
rect 33816 17924 33872 17926
rect 33576 16890 33632 16892
rect 33656 16890 33712 16892
rect 33736 16890 33792 16892
rect 33816 16890 33872 16892
rect 33576 16838 33622 16890
rect 33622 16838 33632 16890
rect 33656 16838 33686 16890
rect 33686 16838 33698 16890
rect 33698 16838 33712 16890
rect 33736 16838 33750 16890
rect 33750 16838 33762 16890
rect 33762 16838 33792 16890
rect 33816 16838 33826 16890
rect 33826 16838 33872 16890
rect 33576 16836 33632 16838
rect 33656 16836 33712 16838
rect 33736 16836 33792 16838
rect 33816 16836 33872 16838
rect 33690 16516 33746 16552
rect 33690 16496 33692 16516
rect 33692 16496 33744 16516
rect 33744 16496 33746 16516
rect 33576 15802 33632 15804
rect 33656 15802 33712 15804
rect 33736 15802 33792 15804
rect 33816 15802 33872 15804
rect 33576 15750 33622 15802
rect 33622 15750 33632 15802
rect 33656 15750 33686 15802
rect 33686 15750 33698 15802
rect 33698 15750 33712 15802
rect 33736 15750 33750 15802
rect 33750 15750 33762 15802
rect 33762 15750 33792 15802
rect 33816 15750 33826 15802
rect 33826 15750 33872 15802
rect 33576 15748 33632 15750
rect 33656 15748 33712 15750
rect 33736 15748 33792 15750
rect 33816 15748 33872 15750
rect 32954 13776 33010 13832
rect 32494 10920 32550 10976
rect 32310 10240 32366 10296
rect 32034 9580 32090 9616
rect 32034 9560 32036 9580
rect 32036 9560 32088 9580
rect 32088 9560 32090 9580
rect 32402 9968 32458 10024
rect 32494 8472 32550 8528
rect 31666 8200 31722 8256
rect 32126 8336 32182 8392
rect 32862 11464 32918 11520
rect 33576 14714 33632 14716
rect 33656 14714 33712 14716
rect 33736 14714 33792 14716
rect 33816 14714 33872 14716
rect 33576 14662 33622 14714
rect 33622 14662 33632 14714
rect 33656 14662 33686 14714
rect 33686 14662 33698 14714
rect 33698 14662 33712 14714
rect 33736 14662 33750 14714
rect 33750 14662 33762 14714
rect 33762 14662 33792 14714
rect 33816 14662 33826 14714
rect 33826 14662 33872 14714
rect 33576 14660 33632 14662
rect 33656 14660 33712 14662
rect 33736 14660 33792 14662
rect 33816 14660 33872 14662
rect 33230 13912 33286 13968
rect 33576 13626 33632 13628
rect 33656 13626 33712 13628
rect 33736 13626 33792 13628
rect 33816 13626 33872 13628
rect 33576 13574 33622 13626
rect 33622 13574 33632 13626
rect 33656 13574 33686 13626
rect 33686 13574 33698 13626
rect 33698 13574 33712 13626
rect 33736 13574 33750 13626
rect 33750 13574 33762 13626
rect 33762 13574 33792 13626
rect 33816 13574 33826 13626
rect 33826 13574 33872 13626
rect 33576 13572 33632 13574
rect 33656 13572 33712 13574
rect 33736 13572 33792 13574
rect 33816 13572 33872 13574
rect 33230 12860 33232 12880
rect 33232 12860 33284 12880
rect 33284 12860 33286 12880
rect 33230 12824 33286 12860
rect 33138 12688 33194 12744
rect 33322 12300 33378 12336
rect 33322 12280 33324 12300
rect 33324 12280 33376 12300
rect 33376 12280 33378 12300
rect 32954 10784 33010 10840
rect 32862 10240 32918 10296
rect 33322 10648 33378 10704
rect 32862 6296 32918 6352
rect 32218 5072 32274 5128
rect 29274 4256 29330 4312
rect 26076 2202 26132 2204
rect 26156 2202 26212 2204
rect 26236 2202 26292 2204
rect 26316 2202 26372 2204
rect 26076 2150 26122 2202
rect 26122 2150 26132 2202
rect 26156 2150 26186 2202
rect 26186 2150 26198 2202
rect 26198 2150 26212 2202
rect 26236 2150 26250 2202
rect 26250 2150 26262 2202
rect 26262 2150 26292 2202
rect 26316 2150 26326 2202
rect 26326 2150 26372 2202
rect 26076 2148 26132 2150
rect 26156 2148 26212 2150
rect 26236 2148 26292 2150
rect 26316 2148 26372 2150
rect 26882 2080 26938 2136
rect 26076 1114 26132 1116
rect 26156 1114 26212 1116
rect 26236 1114 26292 1116
rect 26316 1114 26372 1116
rect 26076 1062 26122 1114
rect 26122 1062 26132 1114
rect 26156 1062 26186 1114
rect 26186 1062 26198 1114
rect 26198 1062 26212 1114
rect 26236 1062 26250 1114
rect 26250 1062 26262 1114
rect 26262 1062 26292 1114
rect 26316 1062 26326 1114
rect 26326 1062 26372 1114
rect 26076 1060 26132 1062
rect 26156 1060 26212 1062
rect 26236 1060 26292 1062
rect 26316 1060 26372 1062
rect 27710 2508 27766 2544
rect 27710 2488 27712 2508
rect 27712 2488 27764 2508
rect 27764 2488 27766 2508
rect 28262 3032 28318 3088
rect 28078 2100 28134 2136
rect 28078 2080 28080 2100
rect 28080 2080 28132 2100
rect 28132 2080 28134 2100
rect 28354 2896 28410 2952
rect 28814 3168 28870 3224
rect 28576 2746 28632 2748
rect 28656 2746 28712 2748
rect 28736 2746 28792 2748
rect 28816 2746 28872 2748
rect 28576 2694 28622 2746
rect 28622 2694 28632 2746
rect 28656 2694 28686 2746
rect 28686 2694 28698 2746
rect 28698 2694 28712 2746
rect 28736 2694 28750 2746
rect 28750 2694 28762 2746
rect 28762 2694 28792 2746
rect 28816 2694 28826 2746
rect 28826 2694 28872 2746
rect 28576 2692 28632 2694
rect 28656 2692 28712 2694
rect 28736 2692 28792 2694
rect 28816 2692 28872 2694
rect 29274 3440 29330 3496
rect 28576 1658 28632 1660
rect 28656 1658 28712 1660
rect 28736 1658 28792 1660
rect 28816 1658 28872 1660
rect 28576 1606 28622 1658
rect 28622 1606 28632 1658
rect 28656 1606 28686 1658
rect 28686 1606 28698 1658
rect 28698 1606 28712 1658
rect 28736 1606 28750 1658
rect 28750 1606 28762 1658
rect 28762 1606 28792 1658
rect 28816 1606 28826 1658
rect 28826 1606 28872 1658
rect 28576 1604 28632 1606
rect 28656 1604 28712 1606
rect 28736 1604 28792 1606
rect 28816 1604 28872 1606
rect 31076 4378 31132 4380
rect 31156 4378 31212 4380
rect 31236 4378 31292 4380
rect 31316 4378 31372 4380
rect 31076 4326 31122 4378
rect 31122 4326 31132 4378
rect 31156 4326 31186 4378
rect 31186 4326 31198 4378
rect 31198 4326 31212 4378
rect 31236 4326 31250 4378
rect 31250 4326 31262 4378
rect 31262 4326 31292 4378
rect 31316 4326 31326 4378
rect 31326 4326 31372 4378
rect 31076 4324 31132 4326
rect 31156 4324 31212 4326
rect 31236 4324 31292 4326
rect 31316 4324 31372 4326
rect 30286 3168 30342 3224
rect 30378 2896 30434 2952
rect 33230 8780 33232 8800
rect 33232 8780 33284 8800
rect 33284 8780 33286 8800
rect 33230 8744 33286 8780
rect 33576 12538 33632 12540
rect 33656 12538 33712 12540
rect 33736 12538 33792 12540
rect 33816 12538 33872 12540
rect 33576 12486 33622 12538
rect 33622 12486 33632 12538
rect 33656 12486 33686 12538
rect 33686 12486 33698 12538
rect 33698 12486 33712 12538
rect 33736 12486 33750 12538
rect 33750 12486 33762 12538
rect 33762 12486 33792 12538
rect 33816 12486 33826 12538
rect 33826 12486 33872 12538
rect 33576 12484 33632 12486
rect 33656 12484 33712 12486
rect 33736 12484 33792 12486
rect 33816 12484 33872 12486
rect 34702 20848 34758 20904
rect 35438 22108 35440 22128
rect 35440 22108 35492 22128
rect 35492 22108 35494 22128
rect 35438 22072 35494 22108
rect 35162 18808 35218 18864
rect 36076 21786 36132 21788
rect 36156 21786 36212 21788
rect 36236 21786 36292 21788
rect 36316 21786 36372 21788
rect 36076 21734 36122 21786
rect 36122 21734 36132 21786
rect 36156 21734 36186 21786
rect 36186 21734 36198 21786
rect 36198 21734 36212 21786
rect 36236 21734 36250 21786
rect 36250 21734 36262 21786
rect 36262 21734 36292 21786
rect 36316 21734 36326 21786
rect 36326 21734 36372 21786
rect 36076 21732 36132 21734
rect 36156 21732 36212 21734
rect 36236 21732 36292 21734
rect 36316 21732 36372 21734
rect 36634 21528 36690 21584
rect 36076 20698 36132 20700
rect 36156 20698 36212 20700
rect 36236 20698 36292 20700
rect 36316 20698 36372 20700
rect 36076 20646 36122 20698
rect 36122 20646 36132 20698
rect 36156 20646 36186 20698
rect 36186 20646 36198 20698
rect 36198 20646 36212 20698
rect 36236 20646 36250 20698
rect 36250 20646 36262 20698
rect 36262 20646 36292 20698
rect 36316 20646 36326 20698
rect 36326 20646 36372 20698
rect 36076 20644 36132 20646
rect 36156 20644 36212 20646
rect 36236 20644 36292 20646
rect 36316 20644 36372 20646
rect 36076 19610 36132 19612
rect 36156 19610 36212 19612
rect 36236 19610 36292 19612
rect 36316 19610 36372 19612
rect 36076 19558 36122 19610
rect 36122 19558 36132 19610
rect 36156 19558 36186 19610
rect 36186 19558 36198 19610
rect 36198 19558 36212 19610
rect 36236 19558 36250 19610
rect 36250 19558 36262 19610
rect 36262 19558 36292 19610
rect 36316 19558 36326 19610
rect 36326 19558 36372 19610
rect 36076 19556 36132 19558
rect 36156 19556 36212 19558
rect 36236 19556 36292 19558
rect 36316 19556 36372 19558
rect 36076 18522 36132 18524
rect 36156 18522 36212 18524
rect 36236 18522 36292 18524
rect 36316 18522 36372 18524
rect 36076 18470 36122 18522
rect 36122 18470 36132 18522
rect 36156 18470 36186 18522
rect 36186 18470 36198 18522
rect 36198 18470 36212 18522
rect 36236 18470 36250 18522
rect 36250 18470 36262 18522
rect 36262 18470 36292 18522
rect 36316 18470 36326 18522
rect 36326 18470 36372 18522
rect 36076 18468 36132 18470
rect 36156 18468 36212 18470
rect 36236 18468 36292 18470
rect 36316 18468 36372 18470
rect 33506 11736 33562 11792
rect 33576 11450 33632 11452
rect 33656 11450 33712 11452
rect 33736 11450 33792 11452
rect 33816 11450 33872 11452
rect 33576 11398 33622 11450
rect 33622 11398 33632 11450
rect 33656 11398 33686 11450
rect 33686 11398 33698 11450
rect 33698 11398 33712 11450
rect 33736 11398 33750 11450
rect 33750 11398 33762 11450
rect 33762 11398 33792 11450
rect 33816 11398 33826 11450
rect 33826 11398 33872 11450
rect 33576 11396 33632 11398
rect 33656 11396 33712 11398
rect 33736 11396 33792 11398
rect 33816 11396 33872 11398
rect 33966 10920 34022 10976
rect 33576 10362 33632 10364
rect 33656 10362 33712 10364
rect 33736 10362 33792 10364
rect 33816 10362 33872 10364
rect 33576 10310 33622 10362
rect 33622 10310 33632 10362
rect 33656 10310 33686 10362
rect 33686 10310 33698 10362
rect 33698 10310 33712 10362
rect 33736 10310 33750 10362
rect 33750 10310 33762 10362
rect 33762 10310 33792 10362
rect 33816 10310 33826 10362
rect 33826 10310 33872 10362
rect 33576 10308 33632 10310
rect 33656 10308 33712 10310
rect 33736 10308 33792 10310
rect 33816 10308 33872 10310
rect 33506 10104 33562 10160
rect 33598 9968 33654 10024
rect 37830 21392 37886 21448
rect 37830 20984 37886 21040
rect 38014 20440 38070 20496
rect 38576 22330 38632 22332
rect 38656 22330 38712 22332
rect 38736 22330 38792 22332
rect 38816 22330 38872 22332
rect 38576 22278 38622 22330
rect 38622 22278 38632 22330
rect 38656 22278 38686 22330
rect 38686 22278 38698 22330
rect 38698 22278 38712 22330
rect 38736 22278 38750 22330
rect 38750 22278 38762 22330
rect 38762 22278 38792 22330
rect 38816 22278 38826 22330
rect 38826 22278 38872 22330
rect 38576 22276 38632 22278
rect 38656 22276 38712 22278
rect 38736 22276 38792 22278
rect 38816 22276 38872 22278
rect 38576 21242 38632 21244
rect 38656 21242 38712 21244
rect 38736 21242 38792 21244
rect 38816 21242 38872 21244
rect 38576 21190 38622 21242
rect 38622 21190 38632 21242
rect 38656 21190 38686 21242
rect 38686 21190 38698 21242
rect 38698 21190 38712 21242
rect 38736 21190 38750 21242
rect 38750 21190 38762 21242
rect 38762 21190 38792 21242
rect 38816 21190 38826 21242
rect 38826 21190 38872 21242
rect 38576 21188 38632 21190
rect 38656 21188 38712 21190
rect 38736 21188 38792 21190
rect 38816 21188 38872 21190
rect 38576 20154 38632 20156
rect 38656 20154 38712 20156
rect 38736 20154 38792 20156
rect 38816 20154 38872 20156
rect 38576 20102 38622 20154
rect 38622 20102 38632 20154
rect 38656 20102 38686 20154
rect 38686 20102 38698 20154
rect 38698 20102 38712 20154
rect 38736 20102 38750 20154
rect 38750 20102 38762 20154
rect 38762 20102 38792 20154
rect 38816 20102 38826 20154
rect 38826 20102 38872 20154
rect 38576 20100 38632 20102
rect 38656 20100 38712 20102
rect 38736 20100 38792 20102
rect 38816 20100 38872 20102
rect 38750 19796 38752 19816
rect 38752 19796 38804 19816
rect 38804 19796 38806 19816
rect 38750 19760 38806 19796
rect 38934 19216 38990 19272
rect 38576 19066 38632 19068
rect 38656 19066 38712 19068
rect 38736 19066 38792 19068
rect 38816 19066 38872 19068
rect 38576 19014 38622 19066
rect 38622 19014 38632 19066
rect 38656 19014 38686 19066
rect 38686 19014 38698 19066
rect 38698 19014 38712 19066
rect 38736 19014 38750 19066
rect 38750 19014 38762 19066
rect 38762 19014 38792 19066
rect 38816 19014 38826 19066
rect 38826 19014 38872 19066
rect 38576 19012 38632 19014
rect 38656 19012 38712 19014
rect 38736 19012 38792 19014
rect 38816 19012 38872 19014
rect 37738 17720 37794 17776
rect 36076 17434 36132 17436
rect 36156 17434 36212 17436
rect 36236 17434 36292 17436
rect 36316 17434 36372 17436
rect 36076 17382 36122 17434
rect 36122 17382 36132 17434
rect 36156 17382 36186 17434
rect 36186 17382 36198 17434
rect 36198 17382 36212 17434
rect 36236 17382 36250 17434
rect 36250 17382 36262 17434
rect 36262 17382 36292 17434
rect 36316 17382 36326 17434
rect 36326 17382 36372 17434
rect 36076 17380 36132 17382
rect 36156 17380 36212 17382
rect 36236 17380 36292 17382
rect 36316 17380 36372 17382
rect 34242 12144 34298 12200
rect 34886 13232 34942 13288
rect 33598 9424 33654 9480
rect 33576 9274 33632 9276
rect 33656 9274 33712 9276
rect 33736 9274 33792 9276
rect 33816 9274 33872 9276
rect 33576 9222 33622 9274
rect 33622 9222 33632 9274
rect 33656 9222 33686 9274
rect 33686 9222 33698 9274
rect 33698 9222 33712 9274
rect 33736 9222 33750 9274
rect 33750 9222 33762 9274
rect 33762 9222 33792 9274
rect 33816 9222 33826 9274
rect 33826 9222 33872 9274
rect 33576 9220 33632 9222
rect 33656 9220 33712 9222
rect 33736 9220 33792 9222
rect 33816 9220 33872 9222
rect 34058 9152 34114 9208
rect 33506 8880 33562 8936
rect 33322 8336 33378 8392
rect 33576 8186 33632 8188
rect 33656 8186 33712 8188
rect 33736 8186 33792 8188
rect 33816 8186 33872 8188
rect 33576 8134 33622 8186
rect 33622 8134 33632 8186
rect 33656 8134 33686 8186
rect 33686 8134 33698 8186
rect 33698 8134 33712 8186
rect 33736 8134 33750 8186
rect 33750 8134 33762 8186
rect 33762 8134 33792 8186
rect 33816 8134 33826 8186
rect 33826 8134 33872 8186
rect 33576 8132 33632 8134
rect 33656 8132 33712 8134
rect 33736 8132 33792 8134
rect 33816 8132 33872 8134
rect 33576 7098 33632 7100
rect 33656 7098 33712 7100
rect 33736 7098 33792 7100
rect 33816 7098 33872 7100
rect 33576 7046 33622 7098
rect 33622 7046 33632 7098
rect 33656 7046 33686 7098
rect 33686 7046 33698 7098
rect 33698 7046 33712 7098
rect 33736 7046 33750 7098
rect 33750 7046 33762 7098
rect 33762 7046 33792 7098
rect 33816 7046 33826 7098
rect 33826 7046 33872 7098
rect 33576 7044 33632 7046
rect 33656 7044 33712 7046
rect 33736 7044 33792 7046
rect 33816 7044 33872 7046
rect 34334 8628 34390 8664
rect 34334 8608 34336 8628
rect 34336 8608 34388 8628
rect 34388 8608 34390 8628
rect 34426 8336 34482 8392
rect 33782 6296 33838 6352
rect 33230 5616 33286 5672
rect 33576 6010 33632 6012
rect 33656 6010 33712 6012
rect 33736 6010 33792 6012
rect 33816 6010 33872 6012
rect 33576 5958 33622 6010
rect 33622 5958 33632 6010
rect 33656 5958 33686 6010
rect 33686 5958 33698 6010
rect 33698 5958 33712 6010
rect 33736 5958 33750 6010
rect 33750 5958 33762 6010
rect 33762 5958 33792 6010
rect 33816 5958 33826 6010
rect 33826 5958 33872 6010
rect 33576 5956 33632 5958
rect 33656 5956 33712 5958
rect 33736 5956 33792 5958
rect 33816 5956 33872 5958
rect 34702 11600 34758 11656
rect 34794 10784 34850 10840
rect 34702 9560 34758 9616
rect 36076 16346 36132 16348
rect 36156 16346 36212 16348
rect 36236 16346 36292 16348
rect 36316 16346 36372 16348
rect 36076 16294 36122 16346
rect 36122 16294 36132 16346
rect 36156 16294 36186 16346
rect 36186 16294 36198 16346
rect 36198 16294 36212 16346
rect 36236 16294 36250 16346
rect 36250 16294 36262 16346
rect 36262 16294 36292 16346
rect 36316 16294 36326 16346
rect 36326 16294 36372 16346
rect 36076 16292 36132 16294
rect 36156 16292 36212 16294
rect 36236 16292 36292 16294
rect 36316 16292 36372 16294
rect 36076 15258 36132 15260
rect 36156 15258 36212 15260
rect 36236 15258 36292 15260
rect 36316 15258 36372 15260
rect 36076 15206 36122 15258
rect 36122 15206 36132 15258
rect 36156 15206 36186 15258
rect 36186 15206 36198 15258
rect 36198 15206 36212 15258
rect 36236 15206 36250 15258
rect 36250 15206 36262 15258
rect 36262 15206 36292 15258
rect 36316 15206 36326 15258
rect 36326 15206 36372 15258
rect 36076 15204 36132 15206
rect 36156 15204 36212 15206
rect 36236 15204 36292 15206
rect 36316 15204 36372 15206
rect 36818 14884 36874 14920
rect 36818 14864 36820 14884
rect 36820 14864 36872 14884
rect 36872 14864 36874 14884
rect 37278 15408 37334 15464
rect 37830 15408 37886 15464
rect 36076 14170 36132 14172
rect 36156 14170 36212 14172
rect 36236 14170 36292 14172
rect 36316 14170 36372 14172
rect 36076 14118 36122 14170
rect 36122 14118 36132 14170
rect 36156 14118 36186 14170
rect 36186 14118 36198 14170
rect 36198 14118 36212 14170
rect 36236 14118 36250 14170
rect 36250 14118 36262 14170
rect 36262 14118 36292 14170
rect 36316 14118 36326 14170
rect 36326 14118 36372 14170
rect 36076 14116 36132 14118
rect 36156 14116 36212 14118
rect 36236 14116 36292 14118
rect 36316 14116 36372 14118
rect 36076 13082 36132 13084
rect 36156 13082 36212 13084
rect 36236 13082 36292 13084
rect 36316 13082 36372 13084
rect 36076 13030 36122 13082
rect 36122 13030 36132 13082
rect 36156 13030 36186 13082
rect 36186 13030 36198 13082
rect 36198 13030 36212 13082
rect 36236 13030 36250 13082
rect 36250 13030 36262 13082
rect 36262 13030 36292 13082
rect 36316 13030 36326 13082
rect 36326 13030 36372 13082
rect 36076 13028 36132 13030
rect 36156 13028 36212 13030
rect 36236 13028 36292 13030
rect 36316 13028 36372 13030
rect 36634 12144 36690 12200
rect 36076 11994 36132 11996
rect 36156 11994 36212 11996
rect 36236 11994 36292 11996
rect 36316 11994 36372 11996
rect 36076 11942 36122 11994
rect 36122 11942 36132 11994
rect 36156 11942 36186 11994
rect 36186 11942 36198 11994
rect 36198 11942 36212 11994
rect 36236 11942 36250 11994
rect 36250 11942 36262 11994
rect 36262 11942 36292 11994
rect 36316 11942 36326 11994
rect 36326 11942 36372 11994
rect 36076 11940 36132 11942
rect 36156 11940 36212 11942
rect 36236 11940 36292 11942
rect 36316 11940 36372 11942
rect 36076 10906 36132 10908
rect 36156 10906 36212 10908
rect 36236 10906 36292 10908
rect 36316 10906 36372 10908
rect 36076 10854 36122 10906
rect 36122 10854 36132 10906
rect 36156 10854 36186 10906
rect 36186 10854 36198 10906
rect 36198 10854 36212 10906
rect 36236 10854 36250 10906
rect 36250 10854 36262 10906
rect 36262 10854 36292 10906
rect 36316 10854 36326 10906
rect 36326 10854 36372 10906
rect 36076 10852 36132 10854
rect 36156 10852 36212 10854
rect 36236 10852 36292 10854
rect 36316 10852 36372 10854
rect 37462 12280 37518 12336
rect 36818 10648 36874 10704
rect 36076 9818 36132 9820
rect 36156 9818 36212 9820
rect 36236 9818 36292 9820
rect 36316 9818 36372 9820
rect 36076 9766 36122 9818
rect 36122 9766 36132 9818
rect 36156 9766 36186 9818
rect 36186 9766 36198 9818
rect 36198 9766 36212 9818
rect 36236 9766 36250 9818
rect 36250 9766 36262 9818
rect 36262 9766 36292 9818
rect 36316 9766 36326 9818
rect 36326 9766 36372 9818
rect 36076 9764 36132 9766
rect 36156 9764 36212 9766
rect 36236 9764 36292 9766
rect 36316 9764 36372 9766
rect 31850 3576 31906 3632
rect 31298 3440 31354 3496
rect 31076 3290 31132 3292
rect 31156 3290 31212 3292
rect 31236 3290 31292 3292
rect 31316 3290 31372 3292
rect 31076 3238 31122 3290
rect 31122 3238 31132 3290
rect 31156 3238 31186 3290
rect 31186 3238 31198 3290
rect 31198 3238 31212 3290
rect 31236 3238 31250 3290
rect 31250 3238 31262 3290
rect 31262 3238 31292 3290
rect 31316 3238 31326 3290
rect 31326 3238 31372 3290
rect 31076 3236 31132 3238
rect 31156 3236 31212 3238
rect 31236 3236 31292 3238
rect 31316 3236 31372 3238
rect 31206 2624 31262 2680
rect 31390 2372 31446 2408
rect 31390 2352 31392 2372
rect 31392 2352 31444 2372
rect 31444 2352 31446 2372
rect 31076 2202 31132 2204
rect 31156 2202 31212 2204
rect 31236 2202 31292 2204
rect 31316 2202 31372 2204
rect 31076 2150 31122 2202
rect 31122 2150 31132 2202
rect 31156 2150 31186 2202
rect 31186 2150 31198 2202
rect 31198 2150 31212 2202
rect 31236 2150 31250 2202
rect 31250 2150 31262 2202
rect 31262 2150 31292 2202
rect 31316 2150 31326 2202
rect 31326 2150 31372 2202
rect 31076 2148 31132 2150
rect 31156 2148 31212 2150
rect 31236 2148 31292 2150
rect 31316 2148 31372 2150
rect 30470 1400 30526 1456
rect 31942 2624 31998 2680
rect 32034 2352 32090 2408
rect 31942 1964 31998 2000
rect 31942 1944 31944 1964
rect 31944 1944 31996 1964
rect 31996 1944 31998 1964
rect 31076 1114 31132 1116
rect 31156 1114 31212 1116
rect 31236 1114 31292 1116
rect 31316 1114 31372 1116
rect 31076 1062 31122 1114
rect 31122 1062 31132 1114
rect 31156 1062 31186 1114
rect 31186 1062 31198 1114
rect 31198 1062 31212 1114
rect 31236 1062 31250 1114
rect 31250 1062 31262 1114
rect 31262 1062 31292 1114
rect 31316 1062 31326 1114
rect 31326 1062 31372 1114
rect 31076 1060 31132 1062
rect 31156 1060 31212 1062
rect 31236 1060 31292 1062
rect 31316 1060 31372 1062
rect 33576 4922 33632 4924
rect 33656 4922 33712 4924
rect 33736 4922 33792 4924
rect 33816 4922 33872 4924
rect 33576 4870 33622 4922
rect 33622 4870 33632 4922
rect 33656 4870 33686 4922
rect 33686 4870 33698 4922
rect 33698 4870 33712 4922
rect 33736 4870 33750 4922
rect 33750 4870 33762 4922
rect 33762 4870 33792 4922
rect 33816 4870 33826 4922
rect 33826 4870 33872 4922
rect 33576 4868 33632 4870
rect 33656 4868 33712 4870
rect 33736 4868 33792 4870
rect 33816 4868 33872 4870
rect 33966 4800 34022 4856
rect 35530 9036 35586 9072
rect 35530 9016 35532 9036
rect 35532 9016 35584 9036
rect 35584 9016 35586 9036
rect 36082 9152 36138 9208
rect 34886 8744 34942 8800
rect 34886 8608 34942 8664
rect 35346 8336 35402 8392
rect 33576 3834 33632 3836
rect 33656 3834 33712 3836
rect 33736 3834 33792 3836
rect 33816 3834 33872 3836
rect 33576 3782 33622 3834
rect 33622 3782 33632 3834
rect 33656 3782 33686 3834
rect 33686 3782 33698 3834
rect 33698 3782 33712 3834
rect 33736 3782 33750 3834
rect 33750 3782 33762 3834
rect 33762 3782 33792 3834
rect 33816 3782 33826 3834
rect 33826 3782 33872 3834
rect 33576 3780 33632 3782
rect 33656 3780 33712 3782
rect 33736 3780 33792 3782
rect 33816 3780 33872 3782
rect 32586 2896 32642 2952
rect 32494 2624 32550 2680
rect 33690 3460 33746 3496
rect 33690 3440 33692 3460
rect 33692 3440 33744 3460
rect 33744 3440 33746 3460
rect 32770 2352 32826 2408
rect 33576 2746 33632 2748
rect 33656 2746 33712 2748
rect 33736 2746 33792 2748
rect 33816 2746 33872 2748
rect 33576 2694 33622 2746
rect 33622 2694 33632 2746
rect 33656 2694 33686 2746
rect 33686 2694 33698 2746
rect 33698 2694 33712 2746
rect 33736 2694 33750 2746
rect 33750 2694 33762 2746
rect 33762 2694 33792 2746
rect 33816 2694 33826 2746
rect 33826 2694 33872 2746
rect 33576 2692 33632 2694
rect 33656 2692 33712 2694
rect 33736 2692 33792 2694
rect 33816 2692 33872 2694
rect 33782 1964 33838 2000
rect 33782 1944 33784 1964
rect 33784 1944 33836 1964
rect 33836 1944 33838 1964
rect 33576 1658 33632 1660
rect 33656 1658 33712 1660
rect 33736 1658 33792 1660
rect 33816 1658 33872 1660
rect 33576 1606 33622 1658
rect 33622 1606 33632 1658
rect 33656 1606 33686 1658
rect 33686 1606 33698 1658
rect 33698 1606 33712 1658
rect 33736 1606 33750 1658
rect 33750 1606 33762 1658
rect 33762 1606 33792 1658
rect 33816 1606 33826 1658
rect 33826 1606 33872 1658
rect 33576 1604 33632 1606
rect 33656 1604 33712 1606
rect 33736 1604 33792 1606
rect 33816 1604 33872 1606
rect 35162 7384 35218 7440
rect 33874 1300 33876 1320
rect 33876 1300 33928 1320
rect 33928 1300 33930 1320
rect 33874 1264 33930 1300
rect 35254 2760 35310 2816
rect 36174 8900 36230 8936
rect 36174 8880 36176 8900
rect 36176 8880 36228 8900
rect 36228 8880 36230 8900
rect 36076 8730 36132 8732
rect 36156 8730 36212 8732
rect 36236 8730 36292 8732
rect 36316 8730 36372 8732
rect 36076 8678 36122 8730
rect 36122 8678 36132 8730
rect 36156 8678 36186 8730
rect 36186 8678 36198 8730
rect 36198 8678 36212 8730
rect 36236 8678 36250 8730
rect 36250 8678 36262 8730
rect 36262 8678 36292 8730
rect 36316 8678 36326 8730
rect 36326 8678 36372 8730
rect 36076 8676 36132 8678
rect 36156 8676 36212 8678
rect 36236 8676 36292 8678
rect 36316 8676 36372 8678
rect 35714 6704 35770 6760
rect 36542 8472 36598 8528
rect 36174 8336 36230 8392
rect 37738 10512 37794 10568
rect 36634 7928 36690 7984
rect 36076 7642 36132 7644
rect 36156 7642 36212 7644
rect 36236 7642 36292 7644
rect 36316 7642 36372 7644
rect 36076 7590 36122 7642
rect 36122 7590 36132 7642
rect 36156 7590 36186 7642
rect 36186 7590 36198 7642
rect 36198 7590 36212 7642
rect 36236 7590 36250 7642
rect 36250 7590 36262 7642
rect 36262 7590 36292 7642
rect 36316 7590 36326 7642
rect 36326 7590 36372 7642
rect 36076 7588 36132 7590
rect 36156 7588 36212 7590
rect 36236 7588 36292 7590
rect 36316 7588 36372 7590
rect 35898 7248 35954 7304
rect 35990 6740 35992 6760
rect 35992 6740 36044 6760
rect 36044 6740 36046 6760
rect 35990 6704 36046 6740
rect 37738 7928 37794 7984
rect 41076 22874 41132 22876
rect 41156 22874 41212 22876
rect 41236 22874 41292 22876
rect 41316 22874 41372 22876
rect 41076 22822 41122 22874
rect 41122 22822 41132 22874
rect 41156 22822 41186 22874
rect 41186 22822 41198 22874
rect 41198 22822 41212 22874
rect 41236 22822 41250 22874
rect 41250 22822 41262 22874
rect 41262 22822 41292 22874
rect 41316 22822 41326 22874
rect 41326 22822 41372 22874
rect 41076 22820 41132 22822
rect 41156 22820 41212 22822
rect 41236 22820 41292 22822
rect 41316 22820 41372 22822
rect 41076 21786 41132 21788
rect 41156 21786 41212 21788
rect 41236 21786 41292 21788
rect 41316 21786 41372 21788
rect 41076 21734 41122 21786
rect 41122 21734 41132 21786
rect 41156 21734 41186 21786
rect 41186 21734 41198 21786
rect 41198 21734 41212 21786
rect 41236 21734 41250 21786
rect 41250 21734 41262 21786
rect 41262 21734 41292 21786
rect 41316 21734 41326 21786
rect 41326 21734 41372 21786
rect 41076 21732 41132 21734
rect 41156 21732 41212 21734
rect 41236 21732 41292 21734
rect 41316 21732 41372 21734
rect 38576 17978 38632 17980
rect 38656 17978 38712 17980
rect 38736 17978 38792 17980
rect 38816 17978 38872 17980
rect 38576 17926 38622 17978
rect 38622 17926 38632 17978
rect 38656 17926 38686 17978
rect 38686 17926 38698 17978
rect 38698 17926 38712 17978
rect 38736 17926 38750 17978
rect 38750 17926 38762 17978
rect 38762 17926 38792 17978
rect 38816 17926 38826 17978
rect 38826 17926 38872 17978
rect 38576 17924 38632 17926
rect 38656 17924 38712 17926
rect 38736 17924 38792 17926
rect 38816 17924 38872 17926
rect 41076 20698 41132 20700
rect 41156 20698 41212 20700
rect 41236 20698 41292 20700
rect 41316 20698 41372 20700
rect 41076 20646 41122 20698
rect 41122 20646 41132 20698
rect 41156 20646 41186 20698
rect 41186 20646 41198 20698
rect 41198 20646 41212 20698
rect 41236 20646 41250 20698
rect 41250 20646 41262 20698
rect 41262 20646 41292 20698
rect 41316 20646 41326 20698
rect 41326 20646 41372 20698
rect 41076 20644 41132 20646
rect 41156 20644 41212 20646
rect 41236 20644 41292 20646
rect 41316 20644 41372 20646
rect 41076 19610 41132 19612
rect 41156 19610 41212 19612
rect 41236 19610 41292 19612
rect 41316 19610 41372 19612
rect 41076 19558 41122 19610
rect 41122 19558 41132 19610
rect 41156 19558 41186 19610
rect 41186 19558 41198 19610
rect 41198 19558 41212 19610
rect 41236 19558 41250 19610
rect 41250 19558 41262 19610
rect 41262 19558 41292 19610
rect 41316 19558 41326 19610
rect 41326 19558 41372 19610
rect 41076 19556 41132 19558
rect 41156 19556 41212 19558
rect 41236 19556 41292 19558
rect 41316 19556 41372 19558
rect 41878 20848 41934 20904
rect 41076 18522 41132 18524
rect 41156 18522 41212 18524
rect 41236 18522 41292 18524
rect 41316 18522 41372 18524
rect 41076 18470 41122 18522
rect 41122 18470 41132 18522
rect 41156 18470 41186 18522
rect 41186 18470 41198 18522
rect 41198 18470 41212 18522
rect 41236 18470 41250 18522
rect 41250 18470 41262 18522
rect 41262 18470 41292 18522
rect 41316 18470 41326 18522
rect 41326 18470 41372 18522
rect 41076 18468 41132 18470
rect 41156 18468 41212 18470
rect 41236 18468 41292 18470
rect 41316 18468 41372 18470
rect 40038 17720 40094 17776
rect 38576 16890 38632 16892
rect 38656 16890 38712 16892
rect 38736 16890 38792 16892
rect 38816 16890 38872 16892
rect 38576 16838 38622 16890
rect 38622 16838 38632 16890
rect 38656 16838 38686 16890
rect 38686 16838 38698 16890
rect 38698 16838 38712 16890
rect 38736 16838 38750 16890
rect 38750 16838 38762 16890
rect 38762 16838 38792 16890
rect 38816 16838 38826 16890
rect 38826 16838 38872 16890
rect 38576 16836 38632 16838
rect 38656 16836 38712 16838
rect 38736 16836 38792 16838
rect 38816 16836 38872 16838
rect 39118 16532 39120 16552
rect 39120 16532 39172 16552
rect 39172 16532 39174 16552
rect 39118 16496 39174 16532
rect 38576 15802 38632 15804
rect 38656 15802 38712 15804
rect 38736 15802 38792 15804
rect 38816 15802 38872 15804
rect 38576 15750 38622 15802
rect 38622 15750 38632 15802
rect 38656 15750 38686 15802
rect 38686 15750 38698 15802
rect 38698 15750 38712 15802
rect 38736 15750 38750 15802
rect 38750 15750 38762 15802
rect 38762 15750 38792 15802
rect 38816 15750 38826 15802
rect 38826 15750 38872 15802
rect 38576 15748 38632 15750
rect 38656 15748 38712 15750
rect 38736 15748 38792 15750
rect 38816 15748 38872 15750
rect 38576 14714 38632 14716
rect 38656 14714 38712 14716
rect 38736 14714 38792 14716
rect 38816 14714 38872 14716
rect 38576 14662 38622 14714
rect 38622 14662 38632 14714
rect 38656 14662 38686 14714
rect 38686 14662 38698 14714
rect 38698 14662 38712 14714
rect 38736 14662 38750 14714
rect 38750 14662 38762 14714
rect 38762 14662 38792 14714
rect 38816 14662 38826 14714
rect 38826 14662 38872 14714
rect 38576 14660 38632 14662
rect 38656 14660 38712 14662
rect 38736 14660 38792 14662
rect 38816 14660 38872 14662
rect 38576 13626 38632 13628
rect 38656 13626 38712 13628
rect 38736 13626 38792 13628
rect 38816 13626 38872 13628
rect 38576 13574 38622 13626
rect 38622 13574 38632 13626
rect 38656 13574 38686 13626
rect 38686 13574 38698 13626
rect 38698 13574 38712 13626
rect 38736 13574 38750 13626
rect 38750 13574 38762 13626
rect 38762 13574 38792 13626
rect 38816 13574 38826 13626
rect 38826 13574 38872 13626
rect 38576 13572 38632 13574
rect 38656 13572 38712 13574
rect 38736 13572 38792 13574
rect 38816 13572 38872 13574
rect 38576 12538 38632 12540
rect 38656 12538 38712 12540
rect 38736 12538 38792 12540
rect 38816 12538 38872 12540
rect 38576 12486 38622 12538
rect 38622 12486 38632 12538
rect 38656 12486 38686 12538
rect 38686 12486 38698 12538
rect 38698 12486 38712 12538
rect 38736 12486 38750 12538
rect 38750 12486 38762 12538
rect 38762 12486 38792 12538
rect 38816 12486 38826 12538
rect 38826 12486 38872 12538
rect 38576 12484 38632 12486
rect 38656 12484 38712 12486
rect 38736 12484 38792 12486
rect 38816 12484 38872 12486
rect 38576 11450 38632 11452
rect 38656 11450 38712 11452
rect 38736 11450 38792 11452
rect 38816 11450 38872 11452
rect 38576 11398 38622 11450
rect 38622 11398 38632 11450
rect 38656 11398 38686 11450
rect 38686 11398 38698 11450
rect 38698 11398 38712 11450
rect 38736 11398 38750 11450
rect 38750 11398 38762 11450
rect 38762 11398 38792 11450
rect 38816 11398 38826 11450
rect 38826 11398 38872 11450
rect 38576 11396 38632 11398
rect 38656 11396 38712 11398
rect 38736 11396 38792 11398
rect 38816 11396 38872 11398
rect 38576 10362 38632 10364
rect 38656 10362 38712 10364
rect 38736 10362 38792 10364
rect 38816 10362 38872 10364
rect 38576 10310 38622 10362
rect 38622 10310 38632 10362
rect 38656 10310 38686 10362
rect 38686 10310 38698 10362
rect 38698 10310 38712 10362
rect 38736 10310 38750 10362
rect 38750 10310 38762 10362
rect 38762 10310 38792 10362
rect 38816 10310 38826 10362
rect 38826 10310 38872 10362
rect 38576 10308 38632 10310
rect 38656 10308 38712 10310
rect 38736 10308 38792 10310
rect 38816 10308 38872 10310
rect 41076 17434 41132 17436
rect 41156 17434 41212 17436
rect 41236 17434 41292 17436
rect 41316 17434 41372 17436
rect 41076 17382 41122 17434
rect 41122 17382 41132 17434
rect 41156 17382 41186 17434
rect 41186 17382 41198 17434
rect 41198 17382 41212 17434
rect 41236 17382 41250 17434
rect 41250 17382 41262 17434
rect 41262 17382 41292 17434
rect 41316 17382 41326 17434
rect 41326 17382 41372 17434
rect 41076 17380 41132 17382
rect 41156 17380 41212 17382
rect 41236 17380 41292 17382
rect 41316 17380 41372 17382
rect 40958 16532 40960 16552
rect 40960 16532 41012 16552
rect 41012 16532 41014 16552
rect 40958 16496 41014 16532
rect 41076 16346 41132 16348
rect 41156 16346 41212 16348
rect 41236 16346 41292 16348
rect 41316 16346 41372 16348
rect 41076 16294 41122 16346
rect 41122 16294 41132 16346
rect 41156 16294 41186 16346
rect 41186 16294 41198 16346
rect 41198 16294 41212 16346
rect 41236 16294 41250 16346
rect 41250 16294 41262 16346
rect 41262 16294 41292 16346
rect 41316 16294 41326 16346
rect 41326 16294 41372 16346
rect 41076 16292 41132 16294
rect 41156 16292 41212 16294
rect 41236 16292 41292 16294
rect 41316 16292 41372 16294
rect 41076 15258 41132 15260
rect 41156 15258 41212 15260
rect 41236 15258 41292 15260
rect 41316 15258 41372 15260
rect 41076 15206 41122 15258
rect 41122 15206 41132 15258
rect 41156 15206 41186 15258
rect 41186 15206 41198 15258
rect 41198 15206 41212 15258
rect 41236 15206 41250 15258
rect 41250 15206 41262 15258
rect 41262 15206 41292 15258
rect 41316 15206 41326 15258
rect 41326 15206 41372 15258
rect 41076 15204 41132 15206
rect 41156 15204 41212 15206
rect 41236 15204 41292 15206
rect 41316 15204 41372 15206
rect 41076 14170 41132 14172
rect 41156 14170 41212 14172
rect 41236 14170 41292 14172
rect 41316 14170 41372 14172
rect 41076 14118 41122 14170
rect 41122 14118 41132 14170
rect 41156 14118 41186 14170
rect 41186 14118 41198 14170
rect 41198 14118 41212 14170
rect 41236 14118 41250 14170
rect 41250 14118 41262 14170
rect 41262 14118 41292 14170
rect 41316 14118 41326 14170
rect 41326 14118 41372 14170
rect 41076 14116 41132 14118
rect 41156 14116 41212 14118
rect 41236 14116 41292 14118
rect 41316 14116 41372 14118
rect 38576 9274 38632 9276
rect 38656 9274 38712 9276
rect 38736 9274 38792 9276
rect 38816 9274 38872 9276
rect 38576 9222 38622 9274
rect 38622 9222 38632 9274
rect 38656 9222 38686 9274
rect 38686 9222 38698 9274
rect 38698 9222 38712 9274
rect 38736 9222 38750 9274
rect 38750 9222 38762 9274
rect 38762 9222 38792 9274
rect 38816 9222 38826 9274
rect 38826 9222 38872 9274
rect 38576 9220 38632 9222
rect 38656 9220 38712 9222
rect 38736 9220 38792 9222
rect 38816 9220 38872 9222
rect 38750 8472 38806 8528
rect 38576 8186 38632 8188
rect 38656 8186 38712 8188
rect 38736 8186 38792 8188
rect 38816 8186 38872 8188
rect 38576 8134 38622 8186
rect 38622 8134 38632 8186
rect 38656 8134 38686 8186
rect 38686 8134 38698 8186
rect 38698 8134 38712 8186
rect 38736 8134 38750 8186
rect 38750 8134 38762 8186
rect 38762 8134 38792 8186
rect 38816 8134 38826 8186
rect 38826 8134 38872 8186
rect 38576 8132 38632 8134
rect 38656 8132 38712 8134
rect 38736 8132 38792 8134
rect 38816 8132 38872 8134
rect 40038 8508 40040 8528
rect 40040 8508 40092 8528
rect 40092 8508 40094 8528
rect 40038 8472 40094 8508
rect 41076 13082 41132 13084
rect 41156 13082 41212 13084
rect 41236 13082 41292 13084
rect 41316 13082 41372 13084
rect 41076 13030 41122 13082
rect 41122 13030 41132 13082
rect 41156 13030 41186 13082
rect 41186 13030 41198 13082
rect 41198 13030 41212 13082
rect 41236 13030 41250 13082
rect 41250 13030 41262 13082
rect 41262 13030 41292 13082
rect 41316 13030 41326 13082
rect 41326 13030 41372 13082
rect 41076 13028 41132 13030
rect 41156 13028 41212 13030
rect 41236 13028 41292 13030
rect 41316 13028 41372 13030
rect 41076 11994 41132 11996
rect 41156 11994 41212 11996
rect 41236 11994 41292 11996
rect 41316 11994 41372 11996
rect 41076 11942 41122 11994
rect 41122 11942 41132 11994
rect 41156 11942 41186 11994
rect 41186 11942 41198 11994
rect 41198 11942 41212 11994
rect 41236 11942 41250 11994
rect 41250 11942 41262 11994
rect 41262 11942 41292 11994
rect 41316 11942 41326 11994
rect 41326 11942 41372 11994
rect 41076 11940 41132 11942
rect 41156 11940 41212 11942
rect 41236 11940 41292 11942
rect 41316 11940 41372 11942
rect 41076 10906 41132 10908
rect 41156 10906 41212 10908
rect 41236 10906 41292 10908
rect 41316 10906 41372 10908
rect 41076 10854 41122 10906
rect 41122 10854 41132 10906
rect 41156 10854 41186 10906
rect 41186 10854 41198 10906
rect 41198 10854 41212 10906
rect 41236 10854 41250 10906
rect 41250 10854 41262 10906
rect 41262 10854 41292 10906
rect 41316 10854 41326 10906
rect 41326 10854 41372 10906
rect 41076 10852 41132 10854
rect 41156 10852 41212 10854
rect 41236 10852 41292 10854
rect 41316 10852 41372 10854
rect 41076 9818 41132 9820
rect 41156 9818 41212 9820
rect 41236 9818 41292 9820
rect 41316 9818 41372 9820
rect 41076 9766 41122 9818
rect 41122 9766 41132 9818
rect 41156 9766 41186 9818
rect 41186 9766 41198 9818
rect 41198 9766 41212 9818
rect 41236 9766 41250 9818
rect 41250 9766 41262 9818
rect 41262 9766 41292 9818
rect 41316 9766 41326 9818
rect 41326 9766 41372 9818
rect 41076 9764 41132 9766
rect 41156 9764 41212 9766
rect 41236 9764 41292 9766
rect 41316 9764 41372 9766
rect 36726 6740 36728 6760
rect 36728 6740 36780 6760
rect 36780 6740 36782 6760
rect 36726 6704 36782 6740
rect 36076 6554 36132 6556
rect 36156 6554 36212 6556
rect 36236 6554 36292 6556
rect 36316 6554 36372 6556
rect 36076 6502 36122 6554
rect 36122 6502 36132 6554
rect 36156 6502 36186 6554
rect 36186 6502 36198 6554
rect 36198 6502 36212 6554
rect 36236 6502 36250 6554
rect 36250 6502 36262 6554
rect 36262 6502 36292 6554
rect 36316 6502 36326 6554
rect 36326 6502 36372 6554
rect 36076 6500 36132 6502
rect 36156 6500 36212 6502
rect 36236 6500 36292 6502
rect 36316 6500 36372 6502
rect 36076 5466 36132 5468
rect 36156 5466 36212 5468
rect 36236 5466 36292 5468
rect 36316 5466 36372 5468
rect 36076 5414 36122 5466
rect 36122 5414 36132 5466
rect 36156 5414 36186 5466
rect 36186 5414 36198 5466
rect 36198 5414 36212 5466
rect 36236 5414 36250 5466
rect 36250 5414 36262 5466
rect 36262 5414 36292 5466
rect 36316 5414 36326 5466
rect 36326 5414 36372 5466
rect 36076 5412 36132 5414
rect 36156 5412 36212 5414
rect 36236 5412 36292 5414
rect 36316 5412 36372 5414
rect 37002 6160 37058 6216
rect 38106 6840 38162 6896
rect 36076 4378 36132 4380
rect 36156 4378 36212 4380
rect 36236 4378 36292 4380
rect 36316 4378 36372 4380
rect 36076 4326 36122 4378
rect 36122 4326 36132 4378
rect 36156 4326 36186 4378
rect 36186 4326 36198 4378
rect 36198 4326 36212 4378
rect 36236 4326 36250 4378
rect 36250 4326 36262 4378
rect 36262 4326 36292 4378
rect 36316 4326 36326 4378
rect 36326 4326 36372 4378
rect 36076 4324 36132 4326
rect 36156 4324 36212 4326
rect 36236 4324 36292 4326
rect 36316 4324 36372 4326
rect 36818 4004 36874 4040
rect 36818 3984 36820 4004
rect 36820 3984 36872 4004
rect 36872 3984 36874 4004
rect 36076 3290 36132 3292
rect 36156 3290 36212 3292
rect 36236 3290 36292 3292
rect 36316 3290 36372 3292
rect 36076 3238 36122 3290
rect 36122 3238 36132 3290
rect 36156 3238 36186 3290
rect 36186 3238 36198 3290
rect 36198 3238 36212 3290
rect 36236 3238 36250 3290
rect 36250 3238 36262 3290
rect 36262 3238 36292 3290
rect 36316 3238 36326 3290
rect 36326 3238 36372 3290
rect 36076 3236 36132 3238
rect 36156 3236 36212 3238
rect 36236 3236 36292 3238
rect 36316 3236 36372 3238
rect 35714 2624 35770 2680
rect 35898 2760 35954 2816
rect 36076 2202 36132 2204
rect 36156 2202 36212 2204
rect 36236 2202 36292 2204
rect 36316 2202 36372 2204
rect 36076 2150 36122 2202
rect 36122 2150 36132 2202
rect 36156 2150 36186 2202
rect 36186 2150 36198 2202
rect 36198 2150 36212 2202
rect 36236 2150 36250 2202
rect 36250 2150 36262 2202
rect 36262 2150 36292 2202
rect 36316 2150 36326 2202
rect 36326 2150 36372 2202
rect 36076 2148 36132 2150
rect 36156 2148 36212 2150
rect 36236 2148 36292 2150
rect 36316 2148 36372 2150
rect 36726 3032 36782 3088
rect 38106 6296 38162 6352
rect 38576 7098 38632 7100
rect 38656 7098 38712 7100
rect 38736 7098 38792 7100
rect 38816 7098 38872 7100
rect 38576 7046 38622 7098
rect 38622 7046 38632 7098
rect 38656 7046 38686 7098
rect 38686 7046 38698 7098
rect 38698 7046 38712 7098
rect 38736 7046 38750 7098
rect 38750 7046 38762 7098
rect 38762 7046 38792 7098
rect 38816 7046 38826 7098
rect 38826 7046 38872 7098
rect 38576 7044 38632 7046
rect 38656 7044 38712 7046
rect 38736 7044 38792 7046
rect 38816 7044 38872 7046
rect 38576 6010 38632 6012
rect 38656 6010 38712 6012
rect 38736 6010 38792 6012
rect 38816 6010 38872 6012
rect 38576 5958 38622 6010
rect 38622 5958 38632 6010
rect 38656 5958 38686 6010
rect 38686 5958 38698 6010
rect 38698 5958 38712 6010
rect 38736 5958 38750 6010
rect 38750 5958 38762 6010
rect 38762 5958 38792 6010
rect 38816 5958 38826 6010
rect 38826 5958 38872 6010
rect 38576 5956 38632 5958
rect 38656 5956 38712 5958
rect 38736 5956 38792 5958
rect 38816 5956 38872 5958
rect 38382 4820 38438 4856
rect 38382 4800 38384 4820
rect 38384 4800 38436 4820
rect 38436 4800 38438 4820
rect 37738 4548 37794 4584
rect 37738 4528 37740 4548
rect 37740 4528 37792 4548
rect 37792 4528 37794 4548
rect 36082 1400 36138 1456
rect 36174 1300 36176 1320
rect 36176 1300 36228 1320
rect 36228 1300 36230 1320
rect 36174 1264 36230 1300
rect 35898 1128 35954 1184
rect 36076 1114 36132 1116
rect 36156 1114 36212 1116
rect 36236 1114 36292 1116
rect 36316 1114 36372 1116
rect 36076 1062 36122 1114
rect 36122 1062 36132 1114
rect 36156 1062 36186 1114
rect 36186 1062 36198 1114
rect 36198 1062 36212 1114
rect 36236 1062 36250 1114
rect 36250 1062 36262 1114
rect 36262 1062 36292 1114
rect 36316 1062 36326 1114
rect 36326 1062 36372 1114
rect 36076 1060 36132 1062
rect 36156 1060 36212 1062
rect 36236 1060 36292 1062
rect 36316 1060 36372 1062
rect 37922 3576 37978 3632
rect 38014 3168 38070 3224
rect 37646 2896 37702 2952
rect 38290 2624 38346 2680
rect 43576 22330 43632 22332
rect 43656 22330 43712 22332
rect 43736 22330 43792 22332
rect 43816 22330 43872 22332
rect 43576 22278 43622 22330
rect 43622 22278 43632 22330
rect 43656 22278 43686 22330
rect 43686 22278 43698 22330
rect 43698 22278 43712 22330
rect 43736 22278 43750 22330
rect 43750 22278 43762 22330
rect 43762 22278 43792 22330
rect 43816 22278 43826 22330
rect 43826 22278 43872 22330
rect 43576 22276 43632 22278
rect 43656 22276 43712 22278
rect 43736 22276 43792 22278
rect 43816 22276 43872 22278
rect 43576 21242 43632 21244
rect 43656 21242 43712 21244
rect 43736 21242 43792 21244
rect 43816 21242 43872 21244
rect 43576 21190 43622 21242
rect 43622 21190 43632 21242
rect 43656 21190 43686 21242
rect 43686 21190 43698 21242
rect 43698 21190 43712 21242
rect 43736 21190 43750 21242
rect 43750 21190 43762 21242
rect 43762 21190 43792 21242
rect 43816 21190 43826 21242
rect 43826 21190 43872 21242
rect 43576 21188 43632 21190
rect 43656 21188 43712 21190
rect 43736 21188 43792 21190
rect 43816 21188 43872 21190
rect 43810 20324 43866 20360
rect 43810 20304 43812 20324
rect 43812 20304 43864 20324
rect 43864 20304 43866 20324
rect 43576 20154 43632 20156
rect 43656 20154 43712 20156
rect 43736 20154 43792 20156
rect 43816 20154 43872 20156
rect 43576 20102 43622 20154
rect 43622 20102 43632 20154
rect 43656 20102 43686 20154
rect 43686 20102 43698 20154
rect 43698 20102 43712 20154
rect 43736 20102 43750 20154
rect 43750 20102 43762 20154
rect 43762 20102 43792 20154
rect 43816 20102 43826 20154
rect 43826 20102 43872 20154
rect 43576 20100 43632 20102
rect 43656 20100 43712 20102
rect 43736 20100 43792 20102
rect 43816 20100 43872 20102
rect 43576 19066 43632 19068
rect 43656 19066 43712 19068
rect 43736 19066 43792 19068
rect 43816 19066 43872 19068
rect 43576 19014 43622 19066
rect 43622 19014 43632 19066
rect 43656 19014 43686 19066
rect 43686 19014 43698 19066
rect 43698 19014 43712 19066
rect 43736 19014 43750 19066
rect 43750 19014 43762 19066
rect 43762 19014 43792 19066
rect 43816 19014 43826 19066
rect 43826 19014 43872 19066
rect 43576 19012 43632 19014
rect 43656 19012 43712 19014
rect 43736 19012 43792 19014
rect 43816 19012 43872 19014
rect 43576 17978 43632 17980
rect 43656 17978 43712 17980
rect 43736 17978 43792 17980
rect 43816 17978 43872 17980
rect 43576 17926 43622 17978
rect 43622 17926 43632 17978
rect 43656 17926 43686 17978
rect 43686 17926 43698 17978
rect 43698 17926 43712 17978
rect 43736 17926 43750 17978
rect 43750 17926 43762 17978
rect 43762 17926 43792 17978
rect 43816 17926 43826 17978
rect 43826 17926 43872 17978
rect 43576 17924 43632 17926
rect 43656 17924 43712 17926
rect 43736 17924 43792 17926
rect 43816 17924 43872 17926
rect 43576 16890 43632 16892
rect 43656 16890 43712 16892
rect 43736 16890 43792 16892
rect 43816 16890 43872 16892
rect 43576 16838 43622 16890
rect 43622 16838 43632 16890
rect 43656 16838 43686 16890
rect 43686 16838 43698 16890
rect 43698 16838 43712 16890
rect 43736 16838 43750 16890
rect 43750 16838 43762 16890
rect 43762 16838 43792 16890
rect 43816 16838 43826 16890
rect 43826 16838 43872 16890
rect 43576 16836 43632 16838
rect 43656 16836 43712 16838
rect 43736 16836 43792 16838
rect 43816 16836 43872 16838
rect 43576 15802 43632 15804
rect 43656 15802 43712 15804
rect 43736 15802 43792 15804
rect 43816 15802 43872 15804
rect 43576 15750 43622 15802
rect 43622 15750 43632 15802
rect 43656 15750 43686 15802
rect 43686 15750 43698 15802
rect 43698 15750 43712 15802
rect 43736 15750 43750 15802
rect 43750 15750 43762 15802
rect 43762 15750 43792 15802
rect 43816 15750 43826 15802
rect 43826 15750 43872 15802
rect 43576 15748 43632 15750
rect 43656 15748 43712 15750
rect 43736 15748 43792 15750
rect 43816 15748 43872 15750
rect 43576 14714 43632 14716
rect 43656 14714 43712 14716
rect 43736 14714 43792 14716
rect 43816 14714 43872 14716
rect 43576 14662 43622 14714
rect 43622 14662 43632 14714
rect 43656 14662 43686 14714
rect 43686 14662 43698 14714
rect 43698 14662 43712 14714
rect 43736 14662 43750 14714
rect 43750 14662 43762 14714
rect 43762 14662 43792 14714
rect 43816 14662 43826 14714
rect 43826 14662 43872 14714
rect 43576 14660 43632 14662
rect 43656 14660 43712 14662
rect 43736 14660 43792 14662
rect 43816 14660 43872 14662
rect 42522 9560 42578 9616
rect 41970 9016 42026 9072
rect 45190 20712 45246 20768
rect 43576 13626 43632 13628
rect 43656 13626 43712 13628
rect 43736 13626 43792 13628
rect 43816 13626 43872 13628
rect 43576 13574 43622 13626
rect 43622 13574 43632 13626
rect 43656 13574 43686 13626
rect 43686 13574 43698 13626
rect 43698 13574 43712 13626
rect 43736 13574 43750 13626
rect 43750 13574 43762 13626
rect 43762 13574 43792 13626
rect 43816 13574 43826 13626
rect 43826 13574 43872 13626
rect 43576 13572 43632 13574
rect 43656 13572 43712 13574
rect 43736 13572 43792 13574
rect 43816 13572 43872 13574
rect 43576 12538 43632 12540
rect 43656 12538 43712 12540
rect 43736 12538 43792 12540
rect 43816 12538 43872 12540
rect 43576 12486 43622 12538
rect 43622 12486 43632 12538
rect 43656 12486 43686 12538
rect 43686 12486 43698 12538
rect 43698 12486 43712 12538
rect 43736 12486 43750 12538
rect 43750 12486 43762 12538
rect 43762 12486 43792 12538
rect 43816 12486 43826 12538
rect 43826 12486 43872 12538
rect 43576 12484 43632 12486
rect 43656 12484 43712 12486
rect 43736 12484 43792 12486
rect 43816 12484 43872 12486
rect 43576 11450 43632 11452
rect 43656 11450 43712 11452
rect 43736 11450 43792 11452
rect 43816 11450 43872 11452
rect 43576 11398 43622 11450
rect 43622 11398 43632 11450
rect 43656 11398 43686 11450
rect 43686 11398 43698 11450
rect 43698 11398 43712 11450
rect 43736 11398 43750 11450
rect 43750 11398 43762 11450
rect 43762 11398 43792 11450
rect 43816 11398 43826 11450
rect 43826 11398 43872 11450
rect 43576 11396 43632 11398
rect 43656 11396 43712 11398
rect 43736 11396 43792 11398
rect 43816 11396 43872 11398
rect 43576 10362 43632 10364
rect 43656 10362 43712 10364
rect 43736 10362 43792 10364
rect 43816 10362 43872 10364
rect 43576 10310 43622 10362
rect 43622 10310 43632 10362
rect 43656 10310 43686 10362
rect 43686 10310 43698 10362
rect 43698 10310 43712 10362
rect 43736 10310 43750 10362
rect 43750 10310 43762 10362
rect 43762 10310 43792 10362
rect 43816 10310 43826 10362
rect 43826 10310 43872 10362
rect 43576 10308 43632 10310
rect 43656 10308 43712 10310
rect 43736 10308 43792 10310
rect 43816 10308 43872 10310
rect 45190 14728 45246 14784
rect 44822 11192 44878 11248
rect 41076 8730 41132 8732
rect 41156 8730 41212 8732
rect 41236 8730 41292 8732
rect 41316 8730 41372 8732
rect 41076 8678 41122 8730
rect 41122 8678 41132 8730
rect 41156 8678 41186 8730
rect 41186 8678 41198 8730
rect 41198 8678 41212 8730
rect 41236 8678 41250 8730
rect 41250 8678 41262 8730
rect 41262 8678 41292 8730
rect 41316 8678 41326 8730
rect 41326 8678 41372 8730
rect 41076 8676 41132 8678
rect 41156 8676 41212 8678
rect 41236 8676 41292 8678
rect 41316 8676 41372 8678
rect 40866 7928 40922 7984
rect 41076 7642 41132 7644
rect 41156 7642 41212 7644
rect 41236 7642 41292 7644
rect 41316 7642 41372 7644
rect 41076 7590 41122 7642
rect 41122 7590 41132 7642
rect 41156 7590 41186 7642
rect 41186 7590 41198 7642
rect 41198 7590 41212 7642
rect 41236 7590 41250 7642
rect 41250 7590 41262 7642
rect 41262 7590 41292 7642
rect 41316 7590 41326 7642
rect 41326 7590 41372 7642
rect 41076 7588 41132 7590
rect 41156 7588 41212 7590
rect 41236 7588 41292 7590
rect 41316 7588 41372 7590
rect 38576 4922 38632 4924
rect 38656 4922 38712 4924
rect 38736 4922 38792 4924
rect 38816 4922 38872 4924
rect 38576 4870 38622 4922
rect 38622 4870 38632 4922
rect 38656 4870 38686 4922
rect 38686 4870 38698 4922
rect 38698 4870 38712 4922
rect 38736 4870 38750 4922
rect 38750 4870 38762 4922
rect 38762 4870 38792 4922
rect 38816 4870 38826 4922
rect 38826 4870 38872 4922
rect 38576 4868 38632 4870
rect 38656 4868 38712 4870
rect 38736 4868 38792 4870
rect 38816 4868 38872 4870
rect 38576 3834 38632 3836
rect 38656 3834 38712 3836
rect 38736 3834 38792 3836
rect 38816 3834 38872 3836
rect 38576 3782 38622 3834
rect 38622 3782 38632 3834
rect 38656 3782 38686 3834
rect 38686 3782 38698 3834
rect 38698 3782 38712 3834
rect 38736 3782 38750 3834
rect 38750 3782 38762 3834
rect 38762 3782 38792 3834
rect 38816 3782 38826 3834
rect 38826 3782 38872 3834
rect 38576 3780 38632 3782
rect 38656 3780 38712 3782
rect 38736 3780 38792 3782
rect 38816 3780 38872 3782
rect 40774 6180 40830 6216
rect 40774 6160 40776 6180
rect 40776 6160 40828 6180
rect 40828 6160 40830 6180
rect 41076 6554 41132 6556
rect 41156 6554 41212 6556
rect 41236 6554 41292 6556
rect 41316 6554 41372 6556
rect 41076 6502 41122 6554
rect 41122 6502 41132 6554
rect 41156 6502 41186 6554
rect 41186 6502 41198 6554
rect 41198 6502 41212 6554
rect 41236 6502 41250 6554
rect 41250 6502 41262 6554
rect 41262 6502 41292 6554
rect 41316 6502 41326 6554
rect 41326 6502 41372 6554
rect 41076 6500 41132 6502
rect 41156 6500 41212 6502
rect 41236 6500 41292 6502
rect 41316 6500 41372 6502
rect 44730 9560 44786 9616
rect 43576 9274 43632 9276
rect 43656 9274 43712 9276
rect 43736 9274 43792 9276
rect 43816 9274 43872 9276
rect 43576 9222 43622 9274
rect 43622 9222 43632 9274
rect 43656 9222 43686 9274
rect 43686 9222 43698 9274
rect 43698 9222 43712 9274
rect 43736 9222 43750 9274
rect 43750 9222 43762 9274
rect 43762 9222 43792 9274
rect 43816 9222 43826 9274
rect 43826 9222 43872 9274
rect 43576 9220 43632 9222
rect 43656 9220 43712 9222
rect 43736 9220 43792 9222
rect 43816 9220 43872 9222
rect 44638 8744 44694 8800
rect 42890 7792 42946 7848
rect 42706 6840 42762 6896
rect 43576 8186 43632 8188
rect 43656 8186 43712 8188
rect 43736 8186 43792 8188
rect 43816 8186 43872 8188
rect 43576 8134 43622 8186
rect 43622 8134 43632 8186
rect 43656 8134 43686 8186
rect 43686 8134 43698 8186
rect 43698 8134 43712 8186
rect 43736 8134 43750 8186
rect 43750 8134 43762 8186
rect 43762 8134 43792 8186
rect 43816 8134 43826 8186
rect 43826 8134 43872 8186
rect 43576 8132 43632 8134
rect 43656 8132 43712 8134
rect 43736 8132 43792 8134
rect 43816 8132 43872 8134
rect 38576 2746 38632 2748
rect 38656 2746 38712 2748
rect 38736 2746 38792 2748
rect 38816 2746 38872 2748
rect 38576 2694 38622 2746
rect 38622 2694 38632 2746
rect 38656 2694 38686 2746
rect 38686 2694 38698 2746
rect 38698 2694 38712 2746
rect 38736 2694 38750 2746
rect 38750 2694 38762 2746
rect 38762 2694 38792 2746
rect 38816 2694 38826 2746
rect 38826 2694 38872 2746
rect 38576 2692 38632 2694
rect 38656 2692 38712 2694
rect 38736 2692 38792 2694
rect 38816 2692 38872 2694
rect 38576 1658 38632 1660
rect 38656 1658 38712 1660
rect 38736 1658 38792 1660
rect 38816 1658 38872 1660
rect 38576 1606 38622 1658
rect 38622 1606 38632 1658
rect 38656 1606 38686 1658
rect 38686 1606 38698 1658
rect 38698 1606 38712 1658
rect 38736 1606 38750 1658
rect 38750 1606 38762 1658
rect 38762 1606 38792 1658
rect 38816 1606 38826 1658
rect 38826 1606 38872 1658
rect 38576 1604 38632 1606
rect 38656 1604 38712 1606
rect 38736 1604 38792 1606
rect 38816 1604 38872 1606
rect 41076 5466 41132 5468
rect 41156 5466 41212 5468
rect 41236 5466 41292 5468
rect 41316 5466 41372 5468
rect 41076 5414 41122 5466
rect 41122 5414 41132 5466
rect 41156 5414 41186 5466
rect 41186 5414 41198 5466
rect 41198 5414 41212 5466
rect 41236 5414 41250 5466
rect 41250 5414 41262 5466
rect 41262 5414 41292 5466
rect 41316 5414 41326 5466
rect 41326 5414 41372 5466
rect 41076 5412 41132 5414
rect 41156 5412 41212 5414
rect 41236 5412 41292 5414
rect 41316 5412 41372 5414
rect 41076 4378 41132 4380
rect 41156 4378 41212 4380
rect 41236 4378 41292 4380
rect 41316 4378 41372 4380
rect 41076 4326 41122 4378
rect 41122 4326 41132 4378
rect 41156 4326 41186 4378
rect 41186 4326 41198 4378
rect 41198 4326 41212 4378
rect 41236 4326 41250 4378
rect 41250 4326 41262 4378
rect 41262 4326 41292 4378
rect 41316 4326 41326 4378
rect 41326 4326 41372 4378
rect 41076 4324 41132 4326
rect 41156 4324 41212 4326
rect 41236 4324 41292 4326
rect 41316 4324 41372 4326
rect 40682 3032 40738 3088
rect 41970 4664 42026 4720
rect 41510 4120 41566 4176
rect 41076 3290 41132 3292
rect 41156 3290 41212 3292
rect 41236 3290 41292 3292
rect 41316 3290 41372 3292
rect 41076 3238 41122 3290
rect 41122 3238 41132 3290
rect 41156 3238 41186 3290
rect 41186 3238 41198 3290
rect 41198 3238 41212 3290
rect 41236 3238 41250 3290
rect 41250 3238 41262 3290
rect 41262 3238 41292 3290
rect 41316 3238 41326 3290
rect 41326 3238 41372 3290
rect 41076 3236 41132 3238
rect 41156 3236 41212 3238
rect 41236 3236 41292 3238
rect 41316 3236 41372 3238
rect 40866 2352 40922 2408
rect 41076 2202 41132 2204
rect 41156 2202 41212 2204
rect 41236 2202 41292 2204
rect 41316 2202 41372 2204
rect 41076 2150 41122 2202
rect 41122 2150 41132 2202
rect 41156 2150 41186 2202
rect 41186 2150 41198 2202
rect 41198 2150 41212 2202
rect 41236 2150 41250 2202
rect 41250 2150 41262 2202
rect 41262 2150 41292 2202
rect 41316 2150 41326 2202
rect 41326 2150 41372 2202
rect 41076 2148 41132 2150
rect 41156 2148 41212 2150
rect 41236 2148 41292 2150
rect 41316 2148 41372 2150
rect 40498 1264 40554 1320
rect 41510 2488 41566 2544
rect 41076 1114 41132 1116
rect 41156 1114 41212 1116
rect 41236 1114 41292 1116
rect 41316 1114 41372 1116
rect 41076 1062 41122 1114
rect 41122 1062 41132 1114
rect 41156 1062 41186 1114
rect 41186 1062 41198 1114
rect 41198 1062 41212 1114
rect 41236 1062 41250 1114
rect 41250 1062 41262 1114
rect 41262 1062 41292 1114
rect 41316 1062 41326 1114
rect 41326 1062 41372 1114
rect 41076 1060 41132 1062
rect 41156 1060 41212 1062
rect 41236 1060 41292 1062
rect 41316 1060 41372 1062
rect 44178 7420 44180 7440
rect 44180 7420 44232 7440
rect 44232 7420 44234 7440
rect 44178 7384 44234 7420
rect 43576 7098 43632 7100
rect 43656 7098 43712 7100
rect 43736 7098 43792 7100
rect 43816 7098 43872 7100
rect 43576 7046 43622 7098
rect 43622 7046 43632 7098
rect 43656 7046 43686 7098
rect 43686 7046 43698 7098
rect 43698 7046 43712 7098
rect 43736 7046 43750 7098
rect 43750 7046 43762 7098
rect 43762 7046 43792 7098
rect 43816 7046 43826 7098
rect 43826 7046 43872 7098
rect 43576 7044 43632 7046
rect 43656 7044 43712 7046
rect 43736 7044 43792 7046
rect 43816 7044 43872 7046
rect 43576 6010 43632 6012
rect 43656 6010 43712 6012
rect 43736 6010 43792 6012
rect 43816 6010 43872 6012
rect 43576 5958 43622 6010
rect 43622 5958 43632 6010
rect 43656 5958 43686 6010
rect 43686 5958 43698 6010
rect 43698 5958 43712 6010
rect 43736 5958 43750 6010
rect 43750 5958 43762 6010
rect 43762 5958 43792 6010
rect 43816 5958 43826 6010
rect 43826 5958 43872 6010
rect 43576 5956 43632 5958
rect 43656 5956 43712 5958
rect 43736 5956 43792 5958
rect 43816 5956 43872 5958
rect 43576 4922 43632 4924
rect 43656 4922 43712 4924
rect 43736 4922 43792 4924
rect 43816 4922 43872 4924
rect 43576 4870 43622 4922
rect 43622 4870 43632 4922
rect 43656 4870 43686 4922
rect 43686 4870 43698 4922
rect 43698 4870 43712 4922
rect 43736 4870 43750 4922
rect 43750 4870 43762 4922
rect 43762 4870 43792 4922
rect 43816 4870 43826 4922
rect 43826 4870 43872 4922
rect 43576 4868 43632 4870
rect 43656 4868 43712 4870
rect 43736 4868 43792 4870
rect 43816 4868 43872 4870
rect 43576 3834 43632 3836
rect 43656 3834 43712 3836
rect 43736 3834 43792 3836
rect 43816 3834 43872 3836
rect 43576 3782 43622 3834
rect 43622 3782 43632 3834
rect 43656 3782 43686 3834
rect 43686 3782 43698 3834
rect 43698 3782 43712 3834
rect 43736 3782 43750 3834
rect 43750 3782 43762 3834
rect 43762 3782 43792 3834
rect 43816 3782 43826 3834
rect 43826 3782 43872 3834
rect 43576 3780 43632 3782
rect 43656 3780 43712 3782
rect 43736 3780 43792 3782
rect 43816 3780 43872 3782
rect 43576 2746 43632 2748
rect 43656 2746 43712 2748
rect 43736 2746 43792 2748
rect 43816 2746 43872 2748
rect 43576 2694 43622 2746
rect 43622 2694 43632 2746
rect 43656 2694 43686 2746
rect 43686 2694 43698 2746
rect 43698 2694 43712 2746
rect 43736 2694 43750 2746
rect 43750 2694 43762 2746
rect 43762 2694 43792 2746
rect 43816 2694 43826 2746
rect 43826 2694 43872 2746
rect 43576 2692 43632 2694
rect 43656 2692 43712 2694
rect 43736 2692 43792 2694
rect 43816 2692 43872 2694
rect 43576 1658 43632 1660
rect 43656 1658 43712 1660
rect 43736 1658 43792 1660
rect 43816 1658 43872 1660
rect 43576 1606 43622 1658
rect 43622 1606 43632 1658
rect 43656 1606 43686 1658
rect 43686 1606 43698 1658
rect 43698 1606 43712 1658
rect 43736 1606 43750 1658
rect 43750 1606 43762 1658
rect 43762 1606 43792 1658
rect 43816 1606 43826 1658
rect 43826 1606 43872 1658
rect 43576 1604 43632 1606
rect 43656 1604 43712 1606
rect 43736 1604 43792 1606
rect 43816 1604 43872 1606
rect 44638 2760 44694 2816
<< metal3 >>
rect 6066 22880 6382 22881
rect 6066 22816 6072 22880
rect 6136 22816 6152 22880
rect 6216 22816 6232 22880
rect 6296 22816 6312 22880
rect 6376 22816 6382 22880
rect 6066 22815 6382 22816
rect 11066 22880 11382 22881
rect 11066 22816 11072 22880
rect 11136 22816 11152 22880
rect 11216 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11382 22880
rect 11066 22815 11382 22816
rect 16066 22880 16382 22881
rect 16066 22816 16072 22880
rect 16136 22816 16152 22880
rect 16216 22816 16232 22880
rect 16296 22816 16312 22880
rect 16376 22816 16382 22880
rect 16066 22815 16382 22816
rect 21066 22880 21382 22881
rect 21066 22816 21072 22880
rect 21136 22816 21152 22880
rect 21216 22816 21232 22880
rect 21296 22816 21312 22880
rect 21376 22816 21382 22880
rect 21066 22815 21382 22816
rect 26066 22880 26382 22881
rect 26066 22816 26072 22880
rect 26136 22816 26152 22880
rect 26216 22816 26232 22880
rect 26296 22816 26312 22880
rect 26376 22816 26382 22880
rect 26066 22815 26382 22816
rect 31066 22880 31382 22881
rect 31066 22816 31072 22880
rect 31136 22816 31152 22880
rect 31216 22816 31232 22880
rect 31296 22816 31312 22880
rect 31376 22816 31382 22880
rect 31066 22815 31382 22816
rect 36066 22880 36382 22881
rect 36066 22816 36072 22880
rect 36136 22816 36152 22880
rect 36216 22816 36232 22880
rect 36296 22816 36312 22880
rect 36376 22816 36382 22880
rect 36066 22815 36382 22816
rect 41066 22880 41382 22881
rect 41066 22816 41072 22880
rect 41136 22816 41152 22880
rect 41216 22816 41232 22880
rect 41296 22816 41312 22880
rect 41376 22816 41382 22880
rect 41066 22815 41382 22816
rect 12801 22538 12867 22541
rect 17125 22538 17191 22541
rect 12801 22536 17191 22538
rect 12801 22480 12806 22536
rect 12862 22480 17130 22536
rect 17186 22480 17191 22536
rect 12801 22478 17191 22480
rect 12801 22475 12867 22478
rect 17125 22475 17191 22478
rect 17953 22538 18019 22541
rect 19190 22538 19196 22540
rect 17953 22536 19196 22538
rect 17953 22480 17958 22536
rect 18014 22480 19196 22536
rect 17953 22478 19196 22480
rect 17953 22475 18019 22478
rect 19190 22476 19196 22478
rect 19260 22538 19266 22540
rect 19260 22478 22110 22538
rect 19260 22476 19266 22478
rect 3566 22336 3882 22337
rect 3566 22272 3572 22336
rect 3636 22272 3652 22336
rect 3716 22272 3732 22336
rect 3796 22272 3812 22336
rect 3876 22272 3882 22336
rect 3566 22271 3882 22272
rect 8566 22336 8882 22337
rect 8566 22272 8572 22336
rect 8636 22272 8652 22336
rect 8716 22272 8732 22336
rect 8796 22272 8812 22336
rect 8876 22272 8882 22336
rect 8566 22271 8882 22272
rect 13566 22336 13882 22337
rect 13566 22272 13572 22336
rect 13636 22272 13652 22336
rect 13716 22272 13732 22336
rect 13796 22272 13812 22336
rect 13876 22272 13882 22336
rect 13566 22271 13882 22272
rect 18566 22336 18882 22337
rect 18566 22272 18572 22336
rect 18636 22272 18652 22336
rect 18716 22272 18732 22336
rect 18796 22272 18812 22336
rect 18876 22272 18882 22336
rect 18566 22271 18882 22272
rect 22050 22266 22110 22478
rect 23566 22336 23882 22337
rect 23566 22272 23572 22336
rect 23636 22272 23652 22336
rect 23716 22272 23732 22336
rect 23796 22272 23812 22336
rect 23876 22272 23882 22336
rect 23566 22271 23882 22272
rect 28566 22336 28882 22337
rect 28566 22272 28572 22336
rect 28636 22272 28652 22336
rect 28716 22272 28732 22336
rect 28796 22272 28812 22336
rect 28876 22272 28882 22336
rect 28566 22271 28882 22272
rect 33566 22336 33882 22337
rect 33566 22272 33572 22336
rect 33636 22272 33652 22336
rect 33716 22272 33732 22336
rect 33796 22272 33812 22336
rect 33876 22272 33882 22336
rect 33566 22271 33882 22272
rect 38566 22336 38882 22337
rect 38566 22272 38572 22336
rect 38636 22272 38652 22336
rect 38716 22272 38732 22336
rect 38796 22272 38812 22336
rect 38876 22272 38882 22336
rect 38566 22271 38882 22272
rect 43566 22336 43882 22337
rect 43566 22272 43572 22336
rect 43636 22272 43652 22336
rect 43716 22272 43732 22336
rect 43796 22272 43812 22336
rect 43876 22272 43882 22336
rect 43566 22271 43882 22272
rect 22050 22206 23490 22266
rect 5073 22130 5139 22133
rect 23430 22130 23490 22206
rect 25454 22206 26250 22266
rect 25454 22130 25514 22206
rect 5073 22128 22202 22130
rect 5073 22072 5078 22128
rect 5134 22072 22202 22128
rect 5073 22070 22202 22072
rect 23430 22070 25514 22130
rect 25589 22130 25655 22133
rect 25814 22130 25820 22132
rect 25589 22128 25820 22130
rect 25589 22072 25594 22128
rect 25650 22072 25820 22128
rect 25589 22070 25820 22072
rect 5073 22067 5139 22070
rect 4429 21994 4495 21997
rect 5349 21994 5415 21997
rect 18321 21994 18387 21997
rect 19793 21994 19859 21997
rect 4429 21992 17234 21994
rect 4429 21936 4434 21992
rect 4490 21936 5354 21992
rect 5410 21936 17234 21992
rect 4429 21934 17234 21936
rect 4429 21931 4495 21934
rect 5349 21931 5415 21934
rect 17174 21858 17234 21934
rect 18321 21992 19859 21994
rect 18321 21936 18326 21992
rect 18382 21936 19798 21992
rect 19854 21936 19859 21992
rect 18321 21934 19859 21936
rect 22142 21994 22202 22070
rect 25589 22067 25655 22070
rect 25814 22068 25820 22070
rect 25884 22068 25890 22132
rect 26190 21994 26250 22206
rect 28206 22068 28212 22132
rect 28276 22130 28282 22132
rect 32397 22130 32463 22133
rect 28276 22128 32463 22130
rect 28276 22072 32402 22128
rect 32458 22072 32463 22128
rect 28276 22070 32463 22072
rect 28276 22068 28282 22070
rect 32397 22067 32463 22070
rect 32949 22130 33015 22133
rect 35433 22130 35499 22133
rect 32949 22128 35499 22130
rect 32949 22072 32954 22128
rect 33010 22072 35438 22128
rect 35494 22072 35499 22128
rect 32949 22070 35499 22072
rect 32949 22067 33015 22070
rect 35433 22067 35499 22070
rect 27613 21994 27679 21997
rect 22142 21934 22386 21994
rect 26190 21992 27679 21994
rect 26190 21936 27618 21992
rect 27674 21936 27679 21992
rect 26190 21934 27679 21936
rect 18321 21931 18387 21934
rect 19793 21931 19859 21934
rect 20253 21858 20319 21861
rect 17174 21856 20319 21858
rect 17174 21800 20258 21856
rect 20314 21800 20319 21856
rect 17174 21798 20319 21800
rect 20253 21795 20319 21798
rect 6066 21792 6382 21793
rect 6066 21728 6072 21792
rect 6136 21728 6152 21792
rect 6216 21728 6232 21792
rect 6296 21728 6312 21792
rect 6376 21728 6382 21792
rect 6066 21727 6382 21728
rect 11066 21792 11382 21793
rect 11066 21728 11072 21792
rect 11136 21728 11152 21792
rect 11216 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11382 21792
rect 11066 21727 11382 21728
rect 16066 21792 16382 21793
rect 16066 21728 16072 21792
rect 16136 21728 16152 21792
rect 16216 21728 16232 21792
rect 16296 21728 16312 21792
rect 16376 21728 16382 21792
rect 16066 21727 16382 21728
rect 21066 21792 21382 21793
rect 21066 21728 21072 21792
rect 21136 21728 21152 21792
rect 21216 21728 21232 21792
rect 21296 21728 21312 21792
rect 21376 21728 21382 21792
rect 21066 21727 21382 21728
rect 19517 21722 19583 21725
rect 19926 21722 19932 21724
rect 19517 21720 19932 21722
rect 19517 21664 19522 21720
rect 19578 21664 19932 21720
rect 19517 21662 19932 21664
rect 19517 21659 19583 21662
rect 19926 21660 19932 21662
rect 19996 21660 20002 21724
rect 22326 21722 22386 21934
rect 27613 21931 27679 21934
rect 28349 21994 28415 21997
rect 33409 21994 33475 21997
rect 28349 21992 33475 21994
rect 28349 21936 28354 21992
rect 28410 21936 33414 21992
rect 33470 21936 33475 21992
rect 28349 21934 33475 21936
rect 28349 21931 28415 21934
rect 33409 21931 33475 21934
rect 26066 21792 26382 21793
rect 26066 21728 26072 21792
rect 26136 21728 26152 21792
rect 26216 21728 26232 21792
rect 26296 21728 26312 21792
rect 26376 21728 26382 21792
rect 26066 21727 26382 21728
rect 31066 21792 31382 21793
rect 31066 21728 31072 21792
rect 31136 21728 31152 21792
rect 31216 21728 31232 21792
rect 31296 21728 31312 21792
rect 31376 21728 31382 21792
rect 31066 21727 31382 21728
rect 36066 21792 36382 21793
rect 36066 21728 36072 21792
rect 36136 21728 36152 21792
rect 36216 21728 36232 21792
rect 36296 21728 36312 21792
rect 36376 21728 36382 21792
rect 36066 21727 36382 21728
rect 41066 21792 41382 21793
rect 41066 21728 41072 21792
rect 41136 21728 41152 21792
rect 41216 21728 41232 21792
rect 41296 21728 41312 21792
rect 41376 21728 41382 21792
rect 41066 21727 41382 21728
rect 25681 21722 25747 21725
rect 22326 21720 25747 21722
rect 22326 21664 25686 21720
rect 25742 21664 25747 21720
rect 22326 21662 25747 21664
rect 25681 21659 25747 21662
rect 26734 21660 26740 21724
rect 26804 21722 26810 21724
rect 27705 21722 27771 21725
rect 26804 21720 27771 21722
rect 26804 21664 27710 21720
rect 27766 21664 27771 21720
rect 26804 21662 27771 21664
rect 26804 21660 26810 21662
rect 27705 21659 27771 21662
rect 6453 21586 6519 21589
rect 23289 21586 23355 21589
rect 6453 21584 23355 21586
rect 6453 21528 6458 21584
rect 6514 21528 23294 21584
rect 23350 21528 23355 21584
rect 6453 21526 23355 21528
rect 6453 21523 6519 21526
rect 23289 21523 23355 21526
rect 23657 21586 23723 21589
rect 30005 21586 30071 21589
rect 23657 21584 30071 21586
rect 23657 21528 23662 21584
rect 23718 21528 30010 21584
rect 30066 21528 30071 21584
rect 23657 21526 30071 21528
rect 23657 21523 23723 21526
rect 30005 21523 30071 21526
rect 30741 21586 30807 21589
rect 36629 21586 36695 21589
rect 30741 21584 36695 21586
rect 30741 21528 30746 21584
rect 30802 21528 36634 21584
rect 36690 21528 36695 21584
rect 30741 21526 36695 21528
rect 30741 21523 30807 21526
rect 36629 21523 36695 21526
rect 11697 21450 11763 21453
rect 17309 21450 17375 21453
rect 11697 21448 17375 21450
rect 11697 21392 11702 21448
rect 11758 21392 17314 21448
rect 17370 21392 17375 21448
rect 11697 21390 17375 21392
rect 11697 21387 11763 21390
rect 17309 21387 17375 21390
rect 18137 21450 18203 21453
rect 20253 21450 20319 21453
rect 23013 21450 23079 21453
rect 23381 21450 23447 21453
rect 26693 21450 26759 21453
rect 18137 21448 20178 21450
rect 18137 21392 18142 21448
rect 18198 21392 20178 21448
rect 18137 21390 20178 21392
rect 18137 21387 18203 21390
rect 14273 21314 14339 21317
rect 17493 21314 17559 21317
rect 14273 21312 17559 21314
rect 14273 21256 14278 21312
rect 14334 21256 17498 21312
rect 17554 21256 17559 21312
rect 14273 21254 17559 21256
rect 20118 21314 20178 21390
rect 20253 21448 23079 21450
rect 20253 21392 20258 21448
rect 20314 21392 23018 21448
rect 23074 21392 23079 21448
rect 20253 21390 23079 21392
rect 20253 21387 20319 21390
rect 23013 21387 23079 21390
rect 23246 21448 26759 21450
rect 23246 21392 23386 21448
rect 23442 21392 26698 21448
rect 26754 21392 26759 21448
rect 23246 21390 26759 21392
rect 23246 21314 23306 21390
rect 23381 21387 23447 21390
rect 26693 21387 26759 21390
rect 31109 21450 31175 21453
rect 37825 21450 37891 21453
rect 31109 21448 37891 21450
rect 31109 21392 31114 21448
rect 31170 21392 37830 21448
rect 37886 21392 37891 21448
rect 31109 21390 37891 21392
rect 31109 21387 31175 21390
rect 37825 21387 37891 21390
rect 20118 21254 23306 21314
rect 14273 21251 14339 21254
rect 17493 21251 17559 21254
rect 3566 21248 3882 21249
rect 3566 21184 3572 21248
rect 3636 21184 3652 21248
rect 3716 21184 3732 21248
rect 3796 21184 3812 21248
rect 3876 21184 3882 21248
rect 3566 21183 3882 21184
rect 8566 21248 8882 21249
rect 8566 21184 8572 21248
rect 8636 21184 8652 21248
rect 8716 21184 8732 21248
rect 8796 21184 8812 21248
rect 8876 21184 8882 21248
rect 8566 21183 8882 21184
rect 13566 21248 13882 21249
rect 13566 21184 13572 21248
rect 13636 21184 13652 21248
rect 13716 21184 13732 21248
rect 13796 21184 13812 21248
rect 13876 21184 13882 21248
rect 13566 21183 13882 21184
rect 18566 21248 18882 21249
rect 18566 21184 18572 21248
rect 18636 21184 18652 21248
rect 18716 21184 18732 21248
rect 18796 21184 18812 21248
rect 18876 21184 18882 21248
rect 18566 21183 18882 21184
rect 23566 21248 23882 21249
rect 23566 21184 23572 21248
rect 23636 21184 23652 21248
rect 23716 21184 23732 21248
rect 23796 21184 23812 21248
rect 23876 21184 23882 21248
rect 23566 21183 23882 21184
rect 28566 21248 28882 21249
rect 28566 21184 28572 21248
rect 28636 21184 28652 21248
rect 28716 21184 28732 21248
rect 28796 21184 28812 21248
rect 28876 21184 28882 21248
rect 28566 21183 28882 21184
rect 33566 21248 33882 21249
rect 33566 21184 33572 21248
rect 33636 21184 33652 21248
rect 33716 21184 33732 21248
rect 33796 21184 33812 21248
rect 33876 21184 33882 21248
rect 33566 21183 33882 21184
rect 38566 21248 38882 21249
rect 38566 21184 38572 21248
rect 38636 21184 38652 21248
rect 38716 21184 38732 21248
rect 38796 21184 38812 21248
rect 38876 21184 38882 21248
rect 38566 21183 38882 21184
rect 43566 21248 43882 21249
rect 43566 21184 43572 21248
rect 43636 21184 43652 21248
rect 43716 21184 43732 21248
rect 43796 21184 43812 21248
rect 43876 21184 43882 21248
rect 43566 21183 43882 21184
rect 13997 21178 14063 21181
rect 18229 21178 18295 21181
rect 13997 21176 18295 21178
rect 13997 21120 14002 21176
rect 14058 21120 18234 21176
rect 18290 21120 18295 21176
rect 13997 21118 18295 21120
rect 13997 21115 14063 21118
rect 18229 21115 18295 21118
rect 18965 21178 19031 21181
rect 21173 21178 21239 21181
rect 21633 21178 21699 21181
rect 18965 21176 21699 21178
rect 18965 21120 18970 21176
rect 19026 21120 21178 21176
rect 21234 21120 21638 21176
rect 21694 21120 21699 21176
rect 18965 21118 21699 21120
rect 18965 21115 19031 21118
rect 21173 21115 21239 21118
rect 21633 21115 21699 21118
rect 25681 21178 25747 21181
rect 27654 21178 27660 21180
rect 25681 21176 27660 21178
rect 25681 21120 25686 21176
rect 25742 21120 27660 21176
rect 25681 21118 27660 21120
rect 25681 21115 25747 21118
rect 27654 21116 27660 21118
rect 27724 21116 27730 21180
rect 30373 21178 30439 21181
rect 30373 21176 33426 21178
rect 30373 21120 30378 21176
rect 30434 21120 33426 21176
rect 30373 21118 33426 21120
rect 30373 21115 30439 21118
rect 12617 21042 12683 21045
rect 17861 21042 17927 21045
rect 12617 21040 17927 21042
rect 12617 20984 12622 21040
rect 12678 20984 17866 21040
rect 17922 20984 17927 21040
rect 12617 20982 17927 20984
rect 12617 20979 12683 20982
rect 17861 20979 17927 20982
rect 19057 21042 19123 21045
rect 19517 21042 19583 21045
rect 27153 21042 27219 21045
rect 32121 21042 32187 21045
rect 19057 21040 19583 21042
rect 19057 20984 19062 21040
rect 19118 20984 19522 21040
rect 19578 20984 19583 21040
rect 19057 20982 19583 20984
rect 19057 20979 19123 20982
rect 19517 20979 19583 20982
rect 22050 21040 32187 21042
rect 22050 20984 27158 21040
rect 27214 20984 32126 21040
rect 32182 20984 32187 21040
rect 22050 20982 32187 20984
rect 15285 20906 15351 20909
rect 16297 20906 16363 20909
rect 15285 20904 16363 20906
rect 15285 20848 15290 20904
rect 15346 20848 16302 20904
rect 16358 20848 16363 20904
rect 15285 20846 16363 20848
rect 15285 20843 15351 20846
rect 16297 20843 16363 20846
rect 16481 20906 16547 20909
rect 17401 20906 17467 20909
rect 18045 20906 18111 20909
rect 16481 20904 18111 20906
rect 16481 20848 16486 20904
rect 16542 20848 17406 20904
rect 17462 20848 18050 20904
rect 18106 20848 18111 20904
rect 16481 20846 18111 20848
rect 16481 20843 16547 20846
rect 17401 20843 17467 20846
rect 18045 20843 18111 20846
rect 18229 20906 18295 20909
rect 22050 20906 22110 20982
rect 27153 20979 27219 20982
rect 32121 20979 32187 20982
rect 32581 21042 32647 21045
rect 33225 21042 33291 21045
rect 32581 21040 33291 21042
rect 32581 20984 32586 21040
rect 32642 20984 33230 21040
rect 33286 20984 33291 21040
rect 32581 20982 33291 20984
rect 33366 21042 33426 21118
rect 37825 21042 37891 21045
rect 33366 21040 37891 21042
rect 33366 20984 37830 21040
rect 37886 20984 37891 21040
rect 33366 20982 37891 20984
rect 32581 20979 32647 20982
rect 33225 20979 33291 20982
rect 37825 20979 37891 20982
rect 18229 20904 22110 20906
rect 18229 20848 18234 20904
rect 18290 20848 22110 20904
rect 18229 20846 22110 20848
rect 23013 20906 23079 20909
rect 26734 20906 26740 20908
rect 23013 20904 26740 20906
rect 23013 20848 23018 20904
rect 23074 20848 26740 20904
rect 23013 20846 26740 20848
rect 18229 20843 18295 20846
rect 23013 20843 23079 20846
rect 26734 20844 26740 20846
rect 26804 20844 26810 20908
rect 29913 20906 29979 20909
rect 34697 20906 34763 20909
rect 41873 20906 41939 20909
rect 29913 20904 34763 20906
rect 29913 20848 29918 20904
rect 29974 20848 34702 20904
rect 34758 20848 34763 20904
rect 29913 20846 34763 20848
rect 29913 20843 29979 20846
rect 34697 20843 34763 20846
rect 34838 20904 41939 20906
rect 34838 20848 41878 20904
rect 41934 20848 41939 20904
rect 34838 20846 41939 20848
rect -300 20770 160 20800
rect 933 20770 999 20773
rect -300 20768 999 20770
rect -300 20712 938 20768
rect 994 20712 999 20768
rect -300 20710 999 20712
rect -300 20680 160 20710
rect 933 20707 999 20710
rect 8937 20770 9003 20773
rect 9254 20770 9260 20772
rect 8937 20768 9260 20770
rect 8937 20712 8942 20768
rect 8998 20712 9260 20768
rect 8937 20710 9260 20712
rect 8937 20707 9003 20710
rect 9254 20708 9260 20710
rect 9324 20708 9330 20772
rect 16982 20708 16988 20772
rect 17052 20770 17058 20772
rect 17125 20770 17191 20773
rect 17493 20772 17559 20773
rect 19793 20772 19859 20773
rect 17493 20770 17540 20772
rect 17052 20768 17191 20770
rect 17052 20712 17130 20768
rect 17186 20712 17191 20768
rect 17052 20710 17191 20712
rect 17448 20768 17540 20770
rect 17448 20712 17498 20768
rect 17448 20710 17540 20712
rect 17052 20708 17058 20710
rect 17125 20707 17191 20710
rect 17493 20708 17540 20710
rect 17604 20708 17610 20772
rect 19742 20708 19748 20772
rect 19812 20770 19859 20772
rect 19812 20768 19904 20770
rect 19854 20712 19904 20768
rect 19812 20710 19904 20712
rect 19812 20708 19859 20710
rect 21582 20708 21588 20772
rect 21652 20770 21658 20772
rect 22369 20770 22435 20773
rect 23289 20772 23355 20773
rect 21652 20768 22435 20770
rect 21652 20712 22374 20768
rect 22430 20712 22435 20768
rect 21652 20710 22435 20712
rect 21652 20708 21658 20710
rect 17493 20707 17559 20708
rect 19793 20707 19859 20708
rect 22369 20707 22435 20710
rect 23238 20708 23244 20772
rect 23308 20770 23355 20772
rect 24853 20770 24919 20773
rect 25446 20770 25452 20772
rect 23308 20768 23400 20770
rect 23350 20712 23400 20768
rect 23308 20710 23400 20712
rect 24853 20768 25452 20770
rect 24853 20712 24858 20768
rect 24914 20712 25452 20768
rect 24853 20710 25452 20712
rect 23308 20708 23355 20710
rect 23289 20707 23355 20708
rect 24853 20707 24919 20710
rect 25446 20708 25452 20710
rect 25516 20708 25522 20772
rect 27654 20708 27660 20772
rect 27724 20770 27730 20772
rect 29085 20770 29151 20773
rect 27724 20768 29151 20770
rect 27724 20712 29090 20768
rect 29146 20712 29151 20768
rect 27724 20710 29151 20712
rect 27724 20708 27730 20710
rect 29085 20707 29151 20710
rect 31886 20708 31892 20772
rect 31956 20770 31962 20772
rect 32949 20770 33015 20773
rect 31956 20768 33015 20770
rect 31956 20712 32954 20768
rect 33010 20712 33015 20768
rect 31956 20710 33015 20712
rect 31956 20708 31962 20710
rect 32949 20707 33015 20710
rect 6066 20704 6382 20705
rect 6066 20640 6072 20704
rect 6136 20640 6152 20704
rect 6216 20640 6232 20704
rect 6296 20640 6312 20704
rect 6376 20640 6382 20704
rect 6066 20639 6382 20640
rect 11066 20704 11382 20705
rect 11066 20640 11072 20704
rect 11136 20640 11152 20704
rect 11216 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11382 20704
rect 11066 20639 11382 20640
rect 16066 20704 16382 20705
rect 16066 20640 16072 20704
rect 16136 20640 16152 20704
rect 16216 20640 16232 20704
rect 16296 20640 16312 20704
rect 16376 20640 16382 20704
rect 16066 20639 16382 20640
rect 21066 20704 21382 20705
rect 21066 20640 21072 20704
rect 21136 20640 21152 20704
rect 21216 20640 21232 20704
rect 21296 20640 21312 20704
rect 21376 20640 21382 20704
rect 21066 20639 21382 20640
rect 26066 20704 26382 20705
rect 26066 20640 26072 20704
rect 26136 20640 26152 20704
rect 26216 20640 26232 20704
rect 26296 20640 26312 20704
rect 26376 20640 26382 20704
rect 26066 20639 26382 20640
rect 31066 20704 31382 20705
rect 31066 20640 31072 20704
rect 31136 20640 31152 20704
rect 31216 20640 31232 20704
rect 31296 20640 31312 20704
rect 31376 20640 31382 20704
rect 31066 20639 31382 20640
rect 30741 20634 30807 20637
rect 28950 20632 30807 20634
rect 28950 20576 30746 20632
rect 30802 20576 30807 20632
rect 28950 20574 30807 20576
rect 14273 20498 14339 20501
rect 14457 20498 14523 20501
rect 15745 20498 15811 20501
rect 16573 20498 16639 20501
rect 14273 20496 16639 20498
rect 14273 20440 14278 20496
rect 14334 20440 14462 20496
rect 14518 20440 15750 20496
rect 15806 20440 16578 20496
rect 16634 20440 16639 20496
rect 14273 20438 16639 20440
rect 14273 20435 14339 20438
rect 14457 20435 14523 20438
rect 15745 20435 15811 20438
rect 16573 20435 16639 20438
rect 16941 20498 17007 20501
rect 20069 20498 20135 20501
rect 16941 20496 20135 20498
rect 16941 20440 16946 20496
rect 17002 20440 20074 20496
rect 20130 20440 20135 20496
rect 16941 20438 20135 20440
rect 16941 20435 17007 20438
rect 20069 20435 20135 20438
rect 22093 20498 22159 20501
rect 27705 20498 27771 20501
rect 28950 20498 29010 20574
rect 30741 20571 30807 20574
rect 32765 20634 32831 20637
rect 34838 20634 34898 20846
rect 41873 20843 41939 20846
rect 45185 20770 45251 20773
rect 45840 20770 46300 20800
rect 45185 20768 46300 20770
rect 45185 20712 45190 20768
rect 45246 20712 46300 20768
rect 45185 20710 46300 20712
rect 45185 20707 45251 20710
rect 36066 20704 36382 20705
rect 36066 20640 36072 20704
rect 36136 20640 36152 20704
rect 36216 20640 36232 20704
rect 36296 20640 36312 20704
rect 36376 20640 36382 20704
rect 36066 20639 36382 20640
rect 41066 20704 41382 20705
rect 41066 20640 41072 20704
rect 41136 20640 41152 20704
rect 41216 20640 41232 20704
rect 41296 20640 41312 20704
rect 41376 20640 41382 20704
rect 45840 20680 46300 20710
rect 41066 20639 41382 20640
rect 32765 20632 34898 20634
rect 32765 20576 32770 20632
rect 32826 20576 34898 20632
rect 32765 20574 34898 20576
rect 32765 20571 32831 20574
rect 22093 20496 29010 20498
rect 22093 20440 22098 20496
rect 22154 20440 27710 20496
rect 27766 20440 29010 20496
rect 22093 20438 29010 20440
rect 29177 20498 29243 20501
rect 32029 20498 32095 20501
rect 29177 20496 32095 20498
rect 29177 20440 29182 20496
rect 29238 20440 32034 20496
rect 32090 20440 32095 20496
rect 29177 20438 32095 20440
rect 22093 20435 22159 20438
rect 27705 20435 27771 20438
rect 29177 20435 29243 20438
rect 32029 20435 32095 20438
rect 32949 20498 33015 20501
rect 38009 20498 38075 20501
rect 32949 20496 38075 20498
rect 32949 20440 32954 20496
rect 33010 20440 38014 20496
rect 38070 20440 38075 20496
rect 32949 20438 38075 20440
rect 32949 20435 33015 20438
rect 38009 20435 38075 20438
rect 11605 20362 11671 20365
rect 26550 20362 26556 20364
rect 11605 20360 26556 20362
rect 11605 20304 11610 20360
rect 11666 20304 26556 20360
rect 11605 20302 26556 20304
rect 11605 20299 11671 20302
rect 26550 20300 26556 20302
rect 26620 20362 26626 20364
rect 32305 20362 32371 20365
rect 26620 20360 32371 20362
rect 26620 20304 32310 20360
rect 32366 20304 32371 20360
rect 26620 20302 32371 20304
rect 26620 20300 26626 20302
rect 32305 20299 32371 20302
rect 33225 20362 33291 20365
rect 34329 20362 34395 20365
rect 43805 20362 43871 20365
rect 33225 20360 43871 20362
rect 33225 20304 33230 20360
rect 33286 20304 34334 20360
rect 34390 20304 43810 20360
rect 43866 20304 43871 20360
rect 33225 20302 43871 20304
rect 33225 20299 33291 20302
rect 34329 20299 34395 20302
rect 43805 20299 43871 20302
rect 14917 20226 14983 20229
rect 17033 20226 17099 20229
rect 14917 20224 17099 20226
rect 14917 20168 14922 20224
rect 14978 20168 17038 20224
rect 17094 20168 17099 20224
rect 14917 20166 17099 20168
rect 14917 20163 14983 20166
rect 17033 20163 17099 20166
rect 30741 20226 30807 20229
rect 31661 20226 31727 20229
rect 30741 20224 31727 20226
rect 30741 20168 30746 20224
rect 30802 20168 31666 20224
rect 31722 20168 31727 20224
rect 30741 20166 31727 20168
rect 30741 20163 30807 20166
rect 31661 20163 31727 20166
rect 3566 20160 3882 20161
rect 3566 20096 3572 20160
rect 3636 20096 3652 20160
rect 3716 20096 3732 20160
rect 3796 20096 3812 20160
rect 3876 20096 3882 20160
rect 3566 20095 3882 20096
rect 8566 20160 8882 20161
rect 8566 20096 8572 20160
rect 8636 20096 8652 20160
rect 8716 20096 8732 20160
rect 8796 20096 8812 20160
rect 8876 20096 8882 20160
rect 8566 20095 8882 20096
rect 13566 20160 13882 20161
rect 13566 20096 13572 20160
rect 13636 20096 13652 20160
rect 13716 20096 13732 20160
rect 13796 20096 13812 20160
rect 13876 20096 13882 20160
rect 13566 20095 13882 20096
rect 18566 20160 18882 20161
rect 18566 20096 18572 20160
rect 18636 20096 18652 20160
rect 18716 20096 18732 20160
rect 18796 20096 18812 20160
rect 18876 20096 18882 20160
rect 18566 20095 18882 20096
rect 23566 20160 23882 20161
rect 23566 20096 23572 20160
rect 23636 20096 23652 20160
rect 23716 20096 23732 20160
rect 23796 20096 23812 20160
rect 23876 20096 23882 20160
rect 23566 20095 23882 20096
rect 28566 20160 28882 20161
rect 28566 20096 28572 20160
rect 28636 20096 28652 20160
rect 28716 20096 28732 20160
rect 28796 20096 28812 20160
rect 28876 20096 28882 20160
rect 28566 20095 28882 20096
rect 33566 20160 33882 20161
rect 33566 20096 33572 20160
rect 33636 20096 33652 20160
rect 33716 20096 33732 20160
rect 33796 20096 33812 20160
rect 33876 20096 33882 20160
rect 33566 20095 33882 20096
rect 38566 20160 38882 20161
rect 38566 20096 38572 20160
rect 38636 20096 38652 20160
rect 38716 20096 38732 20160
rect 38796 20096 38812 20160
rect 38876 20096 38882 20160
rect 38566 20095 38882 20096
rect 43566 20160 43882 20161
rect 43566 20096 43572 20160
rect 43636 20096 43652 20160
rect 43716 20096 43732 20160
rect 43796 20096 43812 20160
rect 43876 20096 43882 20160
rect 43566 20095 43882 20096
rect 14181 20090 14247 20093
rect 16665 20090 16731 20093
rect 14181 20088 16731 20090
rect 14181 20032 14186 20088
rect 14242 20032 16670 20088
rect 16726 20032 16731 20088
rect 14181 20030 16731 20032
rect 14181 20027 14247 20030
rect 16665 20027 16731 20030
rect 30373 20090 30439 20093
rect 31017 20090 31083 20093
rect 33317 20090 33383 20093
rect 30373 20088 31083 20090
rect 30373 20032 30378 20088
rect 30434 20032 31022 20088
rect 31078 20032 31083 20088
rect 30373 20030 31083 20032
rect 30373 20027 30439 20030
rect 31017 20027 31083 20030
rect 31710 20088 33383 20090
rect 31710 20032 33322 20088
rect 33378 20032 33383 20088
rect 31710 20030 33383 20032
rect 5441 19954 5507 19957
rect 17217 19954 17283 19957
rect 5441 19952 17283 19954
rect 5441 19896 5446 19952
rect 5502 19896 17222 19952
rect 17278 19896 17283 19952
rect 5441 19894 17283 19896
rect 5441 19891 5507 19894
rect 17217 19891 17283 19894
rect 17585 19954 17651 19957
rect 19425 19954 19491 19957
rect 17585 19952 19491 19954
rect 17585 19896 17590 19952
rect 17646 19896 19430 19952
rect 19486 19896 19491 19952
rect 17585 19894 19491 19896
rect 17585 19891 17651 19894
rect 19425 19891 19491 19894
rect 20069 19954 20135 19957
rect 20989 19954 21055 19957
rect 20069 19952 21055 19954
rect 20069 19896 20074 19952
rect 20130 19896 20994 19952
rect 21050 19896 21055 19952
rect 20069 19894 21055 19896
rect 20069 19891 20135 19894
rect 20989 19891 21055 19894
rect 24853 19954 24919 19957
rect 25865 19954 25931 19957
rect 28349 19954 28415 19957
rect 24853 19952 28415 19954
rect 24853 19896 24858 19952
rect 24914 19896 25870 19952
rect 25926 19896 28354 19952
rect 28410 19896 28415 19952
rect 24853 19894 28415 19896
rect 24853 19891 24919 19894
rect 25865 19891 25931 19894
rect 28349 19891 28415 19894
rect 28625 19954 28691 19957
rect 31710 19954 31770 20030
rect 33317 20027 33383 20030
rect 28625 19952 31770 19954
rect 28625 19896 28630 19952
rect 28686 19896 31770 19952
rect 28625 19894 31770 19896
rect 28625 19891 28691 19894
rect 12065 19818 12131 19821
rect 23054 19818 23060 19820
rect 12065 19816 23060 19818
rect 12065 19760 12070 19816
rect 12126 19760 23060 19816
rect 12065 19758 23060 19760
rect 12065 19755 12131 19758
rect 23054 19756 23060 19758
rect 23124 19818 23130 19820
rect 23124 19758 25514 19818
rect 23124 19756 23130 19758
rect 18321 19682 18387 19685
rect 19057 19682 19123 19685
rect 18321 19680 19123 19682
rect 18321 19624 18326 19680
rect 18382 19624 19062 19680
rect 19118 19624 19123 19680
rect 18321 19622 19123 19624
rect 18321 19619 18387 19622
rect 19057 19619 19123 19622
rect 19701 19682 19767 19685
rect 20529 19682 20595 19685
rect 19701 19680 20595 19682
rect 19701 19624 19706 19680
rect 19762 19624 20534 19680
rect 20590 19624 20595 19680
rect 19701 19622 20595 19624
rect 19701 19619 19767 19622
rect 20529 19619 20595 19622
rect 6066 19616 6382 19617
rect 6066 19552 6072 19616
rect 6136 19552 6152 19616
rect 6216 19552 6232 19616
rect 6296 19552 6312 19616
rect 6376 19552 6382 19616
rect 6066 19551 6382 19552
rect 11066 19616 11382 19617
rect 11066 19552 11072 19616
rect 11136 19552 11152 19616
rect 11216 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11382 19616
rect 11066 19551 11382 19552
rect 16066 19616 16382 19617
rect 16066 19552 16072 19616
rect 16136 19552 16152 19616
rect 16216 19552 16232 19616
rect 16296 19552 16312 19616
rect 16376 19552 16382 19616
rect 16066 19551 16382 19552
rect 21066 19616 21382 19617
rect 21066 19552 21072 19616
rect 21136 19552 21152 19616
rect 21216 19552 21232 19616
rect 21296 19552 21312 19616
rect 21376 19552 21382 19616
rect 21066 19551 21382 19552
rect 17217 19410 17283 19413
rect 24342 19410 24348 19412
rect 17217 19408 24348 19410
rect 17217 19352 17222 19408
rect 17278 19352 24348 19408
rect 17217 19350 24348 19352
rect 17217 19347 17283 19350
rect 24342 19348 24348 19350
rect 24412 19410 24418 19412
rect 25313 19410 25379 19413
rect 24412 19408 25379 19410
rect 24412 19352 25318 19408
rect 25374 19352 25379 19408
rect 24412 19350 25379 19352
rect 25454 19410 25514 19758
rect 25630 19756 25636 19820
rect 25700 19818 25706 19820
rect 26141 19818 26207 19821
rect 32489 19818 32555 19821
rect 25700 19816 26207 19818
rect 25700 19760 26146 19816
rect 26202 19760 26207 19816
rect 25700 19758 26207 19760
rect 25700 19756 25706 19758
rect 26141 19755 26207 19758
rect 26558 19816 32555 19818
rect 26558 19760 32494 19816
rect 32550 19760 32555 19816
rect 26558 19758 32555 19760
rect 26066 19616 26382 19617
rect 26066 19552 26072 19616
rect 26136 19552 26152 19616
rect 26216 19552 26232 19616
rect 26296 19552 26312 19616
rect 26376 19552 26382 19616
rect 26066 19551 26382 19552
rect 26558 19410 26618 19758
rect 32489 19755 32555 19758
rect 34145 19818 34211 19821
rect 38745 19818 38811 19821
rect 34145 19816 38811 19818
rect 34145 19760 34150 19816
rect 34206 19760 38750 19816
rect 38806 19760 38811 19816
rect 34145 19758 38811 19760
rect 34145 19755 34211 19758
rect 38745 19755 38811 19758
rect 31066 19616 31382 19617
rect 31066 19552 31072 19616
rect 31136 19552 31152 19616
rect 31216 19552 31232 19616
rect 31296 19552 31312 19616
rect 31376 19552 31382 19616
rect 31066 19551 31382 19552
rect 36066 19616 36382 19617
rect 36066 19552 36072 19616
rect 36136 19552 36152 19616
rect 36216 19552 36232 19616
rect 36296 19552 36312 19616
rect 36376 19552 36382 19616
rect 36066 19551 36382 19552
rect 41066 19616 41382 19617
rect 41066 19552 41072 19616
rect 41136 19552 41152 19616
rect 41216 19552 41232 19616
rect 41296 19552 41312 19616
rect 41376 19552 41382 19616
rect 41066 19551 41382 19552
rect 28073 19546 28139 19549
rect 28625 19546 28691 19549
rect 28073 19544 28691 19546
rect 28073 19488 28078 19544
rect 28134 19488 28630 19544
rect 28686 19488 28691 19544
rect 28073 19486 28691 19488
rect 28073 19483 28139 19486
rect 28625 19483 28691 19486
rect 29637 19546 29703 19549
rect 30925 19546 30991 19549
rect 29637 19544 30991 19546
rect 29637 19488 29642 19544
rect 29698 19488 30930 19544
rect 30986 19488 30991 19544
rect 29637 19486 30991 19488
rect 29637 19483 29703 19486
rect 30925 19483 30991 19486
rect 25454 19350 26618 19410
rect 28257 19410 28323 19413
rect 30465 19410 30531 19413
rect 28257 19408 30531 19410
rect 28257 19352 28262 19408
rect 28318 19352 30470 19408
rect 30526 19352 30531 19408
rect 28257 19350 30531 19352
rect 24412 19348 24418 19350
rect 25313 19347 25379 19350
rect 28257 19347 28323 19350
rect 30465 19347 30531 19350
rect 6729 19274 6795 19277
rect 38929 19274 38995 19277
rect 6729 19272 38995 19274
rect 6729 19216 6734 19272
rect 6790 19216 38934 19272
rect 38990 19216 38995 19272
rect 6729 19214 38995 19216
rect 6729 19211 6795 19214
rect 38929 19211 38995 19214
rect 3566 19072 3882 19073
rect 3566 19008 3572 19072
rect 3636 19008 3652 19072
rect 3716 19008 3732 19072
rect 3796 19008 3812 19072
rect 3876 19008 3882 19072
rect 3566 19007 3882 19008
rect 8566 19072 8882 19073
rect 8566 19008 8572 19072
rect 8636 19008 8652 19072
rect 8716 19008 8732 19072
rect 8796 19008 8812 19072
rect 8876 19008 8882 19072
rect 8566 19007 8882 19008
rect 13566 19072 13882 19073
rect 13566 19008 13572 19072
rect 13636 19008 13652 19072
rect 13716 19008 13732 19072
rect 13796 19008 13812 19072
rect 13876 19008 13882 19072
rect 13566 19007 13882 19008
rect 18566 19072 18882 19073
rect 18566 19008 18572 19072
rect 18636 19008 18652 19072
rect 18716 19008 18732 19072
rect 18796 19008 18812 19072
rect 18876 19008 18882 19072
rect 18566 19007 18882 19008
rect 23566 19072 23882 19073
rect 23566 19008 23572 19072
rect 23636 19008 23652 19072
rect 23716 19008 23732 19072
rect 23796 19008 23812 19072
rect 23876 19008 23882 19072
rect 23566 19007 23882 19008
rect 28566 19072 28882 19073
rect 28566 19008 28572 19072
rect 28636 19008 28652 19072
rect 28716 19008 28732 19072
rect 28796 19008 28812 19072
rect 28876 19008 28882 19072
rect 28566 19007 28882 19008
rect 33566 19072 33882 19073
rect 33566 19008 33572 19072
rect 33636 19008 33652 19072
rect 33716 19008 33732 19072
rect 33796 19008 33812 19072
rect 33876 19008 33882 19072
rect 33566 19007 33882 19008
rect 38566 19072 38882 19073
rect 38566 19008 38572 19072
rect 38636 19008 38652 19072
rect 38716 19008 38732 19072
rect 38796 19008 38812 19072
rect 38876 19008 38882 19072
rect 38566 19007 38882 19008
rect 43566 19072 43882 19073
rect 43566 19008 43572 19072
rect 43636 19008 43652 19072
rect 43716 19008 43732 19072
rect 43796 19008 43812 19072
rect 43876 19008 43882 19072
rect 43566 19007 43882 19008
rect 20253 19002 20319 19005
rect 21173 19002 21239 19005
rect 20253 19000 21239 19002
rect 20253 18944 20258 19000
rect 20314 18944 21178 19000
rect 21234 18944 21239 19000
rect 20253 18942 21239 18944
rect 20253 18939 20319 18942
rect 21173 18939 21239 18942
rect 30741 19002 30807 19005
rect 31569 19002 31635 19005
rect 30741 19000 31635 19002
rect 30741 18944 30746 19000
rect 30802 18944 31574 19000
rect 31630 18944 31635 19000
rect 30741 18942 31635 18944
rect 30741 18939 30807 18942
rect 31569 18939 31635 18942
rect 13997 18866 14063 18869
rect 26877 18866 26943 18869
rect 13997 18864 26943 18866
rect 13997 18808 14002 18864
rect 14058 18808 26882 18864
rect 26938 18808 26943 18864
rect 13997 18806 26943 18808
rect 13997 18803 14063 18806
rect 26877 18803 26943 18806
rect 29821 18866 29887 18869
rect 35157 18866 35223 18869
rect 29821 18864 35223 18866
rect 29821 18808 29826 18864
rect 29882 18808 35162 18864
rect 35218 18808 35223 18864
rect 29821 18806 35223 18808
rect 29821 18803 29887 18806
rect 35157 18803 35223 18806
rect 17953 18730 18019 18733
rect 19057 18730 19123 18733
rect 17953 18728 19123 18730
rect 17953 18672 17958 18728
rect 18014 18672 19062 18728
rect 19118 18672 19123 18728
rect 17953 18670 19123 18672
rect 17953 18667 18019 18670
rect 19057 18667 19123 18670
rect 19425 18730 19491 18733
rect 21950 18730 21956 18732
rect 19425 18728 21956 18730
rect 19425 18672 19430 18728
rect 19486 18672 21956 18728
rect 19425 18670 21956 18672
rect 19425 18667 19491 18670
rect 21950 18668 21956 18670
rect 22020 18730 22026 18732
rect 34237 18730 34303 18733
rect 22020 18728 34303 18730
rect 22020 18672 34242 18728
rect 34298 18672 34303 18728
rect 22020 18670 34303 18672
rect 22020 18668 22026 18670
rect 34237 18667 34303 18670
rect 6066 18528 6382 18529
rect 6066 18464 6072 18528
rect 6136 18464 6152 18528
rect 6216 18464 6232 18528
rect 6296 18464 6312 18528
rect 6376 18464 6382 18528
rect 6066 18463 6382 18464
rect 11066 18528 11382 18529
rect 11066 18464 11072 18528
rect 11136 18464 11152 18528
rect 11216 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11382 18528
rect 11066 18463 11382 18464
rect 16066 18528 16382 18529
rect 16066 18464 16072 18528
rect 16136 18464 16152 18528
rect 16216 18464 16232 18528
rect 16296 18464 16312 18528
rect 16376 18464 16382 18528
rect 16066 18463 16382 18464
rect 21066 18528 21382 18529
rect 21066 18464 21072 18528
rect 21136 18464 21152 18528
rect 21216 18464 21232 18528
rect 21296 18464 21312 18528
rect 21376 18464 21382 18528
rect 21066 18463 21382 18464
rect 26066 18528 26382 18529
rect 26066 18464 26072 18528
rect 26136 18464 26152 18528
rect 26216 18464 26232 18528
rect 26296 18464 26312 18528
rect 26376 18464 26382 18528
rect 26066 18463 26382 18464
rect 31066 18528 31382 18529
rect 31066 18464 31072 18528
rect 31136 18464 31152 18528
rect 31216 18464 31232 18528
rect 31296 18464 31312 18528
rect 31376 18464 31382 18528
rect 31066 18463 31382 18464
rect 36066 18528 36382 18529
rect 36066 18464 36072 18528
rect 36136 18464 36152 18528
rect 36216 18464 36232 18528
rect 36296 18464 36312 18528
rect 36376 18464 36382 18528
rect 36066 18463 36382 18464
rect 41066 18528 41382 18529
rect 41066 18464 41072 18528
rect 41136 18464 41152 18528
rect 41216 18464 41232 18528
rect 41296 18464 41312 18528
rect 41376 18464 41382 18528
rect 41066 18463 41382 18464
rect 23197 18458 23263 18461
rect 23933 18458 23999 18461
rect 25681 18458 25747 18461
rect 23197 18456 25747 18458
rect 23197 18400 23202 18456
rect 23258 18400 23938 18456
rect 23994 18400 25686 18456
rect 25742 18400 25747 18456
rect 23197 18398 25747 18400
rect 23197 18395 23263 18398
rect 23933 18395 23999 18398
rect 25681 18395 25747 18398
rect 16481 18322 16547 18325
rect 17033 18322 17099 18325
rect 17953 18322 18019 18325
rect 16481 18320 17099 18322
rect 16481 18264 16486 18320
rect 16542 18264 17038 18320
rect 17094 18264 17099 18320
rect 16481 18262 17099 18264
rect 16481 18259 16547 18262
rect 17033 18259 17099 18262
rect 17358 18320 18019 18322
rect 17358 18264 17958 18320
rect 18014 18264 18019 18320
rect 17358 18262 18019 18264
rect 15285 18186 15351 18189
rect 17125 18186 17191 18189
rect 17358 18186 17418 18262
rect 17953 18259 18019 18262
rect 24853 18322 24919 18325
rect 25957 18322 26023 18325
rect 24853 18320 26023 18322
rect 24853 18264 24858 18320
rect 24914 18264 25962 18320
rect 26018 18264 26023 18320
rect 24853 18262 26023 18264
rect 24853 18259 24919 18262
rect 25957 18259 26023 18262
rect 29085 18322 29151 18325
rect 34237 18322 34303 18325
rect 29085 18320 34303 18322
rect 29085 18264 29090 18320
rect 29146 18264 34242 18320
rect 34298 18264 34303 18320
rect 29085 18262 34303 18264
rect 29085 18259 29151 18262
rect 34237 18259 34303 18262
rect 15285 18184 17418 18186
rect 15285 18128 15290 18184
rect 15346 18128 17130 18184
rect 17186 18128 17418 18184
rect 15285 18126 17418 18128
rect 17493 18186 17559 18189
rect 17769 18186 17835 18189
rect 17493 18184 17835 18186
rect 17493 18128 17498 18184
rect 17554 18128 17774 18184
rect 17830 18128 17835 18184
rect 17493 18126 17835 18128
rect 15285 18123 15351 18126
rect 17125 18123 17191 18126
rect 17493 18123 17559 18126
rect 17769 18123 17835 18126
rect 31201 18186 31267 18189
rect 32857 18186 32923 18189
rect 31201 18184 32923 18186
rect 31201 18128 31206 18184
rect 31262 18128 32862 18184
rect 32918 18128 32923 18184
rect 31201 18126 32923 18128
rect 31201 18123 31267 18126
rect 32857 18123 32923 18126
rect 16573 18050 16639 18053
rect 17309 18050 17375 18053
rect 16573 18048 17375 18050
rect 16573 17992 16578 18048
rect 16634 17992 17314 18048
rect 17370 17992 17375 18048
rect 16573 17990 17375 17992
rect 16573 17987 16639 17990
rect 17309 17987 17375 17990
rect 3566 17984 3882 17985
rect 3566 17920 3572 17984
rect 3636 17920 3652 17984
rect 3716 17920 3732 17984
rect 3796 17920 3812 17984
rect 3876 17920 3882 17984
rect 3566 17919 3882 17920
rect 8566 17984 8882 17985
rect 8566 17920 8572 17984
rect 8636 17920 8652 17984
rect 8716 17920 8732 17984
rect 8796 17920 8812 17984
rect 8876 17920 8882 17984
rect 8566 17919 8882 17920
rect 13566 17984 13882 17985
rect 13566 17920 13572 17984
rect 13636 17920 13652 17984
rect 13716 17920 13732 17984
rect 13796 17920 13812 17984
rect 13876 17920 13882 17984
rect 13566 17919 13882 17920
rect 18566 17984 18882 17985
rect 18566 17920 18572 17984
rect 18636 17920 18652 17984
rect 18716 17920 18732 17984
rect 18796 17920 18812 17984
rect 18876 17920 18882 17984
rect 18566 17919 18882 17920
rect 23566 17984 23882 17985
rect 23566 17920 23572 17984
rect 23636 17920 23652 17984
rect 23716 17920 23732 17984
rect 23796 17920 23812 17984
rect 23876 17920 23882 17984
rect 23566 17919 23882 17920
rect 28566 17984 28882 17985
rect 28566 17920 28572 17984
rect 28636 17920 28652 17984
rect 28716 17920 28732 17984
rect 28796 17920 28812 17984
rect 28876 17920 28882 17984
rect 28566 17919 28882 17920
rect 33566 17984 33882 17985
rect 33566 17920 33572 17984
rect 33636 17920 33652 17984
rect 33716 17920 33732 17984
rect 33796 17920 33812 17984
rect 33876 17920 33882 17984
rect 33566 17919 33882 17920
rect 38566 17984 38882 17985
rect 38566 17920 38572 17984
rect 38636 17920 38652 17984
rect 38716 17920 38732 17984
rect 38796 17920 38812 17984
rect 38876 17920 38882 17984
rect 38566 17919 38882 17920
rect 43566 17984 43882 17985
rect 43566 17920 43572 17984
rect 43636 17920 43652 17984
rect 43716 17920 43732 17984
rect 43796 17920 43812 17984
rect 43876 17920 43882 17984
rect 43566 17919 43882 17920
rect 16389 17914 16455 17917
rect 17953 17914 18019 17917
rect 16389 17912 18019 17914
rect 16389 17856 16394 17912
rect 16450 17856 17958 17912
rect 18014 17856 18019 17912
rect 16389 17854 18019 17856
rect 16389 17851 16455 17854
rect 17953 17851 18019 17854
rect 16389 17778 16455 17781
rect 18229 17778 18295 17781
rect 37733 17778 37799 17781
rect 40033 17778 40099 17781
rect 16389 17776 18295 17778
rect 16389 17720 16394 17776
rect 16450 17720 18234 17776
rect 18290 17720 18295 17776
rect 16389 17718 18295 17720
rect 16389 17715 16455 17718
rect 18229 17715 18295 17718
rect 22050 17776 40099 17778
rect 22050 17720 37738 17776
rect 37794 17720 40038 17776
rect 40094 17720 40099 17776
rect 22050 17718 40099 17720
rect 19793 17642 19859 17645
rect 22050 17642 22110 17718
rect 37733 17715 37799 17718
rect 40033 17715 40099 17718
rect 19793 17640 22110 17642
rect 19793 17584 19798 17640
rect 19854 17584 22110 17640
rect 19793 17582 22110 17584
rect 29913 17642 29979 17645
rect 31569 17642 31635 17645
rect 29913 17640 31635 17642
rect 29913 17584 29918 17640
rect 29974 17584 31574 17640
rect 31630 17584 31635 17640
rect 29913 17582 31635 17584
rect 19793 17579 19859 17582
rect 29913 17579 29979 17582
rect 31569 17579 31635 17582
rect 30465 17508 30531 17509
rect 30414 17506 30420 17508
rect 30374 17446 30420 17506
rect 30484 17504 30531 17508
rect 30526 17448 30531 17504
rect 30414 17444 30420 17446
rect 30484 17444 30531 17448
rect 30465 17443 30531 17444
rect 6066 17440 6382 17441
rect 6066 17376 6072 17440
rect 6136 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6382 17440
rect 6066 17375 6382 17376
rect 11066 17440 11382 17441
rect 11066 17376 11072 17440
rect 11136 17376 11152 17440
rect 11216 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11382 17440
rect 11066 17375 11382 17376
rect 16066 17440 16382 17441
rect 16066 17376 16072 17440
rect 16136 17376 16152 17440
rect 16216 17376 16232 17440
rect 16296 17376 16312 17440
rect 16376 17376 16382 17440
rect 16066 17375 16382 17376
rect 21066 17440 21382 17441
rect 21066 17376 21072 17440
rect 21136 17376 21152 17440
rect 21216 17376 21232 17440
rect 21296 17376 21312 17440
rect 21376 17376 21382 17440
rect 21066 17375 21382 17376
rect 26066 17440 26382 17441
rect 26066 17376 26072 17440
rect 26136 17376 26152 17440
rect 26216 17376 26232 17440
rect 26296 17376 26312 17440
rect 26376 17376 26382 17440
rect 26066 17375 26382 17376
rect 31066 17440 31382 17441
rect 31066 17376 31072 17440
rect 31136 17376 31152 17440
rect 31216 17376 31232 17440
rect 31296 17376 31312 17440
rect 31376 17376 31382 17440
rect 31066 17375 31382 17376
rect 36066 17440 36382 17441
rect 36066 17376 36072 17440
rect 36136 17376 36152 17440
rect 36216 17376 36232 17440
rect 36296 17376 36312 17440
rect 36376 17376 36382 17440
rect 36066 17375 36382 17376
rect 41066 17440 41382 17441
rect 41066 17376 41072 17440
rect 41136 17376 41152 17440
rect 41216 17376 41232 17440
rect 41296 17376 41312 17440
rect 41376 17376 41382 17440
rect 41066 17375 41382 17376
rect 19701 17370 19767 17373
rect 20437 17370 20503 17373
rect 19701 17368 20503 17370
rect 19701 17312 19706 17368
rect 19762 17312 20442 17368
rect 20498 17312 20503 17368
rect 19701 17310 20503 17312
rect 19701 17307 19767 17310
rect 20437 17307 20503 17310
rect 13077 17234 13143 17237
rect 22870 17234 22876 17236
rect 13077 17232 22876 17234
rect 13077 17176 13082 17232
rect 13138 17176 22876 17232
rect 13077 17174 22876 17176
rect 13077 17171 13143 17174
rect 22870 17172 22876 17174
rect 22940 17234 22946 17236
rect 31753 17234 31819 17237
rect 32857 17236 32923 17237
rect 22940 17232 31819 17234
rect 22940 17176 31758 17232
rect 31814 17176 31819 17232
rect 22940 17174 31819 17176
rect 22940 17172 22946 17174
rect 31753 17171 31819 17174
rect 32806 17172 32812 17236
rect 32876 17234 32923 17236
rect 32876 17232 32968 17234
rect 32918 17176 32968 17232
rect 32876 17174 32968 17176
rect 32876 17172 32923 17174
rect 32857 17171 32923 17172
rect 8201 17098 8267 17101
rect 20897 17098 20963 17101
rect 8201 17096 20963 17098
rect 8201 17040 8206 17096
rect 8262 17040 20902 17096
rect 20958 17040 20963 17096
rect 8201 17038 20963 17040
rect 8201 17035 8267 17038
rect 20897 17035 20963 17038
rect 19333 16962 19399 16965
rect 19885 16962 19951 16965
rect 20529 16962 20595 16965
rect 19333 16960 20595 16962
rect 19333 16904 19338 16960
rect 19394 16904 19890 16960
rect 19946 16904 20534 16960
rect 20590 16904 20595 16960
rect 19333 16902 20595 16904
rect 19333 16899 19399 16902
rect 19885 16899 19951 16902
rect 20529 16899 20595 16902
rect 3566 16896 3882 16897
rect 3566 16832 3572 16896
rect 3636 16832 3652 16896
rect 3716 16832 3732 16896
rect 3796 16832 3812 16896
rect 3876 16832 3882 16896
rect 3566 16831 3882 16832
rect 8566 16896 8882 16897
rect 8566 16832 8572 16896
rect 8636 16832 8652 16896
rect 8716 16832 8732 16896
rect 8796 16832 8812 16896
rect 8876 16832 8882 16896
rect 8566 16831 8882 16832
rect 13566 16896 13882 16897
rect 13566 16832 13572 16896
rect 13636 16832 13652 16896
rect 13716 16832 13732 16896
rect 13796 16832 13812 16896
rect 13876 16832 13882 16896
rect 13566 16831 13882 16832
rect 18566 16896 18882 16897
rect 18566 16832 18572 16896
rect 18636 16832 18652 16896
rect 18716 16832 18732 16896
rect 18796 16832 18812 16896
rect 18876 16832 18882 16896
rect 18566 16831 18882 16832
rect 23566 16896 23882 16897
rect 23566 16832 23572 16896
rect 23636 16832 23652 16896
rect 23716 16832 23732 16896
rect 23796 16832 23812 16896
rect 23876 16832 23882 16896
rect 23566 16831 23882 16832
rect 28566 16896 28882 16897
rect 28566 16832 28572 16896
rect 28636 16832 28652 16896
rect 28716 16832 28732 16896
rect 28796 16832 28812 16896
rect 28876 16832 28882 16896
rect 28566 16831 28882 16832
rect 33566 16896 33882 16897
rect 33566 16832 33572 16896
rect 33636 16832 33652 16896
rect 33716 16832 33732 16896
rect 33796 16832 33812 16896
rect 33876 16832 33882 16896
rect 33566 16831 33882 16832
rect 38566 16896 38882 16897
rect 38566 16832 38572 16896
rect 38636 16832 38652 16896
rect 38716 16832 38732 16896
rect 38796 16832 38812 16896
rect 38876 16832 38882 16896
rect 38566 16831 38882 16832
rect 43566 16896 43882 16897
rect 43566 16832 43572 16896
rect 43636 16832 43652 16896
rect 43716 16832 43732 16896
rect 43796 16832 43812 16896
rect 43876 16832 43882 16896
rect 43566 16831 43882 16832
rect 21725 16690 21791 16693
rect 27889 16690 27955 16693
rect 21725 16688 27955 16690
rect 21725 16632 21730 16688
rect 21786 16632 27894 16688
rect 27950 16632 27955 16688
rect 21725 16630 27955 16632
rect 21725 16627 21791 16630
rect 27889 16627 27955 16630
rect 18965 16554 19031 16557
rect 23749 16554 23815 16557
rect 18965 16552 23815 16554
rect 18965 16496 18970 16552
rect 19026 16496 23754 16552
rect 23810 16496 23815 16552
rect 18965 16494 23815 16496
rect 18965 16491 19031 16494
rect 23749 16491 23815 16494
rect 26877 16554 26943 16557
rect 33174 16554 33180 16556
rect 26877 16552 33180 16554
rect 26877 16496 26882 16552
rect 26938 16496 33180 16552
rect 26877 16494 33180 16496
rect 26877 16491 26943 16494
rect 33174 16492 33180 16494
rect 33244 16554 33250 16556
rect 33685 16554 33751 16557
rect 33244 16552 33751 16554
rect 33244 16496 33690 16552
rect 33746 16496 33751 16552
rect 33244 16494 33751 16496
rect 33244 16492 33250 16494
rect 33685 16491 33751 16494
rect 39113 16554 39179 16557
rect 40953 16554 41019 16557
rect 39113 16552 41019 16554
rect 39113 16496 39118 16552
rect 39174 16496 40958 16552
rect 41014 16496 41019 16552
rect 39113 16494 41019 16496
rect 39113 16491 39179 16494
rect 40953 16491 41019 16494
rect 6066 16352 6382 16353
rect 6066 16288 6072 16352
rect 6136 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6382 16352
rect 6066 16287 6382 16288
rect 11066 16352 11382 16353
rect 11066 16288 11072 16352
rect 11136 16288 11152 16352
rect 11216 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11382 16352
rect 11066 16287 11382 16288
rect 16066 16352 16382 16353
rect 16066 16288 16072 16352
rect 16136 16288 16152 16352
rect 16216 16288 16232 16352
rect 16296 16288 16312 16352
rect 16376 16288 16382 16352
rect 16066 16287 16382 16288
rect 21066 16352 21382 16353
rect 21066 16288 21072 16352
rect 21136 16288 21152 16352
rect 21216 16288 21232 16352
rect 21296 16288 21312 16352
rect 21376 16288 21382 16352
rect 21066 16287 21382 16288
rect 26066 16352 26382 16353
rect 26066 16288 26072 16352
rect 26136 16288 26152 16352
rect 26216 16288 26232 16352
rect 26296 16288 26312 16352
rect 26376 16288 26382 16352
rect 26066 16287 26382 16288
rect 31066 16352 31382 16353
rect 31066 16288 31072 16352
rect 31136 16288 31152 16352
rect 31216 16288 31232 16352
rect 31296 16288 31312 16352
rect 31376 16288 31382 16352
rect 31066 16287 31382 16288
rect 36066 16352 36382 16353
rect 36066 16288 36072 16352
rect 36136 16288 36152 16352
rect 36216 16288 36232 16352
rect 36296 16288 36312 16352
rect 36376 16288 36382 16352
rect 36066 16287 36382 16288
rect 41066 16352 41382 16353
rect 41066 16288 41072 16352
rect 41136 16288 41152 16352
rect 41216 16288 41232 16352
rect 41296 16288 41312 16352
rect 41376 16288 41382 16352
rect 41066 16287 41382 16288
rect 16205 16146 16271 16149
rect 18229 16146 18295 16149
rect 16205 16144 18295 16146
rect 16205 16088 16210 16144
rect 16266 16088 18234 16144
rect 18290 16088 18295 16144
rect 16205 16086 18295 16088
rect 16205 16083 16271 16086
rect 18229 16083 18295 16086
rect 22553 16010 22619 16013
rect 26509 16010 26575 16013
rect 26918 16010 26924 16012
rect 22553 16008 26924 16010
rect 22553 15952 22558 16008
rect 22614 15952 26514 16008
rect 26570 15952 26924 16008
rect 22553 15950 26924 15952
rect 22553 15947 22619 15950
rect 26509 15947 26575 15950
rect 26918 15948 26924 15950
rect 26988 15948 26994 16012
rect 29085 16010 29151 16013
rect 30230 16010 30236 16012
rect 29085 16008 30236 16010
rect 29085 15952 29090 16008
rect 29146 15952 30236 16008
rect 29085 15950 30236 15952
rect 29085 15947 29151 15950
rect 30230 15948 30236 15950
rect 30300 15948 30306 16012
rect 3566 15808 3882 15809
rect 3566 15744 3572 15808
rect 3636 15744 3652 15808
rect 3716 15744 3732 15808
rect 3796 15744 3812 15808
rect 3876 15744 3882 15808
rect 3566 15743 3882 15744
rect 8566 15808 8882 15809
rect 8566 15744 8572 15808
rect 8636 15744 8652 15808
rect 8716 15744 8732 15808
rect 8796 15744 8812 15808
rect 8876 15744 8882 15808
rect 8566 15743 8882 15744
rect 13566 15808 13882 15809
rect 13566 15744 13572 15808
rect 13636 15744 13652 15808
rect 13716 15744 13732 15808
rect 13796 15744 13812 15808
rect 13876 15744 13882 15808
rect 13566 15743 13882 15744
rect 18566 15808 18882 15809
rect 18566 15744 18572 15808
rect 18636 15744 18652 15808
rect 18716 15744 18732 15808
rect 18796 15744 18812 15808
rect 18876 15744 18882 15808
rect 18566 15743 18882 15744
rect 23566 15808 23882 15809
rect 23566 15744 23572 15808
rect 23636 15744 23652 15808
rect 23716 15744 23732 15808
rect 23796 15744 23812 15808
rect 23876 15744 23882 15808
rect 23566 15743 23882 15744
rect 28566 15808 28882 15809
rect 28566 15744 28572 15808
rect 28636 15744 28652 15808
rect 28716 15744 28732 15808
rect 28796 15744 28812 15808
rect 28876 15744 28882 15808
rect 28566 15743 28882 15744
rect 33566 15808 33882 15809
rect 33566 15744 33572 15808
rect 33636 15744 33652 15808
rect 33716 15744 33732 15808
rect 33796 15744 33812 15808
rect 33876 15744 33882 15808
rect 33566 15743 33882 15744
rect 38566 15808 38882 15809
rect 38566 15744 38572 15808
rect 38636 15744 38652 15808
rect 38716 15744 38732 15808
rect 38796 15744 38812 15808
rect 38876 15744 38882 15808
rect 38566 15743 38882 15744
rect 43566 15808 43882 15809
rect 43566 15744 43572 15808
rect 43636 15744 43652 15808
rect 43716 15744 43732 15808
rect 43796 15744 43812 15808
rect 43876 15744 43882 15808
rect 43566 15743 43882 15744
rect 23933 15602 23999 15605
rect 27337 15602 27403 15605
rect 23933 15600 27403 15602
rect 23933 15544 23938 15600
rect 23994 15544 27342 15600
rect 27398 15544 27403 15600
rect 23933 15542 27403 15544
rect 23933 15539 23999 15542
rect 27337 15539 27403 15542
rect 14733 15466 14799 15469
rect 15193 15466 15259 15469
rect 37273 15466 37339 15469
rect 37825 15466 37891 15469
rect 14733 15464 37891 15466
rect 14733 15408 14738 15464
rect 14794 15408 15198 15464
rect 15254 15408 37278 15464
rect 37334 15408 37830 15464
rect 37886 15408 37891 15464
rect 14733 15406 37891 15408
rect 14733 15403 14799 15406
rect 15193 15403 15259 15406
rect 37273 15403 37339 15406
rect 37825 15403 37891 15406
rect 27889 15330 27955 15333
rect 29085 15330 29151 15333
rect 27889 15328 29151 15330
rect 27889 15272 27894 15328
rect 27950 15272 29090 15328
rect 29146 15272 29151 15328
rect 27889 15270 29151 15272
rect 27889 15267 27955 15270
rect 29085 15267 29151 15270
rect 6066 15264 6382 15265
rect 6066 15200 6072 15264
rect 6136 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6382 15264
rect 6066 15199 6382 15200
rect 11066 15264 11382 15265
rect 11066 15200 11072 15264
rect 11136 15200 11152 15264
rect 11216 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11382 15264
rect 11066 15199 11382 15200
rect 16066 15264 16382 15265
rect 16066 15200 16072 15264
rect 16136 15200 16152 15264
rect 16216 15200 16232 15264
rect 16296 15200 16312 15264
rect 16376 15200 16382 15264
rect 16066 15199 16382 15200
rect 21066 15264 21382 15265
rect 21066 15200 21072 15264
rect 21136 15200 21152 15264
rect 21216 15200 21232 15264
rect 21296 15200 21312 15264
rect 21376 15200 21382 15264
rect 21066 15199 21382 15200
rect 26066 15264 26382 15265
rect 26066 15200 26072 15264
rect 26136 15200 26152 15264
rect 26216 15200 26232 15264
rect 26296 15200 26312 15264
rect 26376 15200 26382 15264
rect 26066 15199 26382 15200
rect 31066 15264 31382 15265
rect 31066 15200 31072 15264
rect 31136 15200 31152 15264
rect 31216 15200 31232 15264
rect 31296 15200 31312 15264
rect 31376 15200 31382 15264
rect 31066 15199 31382 15200
rect 36066 15264 36382 15265
rect 36066 15200 36072 15264
rect 36136 15200 36152 15264
rect 36216 15200 36232 15264
rect 36296 15200 36312 15264
rect 36376 15200 36382 15264
rect 36066 15199 36382 15200
rect 41066 15264 41382 15265
rect 41066 15200 41072 15264
rect 41136 15200 41152 15264
rect 41216 15200 41232 15264
rect 41296 15200 41312 15264
rect 41376 15200 41382 15264
rect 41066 15199 41382 15200
rect 16297 15058 16363 15061
rect 24209 15058 24275 15061
rect 31937 15058 32003 15061
rect 16297 15056 22110 15058
rect 16297 15000 16302 15056
rect 16358 15000 22110 15056
rect 16297 14998 22110 15000
rect 16297 14995 16363 14998
rect 22050 14922 22110 14998
rect 24209 15056 32003 15058
rect 24209 15000 24214 15056
rect 24270 15000 31942 15056
rect 31998 15000 32003 15056
rect 24209 14998 32003 15000
rect 24209 14995 24275 14998
rect 31937 14995 32003 14998
rect 29361 14924 29427 14925
rect 22686 14922 22692 14924
rect 22050 14862 22692 14922
rect 22686 14860 22692 14862
rect 22756 14922 22762 14924
rect 29310 14922 29316 14924
rect 22756 14862 29010 14922
rect 29270 14862 29316 14922
rect 29380 14920 29427 14924
rect 31753 14922 31819 14925
rect 29422 14864 29427 14920
rect 22756 14860 22762 14862
rect -300 14786 160 14816
rect 933 14786 999 14789
rect -300 14784 999 14786
rect -300 14728 938 14784
rect 994 14728 999 14784
rect -300 14726 999 14728
rect 28950 14786 29010 14862
rect 29310 14860 29316 14862
rect 29380 14860 29427 14864
rect 29361 14859 29427 14860
rect 31710 14920 31819 14922
rect 31710 14864 31758 14920
rect 31814 14864 31819 14920
rect 31710 14859 31819 14864
rect 32213 14922 32279 14925
rect 36813 14922 36879 14925
rect 32213 14920 36879 14922
rect 32213 14864 32218 14920
rect 32274 14864 36818 14920
rect 36874 14864 36879 14920
rect 32213 14862 36879 14864
rect 32213 14859 32279 14862
rect 36813 14859 36879 14862
rect 31710 14786 31770 14859
rect 28950 14726 31770 14786
rect 45185 14786 45251 14789
rect 45840 14786 46300 14816
rect 45185 14784 46300 14786
rect 45185 14728 45190 14784
rect 45246 14728 46300 14784
rect 45185 14726 46300 14728
rect -300 14696 160 14726
rect 933 14723 999 14726
rect 45185 14723 45251 14726
rect 3566 14720 3882 14721
rect 3566 14656 3572 14720
rect 3636 14656 3652 14720
rect 3716 14656 3732 14720
rect 3796 14656 3812 14720
rect 3876 14656 3882 14720
rect 3566 14655 3882 14656
rect 8566 14720 8882 14721
rect 8566 14656 8572 14720
rect 8636 14656 8652 14720
rect 8716 14656 8732 14720
rect 8796 14656 8812 14720
rect 8876 14656 8882 14720
rect 8566 14655 8882 14656
rect 13566 14720 13882 14721
rect 13566 14656 13572 14720
rect 13636 14656 13652 14720
rect 13716 14656 13732 14720
rect 13796 14656 13812 14720
rect 13876 14656 13882 14720
rect 13566 14655 13882 14656
rect 18566 14720 18882 14721
rect 18566 14656 18572 14720
rect 18636 14656 18652 14720
rect 18716 14656 18732 14720
rect 18796 14656 18812 14720
rect 18876 14656 18882 14720
rect 18566 14655 18882 14656
rect 23566 14720 23882 14721
rect 23566 14656 23572 14720
rect 23636 14656 23652 14720
rect 23716 14656 23732 14720
rect 23796 14656 23812 14720
rect 23876 14656 23882 14720
rect 23566 14655 23882 14656
rect 28566 14720 28882 14721
rect 28566 14656 28572 14720
rect 28636 14656 28652 14720
rect 28716 14656 28732 14720
rect 28796 14656 28812 14720
rect 28876 14656 28882 14720
rect 28566 14655 28882 14656
rect 33566 14720 33882 14721
rect 33566 14656 33572 14720
rect 33636 14656 33652 14720
rect 33716 14656 33732 14720
rect 33796 14656 33812 14720
rect 33876 14656 33882 14720
rect 33566 14655 33882 14656
rect 38566 14720 38882 14721
rect 38566 14656 38572 14720
rect 38636 14656 38652 14720
rect 38716 14656 38732 14720
rect 38796 14656 38812 14720
rect 38876 14656 38882 14720
rect 38566 14655 38882 14656
rect 43566 14720 43882 14721
rect 43566 14656 43572 14720
rect 43636 14656 43652 14720
rect 43716 14656 43732 14720
rect 43796 14656 43812 14720
rect 43876 14656 43882 14720
rect 45840 14696 46300 14726
rect 43566 14655 43882 14656
rect 24577 14650 24643 14653
rect 26233 14650 26299 14653
rect 24577 14648 26299 14650
rect 24577 14592 24582 14648
rect 24638 14592 26238 14648
rect 26294 14592 26299 14648
rect 24577 14590 26299 14592
rect 24577 14587 24643 14590
rect 26233 14587 26299 14590
rect 18965 14516 19031 14517
rect 18965 14514 19012 14516
rect 18920 14512 19012 14514
rect 18920 14456 18970 14512
rect 18920 14454 19012 14456
rect 18965 14452 19012 14454
rect 19076 14452 19082 14516
rect 23381 14514 23447 14517
rect 27429 14514 27495 14517
rect 23381 14512 27495 14514
rect 23381 14456 23386 14512
rect 23442 14456 27434 14512
rect 27490 14456 27495 14512
rect 23381 14454 27495 14456
rect 18965 14451 19031 14452
rect 23381 14451 23447 14454
rect 27429 14451 27495 14454
rect 27061 14378 27127 14381
rect 28073 14378 28139 14381
rect 29729 14378 29795 14381
rect 27061 14376 29795 14378
rect 27061 14320 27066 14376
rect 27122 14320 28078 14376
rect 28134 14320 29734 14376
rect 29790 14320 29795 14376
rect 27061 14318 29795 14320
rect 27061 14315 27127 14318
rect 28073 14315 28139 14318
rect 29729 14315 29795 14318
rect 30782 14316 30788 14380
rect 30852 14378 30858 14380
rect 31109 14378 31175 14381
rect 30852 14376 31175 14378
rect 30852 14320 31114 14376
rect 31170 14320 31175 14376
rect 30852 14318 31175 14320
rect 30852 14316 30858 14318
rect 31109 14315 31175 14318
rect 6066 14176 6382 14177
rect 6066 14112 6072 14176
rect 6136 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6382 14176
rect 6066 14111 6382 14112
rect 11066 14176 11382 14177
rect 11066 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11382 14176
rect 11066 14111 11382 14112
rect 16066 14176 16382 14177
rect 16066 14112 16072 14176
rect 16136 14112 16152 14176
rect 16216 14112 16232 14176
rect 16296 14112 16312 14176
rect 16376 14112 16382 14176
rect 16066 14111 16382 14112
rect 21066 14176 21382 14177
rect 21066 14112 21072 14176
rect 21136 14112 21152 14176
rect 21216 14112 21232 14176
rect 21296 14112 21312 14176
rect 21376 14112 21382 14176
rect 21066 14111 21382 14112
rect 26066 14176 26382 14177
rect 26066 14112 26072 14176
rect 26136 14112 26152 14176
rect 26216 14112 26232 14176
rect 26296 14112 26312 14176
rect 26376 14112 26382 14176
rect 26066 14111 26382 14112
rect 31066 14176 31382 14177
rect 31066 14112 31072 14176
rect 31136 14112 31152 14176
rect 31216 14112 31232 14176
rect 31296 14112 31312 14176
rect 31376 14112 31382 14176
rect 31066 14111 31382 14112
rect 36066 14176 36382 14177
rect 36066 14112 36072 14176
rect 36136 14112 36152 14176
rect 36216 14112 36232 14176
rect 36296 14112 36312 14176
rect 36376 14112 36382 14176
rect 36066 14111 36382 14112
rect 41066 14176 41382 14177
rect 41066 14112 41072 14176
rect 41136 14112 41152 14176
rect 41216 14112 41232 14176
rect 41296 14112 41312 14176
rect 41376 14112 41382 14176
rect 41066 14111 41382 14112
rect 26918 14044 26924 14108
rect 26988 14106 26994 14108
rect 28349 14106 28415 14109
rect 26988 14104 28415 14106
rect 26988 14048 28354 14104
rect 28410 14048 28415 14104
rect 26988 14046 28415 14048
rect 26988 14044 26994 14046
rect 28349 14043 28415 14046
rect 21541 13970 21607 13973
rect 33225 13970 33291 13973
rect 21541 13968 33291 13970
rect 21541 13912 21546 13968
rect 21602 13912 33230 13968
rect 33286 13912 33291 13968
rect 21541 13910 33291 13912
rect 21541 13907 21607 13910
rect 33225 13907 33291 13910
rect 13629 13834 13695 13837
rect 14273 13834 14339 13837
rect 13629 13832 14339 13834
rect 13629 13776 13634 13832
rect 13690 13776 14278 13832
rect 14334 13776 14339 13832
rect 13629 13774 14339 13776
rect 13629 13771 13695 13774
rect 14273 13771 14339 13774
rect 29085 13834 29151 13837
rect 32949 13834 33015 13837
rect 29085 13832 33015 13834
rect 29085 13776 29090 13832
rect 29146 13776 32954 13832
rect 33010 13776 33015 13832
rect 29085 13774 33015 13776
rect 29085 13771 29151 13774
rect 32949 13771 33015 13774
rect 3566 13632 3882 13633
rect 3566 13568 3572 13632
rect 3636 13568 3652 13632
rect 3716 13568 3732 13632
rect 3796 13568 3812 13632
rect 3876 13568 3882 13632
rect 3566 13567 3882 13568
rect 8566 13632 8882 13633
rect 8566 13568 8572 13632
rect 8636 13568 8652 13632
rect 8716 13568 8732 13632
rect 8796 13568 8812 13632
rect 8876 13568 8882 13632
rect 8566 13567 8882 13568
rect 13566 13632 13882 13633
rect 13566 13568 13572 13632
rect 13636 13568 13652 13632
rect 13716 13568 13732 13632
rect 13796 13568 13812 13632
rect 13876 13568 13882 13632
rect 13566 13567 13882 13568
rect 18566 13632 18882 13633
rect 18566 13568 18572 13632
rect 18636 13568 18652 13632
rect 18716 13568 18732 13632
rect 18796 13568 18812 13632
rect 18876 13568 18882 13632
rect 18566 13567 18882 13568
rect 23566 13632 23882 13633
rect 23566 13568 23572 13632
rect 23636 13568 23652 13632
rect 23716 13568 23732 13632
rect 23796 13568 23812 13632
rect 23876 13568 23882 13632
rect 23566 13567 23882 13568
rect 28566 13632 28882 13633
rect 28566 13568 28572 13632
rect 28636 13568 28652 13632
rect 28716 13568 28732 13632
rect 28796 13568 28812 13632
rect 28876 13568 28882 13632
rect 28566 13567 28882 13568
rect 33566 13632 33882 13633
rect 33566 13568 33572 13632
rect 33636 13568 33652 13632
rect 33716 13568 33732 13632
rect 33796 13568 33812 13632
rect 33876 13568 33882 13632
rect 33566 13567 33882 13568
rect 38566 13632 38882 13633
rect 38566 13568 38572 13632
rect 38636 13568 38652 13632
rect 38716 13568 38732 13632
rect 38796 13568 38812 13632
rect 38876 13568 38882 13632
rect 38566 13567 38882 13568
rect 43566 13632 43882 13633
rect 43566 13568 43572 13632
rect 43636 13568 43652 13632
rect 43716 13568 43732 13632
rect 43796 13568 43812 13632
rect 43876 13568 43882 13632
rect 43566 13567 43882 13568
rect 27153 13562 27219 13565
rect 23982 13560 27219 13562
rect 23982 13504 27158 13560
rect 27214 13504 27219 13560
rect 23982 13502 27219 13504
rect 20161 13426 20227 13429
rect 20805 13426 20871 13429
rect 20161 13424 20871 13426
rect 20161 13368 20166 13424
rect 20222 13368 20810 13424
rect 20866 13368 20871 13424
rect 20161 13366 20871 13368
rect 20161 13363 20227 13366
rect 20805 13363 20871 13366
rect 21909 13426 21975 13429
rect 23982 13426 24042 13502
rect 27153 13499 27219 13502
rect 21909 13424 24042 13426
rect 21909 13368 21914 13424
rect 21970 13368 24042 13424
rect 21909 13366 24042 13368
rect 25497 13426 25563 13429
rect 29269 13426 29335 13429
rect 25497 13424 29335 13426
rect 25497 13368 25502 13424
rect 25558 13368 29274 13424
rect 29330 13368 29335 13424
rect 25497 13366 29335 13368
rect 21909 13363 21975 13366
rect 25497 13363 25563 13366
rect 29269 13363 29335 13366
rect 16021 13290 16087 13293
rect 19793 13290 19859 13293
rect 16021 13288 19859 13290
rect 16021 13232 16026 13288
rect 16082 13232 19798 13288
rect 19854 13232 19859 13288
rect 16021 13230 19859 13232
rect 16021 13227 16087 13230
rect 19793 13227 19859 13230
rect 23841 13290 23907 13293
rect 25497 13290 25563 13293
rect 23841 13288 25563 13290
rect 23841 13232 23846 13288
rect 23902 13232 25502 13288
rect 25558 13232 25563 13288
rect 23841 13230 25563 13232
rect 23841 13227 23907 13230
rect 25497 13227 25563 13230
rect 30097 13290 30163 13293
rect 34881 13290 34947 13293
rect 30097 13288 34947 13290
rect 30097 13232 30102 13288
rect 30158 13232 34886 13288
rect 34942 13232 34947 13288
rect 30097 13230 34947 13232
rect 30097 13227 30163 13230
rect 34881 13227 34947 13230
rect 24577 13154 24643 13157
rect 25313 13154 25379 13157
rect 24577 13152 25379 13154
rect 24577 13096 24582 13152
rect 24638 13096 25318 13152
rect 25374 13096 25379 13152
rect 24577 13094 25379 13096
rect 24577 13091 24643 13094
rect 25313 13091 25379 13094
rect 6066 13088 6382 13089
rect 6066 13024 6072 13088
rect 6136 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6382 13088
rect 6066 13023 6382 13024
rect 11066 13088 11382 13089
rect 11066 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11382 13088
rect 11066 13023 11382 13024
rect 16066 13088 16382 13089
rect 16066 13024 16072 13088
rect 16136 13024 16152 13088
rect 16216 13024 16232 13088
rect 16296 13024 16312 13088
rect 16376 13024 16382 13088
rect 16066 13023 16382 13024
rect 21066 13088 21382 13089
rect 21066 13024 21072 13088
rect 21136 13024 21152 13088
rect 21216 13024 21232 13088
rect 21296 13024 21312 13088
rect 21376 13024 21382 13088
rect 21066 13023 21382 13024
rect 26066 13088 26382 13089
rect 26066 13024 26072 13088
rect 26136 13024 26152 13088
rect 26216 13024 26232 13088
rect 26296 13024 26312 13088
rect 26376 13024 26382 13088
rect 26066 13023 26382 13024
rect 31066 13088 31382 13089
rect 31066 13024 31072 13088
rect 31136 13024 31152 13088
rect 31216 13024 31232 13088
rect 31296 13024 31312 13088
rect 31376 13024 31382 13088
rect 31066 13023 31382 13024
rect 36066 13088 36382 13089
rect 36066 13024 36072 13088
rect 36136 13024 36152 13088
rect 36216 13024 36232 13088
rect 36296 13024 36312 13088
rect 36376 13024 36382 13088
rect 36066 13023 36382 13024
rect 41066 13088 41382 13089
rect 41066 13024 41072 13088
rect 41136 13024 41152 13088
rect 41216 13024 41232 13088
rect 41296 13024 41312 13088
rect 41376 13024 41382 13088
rect 41066 13023 41382 13024
rect 22277 13018 22343 13021
rect 23289 13018 23355 13021
rect 27613 13018 27679 13021
rect 28257 13018 28323 13021
rect 22277 13016 25698 13018
rect 22277 12960 22282 13016
rect 22338 12960 23294 13016
rect 23350 12960 25698 13016
rect 22277 12958 25698 12960
rect 22277 12955 22343 12958
rect 23289 12955 23355 12958
rect 9397 12882 9463 12885
rect 12709 12882 12775 12885
rect 9397 12880 12775 12882
rect 9397 12824 9402 12880
rect 9458 12824 12714 12880
rect 12770 12824 12775 12880
rect 9397 12822 12775 12824
rect 9397 12819 9463 12822
rect 12709 12819 12775 12822
rect 20161 12882 20227 12885
rect 23841 12882 23907 12885
rect 25405 12882 25471 12885
rect 20161 12880 22110 12882
rect 20161 12824 20166 12880
rect 20222 12824 22110 12880
rect 20161 12822 22110 12824
rect 20161 12819 20227 12822
rect 22050 12746 22110 12822
rect 23841 12880 25471 12882
rect 23841 12824 23846 12880
rect 23902 12824 25410 12880
rect 25466 12824 25471 12880
rect 23841 12822 25471 12824
rect 25638 12882 25698 12958
rect 27613 13016 28323 13018
rect 27613 12960 27618 13016
rect 27674 12960 28262 13016
rect 28318 12960 28323 13016
rect 27613 12958 28323 12960
rect 27613 12955 27679 12958
rect 28257 12955 28323 12958
rect 26049 12882 26115 12885
rect 28349 12882 28415 12885
rect 25638 12880 28415 12882
rect 25638 12824 26054 12880
rect 26110 12824 28354 12880
rect 28410 12824 28415 12880
rect 25638 12822 28415 12824
rect 23841 12819 23907 12822
rect 25405 12819 25471 12822
rect 26049 12819 26115 12822
rect 28349 12819 28415 12822
rect 29913 12882 29979 12885
rect 33225 12882 33291 12885
rect 29913 12880 33291 12882
rect 29913 12824 29918 12880
rect 29974 12824 33230 12880
rect 33286 12824 33291 12880
rect 29913 12822 33291 12824
rect 29913 12819 29979 12822
rect 33225 12819 33291 12822
rect 25221 12746 25287 12749
rect 22050 12744 25287 12746
rect 22050 12688 25226 12744
rect 25282 12688 25287 12744
rect 22050 12686 25287 12688
rect 25221 12683 25287 12686
rect 26969 12746 27035 12749
rect 30414 12746 30420 12748
rect 26969 12744 30420 12746
rect 26969 12688 26974 12744
rect 27030 12688 30420 12744
rect 26969 12686 30420 12688
rect 26969 12683 27035 12686
rect 30414 12684 30420 12686
rect 30484 12746 30490 12748
rect 31937 12746 32003 12749
rect 33133 12746 33199 12749
rect 30484 12744 33199 12746
rect 30484 12688 31942 12744
rect 31998 12688 33138 12744
rect 33194 12688 33199 12744
rect 30484 12686 33199 12688
rect 30484 12684 30490 12686
rect 31937 12683 32003 12686
rect 33133 12683 33199 12686
rect 3566 12544 3882 12545
rect 3566 12480 3572 12544
rect 3636 12480 3652 12544
rect 3716 12480 3732 12544
rect 3796 12480 3812 12544
rect 3876 12480 3882 12544
rect 3566 12479 3882 12480
rect 8566 12544 8882 12545
rect 8566 12480 8572 12544
rect 8636 12480 8652 12544
rect 8716 12480 8732 12544
rect 8796 12480 8812 12544
rect 8876 12480 8882 12544
rect 8566 12479 8882 12480
rect 13566 12544 13882 12545
rect 13566 12480 13572 12544
rect 13636 12480 13652 12544
rect 13716 12480 13732 12544
rect 13796 12480 13812 12544
rect 13876 12480 13882 12544
rect 13566 12479 13882 12480
rect 18566 12544 18882 12545
rect 18566 12480 18572 12544
rect 18636 12480 18652 12544
rect 18716 12480 18732 12544
rect 18796 12480 18812 12544
rect 18876 12480 18882 12544
rect 18566 12479 18882 12480
rect 23566 12544 23882 12545
rect 23566 12480 23572 12544
rect 23636 12480 23652 12544
rect 23716 12480 23732 12544
rect 23796 12480 23812 12544
rect 23876 12480 23882 12544
rect 23566 12479 23882 12480
rect 28566 12544 28882 12545
rect 28566 12480 28572 12544
rect 28636 12480 28652 12544
rect 28716 12480 28732 12544
rect 28796 12480 28812 12544
rect 28876 12480 28882 12544
rect 28566 12479 28882 12480
rect 33566 12544 33882 12545
rect 33566 12480 33572 12544
rect 33636 12480 33652 12544
rect 33716 12480 33732 12544
rect 33796 12480 33812 12544
rect 33876 12480 33882 12544
rect 33566 12479 33882 12480
rect 38566 12544 38882 12545
rect 38566 12480 38572 12544
rect 38636 12480 38652 12544
rect 38716 12480 38732 12544
rect 38796 12480 38812 12544
rect 38876 12480 38882 12544
rect 38566 12479 38882 12480
rect 43566 12544 43882 12545
rect 43566 12480 43572 12544
rect 43636 12480 43652 12544
rect 43716 12480 43732 12544
rect 43796 12480 43812 12544
rect 43876 12480 43882 12544
rect 43566 12479 43882 12480
rect 20161 12474 20227 12477
rect 20118 12472 20227 12474
rect 20118 12416 20166 12472
rect 20222 12416 20227 12472
rect 20118 12411 20227 12416
rect 24853 12472 24919 12477
rect 24853 12416 24858 12472
rect 24914 12416 24919 12472
rect 24853 12411 24919 12416
rect 17401 12338 17467 12341
rect 20118 12338 20178 12411
rect 17401 12336 20178 12338
rect 17401 12280 17406 12336
rect 17462 12280 20178 12336
rect 17401 12278 20178 12280
rect 20437 12338 20503 12341
rect 24856 12338 24916 12411
rect 20437 12336 24916 12338
rect 20437 12280 20442 12336
rect 20498 12280 24916 12336
rect 20437 12278 24916 12280
rect 26417 12338 26483 12341
rect 30782 12338 30788 12340
rect 26417 12336 30788 12338
rect 26417 12280 26422 12336
rect 26478 12280 30788 12336
rect 26417 12278 30788 12280
rect 17401 12275 17467 12278
rect 20437 12275 20503 12278
rect 26417 12275 26483 12278
rect 30782 12276 30788 12278
rect 30852 12276 30858 12340
rect 33317 12338 33383 12341
rect 37457 12338 37523 12341
rect 33317 12336 37523 12338
rect 33317 12280 33322 12336
rect 33378 12280 37462 12336
rect 37518 12280 37523 12336
rect 33317 12278 37523 12280
rect 33317 12275 33383 12278
rect 37457 12275 37523 12278
rect 17677 12202 17743 12205
rect 19149 12202 19215 12205
rect 17677 12200 19215 12202
rect 17677 12144 17682 12200
rect 17738 12144 19154 12200
rect 19210 12144 19215 12200
rect 17677 12142 19215 12144
rect 17677 12139 17743 12142
rect 19149 12139 19215 12142
rect 24853 12202 24919 12205
rect 29177 12202 29243 12205
rect 34237 12202 34303 12205
rect 36629 12202 36695 12205
rect 24853 12200 36695 12202
rect 24853 12144 24858 12200
rect 24914 12144 29182 12200
rect 29238 12144 34242 12200
rect 34298 12144 36634 12200
rect 36690 12144 36695 12200
rect 24853 12142 36695 12144
rect 24853 12139 24919 12142
rect 29177 12139 29243 12142
rect 34237 12139 34303 12142
rect 36629 12139 36695 12142
rect 18689 12066 18755 12069
rect 20621 12066 20687 12069
rect 18689 12064 20687 12066
rect 18689 12008 18694 12064
rect 18750 12008 20626 12064
rect 20682 12008 20687 12064
rect 18689 12006 20687 12008
rect 18689 12003 18755 12006
rect 20621 12003 20687 12006
rect 6066 12000 6382 12001
rect 6066 11936 6072 12000
rect 6136 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6382 12000
rect 6066 11935 6382 11936
rect 11066 12000 11382 12001
rect 11066 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11382 12000
rect 11066 11935 11382 11936
rect 16066 12000 16382 12001
rect 16066 11936 16072 12000
rect 16136 11936 16152 12000
rect 16216 11936 16232 12000
rect 16296 11936 16312 12000
rect 16376 11936 16382 12000
rect 16066 11935 16382 11936
rect 21066 12000 21382 12001
rect 21066 11936 21072 12000
rect 21136 11936 21152 12000
rect 21216 11936 21232 12000
rect 21296 11936 21312 12000
rect 21376 11936 21382 12000
rect 21066 11935 21382 11936
rect 26066 12000 26382 12001
rect 26066 11936 26072 12000
rect 26136 11936 26152 12000
rect 26216 11936 26232 12000
rect 26296 11936 26312 12000
rect 26376 11936 26382 12000
rect 26066 11935 26382 11936
rect 31066 12000 31382 12001
rect 31066 11936 31072 12000
rect 31136 11936 31152 12000
rect 31216 11936 31232 12000
rect 31296 11936 31312 12000
rect 31376 11936 31382 12000
rect 31066 11935 31382 11936
rect 36066 12000 36382 12001
rect 36066 11936 36072 12000
rect 36136 11936 36152 12000
rect 36216 11936 36232 12000
rect 36296 11936 36312 12000
rect 36376 11936 36382 12000
rect 36066 11935 36382 11936
rect 41066 12000 41382 12001
rect 41066 11936 41072 12000
rect 41136 11936 41152 12000
rect 41216 11936 41232 12000
rect 41296 11936 41312 12000
rect 41376 11936 41382 12000
rect 41066 11935 41382 11936
rect 4981 11930 5047 11933
rect 5533 11930 5599 11933
rect 4981 11928 5599 11930
rect 4981 11872 4986 11928
rect 5042 11872 5538 11928
rect 5594 11872 5599 11928
rect 4981 11870 5599 11872
rect 4981 11867 5047 11870
rect 5533 11867 5599 11870
rect 5165 11794 5231 11797
rect 5717 11794 5783 11797
rect 5165 11792 5783 11794
rect 5165 11736 5170 11792
rect 5226 11736 5722 11792
rect 5778 11736 5783 11792
rect 5165 11734 5783 11736
rect 5165 11731 5231 11734
rect 5717 11731 5783 11734
rect 19425 11794 19491 11797
rect 25313 11794 25379 11797
rect 33501 11794 33567 11797
rect 19425 11792 33567 11794
rect 19425 11736 19430 11792
rect 19486 11736 25318 11792
rect 25374 11736 33506 11792
rect 33562 11736 33567 11792
rect 19425 11734 33567 11736
rect 19425 11731 19491 11734
rect 25313 11731 25379 11734
rect 33501 11731 33567 11734
rect 19977 11658 20043 11661
rect 34697 11658 34763 11661
rect 19977 11656 34763 11658
rect 19977 11600 19982 11656
rect 20038 11600 34702 11656
rect 34758 11600 34763 11656
rect 19977 11598 34763 11600
rect 19977 11595 20043 11598
rect 34697 11595 34763 11598
rect 29821 11522 29887 11525
rect 32857 11522 32923 11525
rect 29821 11520 32923 11522
rect 29821 11464 29826 11520
rect 29882 11464 32862 11520
rect 32918 11464 32923 11520
rect 29821 11462 32923 11464
rect 29821 11459 29887 11462
rect 32857 11459 32923 11462
rect 3566 11456 3882 11457
rect 3566 11392 3572 11456
rect 3636 11392 3652 11456
rect 3716 11392 3732 11456
rect 3796 11392 3812 11456
rect 3876 11392 3882 11456
rect 3566 11391 3882 11392
rect 8566 11456 8882 11457
rect 8566 11392 8572 11456
rect 8636 11392 8652 11456
rect 8716 11392 8732 11456
rect 8796 11392 8812 11456
rect 8876 11392 8882 11456
rect 8566 11391 8882 11392
rect 13566 11456 13882 11457
rect 13566 11392 13572 11456
rect 13636 11392 13652 11456
rect 13716 11392 13732 11456
rect 13796 11392 13812 11456
rect 13876 11392 13882 11456
rect 13566 11391 13882 11392
rect 18566 11456 18882 11457
rect 18566 11392 18572 11456
rect 18636 11392 18652 11456
rect 18716 11392 18732 11456
rect 18796 11392 18812 11456
rect 18876 11392 18882 11456
rect 18566 11391 18882 11392
rect 23566 11456 23882 11457
rect 23566 11392 23572 11456
rect 23636 11392 23652 11456
rect 23716 11392 23732 11456
rect 23796 11392 23812 11456
rect 23876 11392 23882 11456
rect 23566 11391 23882 11392
rect 28566 11456 28882 11457
rect 28566 11392 28572 11456
rect 28636 11392 28652 11456
rect 28716 11392 28732 11456
rect 28796 11392 28812 11456
rect 28876 11392 28882 11456
rect 28566 11391 28882 11392
rect 33566 11456 33882 11457
rect 33566 11392 33572 11456
rect 33636 11392 33652 11456
rect 33716 11392 33732 11456
rect 33796 11392 33812 11456
rect 33876 11392 33882 11456
rect 33566 11391 33882 11392
rect 38566 11456 38882 11457
rect 38566 11392 38572 11456
rect 38636 11392 38652 11456
rect 38716 11392 38732 11456
rect 38796 11392 38812 11456
rect 38876 11392 38882 11456
rect 38566 11391 38882 11392
rect 43566 11456 43882 11457
rect 43566 11392 43572 11456
rect 43636 11392 43652 11456
rect 43716 11392 43732 11456
rect 43796 11392 43812 11456
rect 43876 11392 43882 11456
rect 43566 11391 43882 11392
rect 29453 11386 29519 11389
rect 31753 11386 31819 11389
rect 29453 11384 31819 11386
rect 29453 11328 29458 11384
rect 29514 11328 31758 11384
rect 31814 11328 31819 11384
rect 29453 11326 31819 11328
rect 29453 11323 29519 11326
rect 31753 11323 31819 11326
rect 19057 11252 19123 11253
rect 19006 11250 19012 11252
rect 18966 11190 19012 11250
rect 19076 11248 19123 11252
rect 19118 11192 19123 11248
rect 19006 11188 19012 11190
rect 19076 11188 19123 11192
rect 19057 11187 19123 11188
rect 26877 11250 26943 11253
rect 44817 11250 44883 11253
rect 26877 11248 44883 11250
rect 26877 11192 26882 11248
rect 26938 11192 44822 11248
rect 44878 11192 44883 11248
rect 26877 11190 44883 11192
rect 26877 11187 26943 11190
rect 44817 11187 44883 11190
rect 30833 11116 30899 11117
rect 30782 11052 30788 11116
rect 30852 11114 30899 11116
rect 30852 11112 30944 11114
rect 30894 11056 30944 11112
rect 30852 11054 30944 11056
rect 30852 11052 30899 11054
rect 30833 11051 30899 11052
rect 13721 10978 13787 10981
rect 15101 10978 15167 10981
rect 29361 10980 29427 10981
rect 13721 10976 15167 10978
rect 13721 10920 13726 10976
rect 13782 10920 15106 10976
rect 15162 10920 15167 10976
rect 13721 10918 15167 10920
rect 13721 10915 13787 10918
rect 15101 10915 15167 10918
rect 29310 10916 29316 10980
rect 29380 10978 29427 10980
rect 32489 10978 32555 10981
rect 33961 10978 34027 10981
rect 29380 10976 29472 10978
rect 29422 10920 29472 10976
rect 29380 10918 29472 10920
rect 32489 10976 34027 10978
rect 32489 10920 32494 10976
rect 32550 10920 33966 10976
rect 34022 10920 34027 10976
rect 32489 10918 34027 10920
rect 29380 10916 29427 10918
rect 29361 10915 29427 10916
rect 32489 10915 32555 10918
rect 33961 10915 34027 10918
rect 6066 10912 6382 10913
rect 6066 10848 6072 10912
rect 6136 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6382 10912
rect 6066 10847 6382 10848
rect 11066 10912 11382 10913
rect 11066 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11382 10912
rect 11066 10847 11382 10848
rect 16066 10912 16382 10913
rect 16066 10848 16072 10912
rect 16136 10848 16152 10912
rect 16216 10848 16232 10912
rect 16296 10848 16312 10912
rect 16376 10848 16382 10912
rect 16066 10847 16382 10848
rect 21066 10912 21382 10913
rect 21066 10848 21072 10912
rect 21136 10848 21152 10912
rect 21216 10848 21232 10912
rect 21296 10848 21312 10912
rect 21376 10848 21382 10912
rect 21066 10847 21382 10848
rect 26066 10912 26382 10913
rect 26066 10848 26072 10912
rect 26136 10848 26152 10912
rect 26216 10848 26232 10912
rect 26296 10848 26312 10912
rect 26376 10848 26382 10912
rect 26066 10847 26382 10848
rect 31066 10912 31382 10913
rect 31066 10848 31072 10912
rect 31136 10848 31152 10912
rect 31216 10848 31232 10912
rect 31296 10848 31312 10912
rect 31376 10848 31382 10912
rect 31066 10847 31382 10848
rect 36066 10912 36382 10913
rect 36066 10848 36072 10912
rect 36136 10848 36152 10912
rect 36216 10848 36232 10912
rect 36296 10848 36312 10912
rect 36376 10848 36382 10912
rect 36066 10847 36382 10848
rect 41066 10912 41382 10913
rect 41066 10848 41072 10912
rect 41136 10848 41152 10912
rect 41216 10848 41232 10912
rect 41296 10848 41312 10912
rect 41376 10848 41382 10912
rect 41066 10847 41382 10848
rect 32949 10842 33015 10845
rect 34789 10842 34855 10845
rect 32949 10840 34855 10842
rect 32949 10784 32954 10840
rect 33010 10784 34794 10840
rect 34850 10784 34855 10840
rect 32949 10782 34855 10784
rect 32949 10779 33015 10782
rect 34789 10779 34855 10782
rect 33317 10706 33383 10709
rect 36813 10706 36879 10709
rect 33317 10704 36879 10706
rect 33317 10648 33322 10704
rect 33378 10648 36818 10704
rect 36874 10648 36879 10704
rect 33317 10646 36879 10648
rect 33317 10643 33383 10646
rect 36813 10643 36879 10646
rect 13261 10570 13327 10573
rect 37733 10570 37799 10573
rect 13261 10568 37799 10570
rect 13261 10512 13266 10568
rect 13322 10512 37738 10568
rect 37794 10512 37799 10568
rect 13261 10510 37799 10512
rect 13261 10507 13327 10510
rect 37733 10507 37799 10510
rect 3566 10368 3882 10369
rect 3566 10304 3572 10368
rect 3636 10304 3652 10368
rect 3716 10304 3732 10368
rect 3796 10304 3812 10368
rect 3876 10304 3882 10368
rect 3566 10303 3882 10304
rect 8566 10368 8882 10369
rect 8566 10304 8572 10368
rect 8636 10304 8652 10368
rect 8716 10304 8732 10368
rect 8796 10304 8812 10368
rect 8876 10304 8882 10368
rect 8566 10303 8882 10304
rect 13566 10368 13882 10369
rect 13566 10304 13572 10368
rect 13636 10304 13652 10368
rect 13716 10304 13732 10368
rect 13796 10304 13812 10368
rect 13876 10304 13882 10368
rect 13566 10303 13882 10304
rect 18566 10368 18882 10369
rect 18566 10304 18572 10368
rect 18636 10304 18652 10368
rect 18716 10304 18732 10368
rect 18796 10304 18812 10368
rect 18876 10304 18882 10368
rect 18566 10303 18882 10304
rect 23566 10368 23882 10369
rect 23566 10304 23572 10368
rect 23636 10304 23652 10368
rect 23716 10304 23732 10368
rect 23796 10304 23812 10368
rect 23876 10304 23882 10368
rect 23566 10303 23882 10304
rect 28566 10368 28882 10369
rect 28566 10304 28572 10368
rect 28636 10304 28652 10368
rect 28716 10304 28732 10368
rect 28796 10304 28812 10368
rect 28876 10304 28882 10368
rect 28566 10303 28882 10304
rect 33566 10368 33882 10369
rect 33566 10304 33572 10368
rect 33636 10304 33652 10368
rect 33716 10304 33732 10368
rect 33796 10304 33812 10368
rect 33876 10304 33882 10368
rect 33566 10303 33882 10304
rect 38566 10368 38882 10369
rect 38566 10304 38572 10368
rect 38636 10304 38652 10368
rect 38716 10304 38732 10368
rect 38796 10304 38812 10368
rect 38876 10304 38882 10368
rect 38566 10303 38882 10304
rect 43566 10368 43882 10369
rect 43566 10304 43572 10368
rect 43636 10304 43652 10368
rect 43716 10304 43732 10368
rect 43796 10304 43812 10368
rect 43876 10304 43882 10368
rect 43566 10303 43882 10304
rect 32305 10298 32371 10301
rect 32857 10298 32923 10301
rect 32305 10296 32923 10298
rect 32305 10240 32310 10296
rect 32366 10240 32862 10296
rect 32918 10240 32923 10296
rect 32305 10238 32923 10240
rect 32305 10235 32371 10238
rect 32857 10235 32923 10238
rect 29361 10162 29427 10165
rect 33501 10162 33567 10165
rect 29361 10160 33567 10162
rect 29361 10104 29366 10160
rect 29422 10104 33506 10160
rect 33562 10104 33567 10160
rect 29361 10102 33567 10104
rect 29361 10099 29427 10102
rect 33501 10099 33567 10102
rect 32397 10026 32463 10029
rect 33593 10026 33659 10029
rect 32397 10024 33659 10026
rect 32397 9968 32402 10024
rect 32458 9968 33598 10024
rect 33654 9968 33659 10024
rect 32397 9966 33659 9968
rect 32397 9963 32463 9966
rect 33593 9963 33659 9966
rect 22829 9890 22895 9893
rect 23381 9890 23447 9893
rect 22829 9888 23447 9890
rect 22829 9832 22834 9888
rect 22890 9832 23386 9888
rect 23442 9832 23447 9888
rect 22829 9830 23447 9832
rect 22829 9827 22895 9830
rect 23381 9827 23447 9830
rect 6066 9824 6382 9825
rect 6066 9760 6072 9824
rect 6136 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6382 9824
rect 6066 9759 6382 9760
rect 11066 9824 11382 9825
rect 11066 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11382 9824
rect 11066 9759 11382 9760
rect 16066 9824 16382 9825
rect 16066 9760 16072 9824
rect 16136 9760 16152 9824
rect 16216 9760 16232 9824
rect 16296 9760 16312 9824
rect 16376 9760 16382 9824
rect 16066 9759 16382 9760
rect 21066 9824 21382 9825
rect 21066 9760 21072 9824
rect 21136 9760 21152 9824
rect 21216 9760 21232 9824
rect 21296 9760 21312 9824
rect 21376 9760 21382 9824
rect 21066 9759 21382 9760
rect 26066 9824 26382 9825
rect 26066 9760 26072 9824
rect 26136 9760 26152 9824
rect 26216 9760 26232 9824
rect 26296 9760 26312 9824
rect 26376 9760 26382 9824
rect 26066 9759 26382 9760
rect 31066 9824 31382 9825
rect 31066 9760 31072 9824
rect 31136 9760 31152 9824
rect 31216 9760 31232 9824
rect 31296 9760 31312 9824
rect 31376 9760 31382 9824
rect 31066 9759 31382 9760
rect 36066 9824 36382 9825
rect 36066 9760 36072 9824
rect 36136 9760 36152 9824
rect 36216 9760 36232 9824
rect 36296 9760 36312 9824
rect 36376 9760 36382 9824
rect 36066 9759 36382 9760
rect 41066 9824 41382 9825
rect 41066 9760 41072 9824
rect 41136 9760 41152 9824
rect 41216 9760 41232 9824
rect 41296 9760 41312 9824
rect 41376 9760 41382 9824
rect 41066 9759 41382 9760
rect 30230 9692 30236 9756
rect 30300 9754 30306 9756
rect 30465 9754 30531 9757
rect 30300 9752 30531 9754
rect 30300 9696 30470 9752
rect 30526 9696 30531 9752
rect 30300 9694 30531 9696
rect 30300 9692 30306 9694
rect 30465 9691 30531 9694
rect 28165 9620 28231 9621
rect 28165 9618 28212 9620
rect 28120 9616 28212 9618
rect 28120 9560 28170 9616
rect 28120 9558 28212 9560
rect 28165 9556 28212 9558
rect 28276 9556 28282 9620
rect 32029 9618 32095 9621
rect 32806 9618 32812 9620
rect 32029 9616 32812 9618
rect 32029 9560 32034 9616
rect 32090 9560 32812 9616
rect 32029 9558 32812 9560
rect 28165 9555 28231 9556
rect 32029 9555 32095 9558
rect 32806 9556 32812 9558
rect 32876 9618 32882 9620
rect 34697 9618 34763 9621
rect 32876 9616 34763 9618
rect 32876 9560 34702 9616
rect 34758 9560 34763 9616
rect 32876 9558 34763 9560
rect 32876 9556 32882 9558
rect 34697 9555 34763 9558
rect 42517 9618 42583 9621
rect 44725 9618 44791 9621
rect 42517 9616 44791 9618
rect 42517 9560 42522 9616
rect 42578 9560 44730 9616
rect 44786 9560 44791 9616
rect 42517 9558 44791 9560
rect 42517 9555 42583 9558
rect 44725 9555 44791 9558
rect 21173 9482 21239 9485
rect 23473 9482 23539 9485
rect 33593 9482 33659 9485
rect 21173 9480 23539 9482
rect 21173 9424 21178 9480
rect 21234 9424 23478 9480
rect 23534 9424 23539 9480
rect 21173 9422 23539 9424
rect 21173 9419 21239 9422
rect 23473 9419 23539 9422
rect 33412 9480 33659 9482
rect 33412 9424 33598 9480
rect 33654 9424 33659 9480
rect 33412 9422 33659 9424
rect 3566 9280 3882 9281
rect 3566 9216 3572 9280
rect 3636 9216 3652 9280
rect 3716 9216 3732 9280
rect 3796 9216 3812 9280
rect 3876 9216 3882 9280
rect 3566 9215 3882 9216
rect 8566 9280 8882 9281
rect 8566 9216 8572 9280
rect 8636 9216 8652 9280
rect 8716 9216 8732 9280
rect 8796 9216 8812 9280
rect 8876 9216 8882 9280
rect 8566 9215 8882 9216
rect 13566 9280 13882 9281
rect 13566 9216 13572 9280
rect 13636 9216 13652 9280
rect 13716 9216 13732 9280
rect 13796 9216 13812 9280
rect 13876 9216 13882 9280
rect 13566 9215 13882 9216
rect 18566 9280 18882 9281
rect 18566 9216 18572 9280
rect 18636 9216 18652 9280
rect 18716 9216 18732 9280
rect 18796 9216 18812 9280
rect 18876 9216 18882 9280
rect 18566 9215 18882 9216
rect 23566 9280 23882 9281
rect 23566 9216 23572 9280
rect 23636 9216 23652 9280
rect 23716 9216 23732 9280
rect 23796 9216 23812 9280
rect 23876 9216 23882 9280
rect 23566 9215 23882 9216
rect 28566 9280 28882 9281
rect 28566 9216 28572 9280
rect 28636 9216 28652 9280
rect 28716 9216 28732 9280
rect 28796 9216 28812 9280
rect 28876 9216 28882 9280
rect 28566 9215 28882 9216
rect 11237 9210 11303 9213
rect 13261 9210 13327 9213
rect 11237 9208 13327 9210
rect 11237 9152 11242 9208
rect 11298 9152 13266 9208
rect 13322 9152 13327 9208
rect 11237 9150 13327 9152
rect 11237 9147 11303 9150
rect 13261 9147 13327 9150
rect 13077 9074 13143 9077
rect 13537 9074 13603 9077
rect 13077 9072 13603 9074
rect 13077 9016 13082 9072
rect 13138 9016 13542 9072
rect 13598 9016 13603 9072
rect 13077 9014 13603 9016
rect 13077 9011 13143 9014
rect 13537 9011 13603 9014
rect 22001 9074 22067 9077
rect 25037 9074 25103 9077
rect 22001 9072 25103 9074
rect 22001 9016 22006 9072
rect 22062 9016 25042 9072
rect 25098 9016 25103 9072
rect 22001 9014 25103 9016
rect 22001 9011 22067 9014
rect 25037 9011 25103 9014
rect 29545 9074 29611 9077
rect 31201 9074 31267 9077
rect 29545 9072 31267 9074
rect 29545 9016 29550 9072
rect 29606 9016 31206 9072
rect 31262 9016 31267 9072
rect 29545 9014 31267 9016
rect 33412 9074 33472 9422
rect 33593 9419 33659 9422
rect 33566 9280 33882 9281
rect 33566 9216 33572 9280
rect 33636 9216 33652 9280
rect 33716 9216 33732 9280
rect 33796 9216 33812 9280
rect 33876 9216 33882 9280
rect 33566 9215 33882 9216
rect 38566 9280 38882 9281
rect 38566 9216 38572 9280
rect 38636 9216 38652 9280
rect 38716 9216 38732 9280
rect 38796 9216 38812 9280
rect 38876 9216 38882 9280
rect 38566 9215 38882 9216
rect 43566 9280 43882 9281
rect 43566 9216 43572 9280
rect 43636 9216 43652 9280
rect 43716 9216 43732 9280
rect 43796 9216 43812 9280
rect 43876 9216 43882 9280
rect 43566 9215 43882 9216
rect 34053 9210 34119 9213
rect 36077 9210 36143 9213
rect 34053 9208 36143 9210
rect 34053 9152 34058 9208
rect 34114 9152 36082 9208
rect 36138 9152 36143 9208
rect 34053 9150 36143 9152
rect 34053 9147 34119 9150
rect 36077 9147 36143 9150
rect 35525 9074 35591 9077
rect 41965 9074 42031 9077
rect 33412 9014 33610 9074
rect 29545 9011 29611 9014
rect 31201 9011 31267 9014
rect 33550 8941 33610 9014
rect 35525 9072 42031 9074
rect 35525 9016 35530 9072
rect 35586 9016 41970 9072
rect 42026 9016 42031 9072
rect 35525 9014 42031 9016
rect 35525 9011 35591 9014
rect 41965 9011 42031 9014
rect 11973 8938 12039 8941
rect 13813 8938 13879 8941
rect 11973 8936 13879 8938
rect 11973 8880 11978 8936
rect 12034 8880 13818 8936
rect 13874 8880 13879 8936
rect 11973 8878 13879 8880
rect 11973 8875 12039 8878
rect 13813 8875 13879 8878
rect 15837 8938 15903 8941
rect 26509 8938 26575 8941
rect 15837 8936 26575 8938
rect 15837 8880 15842 8936
rect 15898 8880 26514 8936
rect 26570 8880 26575 8936
rect 15837 8878 26575 8880
rect 15837 8875 15903 8878
rect 26509 8875 26575 8878
rect 30097 8938 30163 8941
rect 30741 8938 30807 8941
rect 33501 8938 33610 8941
rect 36169 8938 36235 8941
rect 30097 8936 36235 8938
rect 30097 8880 30102 8936
rect 30158 8880 30746 8936
rect 30802 8880 33506 8936
rect 33562 8880 36174 8936
rect 36230 8880 36235 8936
rect 30097 8878 36235 8880
rect 30097 8875 30163 8878
rect 30741 8875 30807 8878
rect 33501 8875 33567 8878
rect 36169 8875 36235 8878
rect -300 8802 160 8832
rect 933 8802 999 8805
rect -300 8800 999 8802
rect -300 8744 938 8800
rect 994 8744 999 8800
rect -300 8742 999 8744
rect -300 8712 160 8742
rect 933 8739 999 8742
rect 22369 8802 22435 8805
rect 23381 8802 23447 8805
rect 22369 8800 23447 8802
rect 22369 8744 22374 8800
rect 22430 8744 23386 8800
rect 23442 8744 23447 8800
rect 22369 8742 23447 8744
rect 22369 8739 22435 8742
rect 23381 8739 23447 8742
rect 33225 8802 33291 8805
rect 34881 8802 34947 8805
rect 33225 8800 34947 8802
rect 33225 8744 33230 8800
rect 33286 8744 34886 8800
rect 34942 8744 34947 8800
rect 33225 8742 34947 8744
rect 33225 8739 33291 8742
rect 34881 8739 34947 8742
rect 44633 8802 44699 8805
rect 45840 8802 46300 8832
rect 44633 8800 46300 8802
rect 44633 8744 44638 8800
rect 44694 8744 46300 8800
rect 44633 8742 46300 8744
rect 44633 8739 44699 8742
rect 6066 8736 6382 8737
rect 6066 8672 6072 8736
rect 6136 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6382 8736
rect 6066 8671 6382 8672
rect 11066 8736 11382 8737
rect 11066 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11382 8736
rect 11066 8671 11382 8672
rect 16066 8736 16382 8737
rect 16066 8672 16072 8736
rect 16136 8672 16152 8736
rect 16216 8672 16232 8736
rect 16296 8672 16312 8736
rect 16376 8672 16382 8736
rect 16066 8671 16382 8672
rect 21066 8736 21382 8737
rect 21066 8672 21072 8736
rect 21136 8672 21152 8736
rect 21216 8672 21232 8736
rect 21296 8672 21312 8736
rect 21376 8672 21382 8736
rect 21066 8671 21382 8672
rect 26066 8736 26382 8737
rect 26066 8672 26072 8736
rect 26136 8672 26152 8736
rect 26216 8672 26232 8736
rect 26296 8672 26312 8736
rect 26376 8672 26382 8736
rect 26066 8671 26382 8672
rect 31066 8736 31382 8737
rect 31066 8672 31072 8736
rect 31136 8672 31152 8736
rect 31216 8672 31232 8736
rect 31296 8672 31312 8736
rect 31376 8672 31382 8736
rect 31066 8671 31382 8672
rect 36066 8736 36382 8737
rect 36066 8672 36072 8736
rect 36136 8672 36152 8736
rect 36216 8672 36232 8736
rect 36296 8672 36312 8736
rect 36376 8672 36382 8736
rect 36066 8671 36382 8672
rect 41066 8736 41382 8737
rect 41066 8672 41072 8736
rect 41136 8672 41152 8736
rect 41216 8672 41232 8736
rect 41296 8672 41312 8736
rect 41376 8672 41382 8736
rect 45840 8712 46300 8742
rect 41066 8671 41382 8672
rect 34329 8666 34395 8669
rect 34881 8666 34947 8669
rect 34329 8664 34947 8666
rect 34329 8608 34334 8664
rect 34390 8608 34886 8664
rect 34942 8608 34947 8664
rect 34329 8606 34947 8608
rect 34329 8603 34395 8606
rect 34881 8603 34947 8606
rect 28717 8530 28783 8533
rect 32489 8530 32555 8533
rect 36537 8530 36603 8533
rect 28717 8528 36603 8530
rect 28717 8472 28722 8528
rect 28778 8472 32494 8528
rect 32550 8472 36542 8528
rect 36598 8472 36603 8528
rect 28717 8470 36603 8472
rect 28717 8467 28783 8470
rect 32489 8467 32555 8470
rect 36537 8467 36603 8470
rect 38745 8530 38811 8533
rect 40033 8530 40099 8533
rect 38745 8528 40099 8530
rect 38745 8472 38750 8528
rect 38806 8472 40038 8528
rect 40094 8472 40099 8528
rect 38745 8470 40099 8472
rect 38745 8467 38811 8470
rect 40033 8467 40099 8470
rect 21541 8394 21607 8397
rect 25589 8394 25655 8397
rect 21541 8392 25655 8394
rect 21541 8336 21546 8392
rect 21602 8336 25594 8392
rect 25650 8336 25655 8392
rect 21541 8334 25655 8336
rect 21541 8331 21607 8334
rect 25589 8331 25655 8334
rect 27981 8394 28047 8397
rect 28533 8394 28599 8397
rect 27981 8392 28599 8394
rect 27981 8336 27986 8392
rect 28042 8336 28538 8392
rect 28594 8336 28599 8392
rect 27981 8334 28599 8336
rect 27981 8331 28047 8334
rect 28533 8331 28599 8334
rect 29177 8394 29243 8397
rect 32121 8394 32187 8397
rect 29177 8392 32187 8394
rect 29177 8336 29182 8392
rect 29238 8336 32126 8392
rect 32182 8336 32187 8392
rect 29177 8334 32187 8336
rect 29177 8331 29243 8334
rect 32121 8331 32187 8334
rect 33317 8394 33383 8397
rect 34421 8396 34487 8397
rect 34278 8394 34284 8396
rect 33317 8392 34284 8394
rect 33317 8336 33322 8392
rect 33378 8336 34284 8392
rect 33317 8334 34284 8336
rect 33317 8331 33383 8334
rect 34278 8332 34284 8334
rect 34348 8332 34354 8396
rect 34421 8392 34468 8396
rect 34532 8394 34538 8396
rect 35341 8394 35407 8397
rect 36169 8394 36235 8397
rect 34421 8336 34426 8392
rect 34421 8332 34468 8336
rect 34532 8334 34578 8394
rect 35341 8392 36235 8394
rect 35341 8336 35346 8392
rect 35402 8336 36174 8392
rect 36230 8336 36235 8392
rect 35341 8334 36235 8336
rect 34532 8332 34538 8334
rect 34421 8331 34487 8332
rect 35341 8331 35407 8334
rect 36169 8331 36235 8334
rect 31661 8258 31727 8261
rect 31661 8256 31954 8258
rect 31661 8200 31666 8256
rect 31722 8200 31954 8256
rect 31661 8198 31954 8200
rect 31661 8195 31727 8198
rect 3566 8192 3882 8193
rect 3566 8128 3572 8192
rect 3636 8128 3652 8192
rect 3716 8128 3732 8192
rect 3796 8128 3812 8192
rect 3876 8128 3882 8192
rect 3566 8127 3882 8128
rect 8566 8192 8882 8193
rect 8566 8128 8572 8192
rect 8636 8128 8652 8192
rect 8716 8128 8732 8192
rect 8796 8128 8812 8192
rect 8876 8128 8882 8192
rect 8566 8127 8882 8128
rect 13566 8192 13882 8193
rect 13566 8128 13572 8192
rect 13636 8128 13652 8192
rect 13716 8128 13732 8192
rect 13796 8128 13812 8192
rect 13876 8128 13882 8192
rect 13566 8127 13882 8128
rect 18566 8192 18882 8193
rect 18566 8128 18572 8192
rect 18636 8128 18652 8192
rect 18716 8128 18732 8192
rect 18796 8128 18812 8192
rect 18876 8128 18882 8192
rect 18566 8127 18882 8128
rect 23566 8192 23882 8193
rect 23566 8128 23572 8192
rect 23636 8128 23652 8192
rect 23716 8128 23732 8192
rect 23796 8128 23812 8192
rect 23876 8128 23882 8192
rect 23566 8127 23882 8128
rect 28566 8192 28882 8193
rect 28566 8128 28572 8192
rect 28636 8128 28652 8192
rect 28716 8128 28732 8192
rect 28796 8128 28812 8192
rect 28876 8128 28882 8192
rect 28566 8127 28882 8128
rect 26785 7986 26851 7989
rect 28441 7986 28507 7989
rect 26785 7984 28507 7986
rect 26785 7928 26790 7984
rect 26846 7928 28446 7984
rect 28502 7928 28507 7984
rect 26785 7926 28507 7928
rect 26785 7923 26851 7926
rect 28441 7923 28507 7926
rect 30189 7986 30255 7989
rect 31894 7986 31954 8198
rect 33566 8192 33882 8193
rect 33566 8128 33572 8192
rect 33636 8128 33652 8192
rect 33716 8128 33732 8192
rect 33796 8128 33812 8192
rect 33876 8128 33882 8192
rect 33566 8127 33882 8128
rect 38566 8192 38882 8193
rect 38566 8128 38572 8192
rect 38636 8128 38652 8192
rect 38716 8128 38732 8192
rect 38796 8128 38812 8192
rect 38876 8128 38882 8192
rect 38566 8127 38882 8128
rect 43566 8192 43882 8193
rect 43566 8128 43572 8192
rect 43636 8128 43652 8192
rect 43716 8128 43732 8192
rect 43796 8128 43812 8192
rect 43876 8128 43882 8192
rect 43566 8127 43882 8128
rect 36629 7986 36695 7989
rect 30189 7984 36695 7986
rect 30189 7928 30194 7984
rect 30250 7928 36634 7984
rect 36690 7928 36695 7984
rect 30189 7926 36695 7928
rect 30189 7923 30255 7926
rect 36629 7923 36695 7926
rect 37733 7986 37799 7989
rect 40861 7986 40927 7989
rect 37733 7984 40927 7986
rect 37733 7928 37738 7984
rect 37794 7928 40866 7984
rect 40922 7928 40927 7984
rect 37733 7926 40927 7928
rect 37733 7923 37799 7926
rect 40861 7923 40927 7926
rect 25497 7850 25563 7853
rect 25630 7850 25636 7852
rect 25497 7848 25636 7850
rect 25497 7792 25502 7848
rect 25558 7792 25636 7848
rect 25497 7790 25636 7792
rect 25497 7787 25563 7790
rect 25630 7788 25636 7790
rect 25700 7850 25706 7852
rect 26509 7850 26575 7853
rect 25700 7848 26575 7850
rect 25700 7792 26514 7848
rect 26570 7792 26575 7848
rect 25700 7790 26575 7792
rect 25700 7788 25706 7790
rect 26509 7787 26575 7790
rect 30465 7850 30531 7853
rect 42885 7850 42951 7853
rect 30465 7848 42951 7850
rect 30465 7792 30470 7848
rect 30526 7792 42890 7848
rect 42946 7792 42951 7848
rect 30465 7790 42951 7792
rect 30465 7787 30531 7790
rect 42885 7787 42951 7790
rect 6066 7648 6382 7649
rect 6066 7584 6072 7648
rect 6136 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6382 7648
rect 6066 7583 6382 7584
rect 11066 7648 11382 7649
rect 11066 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11382 7648
rect 11066 7583 11382 7584
rect 16066 7648 16382 7649
rect 16066 7584 16072 7648
rect 16136 7584 16152 7648
rect 16216 7584 16232 7648
rect 16296 7584 16312 7648
rect 16376 7584 16382 7648
rect 16066 7583 16382 7584
rect 21066 7648 21382 7649
rect 21066 7584 21072 7648
rect 21136 7584 21152 7648
rect 21216 7584 21232 7648
rect 21296 7584 21312 7648
rect 21376 7584 21382 7648
rect 21066 7583 21382 7584
rect 26066 7648 26382 7649
rect 26066 7584 26072 7648
rect 26136 7584 26152 7648
rect 26216 7584 26232 7648
rect 26296 7584 26312 7648
rect 26376 7584 26382 7648
rect 26066 7583 26382 7584
rect 31066 7648 31382 7649
rect 31066 7584 31072 7648
rect 31136 7584 31152 7648
rect 31216 7584 31232 7648
rect 31296 7584 31312 7648
rect 31376 7584 31382 7648
rect 31066 7583 31382 7584
rect 36066 7648 36382 7649
rect 36066 7584 36072 7648
rect 36136 7584 36152 7648
rect 36216 7584 36232 7648
rect 36296 7584 36312 7648
rect 36376 7584 36382 7648
rect 36066 7583 36382 7584
rect 41066 7648 41382 7649
rect 41066 7584 41072 7648
rect 41136 7584 41152 7648
rect 41216 7584 41232 7648
rect 41296 7584 41312 7648
rect 41376 7584 41382 7648
rect 41066 7583 41382 7584
rect 27429 7442 27495 7445
rect 31109 7442 31175 7445
rect 27429 7440 31175 7442
rect 27429 7384 27434 7440
rect 27490 7384 31114 7440
rect 31170 7384 31175 7440
rect 27429 7382 31175 7384
rect 27429 7379 27495 7382
rect 31109 7379 31175 7382
rect 35157 7442 35223 7445
rect 44173 7442 44239 7445
rect 35157 7440 44239 7442
rect 35157 7384 35162 7440
rect 35218 7384 44178 7440
rect 44234 7384 44239 7440
rect 35157 7382 44239 7384
rect 35157 7379 35223 7382
rect 44173 7379 44239 7382
rect 22553 7306 22619 7309
rect 24117 7306 24183 7309
rect 22553 7304 24183 7306
rect 22553 7248 22558 7304
rect 22614 7248 24122 7304
rect 24178 7248 24183 7304
rect 22553 7246 24183 7248
rect 22553 7243 22619 7246
rect 24117 7243 24183 7246
rect 25773 7306 25839 7309
rect 30833 7306 30899 7309
rect 31886 7306 31892 7308
rect 25773 7304 31892 7306
rect 25773 7248 25778 7304
rect 25834 7248 30838 7304
rect 30894 7248 31892 7304
rect 25773 7246 31892 7248
rect 25773 7243 25839 7246
rect 30833 7243 30899 7246
rect 31886 7244 31892 7246
rect 31956 7306 31962 7308
rect 35893 7306 35959 7309
rect 31956 7304 35959 7306
rect 31956 7248 35898 7304
rect 35954 7248 35959 7304
rect 31956 7246 35959 7248
rect 31956 7244 31962 7246
rect 35893 7243 35959 7246
rect 3566 7104 3882 7105
rect 3566 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3812 7104
rect 3876 7040 3882 7104
rect 3566 7039 3882 7040
rect 8566 7104 8882 7105
rect 8566 7040 8572 7104
rect 8636 7040 8652 7104
rect 8716 7040 8732 7104
rect 8796 7040 8812 7104
rect 8876 7040 8882 7104
rect 8566 7039 8882 7040
rect 13566 7104 13882 7105
rect 13566 7040 13572 7104
rect 13636 7040 13652 7104
rect 13716 7040 13732 7104
rect 13796 7040 13812 7104
rect 13876 7040 13882 7104
rect 13566 7039 13882 7040
rect 18566 7104 18882 7105
rect 18566 7040 18572 7104
rect 18636 7040 18652 7104
rect 18716 7040 18732 7104
rect 18796 7040 18812 7104
rect 18876 7040 18882 7104
rect 18566 7039 18882 7040
rect 23566 7104 23882 7105
rect 23566 7040 23572 7104
rect 23636 7040 23652 7104
rect 23716 7040 23732 7104
rect 23796 7040 23812 7104
rect 23876 7040 23882 7104
rect 23566 7039 23882 7040
rect 28566 7104 28882 7105
rect 28566 7040 28572 7104
rect 28636 7040 28652 7104
rect 28716 7040 28732 7104
rect 28796 7040 28812 7104
rect 28876 7040 28882 7104
rect 28566 7039 28882 7040
rect 33566 7104 33882 7105
rect 33566 7040 33572 7104
rect 33636 7040 33652 7104
rect 33716 7040 33732 7104
rect 33796 7040 33812 7104
rect 33876 7040 33882 7104
rect 33566 7039 33882 7040
rect 38566 7104 38882 7105
rect 38566 7040 38572 7104
rect 38636 7040 38652 7104
rect 38716 7040 38732 7104
rect 38796 7040 38812 7104
rect 38876 7040 38882 7104
rect 38566 7039 38882 7040
rect 43566 7104 43882 7105
rect 43566 7040 43572 7104
rect 43636 7040 43652 7104
rect 43716 7040 43732 7104
rect 43796 7040 43812 7104
rect 43876 7040 43882 7104
rect 43566 7039 43882 7040
rect 23013 7036 23079 7037
rect 23013 7034 23060 7036
rect 22968 7032 23060 7034
rect 22968 6976 23018 7032
rect 22968 6974 23060 6976
rect 23013 6972 23060 6974
rect 23124 6972 23130 7036
rect 24902 6974 26434 7034
rect 23013 6971 23079 6972
rect 9213 6900 9279 6901
rect 19793 6900 19859 6901
rect 9213 6898 9260 6900
rect 9168 6896 9260 6898
rect 9168 6840 9218 6896
rect 9168 6838 9260 6840
rect 9213 6836 9260 6838
rect 9324 6836 9330 6900
rect 17534 6836 17540 6900
rect 17604 6836 17610 6900
rect 19742 6898 19748 6900
rect 19702 6838 19748 6898
rect 19812 6896 19859 6900
rect 19854 6840 19859 6896
rect 19742 6836 19748 6838
rect 19812 6836 19859 6840
rect 22870 6836 22876 6900
rect 22940 6898 22946 6900
rect 23013 6898 23079 6901
rect 24301 6900 24367 6901
rect 24301 6898 24348 6900
rect 22940 6896 23079 6898
rect 22940 6840 23018 6896
rect 23074 6840 23079 6896
rect 22940 6838 23079 6840
rect 24256 6896 24348 6898
rect 24256 6840 24306 6896
rect 24256 6838 24348 6840
rect 22940 6836 22946 6838
rect 9213 6835 9279 6836
rect 17542 6762 17602 6836
rect 19793 6835 19859 6836
rect 23013 6835 23079 6838
rect 24301 6836 24348 6838
rect 24412 6836 24418 6900
rect 24761 6898 24827 6901
rect 24902 6898 24962 6974
rect 24761 6896 24962 6898
rect 24761 6840 24766 6896
rect 24822 6840 24962 6896
rect 24761 6838 24962 6840
rect 25037 6898 25103 6901
rect 25814 6898 25820 6900
rect 25037 6896 25820 6898
rect 25037 6840 25042 6896
rect 25098 6840 25820 6896
rect 25037 6838 25820 6840
rect 24301 6835 24367 6836
rect 24761 6835 24827 6838
rect 25037 6835 25103 6838
rect 25814 6836 25820 6838
rect 25884 6898 25890 6900
rect 26141 6898 26207 6901
rect 25884 6896 26207 6898
rect 25884 6840 26146 6896
rect 26202 6840 26207 6896
rect 25884 6838 26207 6840
rect 26374 6898 26434 6974
rect 27153 6898 27219 6901
rect 31017 6898 31083 6901
rect 26374 6896 31083 6898
rect 26374 6840 27158 6896
rect 27214 6840 31022 6896
rect 31078 6840 31083 6896
rect 26374 6838 31083 6840
rect 25884 6836 25890 6838
rect 26141 6835 26207 6838
rect 27153 6835 27219 6838
rect 31017 6835 31083 6838
rect 38101 6898 38167 6901
rect 42701 6898 42767 6901
rect 38101 6896 42767 6898
rect 38101 6840 38106 6896
rect 38162 6840 42706 6896
rect 42762 6840 42767 6896
rect 38101 6838 42767 6840
rect 38101 6835 38167 6838
rect 42701 6835 42767 6838
rect 25589 6762 25655 6765
rect 35709 6762 35775 6765
rect 17542 6760 25655 6762
rect 17542 6704 25594 6760
rect 25650 6704 25655 6760
rect 17542 6702 25655 6704
rect 25589 6699 25655 6702
rect 25776 6760 35775 6762
rect 25776 6704 35714 6760
rect 35770 6704 35775 6760
rect 25776 6702 35775 6704
rect 22461 6626 22527 6629
rect 24117 6626 24183 6629
rect 25776 6626 25836 6702
rect 35709 6699 35775 6702
rect 35985 6762 36051 6765
rect 36721 6762 36787 6765
rect 35985 6760 36787 6762
rect 35985 6704 35990 6760
rect 36046 6704 36726 6760
rect 36782 6704 36787 6760
rect 35985 6702 36787 6704
rect 35985 6699 36051 6702
rect 36721 6699 36787 6702
rect 22461 6624 24183 6626
rect 22461 6568 22466 6624
rect 22522 6568 24122 6624
rect 24178 6568 24183 6624
rect 22461 6566 24183 6568
rect 22461 6563 22527 6566
rect 24117 6563 24183 6566
rect 25408 6566 25836 6626
rect 6066 6560 6382 6561
rect 6066 6496 6072 6560
rect 6136 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6382 6560
rect 6066 6495 6382 6496
rect 11066 6560 11382 6561
rect 11066 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11382 6560
rect 11066 6495 11382 6496
rect 16066 6560 16382 6561
rect 16066 6496 16072 6560
rect 16136 6496 16152 6560
rect 16216 6496 16232 6560
rect 16296 6496 16312 6560
rect 16376 6496 16382 6560
rect 16066 6495 16382 6496
rect 21066 6560 21382 6561
rect 21066 6496 21072 6560
rect 21136 6496 21152 6560
rect 21216 6496 21232 6560
rect 21296 6496 21312 6560
rect 21376 6496 21382 6560
rect 21066 6495 21382 6496
rect 25408 6493 25468 6566
rect 26066 6560 26382 6561
rect 26066 6496 26072 6560
rect 26136 6496 26152 6560
rect 26216 6496 26232 6560
rect 26296 6496 26312 6560
rect 26376 6496 26382 6560
rect 26066 6495 26382 6496
rect 31066 6560 31382 6561
rect 31066 6496 31072 6560
rect 31136 6496 31152 6560
rect 31216 6496 31232 6560
rect 31296 6496 31312 6560
rect 31376 6496 31382 6560
rect 31066 6495 31382 6496
rect 36066 6560 36382 6561
rect 36066 6496 36072 6560
rect 36136 6496 36152 6560
rect 36216 6496 36232 6560
rect 36296 6496 36312 6560
rect 36376 6496 36382 6560
rect 36066 6495 36382 6496
rect 41066 6560 41382 6561
rect 41066 6496 41072 6560
rect 41136 6496 41152 6560
rect 41216 6496 41232 6560
rect 41296 6496 41312 6560
rect 41376 6496 41382 6560
rect 41066 6495 41382 6496
rect 16982 6428 16988 6492
rect 17052 6490 17058 6492
rect 20897 6490 20963 6493
rect 25405 6490 25471 6493
rect 17052 6488 20963 6490
rect 17052 6432 20902 6488
rect 20958 6432 20963 6488
rect 17052 6430 20963 6432
rect 17052 6428 17058 6430
rect 20897 6427 20963 6430
rect 23292 6488 25471 6490
rect 23292 6432 25410 6488
rect 25466 6432 25471 6488
rect 23292 6430 25471 6432
rect 13353 6354 13419 6357
rect 23105 6354 23171 6357
rect 13353 6352 23171 6354
rect 13353 6296 13358 6352
rect 13414 6296 23110 6352
rect 23166 6296 23171 6352
rect 13353 6294 23171 6296
rect 13353 6291 13419 6294
rect 23105 6291 23171 6294
rect 13629 6218 13695 6221
rect 23292 6218 23352 6430
rect 25405 6427 25471 6430
rect 25129 6354 25195 6357
rect 32857 6354 32923 6357
rect 25129 6352 32923 6354
rect 25129 6296 25134 6352
rect 25190 6296 32862 6352
rect 32918 6296 32923 6352
rect 25129 6294 32923 6296
rect 25129 6291 25195 6294
rect 32857 6291 32923 6294
rect 33777 6354 33843 6357
rect 38101 6354 38167 6357
rect 33777 6352 38167 6354
rect 33777 6296 33782 6352
rect 33838 6296 38106 6352
rect 38162 6296 38167 6352
rect 33777 6294 38167 6296
rect 33777 6291 33843 6294
rect 38101 6291 38167 6294
rect 25589 6218 25655 6221
rect 13629 6216 23352 6218
rect 13629 6160 13634 6216
rect 13690 6160 23352 6216
rect 13629 6158 23352 6160
rect 23430 6216 25655 6218
rect 23430 6160 25594 6216
rect 25650 6160 25655 6216
rect 23430 6158 25655 6160
rect 13629 6155 13695 6158
rect 16113 6082 16179 6085
rect 16849 6082 16915 6085
rect 16113 6080 16915 6082
rect 16113 6024 16118 6080
rect 16174 6024 16854 6080
rect 16910 6024 16915 6080
rect 16113 6022 16915 6024
rect 16113 6019 16179 6022
rect 16849 6019 16915 6022
rect 19057 6082 19123 6085
rect 23430 6082 23490 6158
rect 25589 6155 25655 6158
rect 36997 6218 37063 6221
rect 40769 6218 40835 6221
rect 36997 6216 40835 6218
rect 36997 6160 37002 6216
rect 37058 6160 40774 6216
rect 40830 6160 40835 6216
rect 36997 6158 40835 6160
rect 36997 6155 37063 6158
rect 40769 6155 40835 6158
rect 19057 6080 23490 6082
rect 19057 6024 19062 6080
rect 19118 6024 23490 6080
rect 19057 6022 23490 6024
rect 24209 6082 24275 6085
rect 26734 6082 26740 6084
rect 24209 6080 26740 6082
rect 24209 6024 24214 6080
rect 24270 6024 26740 6080
rect 24209 6022 26740 6024
rect 19057 6019 19123 6022
rect 24209 6019 24275 6022
rect 26734 6020 26740 6022
rect 26804 6020 26810 6084
rect 3566 6016 3882 6017
rect 3566 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3812 6016
rect 3876 5952 3882 6016
rect 3566 5951 3882 5952
rect 8566 6016 8882 6017
rect 8566 5952 8572 6016
rect 8636 5952 8652 6016
rect 8716 5952 8732 6016
rect 8796 5952 8812 6016
rect 8876 5952 8882 6016
rect 8566 5951 8882 5952
rect 13566 6016 13882 6017
rect 13566 5952 13572 6016
rect 13636 5952 13652 6016
rect 13716 5952 13732 6016
rect 13796 5952 13812 6016
rect 13876 5952 13882 6016
rect 13566 5951 13882 5952
rect 18566 6016 18882 6017
rect 18566 5952 18572 6016
rect 18636 5952 18652 6016
rect 18716 5952 18732 6016
rect 18796 5952 18812 6016
rect 18876 5952 18882 6016
rect 18566 5951 18882 5952
rect 23566 6016 23882 6017
rect 23566 5952 23572 6016
rect 23636 5952 23652 6016
rect 23716 5952 23732 6016
rect 23796 5952 23812 6016
rect 23876 5952 23882 6016
rect 23566 5951 23882 5952
rect 28566 6016 28882 6017
rect 28566 5952 28572 6016
rect 28636 5952 28652 6016
rect 28716 5952 28732 6016
rect 28796 5952 28812 6016
rect 28876 5952 28882 6016
rect 28566 5951 28882 5952
rect 33566 6016 33882 6017
rect 33566 5952 33572 6016
rect 33636 5952 33652 6016
rect 33716 5952 33732 6016
rect 33796 5952 33812 6016
rect 33876 5952 33882 6016
rect 33566 5951 33882 5952
rect 38566 6016 38882 6017
rect 38566 5952 38572 6016
rect 38636 5952 38652 6016
rect 38716 5952 38732 6016
rect 38796 5952 38812 6016
rect 38876 5952 38882 6016
rect 38566 5951 38882 5952
rect 43566 6016 43882 6017
rect 43566 5952 43572 6016
rect 43636 5952 43652 6016
rect 43716 5952 43732 6016
rect 43796 5952 43812 6016
rect 43876 5952 43882 6016
rect 43566 5951 43882 5952
rect 14457 5946 14523 5949
rect 17769 5946 17835 5949
rect 14457 5944 17835 5946
rect 14457 5888 14462 5944
rect 14518 5888 17774 5944
rect 17830 5888 17835 5944
rect 14457 5886 17835 5888
rect 14457 5883 14523 5886
rect 17769 5883 17835 5886
rect 22461 5946 22527 5949
rect 22686 5946 22692 5948
rect 22461 5944 22692 5946
rect 22461 5888 22466 5944
rect 22522 5888 22692 5944
rect 22461 5886 22692 5888
rect 22461 5883 22527 5886
rect 22686 5884 22692 5886
rect 22756 5946 22762 5948
rect 23381 5946 23447 5949
rect 22756 5944 23447 5946
rect 22756 5888 23386 5944
rect 23442 5888 23447 5944
rect 22756 5886 23447 5888
rect 22756 5884 22762 5886
rect 23381 5883 23447 5886
rect 25037 5946 25103 5949
rect 25037 5944 26020 5946
rect 25037 5888 25042 5944
rect 25098 5888 26020 5944
rect 25037 5886 26020 5888
rect 25037 5883 25103 5886
rect 14273 5810 14339 5813
rect 25129 5810 25195 5813
rect 14273 5808 25195 5810
rect 14273 5752 14278 5808
rect 14334 5752 25134 5808
rect 25190 5752 25195 5808
rect 14273 5750 25195 5752
rect 14273 5747 14339 5750
rect 25129 5747 25195 5750
rect 25589 5810 25655 5813
rect 25814 5810 25820 5812
rect 25589 5808 25820 5810
rect 25589 5752 25594 5808
rect 25650 5752 25820 5808
rect 25589 5750 25820 5752
rect 25589 5747 25655 5750
rect 25814 5748 25820 5750
rect 25884 5748 25890 5812
rect 25960 5810 26020 5886
rect 30189 5810 30255 5813
rect 25960 5808 30255 5810
rect 25960 5752 30194 5808
rect 30250 5752 30255 5808
rect 25960 5750 30255 5752
rect 30189 5747 30255 5750
rect 3417 5674 3483 5677
rect 14457 5674 14523 5677
rect 24301 5674 24367 5677
rect 3417 5672 24367 5674
rect 3417 5616 3422 5672
rect 3478 5616 14462 5672
rect 14518 5616 24306 5672
rect 24362 5616 24367 5672
rect 3417 5614 24367 5616
rect 3417 5611 3483 5614
rect 14457 5611 14523 5614
rect 24301 5611 24367 5614
rect 24485 5674 24551 5677
rect 33225 5676 33291 5677
rect 33174 5674 33180 5676
rect 24485 5672 33180 5674
rect 33244 5674 33291 5676
rect 33244 5672 33372 5674
rect 24485 5616 24490 5672
rect 24546 5616 33180 5672
rect 33286 5616 33372 5672
rect 24485 5614 33180 5616
rect 24485 5611 24551 5614
rect 33174 5612 33180 5614
rect 33244 5614 33372 5616
rect 33244 5612 33291 5614
rect 33225 5611 33291 5612
rect 17217 5538 17283 5541
rect 19885 5540 19951 5541
rect 23197 5540 23263 5541
rect 17534 5538 17540 5540
rect 17217 5536 17540 5538
rect 17217 5480 17222 5536
rect 17278 5480 17540 5536
rect 17217 5478 17540 5480
rect 17217 5475 17283 5478
rect 17534 5476 17540 5478
rect 17604 5476 17610 5540
rect 19885 5538 19932 5540
rect 19840 5536 19932 5538
rect 19840 5480 19890 5536
rect 19840 5478 19932 5480
rect 19885 5476 19932 5478
rect 19996 5476 20002 5540
rect 21582 5476 21588 5540
rect 21652 5538 21658 5540
rect 23197 5538 23244 5540
rect 21652 5478 22938 5538
rect 23152 5536 23244 5538
rect 23152 5480 23202 5536
rect 23152 5478 23244 5480
rect 21652 5476 21658 5478
rect 19885 5475 19951 5476
rect 6066 5472 6382 5473
rect 6066 5408 6072 5472
rect 6136 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6382 5472
rect 6066 5407 6382 5408
rect 11066 5472 11382 5473
rect 11066 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11382 5472
rect 11066 5407 11382 5408
rect 16066 5472 16382 5473
rect 16066 5408 16072 5472
rect 16136 5408 16152 5472
rect 16216 5408 16232 5472
rect 16296 5408 16312 5472
rect 16376 5408 16382 5472
rect 16066 5407 16382 5408
rect 21066 5472 21382 5473
rect 21066 5408 21072 5472
rect 21136 5408 21152 5472
rect 21216 5408 21232 5472
rect 21296 5408 21312 5472
rect 21376 5408 21382 5472
rect 21066 5407 21382 5408
rect 20805 5402 20871 5405
rect 22001 5404 22067 5405
rect 21950 5402 21956 5404
rect 16806 5400 20871 5402
rect 16806 5344 20810 5400
rect 20866 5344 20871 5400
rect 16806 5342 20871 5344
rect 21910 5342 21956 5402
rect 22020 5400 22067 5404
rect 22062 5344 22067 5400
rect 13721 5266 13787 5269
rect 16806 5266 16866 5342
rect 20805 5339 20871 5342
rect 21950 5340 21956 5342
rect 22020 5340 22067 5344
rect 22878 5402 22938 5478
rect 23197 5476 23244 5478
rect 23308 5476 23314 5540
rect 24577 5538 24643 5541
rect 25446 5538 25452 5540
rect 24577 5536 25452 5538
rect 24577 5480 24582 5536
rect 24638 5480 25452 5536
rect 24577 5478 25452 5480
rect 23197 5475 23263 5476
rect 24577 5475 24643 5478
rect 25446 5476 25452 5478
rect 25516 5476 25522 5540
rect 26066 5472 26382 5473
rect 26066 5408 26072 5472
rect 26136 5408 26152 5472
rect 26216 5408 26232 5472
rect 26296 5408 26312 5472
rect 26376 5408 26382 5472
rect 26066 5407 26382 5408
rect 31066 5472 31382 5473
rect 31066 5408 31072 5472
rect 31136 5408 31152 5472
rect 31216 5408 31232 5472
rect 31296 5408 31312 5472
rect 31376 5408 31382 5472
rect 31066 5407 31382 5408
rect 36066 5472 36382 5473
rect 36066 5408 36072 5472
rect 36136 5408 36152 5472
rect 36216 5408 36232 5472
rect 36296 5408 36312 5472
rect 36376 5408 36382 5472
rect 36066 5407 36382 5408
rect 41066 5472 41382 5473
rect 41066 5408 41072 5472
rect 41136 5408 41152 5472
rect 41216 5408 41232 5472
rect 41296 5408 41312 5472
rect 41376 5408 41382 5472
rect 41066 5407 41382 5408
rect 25037 5402 25103 5405
rect 22878 5400 25103 5402
rect 22878 5344 25042 5400
rect 25098 5344 25103 5400
rect 22878 5342 25103 5344
rect 22001 5339 22067 5340
rect 25037 5339 25103 5342
rect 13721 5264 16866 5266
rect 13721 5208 13726 5264
rect 13782 5208 16866 5264
rect 13721 5206 16866 5208
rect 13721 5203 13787 5206
rect 19190 5204 19196 5268
rect 19260 5266 19266 5268
rect 23289 5266 23355 5269
rect 19260 5264 23355 5266
rect 19260 5208 23294 5264
rect 23350 5208 23355 5264
rect 19260 5206 23355 5208
rect 19260 5204 19266 5206
rect 23289 5203 23355 5206
rect 25129 5266 25195 5269
rect 26969 5266 27035 5269
rect 25129 5264 34162 5266
rect 25129 5208 25134 5264
rect 25190 5208 26974 5264
rect 27030 5208 34162 5264
rect 25129 5206 34162 5208
rect 25129 5203 25195 5206
rect 26969 5203 27035 5206
rect 13997 5130 14063 5133
rect 24117 5130 24183 5133
rect 13997 5128 24183 5130
rect 13997 5072 14002 5128
rect 14058 5072 24122 5128
rect 24178 5072 24183 5128
rect 13997 5070 24183 5072
rect 13997 5067 14063 5070
rect 24117 5067 24183 5070
rect 24485 5130 24551 5133
rect 26550 5130 26556 5132
rect 24485 5128 26556 5130
rect 24485 5072 24490 5128
rect 24546 5072 26556 5128
rect 24485 5070 26556 5072
rect 24485 5067 24551 5070
rect 26550 5068 26556 5070
rect 26620 5068 26626 5132
rect 32213 5130 32279 5133
rect 26742 5128 32279 5130
rect 26742 5072 32218 5128
rect 32274 5072 32279 5128
rect 26742 5070 32279 5072
rect 22461 4994 22527 4997
rect 19014 4992 22527 4994
rect 19014 4936 22466 4992
rect 22522 4936 22527 4992
rect 19014 4934 22527 4936
rect 3566 4928 3882 4929
rect 3566 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3812 4928
rect 3876 4864 3882 4928
rect 3566 4863 3882 4864
rect 8566 4928 8882 4929
rect 8566 4864 8572 4928
rect 8636 4864 8652 4928
rect 8716 4864 8732 4928
rect 8796 4864 8812 4928
rect 8876 4864 8882 4928
rect 8566 4863 8882 4864
rect 13566 4928 13882 4929
rect 13566 4864 13572 4928
rect 13636 4864 13652 4928
rect 13716 4864 13732 4928
rect 13796 4864 13812 4928
rect 13876 4864 13882 4928
rect 13566 4863 13882 4864
rect 18566 4928 18882 4929
rect 18566 4864 18572 4928
rect 18636 4864 18652 4928
rect 18716 4864 18732 4928
rect 18796 4864 18812 4928
rect 18876 4864 18882 4928
rect 18566 4863 18882 4864
rect 5441 4722 5507 4725
rect 16481 4722 16547 4725
rect 19014 4722 19074 4934
rect 22461 4931 22527 4934
rect 24577 4994 24643 4997
rect 26742 4994 26802 5070
rect 32213 5067 32279 5070
rect 24577 4992 26802 4994
rect 24577 4936 24582 4992
rect 24638 4936 26802 4992
rect 24577 4934 26802 4936
rect 24577 4931 24643 4934
rect 23566 4928 23882 4929
rect 23566 4864 23572 4928
rect 23636 4864 23652 4928
rect 23716 4864 23732 4928
rect 23796 4864 23812 4928
rect 23876 4864 23882 4928
rect 23566 4863 23882 4864
rect 28566 4928 28882 4929
rect 28566 4864 28572 4928
rect 28636 4864 28652 4928
rect 28716 4864 28732 4928
rect 28796 4864 28812 4928
rect 28876 4864 28882 4928
rect 28566 4863 28882 4864
rect 33566 4928 33882 4929
rect 33566 4864 33572 4928
rect 33636 4864 33652 4928
rect 33716 4864 33732 4928
rect 33796 4864 33812 4928
rect 33876 4864 33882 4928
rect 33566 4863 33882 4864
rect 19609 4858 19675 4861
rect 22737 4858 22803 4861
rect 19609 4856 22803 4858
rect 19609 4800 19614 4856
rect 19670 4800 22742 4856
rect 22798 4800 22803 4856
rect 19609 4798 22803 4800
rect 19609 4795 19675 4798
rect 22737 4795 22803 4798
rect 26049 4858 26115 4861
rect 27153 4858 27219 4861
rect 26049 4856 27219 4858
rect 26049 4800 26054 4856
rect 26110 4800 27158 4856
rect 27214 4800 27219 4856
rect 26049 4798 27219 4800
rect 26049 4795 26115 4798
rect 27153 4795 27219 4798
rect 33961 4858 34027 4861
rect 34102 4858 34162 5206
rect 38566 4928 38882 4929
rect 38566 4864 38572 4928
rect 38636 4864 38652 4928
rect 38716 4864 38732 4928
rect 38796 4864 38812 4928
rect 38876 4864 38882 4928
rect 38566 4863 38882 4864
rect 43566 4928 43882 4929
rect 43566 4864 43572 4928
rect 43636 4864 43652 4928
rect 43716 4864 43732 4928
rect 43796 4864 43812 4928
rect 43876 4864 43882 4928
rect 43566 4863 43882 4864
rect 38377 4858 38443 4861
rect 33961 4856 38443 4858
rect 33961 4800 33966 4856
rect 34022 4800 38382 4856
rect 38438 4800 38443 4856
rect 33961 4798 38443 4800
rect 33961 4795 34027 4798
rect 38377 4795 38443 4798
rect 5441 4720 19074 4722
rect 5441 4664 5446 4720
rect 5502 4664 16486 4720
rect 16542 4664 19074 4720
rect 5441 4662 19074 4664
rect 19885 4722 19951 4725
rect 19885 4720 22570 4722
rect 19885 4664 19890 4720
rect 19946 4664 22570 4720
rect 19885 4662 22570 4664
rect 5441 4659 5507 4662
rect 16481 4659 16547 4662
rect 19885 4659 19951 4662
rect 3509 4586 3575 4589
rect 16389 4586 16455 4589
rect 21449 4586 21515 4589
rect 3509 4584 21515 4586
rect 3509 4528 3514 4584
rect 3570 4528 16394 4584
rect 16450 4528 21454 4584
rect 21510 4528 21515 4584
rect 3509 4526 21515 4528
rect 22510 4586 22570 4662
rect 22686 4660 22692 4724
rect 22756 4722 22762 4724
rect 22921 4722 22987 4725
rect 27654 4722 27660 4724
rect 22756 4720 27660 4722
rect 22756 4664 22926 4720
rect 22982 4664 27660 4720
rect 22756 4662 27660 4664
rect 22756 4660 22762 4662
rect 22921 4659 22987 4662
rect 27654 4660 27660 4662
rect 27724 4660 27730 4724
rect 28441 4722 28507 4725
rect 41965 4722 42031 4725
rect 28441 4720 42031 4722
rect 28441 4664 28446 4720
rect 28502 4664 41970 4720
rect 42026 4664 42031 4720
rect 28441 4662 42031 4664
rect 28441 4659 28507 4662
rect 41965 4659 42031 4662
rect 23289 4586 23355 4589
rect 22510 4584 23355 4586
rect 22510 4528 23294 4584
rect 23350 4528 23355 4584
rect 22510 4526 23355 4528
rect 3509 4523 3575 4526
rect 16389 4523 16455 4526
rect 21449 4523 21515 4526
rect 23289 4523 23355 4526
rect 25037 4586 25103 4589
rect 28717 4586 28783 4589
rect 25037 4584 28783 4586
rect 25037 4528 25042 4584
rect 25098 4528 28722 4584
rect 28778 4528 28783 4584
rect 25037 4526 28783 4528
rect 25037 4523 25103 4526
rect 28717 4523 28783 4526
rect 30005 4586 30071 4589
rect 37733 4586 37799 4589
rect 30005 4584 37799 4586
rect 30005 4528 30010 4584
rect 30066 4528 37738 4584
rect 37794 4528 37799 4584
rect 30005 4526 37799 4528
rect 30005 4523 30071 4526
rect 37733 4523 37799 4526
rect 22277 4450 22343 4453
rect 24117 4450 24183 4453
rect 22277 4448 24183 4450
rect 22277 4392 22282 4448
rect 22338 4392 24122 4448
rect 24178 4392 24183 4448
rect 22277 4390 24183 4392
rect 22277 4387 22343 4390
rect 24117 4387 24183 4390
rect 6066 4384 6382 4385
rect 6066 4320 6072 4384
rect 6136 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6382 4384
rect 6066 4319 6382 4320
rect 11066 4384 11382 4385
rect 11066 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11382 4384
rect 11066 4319 11382 4320
rect 16066 4384 16382 4385
rect 16066 4320 16072 4384
rect 16136 4320 16152 4384
rect 16216 4320 16232 4384
rect 16296 4320 16312 4384
rect 16376 4320 16382 4384
rect 16066 4319 16382 4320
rect 21066 4384 21382 4385
rect 21066 4320 21072 4384
rect 21136 4320 21152 4384
rect 21216 4320 21232 4384
rect 21296 4320 21312 4384
rect 21376 4320 21382 4384
rect 21066 4319 21382 4320
rect 26066 4384 26382 4385
rect 26066 4320 26072 4384
rect 26136 4320 26152 4384
rect 26216 4320 26232 4384
rect 26296 4320 26312 4384
rect 26376 4320 26382 4384
rect 26066 4319 26382 4320
rect 31066 4384 31382 4385
rect 31066 4320 31072 4384
rect 31136 4320 31152 4384
rect 31216 4320 31232 4384
rect 31296 4320 31312 4384
rect 31376 4320 31382 4384
rect 31066 4319 31382 4320
rect 36066 4384 36382 4385
rect 36066 4320 36072 4384
rect 36136 4320 36152 4384
rect 36216 4320 36232 4384
rect 36296 4320 36312 4384
rect 36376 4320 36382 4384
rect 36066 4319 36382 4320
rect 41066 4384 41382 4385
rect 41066 4320 41072 4384
rect 41136 4320 41152 4384
rect 41216 4320 41232 4384
rect 41296 4320 41312 4384
rect 41376 4320 41382 4384
rect 41066 4319 41382 4320
rect 29269 4314 29335 4317
rect 29269 4312 29378 4314
rect 29269 4256 29274 4312
rect 29330 4256 29378 4312
rect 29269 4251 29378 4256
rect 14825 4178 14891 4181
rect 23841 4178 23907 4181
rect 27429 4178 27495 4181
rect 14825 4176 23907 4178
rect 14825 4120 14830 4176
rect 14886 4120 23846 4176
rect 23902 4120 23907 4176
rect 14825 4118 23907 4120
rect 14825 4115 14891 4118
rect 23841 4115 23907 4118
rect 25684 4176 27495 4178
rect 25684 4120 27434 4176
rect 27490 4120 27495 4176
rect 25684 4118 27495 4120
rect 29318 4178 29378 4251
rect 41505 4178 41571 4181
rect 29318 4176 41571 4178
rect 29318 4120 41510 4176
rect 41566 4120 41571 4176
rect 29318 4118 41571 4120
rect 19149 4044 19215 4045
rect 19149 4042 19196 4044
rect 19104 4040 19196 4042
rect 19104 3984 19154 4040
rect 19104 3982 19196 3984
rect 19149 3980 19196 3982
rect 19260 3980 19266 4044
rect 20345 4042 20411 4045
rect 21725 4042 21791 4045
rect 25221 4042 25287 4045
rect 25684 4042 25744 4118
rect 27429 4115 27495 4118
rect 41505 4115 41571 4118
rect 20345 4040 25744 4042
rect 20345 3984 20350 4040
rect 20406 3984 21730 4040
rect 21786 3984 25226 4040
rect 25282 3984 25744 4040
rect 20345 3982 25744 3984
rect 19149 3979 19215 3980
rect 20345 3979 20411 3982
rect 21725 3979 21791 3982
rect 25221 3979 25287 3982
rect 25814 3980 25820 4044
rect 25884 4042 25890 4044
rect 36813 4042 36879 4045
rect 25884 4040 36879 4042
rect 25884 3984 36818 4040
rect 36874 3984 36879 4040
rect 25884 3982 36879 3984
rect 25884 3980 25890 3982
rect 36813 3979 36879 3982
rect 3566 3840 3882 3841
rect 3566 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3812 3840
rect 3876 3776 3882 3840
rect 3566 3775 3882 3776
rect 8566 3840 8882 3841
rect 8566 3776 8572 3840
rect 8636 3776 8652 3840
rect 8716 3776 8732 3840
rect 8796 3776 8812 3840
rect 8876 3776 8882 3840
rect 8566 3775 8882 3776
rect 13566 3840 13882 3841
rect 13566 3776 13572 3840
rect 13636 3776 13652 3840
rect 13716 3776 13732 3840
rect 13796 3776 13812 3840
rect 13876 3776 13882 3840
rect 13566 3775 13882 3776
rect 18566 3840 18882 3841
rect 18566 3776 18572 3840
rect 18636 3776 18652 3840
rect 18716 3776 18732 3840
rect 18796 3776 18812 3840
rect 18876 3776 18882 3840
rect 18566 3775 18882 3776
rect 23566 3840 23882 3841
rect 23566 3776 23572 3840
rect 23636 3776 23652 3840
rect 23716 3776 23732 3840
rect 23796 3776 23812 3840
rect 23876 3776 23882 3840
rect 23566 3775 23882 3776
rect 28566 3840 28882 3841
rect 28566 3776 28572 3840
rect 28636 3776 28652 3840
rect 28716 3776 28732 3840
rect 28796 3776 28812 3840
rect 28876 3776 28882 3840
rect 28566 3775 28882 3776
rect 33566 3840 33882 3841
rect 33566 3776 33572 3840
rect 33636 3776 33652 3840
rect 33716 3776 33732 3840
rect 33796 3776 33812 3840
rect 33876 3776 33882 3840
rect 33566 3775 33882 3776
rect 38566 3840 38882 3841
rect 38566 3776 38572 3840
rect 38636 3776 38652 3840
rect 38716 3776 38732 3840
rect 38796 3776 38812 3840
rect 38876 3776 38882 3840
rect 38566 3775 38882 3776
rect 43566 3840 43882 3841
rect 43566 3776 43572 3840
rect 43636 3776 43652 3840
rect 43716 3776 43732 3840
rect 43796 3776 43812 3840
rect 43876 3776 43882 3840
rect 43566 3775 43882 3776
rect 21725 3770 21791 3773
rect 23381 3770 23447 3773
rect 21725 3768 23447 3770
rect 21725 3712 21730 3768
rect 21786 3712 23386 3768
rect 23442 3712 23447 3768
rect 21725 3710 23447 3712
rect 21725 3707 21791 3710
rect 23381 3707 23447 3710
rect 28950 3710 31770 3770
rect 10409 3634 10475 3637
rect 23381 3634 23447 3637
rect 10409 3632 23447 3634
rect 10409 3576 10414 3632
rect 10470 3576 23386 3632
rect 23442 3576 23447 3632
rect 10409 3574 23447 3576
rect 10409 3571 10475 3574
rect 23381 3571 23447 3574
rect 24301 3634 24367 3637
rect 28950 3634 29010 3710
rect 24301 3632 29010 3634
rect 24301 3576 24306 3632
rect 24362 3576 29010 3632
rect 24301 3574 29010 3576
rect 24301 3571 24367 3574
rect 29269 3498 29335 3501
rect 31293 3498 31359 3501
rect 29269 3496 31359 3498
rect 29269 3440 29274 3496
rect 29330 3440 31298 3496
rect 31354 3440 31359 3496
rect 29269 3438 31359 3440
rect 31710 3498 31770 3710
rect 31845 3634 31911 3637
rect 37917 3634 37983 3637
rect 31845 3632 37983 3634
rect 31845 3576 31850 3632
rect 31906 3576 37922 3632
rect 37978 3576 37983 3632
rect 31845 3574 37983 3576
rect 31845 3571 31911 3574
rect 37917 3571 37983 3574
rect 33685 3498 33751 3501
rect 31710 3496 33751 3498
rect 31710 3440 33690 3496
rect 33746 3440 33751 3496
rect 31710 3438 33751 3440
rect 29269 3435 29335 3438
rect 31293 3435 31359 3438
rect 33685 3435 33751 3438
rect 6066 3296 6382 3297
rect 6066 3232 6072 3296
rect 6136 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6382 3296
rect 6066 3231 6382 3232
rect 11066 3296 11382 3297
rect 11066 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11382 3296
rect 11066 3231 11382 3232
rect 16066 3296 16382 3297
rect 16066 3232 16072 3296
rect 16136 3232 16152 3296
rect 16216 3232 16232 3296
rect 16296 3232 16312 3296
rect 16376 3232 16382 3296
rect 16066 3231 16382 3232
rect 21066 3296 21382 3297
rect 21066 3232 21072 3296
rect 21136 3232 21152 3296
rect 21216 3232 21232 3296
rect 21296 3232 21312 3296
rect 21376 3232 21382 3296
rect 21066 3231 21382 3232
rect 26066 3296 26382 3297
rect 26066 3232 26072 3296
rect 26136 3232 26152 3296
rect 26216 3232 26232 3296
rect 26296 3232 26312 3296
rect 26376 3232 26382 3296
rect 26066 3231 26382 3232
rect 31066 3296 31382 3297
rect 31066 3232 31072 3296
rect 31136 3232 31152 3296
rect 31216 3232 31232 3296
rect 31296 3232 31312 3296
rect 31376 3232 31382 3296
rect 31066 3231 31382 3232
rect 36066 3296 36382 3297
rect 36066 3232 36072 3296
rect 36136 3232 36152 3296
rect 36216 3232 36232 3296
rect 36296 3232 36312 3296
rect 36376 3232 36382 3296
rect 36066 3231 36382 3232
rect 41066 3296 41382 3297
rect 41066 3232 41072 3296
rect 41136 3232 41152 3296
rect 41216 3232 41232 3296
rect 41296 3232 41312 3296
rect 41376 3232 41382 3296
rect 41066 3231 41382 3232
rect 19425 3226 19491 3229
rect 19290 3224 19491 3226
rect 19290 3168 19430 3224
rect 19486 3168 19491 3224
rect 19290 3166 19491 3168
rect 11329 3090 11395 3093
rect 19290 3090 19350 3166
rect 19425 3163 19491 3166
rect 28809 3226 28875 3229
rect 30281 3226 30347 3229
rect 28809 3224 30347 3226
rect 28809 3168 28814 3224
rect 28870 3168 30286 3224
rect 30342 3168 30347 3224
rect 28809 3166 30347 3168
rect 28809 3163 28875 3166
rect 30281 3163 30347 3166
rect 38009 3226 38075 3229
rect 39982 3226 39988 3228
rect 38009 3224 39988 3226
rect 38009 3168 38014 3224
rect 38070 3168 39988 3224
rect 38009 3166 39988 3168
rect 38009 3163 38075 3166
rect 39982 3164 39988 3166
rect 40052 3164 40058 3228
rect 11329 3088 19350 3090
rect 11329 3032 11334 3088
rect 11390 3032 19350 3088
rect 11329 3030 19350 3032
rect 21173 3090 21239 3093
rect 25129 3090 25195 3093
rect 21173 3088 25195 3090
rect 21173 3032 21178 3088
rect 21234 3032 25134 3088
rect 25190 3032 25195 3088
rect 21173 3030 25195 3032
rect 11329 3027 11395 3030
rect 21173 3027 21239 3030
rect 25129 3027 25195 3030
rect 28257 3090 28323 3093
rect 28942 3090 28948 3092
rect 28257 3088 28948 3090
rect 28257 3032 28262 3088
rect 28318 3032 28948 3088
rect 28257 3030 28948 3032
rect 28257 3027 28323 3030
rect 28942 3028 28948 3030
rect 29012 3028 29018 3092
rect 36721 3090 36787 3093
rect 40677 3090 40743 3093
rect 36721 3088 40743 3090
rect 36721 3032 36726 3088
rect 36782 3032 40682 3088
rect 40738 3032 40743 3088
rect 36721 3030 40743 3032
rect 36721 3027 36787 3030
rect 40677 3027 40743 3030
rect 8293 2954 8359 2957
rect 16389 2954 16455 2957
rect 16982 2954 16988 2956
rect 8293 2952 16988 2954
rect 8293 2896 8298 2952
rect 8354 2896 16394 2952
rect 16450 2896 16988 2952
rect 8293 2894 16988 2896
rect 8293 2891 8359 2894
rect 16389 2891 16455 2894
rect 16982 2892 16988 2894
rect 17052 2892 17058 2956
rect 28349 2954 28415 2957
rect 30373 2954 30439 2957
rect 28349 2952 30439 2954
rect 28349 2896 28354 2952
rect 28410 2896 30378 2952
rect 30434 2896 30439 2952
rect 28349 2894 30439 2896
rect 28349 2891 28415 2894
rect 30373 2891 30439 2894
rect 32581 2954 32647 2957
rect 37641 2954 37707 2957
rect 32581 2952 37707 2954
rect 32581 2896 32586 2952
rect 32642 2896 37646 2952
rect 37702 2896 37707 2952
rect 32581 2894 37707 2896
rect 32581 2891 32647 2894
rect 37641 2891 37707 2894
rect -300 2818 160 2848
rect 749 2818 815 2821
rect -300 2816 815 2818
rect -300 2760 754 2816
rect 810 2760 815 2816
rect -300 2758 815 2760
rect -300 2728 160 2758
rect 749 2755 815 2758
rect 35249 2818 35315 2821
rect 35893 2818 35959 2821
rect 35249 2816 35959 2818
rect 35249 2760 35254 2816
rect 35310 2760 35898 2816
rect 35954 2760 35959 2816
rect 35249 2758 35959 2760
rect 35249 2755 35315 2758
rect 35893 2755 35959 2758
rect 44633 2818 44699 2821
rect 45840 2818 46300 2848
rect 44633 2816 46300 2818
rect 44633 2760 44638 2816
rect 44694 2760 46300 2816
rect 44633 2758 46300 2760
rect 44633 2755 44699 2758
rect 3566 2752 3882 2753
rect 3566 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3812 2752
rect 3876 2688 3882 2752
rect 3566 2687 3882 2688
rect 8566 2752 8882 2753
rect 8566 2688 8572 2752
rect 8636 2688 8652 2752
rect 8716 2688 8732 2752
rect 8796 2688 8812 2752
rect 8876 2688 8882 2752
rect 8566 2687 8882 2688
rect 13566 2752 13882 2753
rect 13566 2688 13572 2752
rect 13636 2688 13652 2752
rect 13716 2688 13732 2752
rect 13796 2688 13812 2752
rect 13876 2688 13882 2752
rect 13566 2687 13882 2688
rect 18566 2752 18882 2753
rect 18566 2688 18572 2752
rect 18636 2688 18652 2752
rect 18716 2688 18732 2752
rect 18796 2688 18812 2752
rect 18876 2688 18882 2752
rect 18566 2687 18882 2688
rect 23566 2752 23882 2753
rect 23566 2688 23572 2752
rect 23636 2688 23652 2752
rect 23716 2688 23732 2752
rect 23796 2688 23812 2752
rect 23876 2688 23882 2752
rect 23566 2687 23882 2688
rect 28566 2752 28882 2753
rect 28566 2688 28572 2752
rect 28636 2688 28652 2752
rect 28716 2688 28732 2752
rect 28796 2688 28812 2752
rect 28876 2688 28882 2752
rect 28566 2687 28882 2688
rect 33566 2752 33882 2753
rect 33566 2688 33572 2752
rect 33636 2688 33652 2752
rect 33716 2688 33732 2752
rect 33796 2688 33812 2752
rect 33876 2688 33882 2752
rect 33566 2687 33882 2688
rect 38566 2752 38882 2753
rect 38566 2688 38572 2752
rect 38636 2688 38652 2752
rect 38716 2688 38732 2752
rect 38796 2688 38812 2752
rect 38876 2688 38882 2752
rect 38566 2687 38882 2688
rect 43566 2752 43882 2753
rect 43566 2688 43572 2752
rect 43636 2688 43652 2752
rect 43716 2688 43732 2752
rect 43796 2688 43812 2752
rect 43876 2688 43882 2752
rect 45840 2728 46300 2758
rect 43566 2687 43882 2688
rect 31201 2682 31267 2685
rect 31937 2682 32003 2685
rect 32489 2682 32555 2685
rect 31201 2680 32555 2682
rect 31201 2624 31206 2680
rect 31262 2624 31942 2680
rect 31998 2624 32494 2680
rect 32550 2624 32555 2680
rect 31201 2622 32555 2624
rect 31201 2619 31267 2622
rect 31937 2619 32003 2622
rect 32489 2619 32555 2622
rect 35709 2682 35775 2685
rect 38285 2682 38351 2685
rect 35709 2680 38351 2682
rect 35709 2624 35714 2680
rect 35770 2624 38290 2680
rect 38346 2624 38351 2680
rect 35709 2622 38351 2624
rect 35709 2619 35775 2622
rect 38285 2619 38351 2622
rect 27705 2546 27771 2549
rect 41505 2546 41571 2549
rect 27705 2544 41571 2546
rect 27705 2488 27710 2544
rect 27766 2488 41510 2544
rect 41566 2488 41571 2544
rect 27705 2486 41571 2488
rect 27705 2483 27771 2486
rect 41505 2483 41571 2486
rect 19241 2410 19307 2413
rect 22686 2410 22692 2412
rect 19241 2408 22692 2410
rect 19241 2352 19246 2408
rect 19302 2352 22692 2408
rect 19241 2350 22692 2352
rect 19241 2347 19307 2350
rect 22686 2348 22692 2350
rect 22756 2348 22762 2412
rect 31385 2410 31451 2413
rect 32029 2410 32095 2413
rect 31385 2408 32095 2410
rect 31385 2352 31390 2408
rect 31446 2352 32034 2408
rect 32090 2352 32095 2408
rect 31385 2350 32095 2352
rect 31385 2347 31451 2350
rect 32029 2347 32095 2350
rect 32765 2410 32831 2413
rect 40861 2410 40927 2413
rect 32765 2408 40927 2410
rect 32765 2352 32770 2408
rect 32826 2352 40866 2408
rect 40922 2352 40927 2408
rect 32765 2350 40927 2352
rect 32765 2347 32831 2350
rect 40861 2347 40927 2350
rect 6066 2208 6382 2209
rect 6066 2144 6072 2208
rect 6136 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6382 2208
rect 6066 2143 6382 2144
rect 11066 2208 11382 2209
rect 11066 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11382 2208
rect 11066 2143 11382 2144
rect 16066 2208 16382 2209
rect 16066 2144 16072 2208
rect 16136 2144 16152 2208
rect 16216 2144 16232 2208
rect 16296 2144 16312 2208
rect 16376 2144 16382 2208
rect 16066 2143 16382 2144
rect 21066 2208 21382 2209
rect 21066 2144 21072 2208
rect 21136 2144 21152 2208
rect 21216 2144 21232 2208
rect 21296 2144 21312 2208
rect 21376 2144 21382 2208
rect 21066 2143 21382 2144
rect 26066 2208 26382 2209
rect 26066 2144 26072 2208
rect 26136 2144 26152 2208
rect 26216 2144 26232 2208
rect 26296 2144 26312 2208
rect 26376 2144 26382 2208
rect 26066 2143 26382 2144
rect 31066 2208 31382 2209
rect 31066 2144 31072 2208
rect 31136 2144 31152 2208
rect 31216 2144 31232 2208
rect 31296 2144 31312 2208
rect 31376 2144 31382 2208
rect 31066 2143 31382 2144
rect 36066 2208 36382 2209
rect 36066 2144 36072 2208
rect 36136 2144 36152 2208
rect 36216 2144 36232 2208
rect 36296 2144 36312 2208
rect 36376 2144 36382 2208
rect 36066 2143 36382 2144
rect 41066 2208 41382 2209
rect 41066 2144 41072 2208
rect 41136 2144 41152 2208
rect 41216 2144 41232 2208
rect 41296 2144 41312 2208
rect 41376 2144 41382 2208
rect 41066 2143 41382 2144
rect 26877 2138 26943 2141
rect 28073 2138 28139 2141
rect 26877 2136 28139 2138
rect 26877 2080 26882 2136
rect 26938 2080 28078 2136
rect 28134 2080 28139 2136
rect 26877 2078 28139 2080
rect 26877 2075 26943 2078
rect 28073 2075 28139 2078
rect 21541 2004 21607 2005
rect 21541 2000 21588 2004
rect 21652 2002 21658 2004
rect 31937 2002 32003 2005
rect 33777 2002 33843 2005
rect 21541 1944 21546 2000
rect 21541 1940 21588 1944
rect 21652 1942 21698 2002
rect 31937 2000 33843 2002
rect 31937 1944 31942 2000
rect 31998 1944 33782 2000
rect 33838 1944 33843 2000
rect 31937 1942 33843 1944
rect 21652 1940 21658 1942
rect 21541 1939 21607 1940
rect 31937 1939 32003 1942
rect 33777 1939 33843 1942
rect 3566 1664 3882 1665
rect 3566 1600 3572 1664
rect 3636 1600 3652 1664
rect 3716 1600 3732 1664
rect 3796 1600 3812 1664
rect 3876 1600 3882 1664
rect 3566 1599 3882 1600
rect 8566 1664 8882 1665
rect 8566 1600 8572 1664
rect 8636 1600 8652 1664
rect 8716 1600 8732 1664
rect 8796 1600 8812 1664
rect 8876 1600 8882 1664
rect 8566 1599 8882 1600
rect 13566 1664 13882 1665
rect 13566 1600 13572 1664
rect 13636 1600 13652 1664
rect 13716 1600 13732 1664
rect 13796 1600 13812 1664
rect 13876 1600 13882 1664
rect 13566 1599 13882 1600
rect 18566 1664 18882 1665
rect 18566 1600 18572 1664
rect 18636 1600 18652 1664
rect 18716 1600 18732 1664
rect 18796 1600 18812 1664
rect 18876 1600 18882 1664
rect 18566 1599 18882 1600
rect 23566 1664 23882 1665
rect 23566 1600 23572 1664
rect 23636 1600 23652 1664
rect 23716 1600 23732 1664
rect 23796 1600 23812 1664
rect 23876 1600 23882 1664
rect 23566 1599 23882 1600
rect 28566 1664 28882 1665
rect 28566 1600 28572 1664
rect 28636 1600 28652 1664
rect 28716 1600 28732 1664
rect 28796 1600 28812 1664
rect 28876 1600 28882 1664
rect 28566 1599 28882 1600
rect 33566 1664 33882 1665
rect 33566 1600 33572 1664
rect 33636 1600 33652 1664
rect 33716 1600 33732 1664
rect 33796 1600 33812 1664
rect 33876 1600 33882 1664
rect 33566 1599 33882 1600
rect 38566 1664 38882 1665
rect 38566 1600 38572 1664
rect 38636 1600 38652 1664
rect 38716 1600 38732 1664
rect 38796 1600 38812 1664
rect 38876 1600 38882 1664
rect 38566 1599 38882 1600
rect 43566 1664 43882 1665
rect 43566 1600 43572 1664
rect 43636 1600 43652 1664
rect 43716 1600 43732 1664
rect 43796 1600 43812 1664
rect 43876 1600 43882 1664
rect 43566 1599 43882 1600
rect 30465 1458 30531 1461
rect 36077 1458 36143 1461
rect 30465 1456 36143 1458
rect 30465 1400 30470 1456
rect 30526 1400 36082 1456
rect 36138 1400 36143 1456
rect 30465 1398 36143 1400
rect 30465 1395 30531 1398
rect 36077 1395 36143 1398
rect 28942 1260 28948 1324
rect 29012 1322 29018 1324
rect 33869 1322 33935 1325
rect 29012 1320 33935 1322
rect 29012 1264 33874 1320
rect 33930 1264 33935 1320
rect 29012 1262 33935 1264
rect 29012 1260 29018 1262
rect 33869 1259 33935 1262
rect 34278 1260 34284 1324
rect 34348 1322 34354 1324
rect 36169 1322 36235 1325
rect 34348 1320 36235 1322
rect 34348 1264 36174 1320
rect 36230 1264 36235 1320
rect 34348 1262 36235 1264
rect 34348 1260 34354 1262
rect 36169 1259 36235 1262
rect 39982 1260 39988 1324
rect 40052 1322 40058 1324
rect 40493 1322 40559 1325
rect 40052 1320 40559 1322
rect 40052 1264 40498 1320
rect 40554 1264 40559 1320
rect 40052 1262 40559 1264
rect 40052 1260 40058 1262
rect 40493 1259 40559 1262
rect 34462 1124 34468 1188
rect 34532 1186 34538 1188
rect 35893 1186 35959 1189
rect 34532 1184 35959 1186
rect 34532 1128 35898 1184
rect 35954 1128 35959 1184
rect 34532 1126 35959 1128
rect 34532 1124 34538 1126
rect 35893 1123 35959 1126
rect 6066 1120 6382 1121
rect 6066 1056 6072 1120
rect 6136 1056 6152 1120
rect 6216 1056 6232 1120
rect 6296 1056 6312 1120
rect 6376 1056 6382 1120
rect 6066 1055 6382 1056
rect 11066 1120 11382 1121
rect 11066 1056 11072 1120
rect 11136 1056 11152 1120
rect 11216 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11382 1120
rect 11066 1055 11382 1056
rect 16066 1120 16382 1121
rect 16066 1056 16072 1120
rect 16136 1056 16152 1120
rect 16216 1056 16232 1120
rect 16296 1056 16312 1120
rect 16376 1056 16382 1120
rect 16066 1055 16382 1056
rect 21066 1120 21382 1121
rect 21066 1056 21072 1120
rect 21136 1056 21152 1120
rect 21216 1056 21232 1120
rect 21296 1056 21312 1120
rect 21376 1056 21382 1120
rect 21066 1055 21382 1056
rect 26066 1120 26382 1121
rect 26066 1056 26072 1120
rect 26136 1056 26152 1120
rect 26216 1056 26232 1120
rect 26296 1056 26312 1120
rect 26376 1056 26382 1120
rect 26066 1055 26382 1056
rect 31066 1120 31382 1121
rect 31066 1056 31072 1120
rect 31136 1056 31152 1120
rect 31216 1056 31232 1120
rect 31296 1056 31312 1120
rect 31376 1056 31382 1120
rect 31066 1055 31382 1056
rect 36066 1120 36382 1121
rect 36066 1056 36072 1120
rect 36136 1056 36152 1120
rect 36216 1056 36232 1120
rect 36296 1056 36312 1120
rect 36376 1056 36382 1120
rect 36066 1055 36382 1056
rect 41066 1120 41382 1121
rect 41066 1056 41072 1120
rect 41136 1056 41152 1120
rect 41216 1056 41232 1120
rect 41296 1056 41312 1120
rect 41376 1056 41382 1120
rect 41066 1055 41382 1056
<< via3 >>
rect 6072 22876 6136 22880
rect 6072 22820 6076 22876
rect 6076 22820 6132 22876
rect 6132 22820 6136 22876
rect 6072 22816 6136 22820
rect 6152 22876 6216 22880
rect 6152 22820 6156 22876
rect 6156 22820 6212 22876
rect 6212 22820 6216 22876
rect 6152 22816 6216 22820
rect 6232 22876 6296 22880
rect 6232 22820 6236 22876
rect 6236 22820 6292 22876
rect 6292 22820 6296 22876
rect 6232 22816 6296 22820
rect 6312 22876 6376 22880
rect 6312 22820 6316 22876
rect 6316 22820 6372 22876
rect 6372 22820 6376 22876
rect 6312 22816 6376 22820
rect 11072 22876 11136 22880
rect 11072 22820 11076 22876
rect 11076 22820 11132 22876
rect 11132 22820 11136 22876
rect 11072 22816 11136 22820
rect 11152 22876 11216 22880
rect 11152 22820 11156 22876
rect 11156 22820 11212 22876
rect 11212 22820 11216 22876
rect 11152 22816 11216 22820
rect 11232 22876 11296 22880
rect 11232 22820 11236 22876
rect 11236 22820 11292 22876
rect 11292 22820 11296 22876
rect 11232 22816 11296 22820
rect 11312 22876 11376 22880
rect 11312 22820 11316 22876
rect 11316 22820 11372 22876
rect 11372 22820 11376 22876
rect 11312 22816 11376 22820
rect 16072 22876 16136 22880
rect 16072 22820 16076 22876
rect 16076 22820 16132 22876
rect 16132 22820 16136 22876
rect 16072 22816 16136 22820
rect 16152 22876 16216 22880
rect 16152 22820 16156 22876
rect 16156 22820 16212 22876
rect 16212 22820 16216 22876
rect 16152 22816 16216 22820
rect 16232 22876 16296 22880
rect 16232 22820 16236 22876
rect 16236 22820 16292 22876
rect 16292 22820 16296 22876
rect 16232 22816 16296 22820
rect 16312 22876 16376 22880
rect 16312 22820 16316 22876
rect 16316 22820 16372 22876
rect 16372 22820 16376 22876
rect 16312 22816 16376 22820
rect 21072 22876 21136 22880
rect 21072 22820 21076 22876
rect 21076 22820 21132 22876
rect 21132 22820 21136 22876
rect 21072 22816 21136 22820
rect 21152 22876 21216 22880
rect 21152 22820 21156 22876
rect 21156 22820 21212 22876
rect 21212 22820 21216 22876
rect 21152 22816 21216 22820
rect 21232 22876 21296 22880
rect 21232 22820 21236 22876
rect 21236 22820 21292 22876
rect 21292 22820 21296 22876
rect 21232 22816 21296 22820
rect 21312 22876 21376 22880
rect 21312 22820 21316 22876
rect 21316 22820 21372 22876
rect 21372 22820 21376 22876
rect 21312 22816 21376 22820
rect 26072 22876 26136 22880
rect 26072 22820 26076 22876
rect 26076 22820 26132 22876
rect 26132 22820 26136 22876
rect 26072 22816 26136 22820
rect 26152 22876 26216 22880
rect 26152 22820 26156 22876
rect 26156 22820 26212 22876
rect 26212 22820 26216 22876
rect 26152 22816 26216 22820
rect 26232 22876 26296 22880
rect 26232 22820 26236 22876
rect 26236 22820 26292 22876
rect 26292 22820 26296 22876
rect 26232 22816 26296 22820
rect 26312 22876 26376 22880
rect 26312 22820 26316 22876
rect 26316 22820 26372 22876
rect 26372 22820 26376 22876
rect 26312 22816 26376 22820
rect 31072 22876 31136 22880
rect 31072 22820 31076 22876
rect 31076 22820 31132 22876
rect 31132 22820 31136 22876
rect 31072 22816 31136 22820
rect 31152 22876 31216 22880
rect 31152 22820 31156 22876
rect 31156 22820 31212 22876
rect 31212 22820 31216 22876
rect 31152 22816 31216 22820
rect 31232 22876 31296 22880
rect 31232 22820 31236 22876
rect 31236 22820 31292 22876
rect 31292 22820 31296 22876
rect 31232 22816 31296 22820
rect 31312 22876 31376 22880
rect 31312 22820 31316 22876
rect 31316 22820 31372 22876
rect 31372 22820 31376 22876
rect 31312 22816 31376 22820
rect 36072 22876 36136 22880
rect 36072 22820 36076 22876
rect 36076 22820 36132 22876
rect 36132 22820 36136 22876
rect 36072 22816 36136 22820
rect 36152 22876 36216 22880
rect 36152 22820 36156 22876
rect 36156 22820 36212 22876
rect 36212 22820 36216 22876
rect 36152 22816 36216 22820
rect 36232 22876 36296 22880
rect 36232 22820 36236 22876
rect 36236 22820 36292 22876
rect 36292 22820 36296 22876
rect 36232 22816 36296 22820
rect 36312 22876 36376 22880
rect 36312 22820 36316 22876
rect 36316 22820 36372 22876
rect 36372 22820 36376 22876
rect 36312 22816 36376 22820
rect 41072 22876 41136 22880
rect 41072 22820 41076 22876
rect 41076 22820 41132 22876
rect 41132 22820 41136 22876
rect 41072 22816 41136 22820
rect 41152 22876 41216 22880
rect 41152 22820 41156 22876
rect 41156 22820 41212 22876
rect 41212 22820 41216 22876
rect 41152 22816 41216 22820
rect 41232 22876 41296 22880
rect 41232 22820 41236 22876
rect 41236 22820 41292 22876
rect 41292 22820 41296 22876
rect 41232 22816 41296 22820
rect 41312 22876 41376 22880
rect 41312 22820 41316 22876
rect 41316 22820 41372 22876
rect 41372 22820 41376 22876
rect 41312 22816 41376 22820
rect 19196 22476 19260 22540
rect 3572 22332 3636 22336
rect 3572 22276 3576 22332
rect 3576 22276 3632 22332
rect 3632 22276 3636 22332
rect 3572 22272 3636 22276
rect 3652 22332 3716 22336
rect 3652 22276 3656 22332
rect 3656 22276 3712 22332
rect 3712 22276 3716 22332
rect 3652 22272 3716 22276
rect 3732 22332 3796 22336
rect 3732 22276 3736 22332
rect 3736 22276 3792 22332
rect 3792 22276 3796 22332
rect 3732 22272 3796 22276
rect 3812 22332 3876 22336
rect 3812 22276 3816 22332
rect 3816 22276 3872 22332
rect 3872 22276 3876 22332
rect 3812 22272 3876 22276
rect 8572 22332 8636 22336
rect 8572 22276 8576 22332
rect 8576 22276 8632 22332
rect 8632 22276 8636 22332
rect 8572 22272 8636 22276
rect 8652 22332 8716 22336
rect 8652 22276 8656 22332
rect 8656 22276 8712 22332
rect 8712 22276 8716 22332
rect 8652 22272 8716 22276
rect 8732 22332 8796 22336
rect 8732 22276 8736 22332
rect 8736 22276 8792 22332
rect 8792 22276 8796 22332
rect 8732 22272 8796 22276
rect 8812 22332 8876 22336
rect 8812 22276 8816 22332
rect 8816 22276 8872 22332
rect 8872 22276 8876 22332
rect 8812 22272 8876 22276
rect 13572 22332 13636 22336
rect 13572 22276 13576 22332
rect 13576 22276 13632 22332
rect 13632 22276 13636 22332
rect 13572 22272 13636 22276
rect 13652 22332 13716 22336
rect 13652 22276 13656 22332
rect 13656 22276 13712 22332
rect 13712 22276 13716 22332
rect 13652 22272 13716 22276
rect 13732 22332 13796 22336
rect 13732 22276 13736 22332
rect 13736 22276 13792 22332
rect 13792 22276 13796 22332
rect 13732 22272 13796 22276
rect 13812 22332 13876 22336
rect 13812 22276 13816 22332
rect 13816 22276 13872 22332
rect 13872 22276 13876 22332
rect 13812 22272 13876 22276
rect 18572 22332 18636 22336
rect 18572 22276 18576 22332
rect 18576 22276 18632 22332
rect 18632 22276 18636 22332
rect 18572 22272 18636 22276
rect 18652 22332 18716 22336
rect 18652 22276 18656 22332
rect 18656 22276 18712 22332
rect 18712 22276 18716 22332
rect 18652 22272 18716 22276
rect 18732 22332 18796 22336
rect 18732 22276 18736 22332
rect 18736 22276 18792 22332
rect 18792 22276 18796 22332
rect 18732 22272 18796 22276
rect 18812 22332 18876 22336
rect 18812 22276 18816 22332
rect 18816 22276 18872 22332
rect 18872 22276 18876 22332
rect 18812 22272 18876 22276
rect 23572 22332 23636 22336
rect 23572 22276 23576 22332
rect 23576 22276 23632 22332
rect 23632 22276 23636 22332
rect 23572 22272 23636 22276
rect 23652 22332 23716 22336
rect 23652 22276 23656 22332
rect 23656 22276 23712 22332
rect 23712 22276 23716 22332
rect 23652 22272 23716 22276
rect 23732 22332 23796 22336
rect 23732 22276 23736 22332
rect 23736 22276 23792 22332
rect 23792 22276 23796 22332
rect 23732 22272 23796 22276
rect 23812 22332 23876 22336
rect 23812 22276 23816 22332
rect 23816 22276 23872 22332
rect 23872 22276 23876 22332
rect 23812 22272 23876 22276
rect 28572 22332 28636 22336
rect 28572 22276 28576 22332
rect 28576 22276 28632 22332
rect 28632 22276 28636 22332
rect 28572 22272 28636 22276
rect 28652 22332 28716 22336
rect 28652 22276 28656 22332
rect 28656 22276 28712 22332
rect 28712 22276 28716 22332
rect 28652 22272 28716 22276
rect 28732 22332 28796 22336
rect 28732 22276 28736 22332
rect 28736 22276 28792 22332
rect 28792 22276 28796 22332
rect 28732 22272 28796 22276
rect 28812 22332 28876 22336
rect 28812 22276 28816 22332
rect 28816 22276 28872 22332
rect 28872 22276 28876 22332
rect 28812 22272 28876 22276
rect 33572 22332 33636 22336
rect 33572 22276 33576 22332
rect 33576 22276 33632 22332
rect 33632 22276 33636 22332
rect 33572 22272 33636 22276
rect 33652 22332 33716 22336
rect 33652 22276 33656 22332
rect 33656 22276 33712 22332
rect 33712 22276 33716 22332
rect 33652 22272 33716 22276
rect 33732 22332 33796 22336
rect 33732 22276 33736 22332
rect 33736 22276 33792 22332
rect 33792 22276 33796 22332
rect 33732 22272 33796 22276
rect 33812 22332 33876 22336
rect 33812 22276 33816 22332
rect 33816 22276 33872 22332
rect 33872 22276 33876 22332
rect 33812 22272 33876 22276
rect 38572 22332 38636 22336
rect 38572 22276 38576 22332
rect 38576 22276 38632 22332
rect 38632 22276 38636 22332
rect 38572 22272 38636 22276
rect 38652 22332 38716 22336
rect 38652 22276 38656 22332
rect 38656 22276 38712 22332
rect 38712 22276 38716 22332
rect 38652 22272 38716 22276
rect 38732 22332 38796 22336
rect 38732 22276 38736 22332
rect 38736 22276 38792 22332
rect 38792 22276 38796 22332
rect 38732 22272 38796 22276
rect 38812 22332 38876 22336
rect 38812 22276 38816 22332
rect 38816 22276 38872 22332
rect 38872 22276 38876 22332
rect 38812 22272 38876 22276
rect 43572 22332 43636 22336
rect 43572 22276 43576 22332
rect 43576 22276 43632 22332
rect 43632 22276 43636 22332
rect 43572 22272 43636 22276
rect 43652 22332 43716 22336
rect 43652 22276 43656 22332
rect 43656 22276 43712 22332
rect 43712 22276 43716 22332
rect 43652 22272 43716 22276
rect 43732 22332 43796 22336
rect 43732 22276 43736 22332
rect 43736 22276 43792 22332
rect 43792 22276 43796 22332
rect 43732 22272 43796 22276
rect 43812 22332 43876 22336
rect 43812 22276 43816 22332
rect 43816 22276 43872 22332
rect 43872 22276 43876 22332
rect 43812 22272 43876 22276
rect 25820 22068 25884 22132
rect 28212 22068 28276 22132
rect 6072 21788 6136 21792
rect 6072 21732 6076 21788
rect 6076 21732 6132 21788
rect 6132 21732 6136 21788
rect 6072 21728 6136 21732
rect 6152 21788 6216 21792
rect 6152 21732 6156 21788
rect 6156 21732 6212 21788
rect 6212 21732 6216 21788
rect 6152 21728 6216 21732
rect 6232 21788 6296 21792
rect 6232 21732 6236 21788
rect 6236 21732 6292 21788
rect 6292 21732 6296 21788
rect 6232 21728 6296 21732
rect 6312 21788 6376 21792
rect 6312 21732 6316 21788
rect 6316 21732 6372 21788
rect 6372 21732 6376 21788
rect 6312 21728 6376 21732
rect 11072 21788 11136 21792
rect 11072 21732 11076 21788
rect 11076 21732 11132 21788
rect 11132 21732 11136 21788
rect 11072 21728 11136 21732
rect 11152 21788 11216 21792
rect 11152 21732 11156 21788
rect 11156 21732 11212 21788
rect 11212 21732 11216 21788
rect 11152 21728 11216 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 16072 21788 16136 21792
rect 16072 21732 16076 21788
rect 16076 21732 16132 21788
rect 16132 21732 16136 21788
rect 16072 21728 16136 21732
rect 16152 21788 16216 21792
rect 16152 21732 16156 21788
rect 16156 21732 16212 21788
rect 16212 21732 16216 21788
rect 16152 21728 16216 21732
rect 16232 21788 16296 21792
rect 16232 21732 16236 21788
rect 16236 21732 16292 21788
rect 16292 21732 16296 21788
rect 16232 21728 16296 21732
rect 16312 21788 16376 21792
rect 16312 21732 16316 21788
rect 16316 21732 16372 21788
rect 16372 21732 16376 21788
rect 16312 21728 16376 21732
rect 21072 21788 21136 21792
rect 21072 21732 21076 21788
rect 21076 21732 21132 21788
rect 21132 21732 21136 21788
rect 21072 21728 21136 21732
rect 21152 21788 21216 21792
rect 21152 21732 21156 21788
rect 21156 21732 21212 21788
rect 21212 21732 21216 21788
rect 21152 21728 21216 21732
rect 21232 21788 21296 21792
rect 21232 21732 21236 21788
rect 21236 21732 21292 21788
rect 21292 21732 21296 21788
rect 21232 21728 21296 21732
rect 21312 21788 21376 21792
rect 21312 21732 21316 21788
rect 21316 21732 21372 21788
rect 21372 21732 21376 21788
rect 21312 21728 21376 21732
rect 19932 21660 19996 21724
rect 26072 21788 26136 21792
rect 26072 21732 26076 21788
rect 26076 21732 26132 21788
rect 26132 21732 26136 21788
rect 26072 21728 26136 21732
rect 26152 21788 26216 21792
rect 26152 21732 26156 21788
rect 26156 21732 26212 21788
rect 26212 21732 26216 21788
rect 26152 21728 26216 21732
rect 26232 21788 26296 21792
rect 26232 21732 26236 21788
rect 26236 21732 26292 21788
rect 26292 21732 26296 21788
rect 26232 21728 26296 21732
rect 26312 21788 26376 21792
rect 26312 21732 26316 21788
rect 26316 21732 26372 21788
rect 26372 21732 26376 21788
rect 26312 21728 26376 21732
rect 31072 21788 31136 21792
rect 31072 21732 31076 21788
rect 31076 21732 31132 21788
rect 31132 21732 31136 21788
rect 31072 21728 31136 21732
rect 31152 21788 31216 21792
rect 31152 21732 31156 21788
rect 31156 21732 31212 21788
rect 31212 21732 31216 21788
rect 31152 21728 31216 21732
rect 31232 21788 31296 21792
rect 31232 21732 31236 21788
rect 31236 21732 31292 21788
rect 31292 21732 31296 21788
rect 31232 21728 31296 21732
rect 31312 21788 31376 21792
rect 31312 21732 31316 21788
rect 31316 21732 31372 21788
rect 31372 21732 31376 21788
rect 31312 21728 31376 21732
rect 36072 21788 36136 21792
rect 36072 21732 36076 21788
rect 36076 21732 36132 21788
rect 36132 21732 36136 21788
rect 36072 21728 36136 21732
rect 36152 21788 36216 21792
rect 36152 21732 36156 21788
rect 36156 21732 36212 21788
rect 36212 21732 36216 21788
rect 36152 21728 36216 21732
rect 36232 21788 36296 21792
rect 36232 21732 36236 21788
rect 36236 21732 36292 21788
rect 36292 21732 36296 21788
rect 36232 21728 36296 21732
rect 36312 21788 36376 21792
rect 36312 21732 36316 21788
rect 36316 21732 36372 21788
rect 36372 21732 36376 21788
rect 36312 21728 36376 21732
rect 41072 21788 41136 21792
rect 41072 21732 41076 21788
rect 41076 21732 41132 21788
rect 41132 21732 41136 21788
rect 41072 21728 41136 21732
rect 41152 21788 41216 21792
rect 41152 21732 41156 21788
rect 41156 21732 41212 21788
rect 41212 21732 41216 21788
rect 41152 21728 41216 21732
rect 41232 21788 41296 21792
rect 41232 21732 41236 21788
rect 41236 21732 41292 21788
rect 41292 21732 41296 21788
rect 41232 21728 41296 21732
rect 41312 21788 41376 21792
rect 41312 21732 41316 21788
rect 41316 21732 41372 21788
rect 41372 21732 41376 21788
rect 41312 21728 41376 21732
rect 26740 21660 26804 21724
rect 3572 21244 3636 21248
rect 3572 21188 3576 21244
rect 3576 21188 3632 21244
rect 3632 21188 3636 21244
rect 3572 21184 3636 21188
rect 3652 21244 3716 21248
rect 3652 21188 3656 21244
rect 3656 21188 3712 21244
rect 3712 21188 3716 21244
rect 3652 21184 3716 21188
rect 3732 21244 3796 21248
rect 3732 21188 3736 21244
rect 3736 21188 3792 21244
rect 3792 21188 3796 21244
rect 3732 21184 3796 21188
rect 3812 21244 3876 21248
rect 3812 21188 3816 21244
rect 3816 21188 3872 21244
rect 3872 21188 3876 21244
rect 3812 21184 3876 21188
rect 8572 21244 8636 21248
rect 8572 21188 8576 21244
rect 8576 21188 8632 21244
rect 8632 21188 8636 21244
rect 8572 21184 8636 21188
rect 8652 21244 8716 21248
rect 8652 21188 8656 21244
rect 8656 21188 8712 21244
rect 8712 21188 8716 21244
rect 8652 21184 8716 21188
rect 8732 21244 8796 21248
rect 8732 21188 8736 21244
rect 8736 21188 8792 21244
rect 8792 21188 8796 21244
rect 8732 21184 8796 21188
rect 8812 21244 8876 21248
rect 8812 21188 8816 21244
rect 8816 21188 8872 21244
rect 8872 21188 8876 21244
rect 8812 21184 8876 21188
rect 13572 21244 13636 21248
rect 13572 21188 13576 21244
rect 13576 21188 13632 21244
rect 13632 21188 13636 21244
rect 13572 21184 13636 21188
rect 13652 21244 13716 21248
rect 13652 21188 13656 21244
rect 13656 21188 13712 21244
rect 13712 21188 13716 21244
rect 13652 21184 13716 21188
rect 13732 21244 13796 21248
rect 13732 21188 13736 21244
rect 13736 21188 13792 21244
rect 13792 21188 13796 21244
rect 13732 21184 13796 21188
rect 13812 21244 13876 21248
rect 13812 21188 13816 21244
rect 13816 21188 13872 21244
rect 13872 21188 13876 21244
rect 13812 21184 13876 21188
rect 18572 21244 18636 21248
rect 18572 21188 18576 21244
rect 18576 21188 18632 21244
rect 18632 21188 18636 21244
rect 18572 21184 18636 21188
rect 18652 21244 18716 21248
rect 18652 21188 18656 21244
rect 18656 21188 18712 21244
rect 18712 21188 18716 21244
rect 18652 21184 18716 21188
rect 18732 21244 18796 21248
rect 18732 21188 18736 21244
rect 18736 21188 18792 21244
rect 18792 21188 18796 21244
rect 18732 21184 18796 21188
rect 18812 21244 18876 21248
rect 18812 21188 18816 21244
rect 18816 21188 18872 21244
rect 18872 21188 18876 21244
rect 18812 21184 18876 21188
rect 23572 21244 23636 21248
rect 23572 21188 23576 21244
rect 23576 21188 23632 21244
rect 23632 21188 23636 21244
rect 23572 21184 23636 21188
rect 23652 21244 23716 21248
rect 23652 21188 23656 21244
rect 23656 21188 23712 21244
rect 23712 21188 23716 21244
rect 23652 21184 23716 21188
rect 23732 21244 23796 21248
rect 23732 21188 23736 21244
rect 23736 21188 23792 21244
rect 23792 21188 23796 21244
rect 23732 21184 23796 21188
rect 23812 21244 23876 21248
rect 23812 21188 23816 21244
rect 23816 21188 23872 21244
rect 23872 21188 23876 21244
rect 23812 21184 23876 21188
rect 28572 21244 28636 21248
rect 28572 21188 28576 21244
rect 28576 21188 28632 21244
rect 28632 21188 28636 21244
rect 28572 21184 28636 21188
rect 28652 21244 28716 21248
rect 28652 21188 28656 21244
rect 28656 21188 28712 21244
rect 28712 21188 28716 21244
rect 28652 21184 28716 21188
rect 28732 21244 28796 21248
rect 28732 21188 28736 21244
rect 28736 21188 28792 21244
rect 28792 21188 28796 21244
rect 28732 21184 28796 21188
rect 28812 21244 28876 21248
rect 28812 21188 28816 21244
rect 28816 21188 28872 21244
rect 28872 21188 28876 21244
rect 28812 21184 28876 21188
rect 33572 21244 33636 21248
rect 33572 21188 33576 21244
rect 33576 21188 33632 21244
rect 33632 21188 33636 21244
rect 33572 21184 33636 21188
rect 33652 21244 33716 21248
rect 33652 21188 33656 21244
rect 33656 21188 33712 21244
rect 33712 21188 33716 21244
rect 33652 21184 33716 21188
rect 33732 21244 33796 21248
rect 33732 21188 33736 21244
rect 33736 21188 33792 21244
rect 33792 21188 33796 21244
rect 33732 21184 33796 21188
rect 33812 21244 33876 21248
rect 33812 21188 33816 21244
rect 33816 21188 33872 21244
rect 33872 21188 33876 21244
rect 33812 21184 33876 21188
rect 38572 21244 38636 21248
rect 38572 21188 38576 21244
rect 38576 21188 38632 21244
rect 38632 21188 38636 21244
rect 38572 21184 38636 21188
rect 38652 21244 38716 21248
rect 38652 21188 38656 21244
rect 38656 21188 38712 21244
rect 38712 21188 38716 21244
rect 38652 21184 38716 21188
rect 38732 21244 38796 21248
rect 38732 21188 38736 21244
rect 38736 21188 38792 21244
rect 38792 21188 38796 21244
rect 38732 21184 38796 21188
rect 38812 21244 38876 21248
rect 38812 21188 38816 21244
rect 38816 21188 38872 21244
rect 38872 21188 38876 21244
rect 38812 21184 38876 21188
rect 43572 21244 43636 21248
rect 43572 21188 43576 21244
rect 43576 21188 43632 21244
rect 43632 21188 43636 21244
rect 43572 21184 43636 21188
rect 43652 21244 43716 21248
rect 43652 21188 43656 21244
rect 43656 21188 43712 21244
rect 43712 21188 43716 21244
rect 43652 21184 43716 21188
rect 43732 21244 43796 21248
rect 43732 21188 43736 21244
rect 43736 21188 43792 21244
rect 43792 21188 43796 21244
rect 43732 21184 43796 21188
rect 43812 21244 43876 21248
rect 43812 21188 43816 21244
rect 43816 21188 43872 21244
rect 43872 21188 43876 21244
rect 43812 21184 43876 21188
rect 27660 21116 27724 21180
rect 26740 20844 26804 20908
rect 9260 20708 9324 20772
rect 16988 20708 17052 20772
rect 17540 20768 17604 20772
rect 17540 20712 17554 20768
rect 17554 20712 17604 20768
rect 17540 20708 17604 20712
rect 19748 20768 19812 20772
rect 19748 20712 19798 20768
rect 19798 20712 19812 20768
rect 19748 20708 19812 20712
rect 21588 20708 21652 20772
rect 23244 20768 23308 20772
rect 23244 20712 23294 20768
rect 23294 20712 23308 20768
rect 23244 20708 23308 20712
rect 25452 20708 25516 20772
rect 27660 20708 27724 20772
rect 31892 20708 31956 20772
rect 6072 20700 6136 20704
rect 6072 20644 6076 20700
rect 6076 20644 6132 20700
rect 6132 20644 6136 20700
rect 6072 20640 6136 20644
rect 6152 20700 6216 20704
rect 6152 20644 6156 20700
rect 6156 20644 6212 20700
rect 6212 20644 6216 20700
rect 6152 20640 6216 20644
rect 6232 20700 6296 20704
rect 6232 20644 6236 20700
rect 6236 20644 6292 20700
rect 6292 20644 6296 20700
rect 6232 20640 6296 20644
rect 6312 20700 6376 20704
rect 6312 20644 6316 20700
rect 6316 20644 6372 20700
rect 6372 20644 6376 20700
rect 6312 20640 6376 20644
rect 11072 20700 11136 20704
rect 11072 20644 11076 20700
rect 11076 20644 11132 20700
rect 11132 20644 11136 20700
rect 11072 20640 11136 20644
rect 11152 20700 11216 20704
rect 11152 20644 11156 20700
rect 11156 20644 11212 20700
rect 11212 20644 11216 20700
rect 11152 20640 11216 20644
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 16072 20700 16136 20704
rect 16072 20644 16076 20700
rect 16076 20644 16132 20700
rect 16132 20644 16136 20700
rect 16072 20640 16136 20644
rect 16152 20700 16216 20704
rect 16152 20644 16156 20700
rect 16156 20644 16212 20700
rect 16212 20644 16216 20700
rect 16152 20640 16216 20644
rect 16232 20700 16296 20704
rect 16232 20644 16236 20700
rect 16236 20644 16292 20700
rect 16292 20644 16296 20700
rect 16232 20640 16296 20644
rect 16312 20700 16376 20704
rect 16312 20644 16316 20700
rect 16316 20644 16372 20700
rect 16372 20644 16376 20700
rect 16312 20640 16376 20644
rect 21072 20700 21136 20704
rect 21072 20644 21076 20700
rect 21076 20644 21132 20700
rect 21132 20644 21136 20700
rect 21072 20640 21136 20644
rect 21152 20700 21216 20704
rect 21152 20644 21156 20700
rect 21156 20644 21212 20700
rect 21212 20644 21216 20700
rect 21152 20640 21216 20644
rect 21232 20700 21296 20704
rect 21232 20644 21236 20700
rect 21236 20644 21292 20700
rect 21292 20644 21296 20700
rect 21232 20640 21296 20644
rect 21312 20700 21376 20704
rect 21312 20644 21316 20700
rect 21316 20644 21372 20700
rect 21372 20644 21376 20700
rect 21312 20640 21376 20644
rect 26072 20700 26136 20704
rect 26072 20644 26076 20700
rect 26076 20644 26132 20700
rect 26132 20644 26136 20700
rect 26072 20640 26136 20644
rect 26152 20700 26216 20704
rect 26152 20644 26156 20700
rect 26156 20644 26212 20700
rect 26212 20644 26216 20700
rect 26152 20640 26216 20644
rect 26232 20700 26296 20704
rect 26232 20644 26236 20700
rect 26236 20644 26292 20700
rect 26292 20644 26296 20700
rect 26232 20640 26296 20644
rect 26312 20700 26376 20704
rect 26312 20644 26316 20700
rect 26316 20644 26372 20700
rect 26372 20644 26376 20700
rect 26312 20640 26376 20644
rect 31072 20700 31136 20704
rect 31072 20644 31076 20700
rect 31076 20644 31132 20700
rect 31132 20644 31136 20700
rect 31072 20640 31136 20644
rect 31152 20700 31216 20704
rect 31152 20644 31156 20700
rect 31156 20644 31212 20700
rect 31212 20644 31216 20700
rect 31152 20640 31216 20644
rect 31232 20700 31296 20704
rect 31232 20644 31236 20700
rect 31236 20644 31292 20700
rect 31292 20644 31296 20700
rect 31232 20640 31296 20644
rect 31312 20700 31376 20704
rect 31312 20644 31316 20700
rect 31316 20644 31372 20700
rect 31372 20644 31376 20700
rect 31312 20640 31376 20644
rect 36072 20700 36136 20704
rect 36072 20644 36076 20700
rect 36076 20644 36132 20700
rect 36132 20644 36136 20700
rect 36072 20640 36136 20644
rect 36152 20700 36216 20704
rect 36152 20644 36156 20700
rect 36156 20644 36212 20700
rect 36212 20644 36216 20700
rect 36152 20640 36216 20644
rect 36232 20700 36296 20704
rect 36232 20644 36236 20700
rect 36236 20644 36292 20700
rect 36292 20644 36296 20700
rect 36232 20640 36296 20644
rect 36312 20700 36376 20704
rect 36312 20644 36316 20700
rect 36316 20644 36372 20700
rect 36372 20644 36376 20700
rect 36312 20640 36376 20644
rect 41072 20700 41136 20704
rect 41072 20644 41076 20700
rect 41076 20644 41132 20700
rect 41132 20644 41136 20700
rect 41072 20640 41136 20644
rect 41152 20700 41216 20704
rect 41152 20644 41156 20700
rect 41156 20644 41212 20700
rect 41212 20644 41216 20700
rect 41152 20640 41216 20644
rect 41232 20700 41296 20704
rect 41232 20644 41236 20700
rect 41236 20644 41292 20700
rect 41292 20644 41296 20700
rect 41232 20640 41296 20644
rect 41312 20700 41376 20704
rect 41312 20644 41316 20700
rect 41316 20644 41372 20700
rect 41372 20644 41376 20700
rect 41312 20640 41376 20644
rect 26556 20300 26620 20364
rect 3572 20156 3636 20160
rect 3572 20100 3576 20156
rect 3576 20100 3632 20156
rect 3632 20100 3636 20156
rect 3572 20096 3636 20100
rect 3652 20156 3716 20160
rect 3652 20100 3656 20156
rect 3656 20100 3712 20156
rect 3712 20100 3716 20156
rect 3652 20096 3716 20100
rect 3732 20156 3796 20160
rect 3732 20100 3736 20156
rect 3736 20100 3792 20156
rect 3792 20100 3796 20156
rect 3732 20096 3796 20100
rect 3812 20156 3876 20160
rect 3812 20100 3816 20156
rect 3816 20100 3872 20156
rect 3872 20100 3876 20156
rect 3812 20096 3876 20100
rect 8572 20156 8636 20160
rect 8572 20100 8576 20156
rect 8576 20100 8632 20156
rect 8632 20100 8636 20156
rect 8572 20096 8636 20100
rect 8652 20156 8716 20160
rect 8652 20100 8656 20156
rect 8656 20100 8712 20156
rect 8712 20100 8716 20156
rect 8652 20096 8716 20100
rect 8732 20156 8796 20160
rect 8732 20100 8736 20156
rect 8736 20100 8792 20156
rect 8792 20100 8796 20156
rect 8732 20096 8796 20100
rect 8812 20156 8876 20160
rect 8812 20100 8816 20156
rect 8816 20100 8872 20156
rect 8872 20100 8876 20156
rect 8812 20096 8876 20100
rect 13572 20156 13636 20160
rect 13572 20100 13576 20156
rect 13576 20100 13632 20156
rect 13632 20100 13636 20156
rect 13572 20096 13636 20100
rect 13652 20156 13716 20160
rect 13652 20100 13656 20156
rect 13656 20100 13712 20156
rect 13712 20100 13716 20156
rect 13652 20096 13716 20100
rect 13732 20156 13796 20160
rect 13732 20100 13736 20156
rect 13736 20100 13792 20156
rect 13792 20100 13796 20156
rect 13732 20096 13796 20100
rect 13812 20156 13876 20160
rect 13812 20100 13816 20156
rect 13816 20100 13872 20156
rect 13872 20100 13876 20156
rect 13812 20096 13876 20100
rect 18572 20156 18636 20160
rect 18572 20100 18576 20156
rect 18576 20100 18632 20156
rect 18632 20100 18636 20156
rect 18572 20096 18636 20100
rect 18652 20156 18716 20160
rect 18652 20100 18656 20156
rect 18656 20100 18712 20156
rect 18712 20100 18716 20156
rect 18652 20096 18716 20100
rect 18732 20156 18796 20160
rect 18732 20100 18736 20156
rect 18736 20100 18792 20156
rect 18792 20100 18796 20156
rect 18732 20096 18796 20100
rect 18812 20156 18876 20160
rect 18812 20100 18816 20156
rect 18816 20100 18872 20156
rect 18872 20100 18876 20156
rect 18812 20096 18876 20100
rect 23572 20156 23636 20160
rect 23572 20100 23576 20156
rect 23576 20100 23632 20156
rect 23632 20100 23636 20156
rect 23572 20096 23636 20100
rect 23652 20156 23716 20160
rect 23652 20100 23656 20156
rect 23656 20100 23712 20156
rect 23712 20100 23716 20156
rect 23652 20096 23716 20100
rect 23732 20156 23796 20160
rect 23732 20100 23736 20156
rect 23736 20100 23792 20156
rect 23792 20100 23796 20156
rect 23732 20096 23796 20100
rect 23812 20156 23876 20160
rect 23812 20100 23816 20156
rect 23816 20100 23872 20156
rect 23872 20100 23876 20156
rect 23812 20096 23876 20100
rect 28572 20156 28636 20160
rect 28572 20100 28576 20156
rect 28576 20100 28632 20156
rect 28632 20100 28636 20156
rect 28572 20096 28636 20100
rect 28652 20156 28716 20160
rect 28652 20100 28656 20156
rect 28656 20100 28712 20156
rect 28712 20100 28716 20156
rect 28652 20096 28716 20100
rect 28732 20156 28796 20160
rect 28732 20100 28736 20156
rect 28736 20100 28792 20156
rect 28792 20100 28796 20156
rect 28732 20096 28796 20100
rect 28812 20156 28876 20160
rect 28812 20100 28816 20156
rect 28816 20100 28872 20156
rect 28872 20100 28876 20156
rect 28812 20096 28876 20100
rect 33572 20156 33636 20160
rect 33572 20100 33576 20156
rect 33576 20100 33632 20156
rect 33632 20100 33636 20156
rect 33572 20096 33636 20100
rect 33652 20156 33716 20160
rect 33652 20100 33656 20156
rect 33656 20100 33712 20156
rect 33712 20100 33716 20156
rect 33652 20096 33716 20100
rect 33732 20156 33796 20160
rect 33732 20100 33736 20156
rect 33736 20100 33792 20156
rect 33792 20100 33796 20156
rect 33732 20096 33796 20100
rect 33812 20156 33876 20160
rect 33812 20100 33816 20156
rect 33816 20100 33872 20156
rect 33872 20100 33876 20156
rect 33812 20096 33876 20100
rect 38572 20156 38636 20160
rect 38572 20100 38576 20156
rect 38576 20100 38632 20156
rect 38632 20100 38636 20156
rect 38572 20096 38636 20100
rect 38652 20156 38716 20160
rect 38652 20100 38656 20156
rect 38656 20100 38712 20156
rect 38712 20100 38716 20156
rect 38652 20096 38716 20100
rect 38732 20156 38796 20160
rect 38732 20100 38736 20156
rect 38736 20100 38792 20156
rect 38792 20100 38796 20156
rect 38732 20096 38796 20100
rect 38812 20156 38876 20160
rect 38812 20100 38816 20156
rect 38816 20100 38872 20156
rect 38872 20100 38876 20156
rect 38812 20096 38876 20100
rect 43572 20156 43636 20160
rect 43572 20100 43576 20156
rect 43576 20100 43632 20156
rect 43632 20100 43636 20156
rect 43572 20096 43636 20100
rect 43652 20156 43716 20160
rect 43652 20100 43656 20156
rect 43656 20100 43712 20156
rect 43712 20100 43716 20156
rect 43652 20096 43716 20100
rect 43732 20156 43796 20160
rect 43732 20100 43736 20156
rect 43736 20100 43792 20156
rect 43792 20100 43796 20156
rect 43732 20096 43796 20100
rect 43812 20156 43876 20160
rect 43812 20100 43816 20156
rect 43816 20100 43872 20156
rect 43872 20100 43876 20156
rect 43812 20096 43876 20100
rect 23060 19756 23124 19820
rect 6072 19612 6136 19616
rect 6072 19556 6076 19612
rect 6076 19556 6132 19612
rect 6132 19556 6136 19612
rect 6072 19552 6136 19556
rect 6152 19612 6216 19616
rect 6152 19556 6156 19612
rect 6156 19556 6212 19612
rect 6212 19556 6216 19612
rect 6152 19552 6216 19556
rect 6232 19612 6296 19616
rect 6232 19556 6236 19612
rect 6236 19556 6292 19612
rect 6292 19556 6296 19612
rect 6232 19552 6296 19556
rect 6312 19612 6376 19616
rect 6312 19556 6316 19612
rect 6316 19556 6372 19612
rect 6372 19556 6376 19612
rect 6312 19552 6376 19556
rect 11072 19612 11136 19616
rect 11072 19556 11076 19612
rect 11076 19556 11132 19612
rect 11132 19556 11136 19612
rect 11072 19552 11136 19556
rect 11152 19612 11216 19616
rect 11152 19556 11156 19612
rect 11156 19556 11212 19612
rect 11212 19556 11216 19612
rect 11152 19552 11216 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 16072 19612 16136 19616
rect 16072 19556 16076 19612
rect 16076 19556 16132 19612
rect 16132 19556 16136 19612
rect 16072 19552 16136 19556
rect 16152 19612 16216 19616
rect 16152 19556 16156 19612
rect 16156 19556 16212 19612
rect 16212 19556 16216 19612
rect 16152 19552 16216 19556
rect 16232 19612 16296 19616
rect 16232 19556 16236 19612
rect 16236 19556 16292 19612
rect 16292 19556 16296 19612
rect 16232 19552 16296 19556
rect 16312 19612 16376 19616
rect 16312 19556 16316 19612
rect 16316 19556 16372 19612
rect 16372 19556 16376 19612
rect 16312 19552 16376 19556
rect 21072 19612 21136 19616
rect 21072 19556 21076 19612
rect 21076 19556 21132 19612
rect 21132 19556 21136 19612
rect 21072 19552 21136 19556
rect 21152 19612 21216 19616
rect 21152 19556 21156 19612
rect 21156 19556 21212 19612
rect 21212 19556 21216 19612
rect 21152 19552 21216 19556
rect 21232 19612 21296 19616
rect 21232 19556 21236 19612
rect 21236 19556 21292 19612
rect 21292 19556 21296 19612
rect 21232 19552 21296 19556
rect 21312 19612 21376 19616
rect 21312 19556 21316 19612
rect 21316 19556 21372 19612
rect 21372 19556 21376 19612
rect 21312 19552 21376 19556
rect 24348 19348 24412 19412
rect 25636 19756 25700 19820
rect 26072 19612 26136 19616
rect 26072 19556 26076 19612
rect 26076 19556 26132 19612
rect 26132 19556 26136 19612
rect 26072 19552 26136 19556
rect 26152 19612 26216 19616
rect 26152 19556 26156 19612
rect 26156 19556 26212 19612
rect 26212 19556 26216 19612
rect 26152 19552 26216 19556
rect 26232 19612 26296 19616
rect 26232 19556 26236 19612
rect 26236 19556 26292 19612
rect 26292 19556 26296 19612
rect 26232 19552 26296 19556
rect 26312 19612 26376 19616
rect 26312 19556 26316 19612
rect 26316 19556 26372 19612
rect 26372 19556 26376 19612
rect 26312 19552 26376 19556
rect 31072 19612 31136 19616
rect 31072 19556 31076 19612
rect 31076 19556 31132 19612
rect 31132 19556 31136 19612
rect 31072 19552 31136 19556
rect 31152 19612 31216 19616
rect 31152 19556 31156 19612
rect 31156 19556 31212 19612
rect 31212 19556 31216 19612
rect 31152 19552 31216 19556
rect 31232 19612 31296 19616
rect 31232 19556 31236 19612
rect 31236 19556 31292 19612
rect 31292 19556 31296 19612
rect 31232 19552 31296 19556
rect 31312 19612 31376 19616
rect 31312 19556 31316 19612
rect 31316 19556 31372 19612
rect 31372 19556 31376 19612
rect 31312 19552 31376 19556
rect 36072 19612 36136 19616
rect 36072 19556 36076 19612
rect 36076 19556 36132 19612
rect 36132 19556 36136 19612
rect 36072 19552 36136 19556
rect 36152 19612 36216 19616
rect 36152 19556 36156 19612
rect 36156 19556 36212 19612
rect 36212 19556 36216 19612
rect 36152 19552 36216 19556
rect 36232 19612 36296 19616
rect 36232 19556 36236 19612
rect 36236 19556 36292 19612
rect 36292 19556 36296 19612
rect 36232 19552 36296 19556
rect 36312 19612 36376 19616
rect 36312 19556 36316 19612
rect 36316 19556 36372 19612
rect 36372 19556 36376 19612
rect 36312 19552 36376 19556
rect 41072 19612 41136 19616
rect 41072 19556 41076 19612
rect 41076 19556 41132 19612
rect 41132 19556 41136 19612
rect 41072 19552 41136 19556
rect 41152 19612 41216 19616
rect 41152 19556 41156 19612
rect 41156 19556 41212 19612
rect 41212 19556 41216 19612
rect 41152 19552 41216 19556
rect 41232 19612 41296 19616
rect 41232 19556 41236 19612
rect 41236 19556 41292 19612
rect 41292 19556 41296 19612
rect 41232 19552 41296 19556
rect 41312 19612 41376 19616
rect 41312 19556 41316 19612
rect 41316 19556 41372 19612
rect 41372 19556 41376 19612
rect 41312 19552 41376 19556
rect 3572 19068 3636 19072
rect 3572 19012 3576 19068
rect 3576 19012 3632 19068
rect 3632 19012 3636 19068
rect 3572 19008 3636 19012
rect 3652 19068 3716 19072
rect 3652 19012 3656 19068
rect 3656 19012 3712 19068
rect 3712 19012 3716 19068
rect 3652 19008 3716 19012
rect 3732 19068 3796 19072
rect 3732 19012 3736 19068
rect 3736 19012 3792 19068
rect 3792 19012 3796 19068
rect 3732 19008 3796 19012
rect 3812 19068 3876 19072
rect 3812 19012 3816 19068
rect 3816 19012 3872 19068
rect 3872 19012 3876 19068
rect 3812 19008 3876 19012
rect 8572 19068 8636 19072
rect 8572 19012 8576 19068
rect 8576 19012 8632 19068
rect 8632 19012 8636 19068
rect 8572 19008 8636 19012
rect 8652 19068 8716 19072
rect 8652 19012 8656 19068
rect 8656 19012 8712 19068
rect 8712 19012 8716 19068
rect 8652 19008 8716 19012
rect 8732 19068 8796 19072
rect 8732 19012 8736 19068
rect 8736 19012 8792 19068
rect 8792 19012 8796 19068
rect 8732 19008 8796 19012
rect 8812 19068 8876 19072
rect 8812 19012 8816 19068
rect 8816 19012 8872 19068
rect 8872 19012 8876 19068
rect 8812 19008 8876 19012
rect 13572 19068 13636 19072
rect 13572 19012 13576 19068
rect 13576 19012 13632 19068
rect 13632 19012 13636 19068
rect 13572 19008 13636 19012
rect 13652 19068 13716 19072
rect 13652 19012 13656 19068
rect 13656 19012 13712 19068
rect 13712 19012 13716 19068
rect 13652 19008 13716 19012
rect 13732 19068 13796 19072
rect 13732 19012 13736 19068
rect 13736 19012 13792 19068
rect 13792 19012 13796 19068
rect 13732 19008 13796 19012
rect 13812 19068 13876 19072
rect 13812 19012 13816 19068
rect 13816 19012 13872 19068
rect 13872 19012 13876 19068
rect 13812 19008 13876 19012
rect 18572 19068 18636 19072
rect 18572 19012 18576 19068
rect 18576 19012 18632 19068
rect 18632 19012 18636 19068
rect 18572 19008 18636 19012
rect 18652 19068 18716 19072
rect 18652 19012 18656 19068
rect 18656 19012 18712 19068
rect 18712 19012 18716 19068
rect 18652 19008 18716 19012
rect 18732 19068 18796 19072
rect 18732 19012 18736 19068
rect 18736 19012 18792 19068
rect 18792 19012 18796 19068
rect 18732 19008 18796 19012
rect 18812 19068 18876 19072
rect 18812 19012 18816 19068
rect 18816 19012 18872 19068
rect 18872 19012 18876 19068
rect 18812 19008 18876 19012
rect 23572 19068 23636 19072
rect 23572 19012 23576 19068
rect 23576 19012 23632 19068
rect 23632 19012 23636 19068
rect 23572 19008 23636 19012
rect 23652 19068 23716 19072
rect 23652 19012 23656 19068
rect 23656 19012 23712 19068
rect 23712 19012 23716 19068
rect 23652 19008 23716 19012
rect 23732 19068 23796 19072
rect 23732 19012 23736 19068
rect 23736 19012 23792 19068
rect 23792 19012 23796 19068
rect 23732 19008 23796 19012
rect 23812 19068 23876 19072
rect 23812 19012 23816 19068
rect 23816 19012 23872 19068
rect 23872 19012 23876 19068
rect 23812 19008 23876 19012
rect 28572 19068 28636 19072
rect 28572 19012 28576 19068
rect 28576 19012 28632 19068
rect 28632 19012 28636 19068
rect 28572 19008 28636 19012
rect 28652 19068 28716 19072
rect 28652 19012 28656 19068
rect 28656 19012 28712 19068
rect 28712 19012 28716 19068
rect 28652 19008 28716 19012
rect 28732 19068 28796 19072
rect 28732 19012 28736 19068
rect 28736 19012 28792 19068
rect 28792 19012 28796 19068
rect 28732 19008 28796 19012
rect 28812 19068 28876 19072
rect 28812 19012 28816 19068
rect 28816 19012 28872 19068
rect 28872 19012 28876 19068
rect 28812 19008 28876 19012
rect 33572 19068 33636 19072
rect 33572 19012 33576 19068
rect 33576 19012 33632 19068
rect 33632 19012 33636 19068
rect 33572 19008 33636 19012
rect 33652 19068 33716 19072
rect 33652 19012 33656 19068
rect 33656 19012 33712 19068
rect 33712 19012 33716 19068
rect 33652 19008 33716 19012
rect 33732 19068 33796 19072
rect 33732 19012 33736 19068
rect 33736 19012 33792 19068
rect 33792 19012 33796 19068
rect 33732 19008 33796 19012
rect 33812 19068 33876 19072
rect 33812 19012 33816 19068
rect 33816 19012 33872 19068
rect 33872 19012 33876 19068
rect 33812 19008 33876 19012
rect 38572 19068 38636 19072
rect 38572 19012 38576 19068
rect 38576 19012 38632 19068
rect 38632 19012 38636 19068
rect 38572 19008 38636 19012
rect 38652 19068 38716 19072
rect 38652 19012 38656 19068
rect 38656 19012 38712 19068
rect 38712 19012 38716 19068
rect 38652 19008 38716 19012
rect 38732 19068 38796 19072
rect 38732 19012 38736 19068
rect 38736 19012 38792 19068
rect 38792 19012 38796 19068
rect 38732 19008 38796 19012
rect 38812 19068 38876 19072
rect 38812 19012 38816 19068
rect 38816 19012 38872 19068
rect 38872 19012 38876 19068
rect 38812 19008 38876 19012
rect 43572 19068 43636 19072
rect 43572 19012 43576 19068
rect 43576 19012 43632 19068
rect 43632 19012 43636 19068
rect 43572 19008 43636 19012
rect 43652 19068 43716 19072
rect 43652 19012 43656 19068
rect 43656 19012 43712 19068
rect 43712 19012 43716 19068
rect 43652 19008 43716 19012
rect 43732 19068 43796 19072
rect 43732 19012 43736 19068
rect 43736 19012 43792 19068
rect 43792 19012 43796 19068
rect 43732 19008 43796 19012
rect 43812 19068 43876 19072
rect 43812 19012 43816 19068
rect 43816 19012 43872 19068
rect 43872 19012 43876 19068
rect 43812 19008 43876 19012
rect 21956 18668 22020 18732
rect 6072 18524 6136 18528
rect 6072 18468 6076 18524
rect 6076 18468 6132 18524
rect 6132 18468 6136 18524
rect 6072 18464 6136 18468
rect 6152 18524 6216 18528
rect 6152 18468 6156 18524
rect 6156 18468 6212 18524
rect 6212 18468 6216 18524
rect 6152 18464 6216 18468
rect 6232 18524 6296 18528
rect 6232 18468 6236 18524
rect 6236 18468 6292 18524
rect 6292 18468 6296 18524
rect 6232 18464 6296 18468
rect 6312 18524 6376 18528
rect 6312 18468 6316 18524
rect 6316 18468 6372 18524
rect 6372 18468 6376 18524
rect 6312 18464 6376 18468
rect 11072 18524 11136 18528
rect 11072 18468 11076 18524
rect 11076 18468 11132 18524
rect 11132 18468 11136 18524
rect 11072 18464 11136 18468
rect 11152 18524 11216 18528
rect 11152 18468 11156 18524
rect 11156 18468 11212 18524
rect 11212 18468 11216 18524
rect 11152 18464 11216 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 16072 18524 16136 18528
rect 16072 18468 16076 18524
rect 16076 18468 16132 18524
rect 16132 18468 16136 18524
rect 16072 18464 16136 18468
rect 16152 18524 16216 18528
rect 16152 18468 16156 18524
rect 16156 18468 16212 18524
rect 16212 18468 16216 18524
rect 16152 18464 16216 18468
rect 16232 18524 16296 18528
rect 16232 18468 16236 18524
rect 16236 18468 16292 18524
rect 16292 18468 16296 18524
rect 16232 18464 16296 18468
rect 16312 18524 16376 18528
rect 16312 18468 16316 18524
rect 16316 18468 16372 18524
rect 16372 18468 16376 18524
rect 16312 18464 16376 18468
rect 21072 18524 21136 18528
rect 21072 18468 21076 18524
rect 21076 18468 21132 18524
rect 21132 18468 21136 18524
rect 21072 18464 21136 18468
rect 21152 18524 21216 18528
rect 21152 18468 21156 18524
rect 21156 18468 21212 18524
rect 21212 18468 21216 18524
rect 21152 18464 21216 18468
rect 21232 18524 21296 18528
rect 21232 18468 21236 18524
rect 21236 18468 21292 18524
rect 21292 18468 21296 18524
rect 21232 18464 21296 18468
rect 21312 18524 21376 18528
rect 21312 18468 21316 18524
rect 21316 18468 21372 18524
rect 21372 18468 21376 18524
rect 21312 18464 21376 18468
rect 26072 18524 26136 18528
rect 26072 18468 26076 18524
rect 26076 18468 26132 18524
rect 26132 18468 26136 18524
rect 26072 18464 26136 18468
rect 26152 18524 26216 18528
rect 26152 18468 26156 18524
rect 26156 18468 26212 18524
rect 26212 18468 26216 18524
rect 26152 18464 26216 18468
rect 26232 18524 26296 18528
rect 26232 18468 26236 18524
rect 26236 18468 26292 18524
rect 26292 18468 26296 18524
rect 26232 18464 26296 18468
rect 26312 18524 26376 18528
rect 26312 18468 26316 18524
rect 26316 18468 26372 18524
rect 26372 18468 26376 18524
rect 26312 18464 26376 18468
rect 31072 18524 31136 18528
rect 31072 18468 31076 18524
rect 31076 18468 31132 18524
rect 31132 18468 31136 18524
rect 31072 18464 31136 18468
rect 31152 18524 31216 18528
rect 31152 18468 31156 18524
rect 31156 18468 31212 18524
rect 31212 18468 31216 18524
rect 31152 18464 31216 18468
rect 31232 18524 31296 18528
rect 31232 18468 31236 18524
rect 31236 18468 31292 18524
rect 31292 18468 31296 18524
rect 31232 18464 31296 18468
rect 31312 18524 31376 18528
rect 31312 18468 31316 18524
rect 31316 18468 31372 18524
rect 31372 18468 31376 18524
rect 31312 18464 31376 18468
rect 36072 18524 36136 18528
rect 36072 18468 36076 18524
rect 36076 18468 36132 18524
rect 36132 18468 36136 18524
rect 36072 18464 36136 18468
rect 36152 18524 36216 18528
rect 36152 18468 36156 18524
rect 36156 18468 36212 18524
rect 36212 18468 36216 18524
rect 36152 18464 36216 18468
rect 36232 18524 36296 18528
rect 36232 18468 36236 18524
rect 36236 18468 36292 18524
rect 36292 18468 36296 18524
rect 36232 18464 36296 18468
rect 36312 18524 36376 18528
rect 36312 18468 36316 18524
rect 36316 18468 36372 18524
rect 36372 18468 36376 18524
rect 36312 18464 36376 18468
rect 41072 18524 41136 18528
rect 41072 18468 41076 18524
rect 41076 18468 41132 18524
rect 41132 18468 41136 18524
rect 41072 18464 41136 18468
rect 41152 18524 41216 18528
rect 41152 18468 41156 18524
rect 41156 18468 41212 18524
rect 41212 18468 41216 18524
rect 41152 18464 41216 18468
rect 41232 18524 41296 18528
rect 41232 18468 41236 18524
rect 41236 18468 41292 18524
rect 41292 18468 41296 18524
rect 41232 18464 41296 18468
rect 41312 18524 41376 18528
rect 41312 18468 41316 18524
rect 41316 18468 41372 18524
rect 41372 18468 41376 18524
rect 41312 18464 41376 18468
rect 3572 17980 3636 17984
rect 3572 17924 3576 17980
rect 3576 17924 3632 17980
rect 3632 17924 3636 17980
rect 3572 17920 3636 17924
rect 3652 17980 3716 17984
rect 3652 17924 3656 17980
rect 3656 17924 3712 17980
rect 3712 17924 3716 17980
rect 3652 17920 3716 17924
rect 3732 17980 3796 17984
rect 3732 17924 3736 17980
rect 3736 17924 3792 17980
rect 3792 17924 3796 17980
rect 3732 17920 3796 17924
rect 3812 17980 3876 17984
rect 3812 17924 3816 17980
rect 3816 17924 3872 17980
rect 3872 17924 3876 17980
rect 3812 17920 3876 17924
rect 8572 17980 8636 17984
rect 8572 17924 8576 17980
rect 8576 17924 8632 17980
rect 8632 17924 8636 17980
rect 8572 17920 8636 17924
rect 8652 17980 8716 17984
rect 8652 17924 8656 17980
rect 8656 17924 8712 17980
rect 8712 17924 8716 17980
rect 8652 17920 8716 17924
rect 8732 17980 8796 17984
rect 8732 17924 8736 17980
rect 8736 17924 8792 17980
rect 8792 17924 8796 17980
rect 8732 17920 8796 17924
rect 8812 17980 8876 17984
rect 8812 17924 8816 17980
rect 8816 17924 8872 17980
rect 8872 17924 8876 17980
rect 8812 17920 8876 17924
rect 13572 17980 13636 17984
rect 13572 17924 13576 17980
rect 13576 17924 13632 17980
rect 13632 17924 13636 17980
rect 13572 17920 13636 17924
rect 13652 17980 13716 17984
rect 13652 17924 13656 17980
rect 13656 17924 13712 17980
rect 13712 17924 13716 17980
rect 13652 17920 13716 17924
rect 13732 17980 13796 17984
rect 13732 17924 13736 17980
rect 13736 17924 13792 17980
rect 13792 17924 13796 17980
rect 13732 17920 13796 17924
rect 13812 17980 13876 17984
rect 13812 17924 13816 17980
rect 13816 17924 13872 17980
rect 13872 17924 13876 17980
rect 13812 17920 13876 17924
rect 18572 17980 18636 17984
rect 18572 17924 18576 17980
rect 18576 17924 18632 17980
rect 18632 17924 18636 17980
rect 18572 17920 18636 17924
rect 18652 17980 18716 17984
rect 18652 17924 18656 17980
rect 18656 17924 18712 17980
rect 18712 17924 18716 17980
rect 18652 17920 18716 17924
rect 18732 17980 18796 17984
rect 18732 17924 18736 17980
rect 18736 17924 18792 17980
rect 18792 17924 18796 17980
rect 18732 17920 18796 17924
rect 18812 17980 18876 17984
rect 18812 17924 18816 17980
rect 18816 17924 18872 17980
rect 18872 17924 18876 17980
rect 18812 17920 18876 17924
rect 23572 17980 23636 17984
rect 23572 17924 23576 17980
rect 23576 17924 23632 17980
rect 23632 17924 23636 17980
rect 23572 17920 23636 17924
rect 23652 17980 23716 17984
rect 23652 17924 23656 17980
rect 23656 17924 23712 17980
rect 23712 17924 23716 17980
rect 23652 17920 23716 17924
rect 23732 17980 23796 17984
rect 23732 17924 23736 17980
rect 23736 17924 23792 17980
rect 23792 17924 23796 17980
rect 23732 17920 23796 17924
rect 23812 17980 23876 17984
rect 23812 17924 23816 17980
rect 23816 17924 23872 17980
rect 23872 17924 23876 17980
rect 23812 17920 23876 17924
rect 28572 17980 28636 17984
rect 28572 17924 28576 17980
rect 28576 17924 28632 17980
rect 28632 17924 28636 17980
rect 28572 17920 28636 17924
rect 28652 17980 28716 17984
rect 28652 17924 28656 17980
rect 28656 17924 28712 17980
rect 28712 17924 28716 17980
rect 28652 17920 28716 17924
rect 28732 17980 28796 17984
rect 28732 17924 28736 17980
rect 28736 17924 28792 17980
rect 28792 17924 28796 17980
rect 28732 17920 28796 17924
rect 28812 17980 28876 17984
rect 28812 17924 28816 17980
rect 28816 17924 28872 17980
rect 28872 17924 28876 17980
rect 28812 17920 28876 17924
rect 33572 17980 33636 17984
rect 33572 17924 33576 17980
rect 33576 17924 33632 17980
rect 33632 17924 33636 17980
rect 33572 17920 33636 17924
rect 33652 17980 33716 17984
rect 33652 17924 33656 17980
rect 33656 17924 33712 17980
rect 33712 17924 33716 17980
rect 33652 17920 33716 17924
rect 33732 17980 33796 17984
rect 33732 17924 33736 17980
rect 33736 17924 33792 17980
rect 33792 17924 33796 17980
rect 33732 17920 33796 17924
rect 33812 17980 33876 17984
rect 33812 17924 33816 17980
rect 33816 17924 33872 17980
rect 33872 17924 33876 17980
rect 33812 17920 33876 17924
rect 38572 17980 38636 17984
rect 38572 17924 38576 17980
rect 38576 17924 38632 17980
rect 38632 17924 38636 17980
rect 38572 17920 38636 17924
rect 38652 17980 38716 17984
rect 38652 17924 38656 17980
rect 38656 17924 38712 17980
rect 38712 17924 38716 17980
rect 38652 17920 38716 17924
rect 38732 17980 38796 17984
rect 38732 17924 38736 17980
rect 38736 17924 38792 17980
rect 38792 17924 38796 17980
rect 38732 17920 38796 17924
rect 38812 17980 38876 17984
rect 38812 17924 38816 17980
rect 38816 17924 38872 17980
rect 38872 17924 38876 17980
rect 38812 17920 38876 17924
rect 43572 17980 43636 17984
rect 43572 17924 43576 17980
rect 43576 17924 43632 17980
rect 43632 17924 43636 17980
rect 43572 17920 43636 17924
rect 43652 17980 43716 17984
rect 43652 17924 43656 17980
rect 43656 17924 43712 17980
rect 43712 17924 43716 17980
rect 43652 17920 43716 17924
rect 43732 17980 43796 17984
rect 43732 17924 43736 17980
rect 43736 17924 43792 17980
rect 43792 17924 43796 17980
rect 43732 17920 43796 17924
rect 43812 17980 43876 17984
rect 43812 17924 43816 17980
rect 43816 17924 43872 17980
rect 43872 17924 43876 17980
rect 43812 17920 43876 17924
rect 30420 17504 30484 17508
rect 30420 17448 30470 17504
rect 30470 17448 30484 17504
rect 30420 17444 30484 17448
rect 6072 17436 6136 17440
rect 6072 17380 6076 17436
rect 6076 17380 6132 17436
rect 6132 17380 6136 17436
rect 6072 17376 6136 17380
rect 6152 17436 6216 17440
rect 6152 17380 6156 17436
rect 6156 17380 6212 17436
rect 6212 17380 6216 17436
rect 6152 17376 6216 17380
rect 6232 17436 6296 17440
rect 6232 17380 6236 17436
rect 6236 17380 6292 17436
rect 6292 17380 6296 17436
rect 6232 17376 6296 17380
rect 6312 17436 6376 17440
rect 6312 17380 6316 17436
rect 6316 17380 6372 17436
rect 6372 17380 6376 17436
rect 6312 17376 6376 17380
rect 11072 17436 11136 17440
rect 11072 17380 11076 17436
rect 11076 17380 11132 17436
rect 11132 17380 11136 17436
rect 11072 17376 11136 17380
rect 11152 17436 11216 17440
rect 11152 17380 11156 17436
rect 11156 17380 11212 17436
rect 11212 17380 11216 17436
rect 11152 17376 11216 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 16072 17436 16136 17440
rect 16072 17380 16076 17436
rect 16076 17380 16132 17436
rect 16132 17380 16136 17436
rect 16072 17376 16136 17380
rect 16152 17436 16216 17440
rect 16152 17380 16156 17436
rect 16156 17380 16212 17436
rect 16212 17380 16216 17436
rect 16152 17376 16216 17380
rect 16232 17436 16296 17440
rect 16232 17380 16236 17436
rect 16236 17380 16292 17436
rect 16292 17380 16296 17436
rect 16232 17376 16296 17380
rect 16312 17436 16376 17440
rect 16312 17380 16316 17436
rect 16316 17380 16372 17436
rect 16372 17380 16376 17436
rect 16312 17376 16376 17380
rect 21072 17436 21136 17440
rect 21072 17380 21076 17436
rect 21076 17380 21132 17436
rect 21132 17380 21136 17436
rect 21072 17376 21136 17380
rect 21152 17436 21216 17440
rect 21152 17380 21156 17436
rect 21156 17380 21212 17436
rect 21212 17380 21216 17436
rect 21152 17376 21216 17380
rect 21232 17436 21296 17440
rect 21232 17380 21236 17436
rect 21236 17380 21292 17436
rect 21292 17380 21296 17436
rect 21232 17376 21296 17380
rect 21312 17436 21376 17440
rect 21312 17380 21316 17436
rect 21316 17380 21372 17436
rect 21372 17380 21376 17436
rect 21312 17376 21376 17380
rect 26072 17436 26136 17440
rect 26072 17380 26076 17436
rect 26076 17380 26132 17436
rect 26132 17380 26136 17436
rect 26072 17376 26136 17380
rect 26152 17436 26216 17440
rect 26152 17380 26156 17436
rect 26156 17380 26212 17436
rect 26212 17380 26216 17436
rect 26152 17376 26216 17380
rect 26232 17436 26296 17440
rect 26232 17380 26236 17436
rect 26236 17380 26292 17436
rect 26292 17380 26296 17436
rect 26232 17376 26296 17380
rect 26312 17436 26376 17440
rect 26312 17380 26316 17436
rect 26316 17380 26372 17436
rect 26372 17380 26376 17436
rect 26312 17376 26376 17380
rect 31072 17436 31136 17440
rect 31072 17380 31076 17436
rect 31076 17380 31132 17436
rect 31132 17380 31136 17436
rect 31072 17376 31136 17380
rect 31152 17436 31216 17440
rect 31152 17380 31156 17436
rect 31156 17380 31212 17436
rect 31212 17380 31216 17436
rect 31152 17376 31216 17380
rect 31232 17436 31296 17440
rect 31232 17380 31236 17436
rect 31236 17380 31292 17436
rect 31292 17380 31296 17436
rect 31232 17376 31296 17380
rect 31312 17436 31376 17440
rect 31312 17380 31316 17436
rect 31316 17380 31372 17436
rect 31372 17380 31376 17436
rect 31312 17376 31376 17380
rect 36072 17436 36136 17440
rect 36072 17380 36076 17436
rect 36076 17380 36132 17436
rect 36132 17380 36136 17436
rect 36072 17376 36136 17380
rect 36152 17436 36216 17440
rect 36152 17380 36156 17436
rect 36156 17380 36212 17436
rect 36212 17380 36216 17436
rect 36152 17376 36216 17380
rect 36232 17436 36296 17440
rect 36232 17380 36236 17436
rect 36236 17380 36292 17436
rect 36292 17380 36296 17436
rect 36232 17376 36296 17380
rect 36312 17436 36376 17440
rect 36312 17380 36316 17436
rect 36316 17380 36372 17436
rect 36372 17380 36376 17436
rect 36312 17376 36376 17380
rect 41072 17436 41136 17440
rect 41072 17380 41076 17436
rect 41076 17380 41132 17436
rect 41132 17380 41136 17436
rect 41072 17376 41136 17380
rect 41152 17436 41216 17440
rect 41152 17380 41156 17436
rect 41156 17380 41212 17436
rect 41212 17380 41216 17436
rect 41152 17376 41216 17380
rect 41232 17436 41296 17440
rect 41232 17380 41236 17436
rect 41236 17380 41292 17436
rect 41292 17380 41296 17436
rect 41232 17376 41296 17380
rect 41312 17436 41376 17440
rect 41312 17380 41316 17436
rect 41316 17380 41372 17436
rect 41372 17380 41376 17436
rect 41312 17376 41376 17380
rect 22876 17172 22940 17236
rect 32812 17232 32876 17236
rect 32812 17176 32862 17232
rect 32862 17176 32876 17232
rect 32812 17172 32876 17176
rect 3572 16892 3636 16896
rect 3572 16836 3576 16892
rect 3576 16836 3632 16892
rect 3632 16836 3636 16892
rect 3572 16832 3636 16836
rect 3652 16892 3716 16896
rect 3652 16836 3656 16892
rect 3656 16836 3712 16892
rect 3712 16836 3716 16892
rect 3652 16832 3716 16836
rect 3732 16892 3796 16896
rect 3732 16836 3736 16892
rect 3736 16836 3792 16892
rect 3792 16836 3796 16892
rect 3732 16832 3796 16836
rect 3812 16892 3876 16896
rect 3812 16836 3816 16892
rect 3816 16836 3872 16892
rect 3872 16836 3876 16892
rect 3812 16832 3876 16836
rect 8572 16892 8636 16896
rect 8572 16836 8576 16892
rect 8576 16836 8632 16892
rect 8632 16836 8636 16892
rect 8572 16832 8636 16836
rect 8652 16892 8716 16896
rect 8652 16836 8656 16892
rect 8656 16836 8712 16892
rect 8712 16836 8716 16892
rect 8652 16832 8716 16836
rect 8732 16892 8796 16896
rect 8732 16836 8736 16892
rect 8736 16836 8792 16892
rect 8792 16836 8796 16892
rect 8732 16832 8796 16836
rect 8812 16892 8876 16896
rect 8812 16836 8816 16892
rect 8816 16836 8872 16892
rect 8872 16836 8876 16892
rect 8812 16832 8876 16836
rect 13572 16892 13636 16896
rect 13572 16836 13576 16892
rect 13576 16836 13632 16892
rect 13632 16836 13636 16892
rect 13572 16832 13636 16836
rect 13652 16892 13716 16896
rect 13652 16836 13656 16892
rect 13656 16836 13712 16892
rect 13712 16836 13716 16892
rect 13652 16832 13716 16836
rect 13732 16892 13796 16896
rect 13732 16836 13736 16892
rect 13736 16836 13792 16892
rect 13792 16836 13796 16892
rect 13732 16832 13796 16836
rect 13812 16892 13876 16896
rect 13812 16836 13816 16892
rect 13816 16836 13872 16892
rect 13872 16836 13876 16892
rect 13812 16832 13876 16836
rect 18572 16892 18636 16896
rect 18572 16836 18576 16892
rect 18576 16836 18632 16892
rect 18632 16836 18636 16892
rect 18572 16832 18636 16836
rect 18652 16892 18716 16896
rect 18652 16836 18656 16892
rect 18656 16836 18712 16892
rect 18712 16836 18716 16892
rect 18652 16832 18716 16836
rect 18732 16892 18796 16896
rect 18732 16836 18736 16892
rect 18736 16836 18792 16892
rect 18792 16836 18796 16892
rect 18732 16832 18796 16836
rect 18812 16892 18876 16896
rect 18812 16836 18816 16892
rect 18816 16836 18872 16892
rect 18872 16836 18876 16892
rect 18812 16832 18876 16836
rect 23572 16892 23636 16896
rect 23572 16836 23576 16892
rect 23576 16836 23632 16892
rect 23632 16836 23636 16892
rect 23572 16832 23636 16836
rect 23652 16892 23716 16896
rect 23652 16836 23656 16892
rect 23656 16836 23712 16892
rect 23712 16836 23716 16892
rect 23652 16832 23716 16836
rect 23732 16892 23796 16896
rect 23732 16836 23736 16892
rect 23736 16836 23792 16892
rect 23792 16836 23796 16892
rect 23732 16832 23796 16836
rect 23812 16892 23876 16896
rect 23812 16836 23816 16892
rect 23816 16836 23872 16892
rect 23872 16836 23876 16892
rect 23812 16832 23876 16836
rect 28572 16892 28636 16896
rect 28572 16836 28576 16892
rect 28576 16836 28632 16892
rect 28632 16836 28636 16892
rect 28572 16832 28636 16836
rect 28652 16892 28716 16896
rect 28652 16836 28656 16892
rect 28656 16836 28712 16892
rect 28712 16836 28716 16892
rect 28652 16832 28716 16836
rect 28732 16892 28796 16896
rect 28732 16836 28736 16892
rect 28736 16836 28792 16892
rect 28792 16836 28796 16892
rect 28732 16832 28796 16836
rect 28812 16892 28876 16896
rect 28812 16836 28816 16892
rect 28816 16836 28872 16892
rect 28872 16836 28876 16892
rect 28812 16832 28876 16836
rect 33572 16892 33636 16896
rect 33572 16836 33576 16892
rect 33576 16836 33632 16892
rect 33632 16836 33636 16892
rect 33572 16832 33636 16836
rect 33652 16892 33716 16896
rect 33652 16836 33656 16892
rect 33656 16836 33712 16892
rect 33712 16836 33716 16892
rect 33652 16832 33716 16836
rect 33732 16892 33796 16896
rect 33732 16836 33736 16892
rect 33736 16836 33792 16892
rect 33792 16836 33796 16892
rect 33732 16832 33796 16836
rect 33812 16892 33876 16896
rect 33812 16836 33816 16892
rect 33816 16836 33872 16892
rect 33872 16836 33876 16892
rect 33812 16832 33876 16836
rect 38572 16892 38636 16896
rect 38572 16836 38576 16892
rect 38576 16836 38632 16892
rect 38632 16836 38636 16892
rect 38572 16832 38636 16836
rect 38652 16892 38716 16896
rect 38652 16836 38656 16892
rect 38656 16836 38712 16892
rect 38712 16836 38716 16892
rect 38652 16832 38716 16836
rect 38732 16892 38796 16896
rect 38732 16836 38736 16892
rect 38736 16836 38792 16892
rect 38792 16836 38796 16892
rect 38732 16832 38796 16836
rect 38812 16892 38876 16896
rect 38812 16836 38816 16892
rect 38816 16836 38872 16892
rect 38872 16836 38876 16892
rect 38812 16832 38876 16836
rect 43572 16892 43636 16896
rect 43572 16836 43576 16892
rect 43576 16836 43632 16892
rect 43632 16836 43636 16892
rect 43572 16832 43636 16836
rect 43652 16892 43716 16896
rect 43652 16836 43656 16892
rect 43656 16836 43712 16892
rect 43712 16836 43716 16892
rect 43652 16832 43716 16836
rect 43732 16892 43796 16896
rect 43732 16836 43736 16892
rect 43736 16836 43792 16892
rect 43792 16836 43796 16892
rect 43732 16832 43796 16836
rect 43812 16892 43876 16896
rect 43812 16836 43816 16892
rect 43816 16836 43872 16892
rect 43872 16836 43876 16892
rect 43812 16832 43876 16836
rect 33180 16492 33244 16556
rect 6072 16348 6136 16352
rect 6072 16292 6076 16348
rect 6076 16292 6132 16348
rect 6132 16292 6136 16348
rect 6072 16288 6136 16292
rect 6152 16348 6216 16352
rect 6152 16292 6156 16348
rect 6156 16292 6212 16348
rect 6212 16292 6216 16348
rect 6152 16288 6216 16292
rect 6232 16348 6296 16352
rect 6232 16292 6236 16348
rect 6236 16292 6292 16348
rect 6292 16292 6296 16348
rect 6232 16288 6296 16292
rect 6312 16348 6376 16352
rect 6312 16292 6316 16348
rect 6316 16292 6372 16348
rect 6372 16292 6376 16348
rect 6312 16288 6376 16292
rect 11072 16348 11136 16352
rect 11072 16292 11076 16348
rect 11076 16292 11132 16348
rect 11132 16292 11136 16348
rect 11072 16288 11136 16292
rect 11152 16348 11216 16352
rect 11152 16292 11156 16348
rect 11156 16292 11212 16348
rect 11212 16292 11216 16348
rect 11152 16288 11216 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 16072 16348 16136 16352
rect 16072 16292 16076 16348
rect 16076 16292 16132 16348
rect 16132 16292 16136 16348
rect 16072 16288 16136 16292
rect 16152 16348 16216 16352
rect 16152 16292 16156 16348
rect 16156 16292 16212 16348
rect 16212 16292 16216 16348
rect 16152 16288 16216 16292
rect 16232 16348 16296 16352
rect 16232 16292 16236 16348
rect 16236 16292 16292 16348
rect 16292 16292 16296 16348
rect 16232 16288 16296 16292
rect 16312 16348 16376 16352
rect 16312 16292 16316 16348
rect 16316 16292 16372 16348
rect 16372 16292 16376 16348
rect 16312 16288 16376 16292
rect 21072 16348 21136 16352
rect 21072 16292 21076 16348
rect 21076 16292 21132 16348
rect 21132 16292 21136 16348
rect 21072 16288 21136 16292
rect 21152 16348 21216 16352
rect 21152 16292 21156 16348
rect 21156 16292 21212 16348
rect 21212 16292 21216 16348
rect 21152 16288 21216 16292
rect 21232 16348 21296 16352
rect 21232 16292 21236 16348
rect 21236 16292 21292 16348
rect 21292 16292 21296 16348
rect 21232 16288 21296 16292
rect 21312 16348 21376 16352
rect 21312 16292 21316 16348
rect 21316 16292 21372 16348
rect 21372 16292 21376 16348
rect 21312 16288 21376 16292
rect 26072 16348 26136 16352
rect 26072 16292 26076 16348
rect 26076 16292 26132 16348
rect 26132 16292 26136 16348
rect 26072 16288 26136 16292
rect 26152 16348 26216 16352
rect 26152 16292 26156 16348
rect 26156 16292 26212 16348
rect 26212 16292 26216 16348
rect 26152 16288 26216 16292
rect 26232 16348 26296 16352
rect 26232 16292 26236 16348
rect 26236 16292 26292 16348
rect 26292 16292 26296 16348
rect 26232 16288 26296 16292
rect 26312 16348 26376 16352
rect 26312 16292 26316 16348
rect 26316 16292 26372 16348
rect 26372 16292 26376 16348
rect 26312 16288 26376 16292
rect 31072 16348 31136 16352
rect 31072 16292 31076 16348
rect 31076 16292 31132 16348
rect 31132 16292 31136 16348
rect 31072 16288 31136 16292
rect 31152 16348 31216 16352
rect 31152 16292 31156 16348
rect 31156 16292 31212 16348
rect 31212 16292 31216 16348
rect 31152 16288 31216 16292
rect 31232 16348 31296 16352
rect 31232 16292 31236 16348
rect 31236 16292 31292 16348
rect 31292 16292 31296 16348
rect 31232 16288 31296 16292
rect 31312 16348 31376 16352
rect 31312 16292 31316 16348
rect 31316 16292 31372 16348
rect 31372 16292 31376 16348
rect 31312 16288 31376 16292
rect 36072 16348 36136 16352
rect 36072 16292 36076 16348
rect 36076 16292 36132 16348
rect 36132 16292 36136 16348
rect 36072 16288 36136 16292
rect 36152 16348 36216 16352
rect 36152 16292 36156 16348
rect 36156 16292 36212 16348
rect 36212 16292 36216 16348
rect 36152 16288 36216 16292
rect 36232 16348 36296 16352
rect 36232 16292 36236 16348
rect 36236 16292 36292 16348
rect 36292 16292 36296 16348
rect 36232 16288 36296 16292
rect 36312 16348 36376 16352
rect 36312 16292 36316 16348
rect 36316 16292 36372 16348
rect 36372 16292 36376 16348
rect 36312 16288 36376 16292
rect 41072 16348 41136 16352
rect 41072 16292 41076 16348
rect 41076 16292 41132 16348
rect 41132 16292 41136 16348
rect 41072 16288 41136 16292
rect 41152 16348 41216 16352
rect 41152 16292 41156 16348
rect 41156 16292 41212 16348
rect 41212 16292 41216 16348
rect 41152 16288 41216 16292
rect 41232 16348 41296 16352
rect 41232 16292 41236 16348
rect 41236 16292 41292 16348
rect 41292 16292 41296 16348
rect 41232 16288 41296 16292
rect 41312 16348 41376 16352
rect 41312 16292 41316 16348
rect 41316 16292 41372 16348
rect 41372 16292 41376 16348
rect 41312 16288 41376 16292
rect 26924 15948 26988 16012
rect 30236 15948 30300 16012
rect 3572 15804 3636 15808
rect 3572 15748 3576 15804
rect 3576 15748 3632 15804
rect 3632 15748 3636 15804
rect 3572 15744 3636 15748
rect 3652 15804 3716 15808
rect 3652 15748 3656 15804
rect 3656 15748 3712 15804
rect 3712 15748 3716 15804
rect 3652 15744 3716 15748
rect 3732 15804 3796 15808
rect 3732 15748 3736 15804
rect 3736 15748 3792 15804
rect 3792 15748 3796 15804
rect 3732 15744 3796 15748
rect 3812 15804 3876 15808
rect 3812 15748 3816 15804
rect 3816 15748 3872 15804
rect 3872 15748 3876 15804
rect 3812 15744 3876 15748
rect 8572 15804 8636 15808
rect 8572 15748 8576 15804
rect 8576 15748 8632 15804
rect 8632 15748 8636 15804
rect 8572 15744 8636 15748
rect 8652 15804 8716 15808
rect 8652 15748 8656 15804
rect 8656 15748 8712 15804
rect 8712 15748 8716 15804
rect 8652 15744 8716 15748
rect 8732 15804 8796 15808
rect 8732 15748 8736 15804
rect 8736 15748 8792 15804
rect 8792 15748 8796 15804
rect 8732 15744 8796 15748
rect 8812 15804 8876 15808
rect 8812 15748 8816 15804
rect 8816 15748 8872 15804
rect 8872 15748 8876 15804
rect 8812 15744 8876 15748
rect 13572 15804 13636 15808
rect 13572 15748 13576 15804
rect 13576 15748 13632 15804
rect 13632 15748 13636 15804
rect 13572 15744 13636 15748
rect 13652 15804 13716 15808
rect 13652 15748 13656 15804
rect 13656 15748 13712 15804
rect 13712 15748 13716 15804
rect 13652 15744 13716 15748
rect 13732 15804 13796 15808
rect 13732 15748 13736 15804
rect 13736 15748 13792 15804
rect 13792 15748 13796 15804
rect 13732 15744 13796 15748
rect 13812 15804 13876 15808
rect 13812 15748 13816 15804
rect 13816 15748 13872 15804
rect 13872 15748 13876 15804
rect 13812 15744 13876 15748
rect 18572 15804 18636 15808
rect 18572 15748 18576 15804
rect 18576 15748 18632 15804
rect 18632 15748 18636 15804
rect 18572 15744 18636 15748
rect 18652 15804 18716 15808
rect 18652 15748 18656 15804
rect 18656 15748 18712 15804
rect 18712 15748 18716 15804
rect 18652 15744 18716 15748
rect 18732 15804 18796 15808
rect 18732 15748 18736 15804
rect 18736 15748 18792 15804
rect 18792 15748 18796 15804
rect 18732 15744 18796 15748
rect 18812 15804 18876 15808
rect 18812 15748 18816 15804
rect 18816 15748 18872 15804
rect 18872 15748 18876 15804
rect 18812 15744 18876 15748
rect 23572 15804 23636 15808
rect 23572 15748 23576 15804
rect 23576 15748 23632 15804
rect 23632 15748 23636 15804
rect 23572 15744 23636 15748
rect 23652 15804 23716 15808
rect 23652 15748 23656 15804
rect 23656 15748 23712 15804
rect 23712 15748 23716 15804
rect 23652 15744 23716 15748
rect 23732 15804 23796 15808
rect 23732 15748 23736 15804
rect 23736 15748 23792 15804
rect 23792 15748 23796 15804
rect 23732 15744 23796 15748
rect 23812 15804 23876 15808
rect 23812 15748 23816 15804
rect 23816 15748 23872 15804
rect 23872 15748 23876 15804
rect 23812 15744 23876 15748
rect 28572 15804 28636 15808
rect 28572 15748 28576 15804
rect 28576 15748 28632 15804
rect 28632 15748 28636 15804
rect 28572 15744 28636 15748
rect 28652 15804 28716 15808
rect 28652 15748 28656 15804
rect 28656 15748 28712 15804
rect 28712 15748 28716 15804
rect 28652 15744 28716 15748
rect 28732 15804 28796 15808
rect 28732 15748 28736 15804
rect 28736 15748 28792 15804
rect 28792 15748 28796 15804
rect 28732 15744 28796 15748
rect 28812 15804 28876 15808
rect 28812 15748 28816 15804
rect 28816 15748 28872 15804
rect 28872 15748 28876 15804
rect 28812 15744 28876 15748
rect 33572 15804 33636 15808
rect 33572 15748 33576 15804
rect 33576 15748 33632 15804
rect 33632 15748 33636 15804
rect 33572 15744 33636 15748
rect 33652 15804 33716 15808
rect 33652 15748 33656 15804
rect 33656 15748 33712 15804
rect 33712 15748 33716 15804
rect 33652 15744 33716 15748
rect 33732 15804 33796 15808
rect 33732 15748 33736 15804
rect 33736 15748 33792 15804
rect 33792 15748 33796 15804
rect 33732 15744 33796 15748
rect 33812 15804 33876 15808
rect 33812 15748 33816 15804
rect 33816 15748 33872 15804
rect 33872 15748 33876 15804
rect 33812 15744 33876 15748
rect 38572 15804 38636 15808
rect 38572 15748 38576 15804
rect 38576 15748 38632 15804
rect 38632 15748 38636 15804
rect 38572 15744 38636 15748
rect 38652 15804 38716 15808
rect 38652 15748 38656 15804
rect 38656 15748 38712 15804
rect 38712 15748 38716 15804
rect 38652 15744 38716 15748
rect 38732 15804 38796 15808
rect 38732 15748 38736 15804
rect 38736 15748 38792 15804
rect 38792 15748 38796 15804
rect 38732 15744 38796 15748
rect 38812 15804 38876 15808
rect 38812 15748 38816 15804
rect 38816 15748 38872 15804
rect 38872 15748 38876 15804
rect 38812 15744 38876 15748
rect 43572 15804 43636 15808
rect 43572 15748 43576 15804
rect 43576 15748 43632 15804
rect 43632 15748 43636 15804
rect 43572 15744 43636 15748
rect 43652 15804 43716 15808
rect 43652 15748 43656 15804
rect 43656 15748 43712 15804
rect 43712 15748 43716 15804
rect 43652 15744 43716 15748
rect 43732 15804 43796 15808
rect 43732 15748 43736 15804
rect 43736 15748 43792 15804
rect 43792 15748 43796 15804
rect 43732 15744 43796 15748
rect 43812 15804 43876 15808
rect 43812 15748 43816 15804
rect 43816 15748 43872 15804
rect 43872 15748 43876 15804
rect 43812 15744 43876 15748
rect 6072 15260 6136 15264
rect 6072 15204 6076 15260
rect 6076 15204 6132 15260
rect 6132 15204 6136 15260
rect 6072 15200 6136 15204
rect 6152 15260 6216 15264
rect 6152 15204 6156 15260
rect 6156 15204 6212 15260
rect 6212 15204 6216 15260
rect 6152 15200 6216 15204
rect 6232 15260 6296 15264
rect 6232 15204 6236 15260
rect 6236 15204 6292 15260
rect 6292 15204 6296 15260
rect 6232 15200 6296 15204
rect 6312 15260 6376 15264
rect 6312 15204 6316 15260
rect 6316 15204 6372 15260
rect 6372 15204 6376 15260
rect 6312 15200 6376 15204
rect 11072 15260 11136 15264
rect 11072 15204 11076 15260
rect 11076 15204 11132 15260
rect 11132 15204 11136 15260
rect 11072 15200 11136 15204
rect 11152 15260 11216 15264
rect 11152 15204 11156 15260
rect 11156 15204 11212 15260
rect 11212 15204 11216 15260
rect 11152 15200 11216 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 16072 15260 16136 15264
rect 16072 15204 16076 15260
rect 16076 15204 16132 15260
rect 16132 15204 16136 15260
rect 16072 15200 16136 15204
rect 16152 15260 16216 15264
rect 16152 15204 16156 15260
rect 16156 15204 16212 15260
rect 16212 15204 16216 15260
rect 16152 15200 16216 15204
rect 16232 15260 16296 15264
rect 16232 15204 16236 15260
rect 16236 15204 16292 15260
rect 16292 15204 16296 15260
rect 16232 15200 16296 15204
rect 16312 15260 16376 15264
rect 16312 15204 16316 15260
rect 16316 15204 16372 15260
rect 16372 15204 16376 15260
rect 16312 15200 16376 15204
rect 21072 15260 21136 15264
rect 21072 15204 21076 15260
rect 21076 15204 21132 15260
rect 21132 15204 21136 15260
rect 21072 15200 21136 15204
rect 21152 15260 21216 15264
rect 21152 15204 21156 15260
rect 21156 15204 21212 15260
rect 21212 15204 21216 15260
rect 21152 15200 21216 15204
rect 21232 15260 21296 15264
rect 21232 15204 21236 15260
rect 21236 15204 21292 15260
rect 21292 15204 21296 15260
rect 21232 15200 21296 15204
rect 21312 15260 21376 15264
rect 21312 15204 21316 15260
rect 21316 15204 21372 15260
rect 21372 15204 21376 15260
rect 21312 15200 21376 15204
rect 26072 15260 26136 15264
rect 26072 15204 26076 15260
rect 26076 15204 26132 15260
rect 26132 15204 26136 15260
rect 26072 15200 26136 15204
rect 26152 15260 26216 15264
rect 26152 15204 26156 15260
rect 26156 15204 26212 15260
rect 26212 15204 26216 15260
rect 26152 15200 26216 15204
rect 26232 15260 26296 15264
rect 26232 15204 26236 15260
rect 26236 15204 26292 15260
rect 26292 15204 26296 15260
rect 26232 15200 26296 15204
rect 26312 15260 26376 15264
rect 26312 15204 26316 15260
rect 26316 15204 26372 15260
rect 26372 15204 26376 15260
rect 26312 15200 26376 15204
rect 31072 15260 31136 15264
rect 31072 15204 31076 15260
rect 31076 15204 31132 15260
rect 31132 15204 31136 15260
rect 31072 15200 31136 15204
rect 31152 15260 31216 15264
rect 31152 15204 31156 15260
rect 31156 15204 31212 15260
rect 31212 15204 31216 15260
rect 31152 15200 31216 15204
rect 31232 15260 31296 15264
rect 31232 15204 31236 15260
rect 31236 15204 31292 15260
rect 31292 15204 31296 15260
rect 31232 15200 31296 15204
rect 31312 15260 31376 15264
rect 31312 15204 31316 15260
rect 31316 15204 31372 15260
rect 31372 15204 31376 15260
rect 31312 15200 31376 15204
rect 36072 15260 36136 15264
rect 36072 15204 36076 15260
rect 36076 15204 36132 15260
rect 36132 15204 36136 15260
rect 36072 15200 36136 15204
rect 36152 15260 36216 15264
rect 36152 15204 36156 15260
rect 36156 15204 36212 15260
rect 36212 15204 36216 15260
rect 36152 15200 36216 15204
rect 36232 15260 36296 15264
rect 36232 15204 36236 15260
rect 36236 15204 36292 15260
rect 36292 15204 36296 15260
rect 36232 15200 36296 15204
rect 36312 15260 36376 15264
rect 36312 15204 36316 15260
rect 36316 15204 36372 15260
rect 36372 15204 36376 15260
rect 36312 15200 36376 15204
rect 41072 15260 41136 15264
rect 41072 15204 41076 15260
rect 41076 15204 41132 15260
rect 41132 15204 41136 15260
rect 41072 15200 41136 15204
rect 41152 15260 41216 15264
rect 41152 15204 41156 15260
rect 41156 15204 41212 15260
rect 41212 15204 41216 15260
rect 41152 15200 41216 15204
rect 41232 15260 41296 15264
rect 41232 15204 41236 15260
rect 41236 15204 41292 15260
rect 41292 15204 41296 15260
rect 41232 15200 41296 15204
rect 41312 15260 41376 15264
rect 41312 15204 41316 15260
rect 41316 15204 41372 15260
rect 41372 15204 41376 15260
rect 41312 15200 41376 15204
rect 22692 14860 22756 14924
rect 29316 14920 29380 14924
rect 29316 14864 29366 14920
rect 29366 14864 29380 14920
rect 29316 14860 29380 14864
rect 3572 14716 3636 14720
rect 3572 14660 3576 14716
rect 3576 14660 3632 14716
rect 3632 14660 3636 14716
rect 3572 14656 3636 14660
rect 3652 14716 3716 14720
rect 3652 14660 3656 14716
rect 3656 14660 3712 14716
rect 3712 14660 3716 14716
rect 3652 14656 3716 14660
rect 3732 14716 3796 14720
rect 3732 14660 3736 14716
rect 3736 14660 3792 14716
rect 3792 14660 3796 14716
rect 3732 14656 3796 14660
rect 3812 14716 3876 14720
rect 3812 14660 3816 14716
rect 3816 14660 3872 14716
rect 3872 14660 3876 14716
rect 3812 14656 3876 14660
rect 8572 14716 8636 14720
rect 8572 14660 8576 14716
rect 8576 14660 8632 14716
rect 8632 14660 8636 14716
rect 8572 14656 8636 14660
rect 8652 14716 8716 14720
rect 8652 14660 8656 14716
rect 8656 14660 8712 14716
rect 8712 14660 8716 14716
rect 8652 14656 8716 14660
rect 8732 14716 8796 14720
rect 8732 14660 8736 14716
rect 8736 14660 8792 14716
rect 8792 14660 8796 14716
rect 8732 14656 8796 14660
rect 8812 14716 8876 14720
rect 8812 14660 8816 14716
rect 8816 14660 8872 14716
rect 8872 14660 8876 14716
rect 8812 14656 8876 14660
rect 13572 14716 13636 14720
rect 13572 14660 13576 14716
rect 13576 14660 13632 14716
rect 13632 14660 13636 14716
rect 13572 14656 13636 14660
rect 13652 14716 13716 14720
rect 13652 14660 13656 14716
rect 13656 14660 13712 14716
rect 13712 14660 13716 14716
rect 13652 14656 13716 14660
rect 13732 14716 13796 14720
rect 13732 14660 13736 14716
rect 13736 14660 13792 14716
rect 13792 14660 13796 14716
rect 13732 14656 13796 14660
rect 13812 14716 13876 14720
rect 13812 14660 13816 14716
rect 13816 14660 13872 14716
rect 13872 14660 13876 14716
rect 13812 14656 13876 14660
rect 18572 14716 18636 14720
rect 18572 14660 18576 14716
rect 18576 14660 18632 14716
rect 18632 14660 18636 14716
rect 18572 14656 18636 14660
rect 18652 14716 18716 14720
rect 18652 14660 18656 14716
rect 18656 14660 18712 14716
rect 18712 14660 18716 14716
rect 18652 14656 18716 14660
rect 18732 14716 18796 14720
rect 18732 14660 18736 14716
rect 18736 14660 18792 14716
rect 18792 14660 18796 14716
rect 18732 14656 18796 14660
rect 18812 14716 18876 14720
rect 18812 14660 18816 14716
rect 18816 14660 18872 14716
rect 18872 14660 18876 14716
rect 18812 14656 18876 14660
rect 23572 14716 23636 14720
rect 23572 14660 23576 14716
rect 23576 14660 23632 14716
rect 23632 14660 23636 14716
rect 23572 14656 23636 14660
rect 23652 14716 23716 14720
rect 23652 14660 23656 14716
rect 23656 14660 23712 14716
rect 23712 14660 23716 14716
rect 23652 14656 23716 14660
rect 23732 14716 23796 14720
rect 23732 14660 23736 14716
rect 23736 14660 23792 14716
rect 23792 14660 23796 14716
rect 23732 14656 23796 14660
rect 23812 14716 23876 14720
rect 23812 14660 23816 14716
rect 23816 14660 23872 14716
rect 23872 14660 23876 14716
rect 23812 14656 23876 14660
rect 28572 14716 28636 14720
rect 28572 14660 28576 14716
rect 28576 14660 28632 14716
rect 28632 14660 28636 14716
rect 28572 14656 28636 14660
rect 28652 14716 28716 14720
rect 28652 14660 28656 14716
rect 28656 14660 28712 14716
rect 28712 14660 28716 14716
rect 28652 14656 28716 14660
rect 28732 14716 28796 14720
rect 28732 14660 28736 14716
rect 28736 14660 28792 14716
rect 28792 14660 28796 14716
rect 28732 14656 28796 14660
rect 28812 14716 28876 14720
rect 28812 14660 28816 14716
rect 28816 14660 28872 14716
rect 28872 14660 28876 14716
rect 28812 14656 28876 14660
rect 33572 14716 33636 14720
rect 33572 14660 33576 14716
rect 33576 14660 33632 14716
rect 33632 14660 33636 14716
rect 33572 14656 33636 14660
rect 33652 14716 33716 14720
rect 33652 14660 33656 14716
rect 33656 14660 33712 14716
rect 33712 14660 33716 14716
rect 33652 14656 33716 14660
rect 33732 14716 33796 14720
rect 33732 14660 33736 14716
rect 33736 14660 33792 14716
rect 33792 14660 33796 14716
rect 33732 14656 33796 14660
rect 33812 14716 33876 14720
rect 33812 14660 33816 14716
rect 33816 14660 33872 14716
rect 33872 14660 33876 14716
rect 33812 14656 33876 14660
rect 38572 14716 38636 14720
rect 38572 14660 38576 14716
rect 38576 14660 38632 14716
rect 38632 14660 38636 14716
rect 38572 14656 38636 14660
rect 38652 14716 38716 14720
rect 38652 14660 38656 14716
rect 38656 14660 38712 14716
rect 38712 14660 38716 14716
rect 38652 14656 38716 14660
rect 38732 14716 38796 14720
rect 38732 14660 38736 14716
rect 38736 14660 38792 14716
rect 38792 14660 38796 14716
rect 38732 14656 38796 14660
rect 38812 14716 38876 14720
rect 38812 14660 38816 14716
rect 38816 14660 38872 14716
rect 38872 14660 38876 14716
rect 38812 14656 38876 14660
rect 43572 14716 43636 14720
rect 43572 14660 43576 14716
rect 43576 14660 43632 14716
rect 43632 14660 43636 14716
rect 43572 14656 43636 14660
rect 43652 14716 43716 14720
rect 43652 14660 43656 14716
rect 43656 14660 43712 14716
rect 43712 14660 43716 14716
rect 43652 14656 43716 14660
rect 43732 14716 43796 14720
rect 43732 14660 43736 14716
rect 43736 14660 43792 14716
rect 43792 14660 43796 14716
rect 43732 14656 43796 14660
rect 43812 14716 43876 14720
rect 43812 14660 43816 14716
rect 43816 14660 43872 14716
rect 43872 14660 43876 14716
rect 43812 14656 43876 14660
rect 19012 14512 19076 14516
rect 19012 14456 19026 14512
rect 19026 14456 19076 14512
rect 19012 14452 19076 14456
rect 30788 14316 30852 14380
rect 6072 14172 6136 14176
rect 6072 14116 6076 14172
rect 6076 14116 6132 14172
rect 6132 14116 6136 14172
rect 6072 14112 6136 14116
rect 6152 14172 6216 14176
rect 6152 14116 6156 14172
rect 6156 14116 6212 14172
rect 6212 14116 6216 14172
rect 6152 14112 6216 14116
rect 6232 14172 6296 14176
rect 6232 14116 6236 14172
rect 6236 14116 6292 14172
rect 6292 14116 6296 14172
rect 6232 14112 6296 14116
rect 6312 14172 6376 14176
rect 6312 14116 6316 14172
rect 6316 14116 6372 14172
rect 6372 14116 6376 14172
rect 6312 14112 6376 14116
rect 11072 14172 11136 14176
rect 11072 14116 11076 14172
rect 11076 14116 11132 14172
rect 11132 14116 11136 14172
rect 11072 14112 11136 14116
rect 11152 14172 11216 14176
rect 11152 14116 11156 14172
rect 11156 14116 11212 14172
rect 11212 14116 11216 14172
rect 11152 14112 11216 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 16072 14172 16136 14176
rect 16072 14116 16076 14172
rect 16076 14116 16132 14172
rect 16132 14116 16136 14172
rect 16072 14112 16136 14116
rect 16152 14172 16216 14176
rect 16152 14116 16156 14172
rect 16156 14116 16212 14172
rect 16212 14116 16216 14172
rect 16152 14112 16216 14116
rect 16232 14172 16296 14176
rect 16232 14116 16236 14172
rect 16236 14116 16292 14172
rect 16292 14116 16296 14172
rect 16232 14112 16296 14116
rect 16312 14172 16376 14176
rect 16312 14116 16316 14172
rect 16316 14116 16372 14172
rect 16372 14116 16376 14172
rect 16312 14112 16376 14116
rect 21072 14172 21136 14176
rect 21072 14116 21076 14172
rect 21076 14116 21132 14172
rect 21132 14116 21136 14172
rect 21072 14112 21136 14116
rect 21152 14172 21216 14176
rect 21152 14116 21156 14172
rect 21156 14116 21212 14172
rect 21212 14116 21216 14172
rect 21152 14112 21216 14116
rect 21232 14172 21296 14176
rect 21232 14116 21236 14172
rect 21236 14116 21292 14172
rect 21292 14116 21296 14172
rect 21232 14112 21296 14116
rect 21312 14172 21376 14176
rect 21312 14116 21316 14172
rect 21316 14116 21372 14172
rect 21372 14116 21376 14172
rect 21312 14112 21376 14116
rect 26072 14172 26136 14176
rect 26072 14116 26076 14172
rect 26076 14116 26132 14172
rect 26132 14116 26136 14172
rect 26072 14112 26136 14116
rect 26152 14172 26216 14176
rect 26152 14116 26156 14172
rect 26156 14116 26212 14172
rect 26212 14116 26216 14172
rect 26152 14112 26216 14116
rect 26232 14172 26296 14176
rect 26232 14116 26236 14172
rect 26236 14116 26292 14172
rect 26292 14116 26296 14172
rect 26232 14112 26296 14116
rect 26312 14172 26376 14176
rect 26312 14116 26316 14172
rect 26316 14116 26372 14172
rect 26372 14116 26376 14172
rect 26312 14112 26376 14116
rect 31072 14172 31136 14176
rect 31072 14116 31076 14172
rect 31076 14116 31132 14172
rect 31132 14116 31136 14172
rect 31072 14112 31136 14116
rect 31152 14172 31216 14176
rect 31152 14116 31156 14172
rect 31156 14116 31212 14172
rect 31212 14116 31216 14172
rect 31152 14112 31216 14116
rect 31232 14172 31296 14176
rect 31232 14116 31236 14172
rect 31236 14116 31292 14172
rect 31292 14116 31296 14172
rect 31232 14112 31296 14116
rect 31312 14172 31376 14176
rect 31312 14116 31316 14172
rect 31316 14116 31372 14172
rect 31372 14116 31376 14172
rect 31312 14112 31376 14116
rect 36072 14172 36136 14176
rect 36072 14116 36076 14172
rect 36076 14116 36132 14172
rect 36132 14116 36136 14172
rect 36072 14112 36136 14116
rect 36152 14172 36216 14176
rect 36152 14116 36156 14172
rect 36156 14116 36212 14172
rect 36212 14116 36216 14172
rect 36152 14112 36216 14116
rect 36232 14172 36296 14176
rect 36232 14116 36236 14172
rect 36236 14116 36292 14172
rect 36292 14116 36296 14172
rect 36232 14112 36296 14116
rect 36312 14172 36376 14176
rect 36312 14116 36316 14172
rect 36316 14116 36372 14172
rect 36372 14116 36376 14172
rect 36312 14112 36376 14116
rect 41072 14172 41136 14176
rect 41072 14116 41076 14172
rect 41076 14116 41132 14172
rect 41132 14116 41136 14172
rect 41072 14112 41136 14116
rect 41152 14172 41216 14176
rect 41152 14116 41156 14172
rect 41156 14116 41212 14172
rect 41212 14116 41216 14172
rect 41152 14112 41216 14116
rect 41232 14172 41296 14176
rect 41232 14116 41236 14172
rect 41236 14116 41292 14172
rect 41292 14116 41296 14172
rect 41232 14112 41296 14116
rect 41312 14172 41376 14176
rect 41312 14116 41316 14172
rect 41316 14116 41372 14172
rect 41372 14116 41376 14172
rect 41312 14112 41376 14116
rect 26924 14044 26988 14108
rect 3572 13628 3636 13632
rect 3572 13572 3576 13628
rect 3576 13572 3632 13628
rect 3632 13572 3636 13628
rect 3572 13568 3636 13572
rect 3652 13628 3716 13632
rect 3652 13572 3656 13628
rect 3656 13572 3712 13628
rect 3712 13572 3716 13628
rect 3652 13568 3716 13572
rect 3732 13628 3796 13632
rect 3732 13572 3736 13628
rect 3736 13572 3792 13628
rect 3792 13572 3796 13628
rect 3732 13568 3796 13572
rect 3812 13628 3876 13632
rect 3812 13572 3816 13628
rect 3816 13572 3872 13628
rect 3872 13572 3876 13628
rect 3812 13568 3876 13572
rect 8572 13628 8636 13632
rect 8572 13572 8576 13628
rect 8576 13572 8632 13628
rect 8632 13572 8636 13628
rect 8572 13568 8636 13572
rect 8652 13628 8716 13632
rect 8652 13572 8656 13628
rect 8656 13572 8712 13628
rect 8712 13572 8716 13628
rect 8652 13568 8716 13572
rect 8732 13628 8796 13632
rect 8732 13572 8736 13628
rect 8736 13572 8792 13628
rect 8792 13572 8796 13628
rect 8732 13568 8796 13572
rect 8812 13628 8876 13632
rect 8812 13572 8816 13628
rect 8816 13572 8872 13628
rect 8872 13572 8876 13628
rect 8812 13568 8876 13572
rect 13572 13628 13636 13632
rect 13572 13572 13576 13628
rect 13576 13572 13632 13628
rect 13632 13572 13636 13628
rect 13572 13568 13636 13572
rect 13652 13628 13716 13632
rect 13652 13572 13656 13628
rect 13656 13572 13712 13628
rect 13712 13572 13716 13628
rect 13652 13568 13716 13572
rect 13732 13628 13796 13632
rect 13732 13572 13736 13628
rect 13736 13572 13792 13628
rect 13792 13572 13796 13628
rect 13732 13568 13796 13572
rect 13812 13628 13876 13632
rect 13812 13572 13816 13628
rect 13816 13572 13872 13628
rect 13872 13572 13876 13628
rect 13812 13568 13876 13572
rect 18572 13628 18636 13632
rect 18572 13572 18576 13628
rect 18576 13572 18632 13628
rect 18632 13572 18636 13628
rect 18572 13568 18636 13572
rect 18652 13628 18716 13632
rect 18652 13572 18656 13628
rect 18656 13572 18712 13628
rect 18712 13572 18716 13628
rect 18652 13568 18716 13572
rect 18732 13628 18796 13632
rect 18732 13572 18736 13628
rect 18736 13572 18792 13628
rect 18792 13572 18796 13628
rect 18732 13568 18796 13572
rect 18812 13628 18876 13632
rect 18812 13572 18816 13628
rect 18816 13572 18872 13628
rect 18872 13572 18876 13628
rect 18812 13568 18876 13572
rect 23572 13628 23636 13632
rect 23572 13572 23576 13628
rect 23576 13572 23632 13628
rect 23632 13572 23636 13628
rect 23572 13568 23636 13572
rect 23652 13628 23716 13632
rect 23652 13572 23656 13628
rect 23656 13572 23712 13628
rect 23712 13572 23716 13628
rect 23652 13568 23716 13572
rect 23732 13628 23796 13632
rect 23732 13572 23736 13628
rect 23736 13572 23792 13628
rect 23792 13572 23796 13628
rect 23732 13568 23796 13572
rect 23812 13628 23876 13632
rect 23812 13572 23816 13628
rect 23816 13572 23872 13628
rect 23872 13572 23876 13628
rect 23812 13568 23876 13572
rect 28572 13628 28636 13632
rect 28572 13572 28576 13628
rect 28576 13572 28632 13628
rect 28632 13572 28636 13628
rect 28572 13568 28636 13572
rect 28652 13628 28716 13632
rect 28652 13572 28656 13628
rect 28656 13572 28712 13628
rect 28712 13572 28716 13628
rect 28652 13568 28716 13572
rect 28732 13628 28796 13632
rect 28732 13572 28736 13628
rect 28736 13572 28792 13628
rect 28792 13572 28796 13628
rect 28732 13568 28796 13572
rect 28812 13628 28876 13632
rect 28812 13572 28816 13628
rect 28816 13572 28872 13628
rect 28872 13572 28876 13628
rect 28812 13568 28876 13572
rect 33572 13628 33636 13632
rect 33572 13572 33576 13628
rect 33576 13572 33632 13628
rect 33632 13572 33636 13628
rect 33572 13568 33636 13572
rect 33652 13628 33716 13632
rect 33652 13572 33656 13628
rect 33656 13572 33712 13628
rect 33712 13572 33716 13628
rect 33652 13568 33716 13572
rect 33732 13628 33796 13632
rect 33732 13572 33736 13628
rect 33736 13572 33792 13628
rect 33792 13572 33796 13628
rect 33732 13568 33796 13572
rect 33812 13628 33876 13632
rect 33812 13572 33816 13628
rect 33816 13572 33872 13628
rect 33872 13572 33876 13628
rect 33812 13568 33876 13572
rect 38572 13628 38636 13632
rect 38572 13572 38576 13628
rect 38576 13572 38632 13628
rect 38632 13572 38636 13628
rect 38572 13568 38636 13572
rect 38652 13628 38716 13632
rect 38652 13572 38656 13628
rect 38656 13572 38712 13628
rect 38712 13572 38716 13628
rect 38652 13568 38716 13572
rect 38732 13628 38796 13632
rect 38732 13572 38736 13628
rect 38736 13572 38792 13628
rect 38792 13572 38796 13628
rect 38732 13568 38796 13572
rect 38812 13628 38876 13632
rect 38812 13572 38816 13628
rect 38816 13572 38872 13628
rect 38872 13572 38876 13628
rect 38812 13568 38876 13572
rect 43572 13628 43636 13632
rect 43572 13572 43576 13628
rect 43576 13572 43632 13628
rect 43632 13572 43636 13628
rect 43572 13568 43636 13572
rect 43652 13628 43716 13632
rect 43652 13572 43656 13628
rect 43656 13572 43712 13628
rect 43712 13572 43716 13628
rect 43652 13568 43716 13572
rect 43732 13628 43796 13632
rect 43732 13572 43736 13628
rect 43736 13572 43792 13628
rect 43792 13572 43796 13628
rect 43732 13568 43796 13572
rect 43812 13628 43876 13632
rect 43812 13572 43816 13628
rect 43816 13572 43872 13628
rect 43872 13572 43876 13628
rect 43812 13568 43876 13572
rect 6072 13084 6136 13088
rect 6072 13028 6076 13084
rect 6076 13028 6132 13084
rect 6132 13028 6136 13084
rect 6072 13024 6136 13028
rect 6152 13084 6216 13088
rect 6152 13028 6156 13084
rect 6156 13028 6212 13084
rect 6212 13028 6216 13084
rect 6152 13024 6216 13028
rect 6232 13084 6296 13088
rect 6232 13028 6236 13084
rect 6236 13028 6292 13084
rect 6292 13028 6296 13084
rect 6232 13024 6296 13028
rect 6312 13084 6376 13088
rect 6312 13028 6316 13084
rect 6316 13028 6372 13084
rect 6372 13028 6376 13084
rect 6312 13024 6376 13028
rect 11072 13084 11136 13088
rect 11072 13028 11076 13084
rect 11076 13028 11132 13084
rect 11132 13028 11136 13084
rect 11072 13024 11136 13028
rect 11152 13084 11216 13088
rect 11152 13028 11156 13084
rect 11156 13028 11212 13084
rect 11212 13028 11216 13084
rect 11152 13024 11216 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 16072 13084 16136 13088
rect 16072 13028 16076 13084
rect 16076 13028 16132 13084
rect 16132 13028 16136 13084
rect 16072 13024 16136 13028
rect 16152 13084 16216 13088
rect 16152 13028 16156 13084
rect 16156 13028 16212 13084
rect 16212 13028 16216 13084
rect 16152 13024 16216 13028
rect 16232 13084 16296 13088
rect 16232 13028 16236 13084
rect 16236 13028 16292 13084
rect 16292 13028 16296 13084
rect 16232 13024 16296 13028
rect 16312 13084 16376 13088
rect 16312 13028 16316 13084
rect 16316 13028 16372 13084
rect 16372 13028 16376 13084
rect 16312 13024 16376 13028
rect 21072 13084 21136 13088
rect 21072 13028 21076 13084
rect 21076 13028 21132 13084
rect 21132 13028 21136 13084
rect 21072 13024 21136 13028
rect 21152 13084 21216 13088
rect 21152 13028 21156 13084
rect 21156 13028 21212 13084
rect 21212 13028 21216 13084
rect 21152 13024 21216 13028
rect 21232 13084 21296 13088
rect 21232 13028 21236 13084
rect 21236 13028 21292 13084
rect 21292 13028 21296 13084
rect 21232 13024 21296 13028
rect 21312 13084 21376 13088
rect 21312 13028 21316 13084
rect 21316 13028 21372 13084
rect 21372 13028 21376 13084
rect 21312 13024 21376 13028
rect 26072 13084 26136 13088
rect 26072 13028 26076 13084
rect 26076 13028 26132 13084
rect 26132 13028 26136 13084
rect 26072 13024 26136 13028
rect 26152 13084 26216 13088
rect 26152 13028 26156 13084
rect 26156 13028 26212 13084
rect 26212 13028 26216 13084
rect 26152 13024 26216 13028
rect 26232 13084 26296 13088
rect 26232 13028 26236 13084
rect 26236 13028 26292 13084
rect 26292 13028 26296 13084
rect 26232 13024 26296 13028
rect 26312 13084 26376 13088
rect 26312 13028 26316 13084
rect 26316 13028 26372 13084
rect 26372 13028 26376 13084
rect 26312 13024 26376 13028
rect 31072 13084 31136 13088
rect 31072 13028 31076 13084
rect 31076 13028 31132 13084
rect 31132 13028 31136 13084
rect 31072 13024 31136 13028
rect 31152 13084 31216 13088
rect 31152 13028 31156 13084
rect 31156 13028 31212 13084
rect 31212 13028 31216 13084
rect 31152 13024 31216 13028
rect 31232 13084 31296 13088
rect 31232 13028 31236 13084
rect 31236 13028 31292 13084
rect 31292 13028 31296 13084
rect 31232 13024 31296 13028
rect 31312 13084 31376 13088
rect 31312 13028 31316 13084
rect 31316 13028 31372 13084
rect 31372 13028 31376 13084
rect 31312 13024 31376 13028
rect 36072 13084 36136 13088
rect 36072 13028 36076 13084
rect 36076 13028 36132 13084
rect 36132 13028 36136 13084
rect 36072 13024 36136 13028
rect 36152 13084 36216 13088
rect 36152 13028 36156 13084
rect 36156 13028 36212 13084
rect 36212 13028 36216 13084
rect 36152 13024 36216 13028
rect 36232 13084 36296 13088
rect 36232 13028 36236 13084
rect 36236 13028 36292 13084
rect 36292 13028 36296 13084
rect 36232 13024 36296 13028
rect 36312 13084 36376 13088
rect 36312 13028 36316 13084
rect 36316 13028 36372 13084
rect 36372 13028 36376 13084
rect 36312 13024 36376 13028
rect 41072 13084 41136 13088
rect 41072 13028 41076 13084
rect 41076 13028 41132 13084
rect 41132 13028 41136 13084
rect 41072 13024 41136 13028
rect 41152 13084 41216 13088
rect 41152 13028 41156 13084
rect 41156 13028 41212 13084
rect 41212 13028 41216 13084
rect 41152 13024 41216 13028
rect 41232 13084 41296 13088
rect 41232 13028 41236 13084
rect 41236 13028 41292 13084
rect 41292 13028 41296 13084
rect 41232 13024 41296 13028
rect 41312 13084 41376 13088
rect 41312 13028 41316 13084
rect 41316 13028 41372 13084
rect 41372 13028 41376 13084
rect 41312 13024 41376 13028
rect 30420 12684 30484 12748
rect 3572 12540 3636 12544
rect 3572 12484 3576 12540
rect 3576 12484 3632 12540
rect 3632 12484 3636 12540
rect 3572 12480 3636 12484
rect 3652 12540 3716 12544
rect 3652 12484 3656 12540
rect 3656 12484 3712 12540
rect 3712 12484 3716 12540
rect 3652 12480 3716 12484
rect 3732 12540 3796 12544
rect 3732 12484 3736 12540
rect 3736 12484 3792 12540
rect 3792 12484 3796 12540
rect 3732 12480 3796 12484
rect 3812 12540 3876 12544
rect 3812 12484 3816 12540
rect 3816 12484 3872 12540
rect 3872 12484 3876 12540
rect 3812 12480 3876 12484
rect 8572 12540 8636 12544
rect 8572 12484 8576 12540
rect 8576 12484 8632 12540
rect 8632 12484 8636 12540
rect 8572 12480 8636 12484
rect 8652 12540 8716 12544
rect 8652 12484 8656 12540
rect 8656 12484 8712 12540
rect 8712 12484 8716 12540
rect 8652 12480 8716 12484
rect 8732 12540 8796 12544
rect 8732 12484 8736 12540
rect 8736 12484 8792 12540
rect 8792 12484 8796 12540
rect 8732 12480 8796 12484
rect 8812 12540 8876 12544
rect 8812 12484 8816 12540
rect 8816 12484 8872 12540
rect 8872 12484 8876 12540
rect 8812 12480 8876 12484
rect 13572 12540 13636 12544
rect 13572 12484 13576 12540
rect 13576 12484 13632 12540
rect 13632 12484 13636 12540
rect 13572 12480 13636 12484
rect 13652 12540 13716 12544
rect 13652 12484 13656 12540
rect 13656 12484 13712 12540
rect 13712 12484 13716 12540
rect 13652 12480 13716 12484
rect 13732 12540 13796 12544
rect 13732 12484 13736 12540
rect 13736 12484 13792 12540
rect 13792 12484 13796 12540
rect 13732 12480 13796 12484
rect 13812 12540 13876 12544
rect 13812 12484 13816 12540
rect 13816 12484 13872 12540
rect 13872 12484 13876 12540
rect 13812 12480 13876 12484
rect 18572 12540 18636 12544
rect 18572 12484 18576 12540
rect 18576 12484 18632 12540
rect 18632 12484 18636 12540
rect 18572 12480 18636 12484
rect 18652 12540 18716 12544
rect 18652 12484 18656 12540
rect 18656 12484 18712 12540
rect 18712 12484 18716 12540
rect 18652 12480 18716 12484
rect 18732 12540 18796 12544
rect 18732 12484 18736 12540
rect 18736 12484 18792 12540
rect 18792 12484 18796 12540
rect 18732 12480 18796 12484
rect 18812 12540 18876 12544
rect 18812 12484 18816 12540
rect 18816 12484 18872 12540
rect 18872 12484 18876 12540
rect 18812 12480 18876 12484
rect 23572 12540 23636 12544
rect 23572 12484 23576 12540
rect 23576 12484 23632 12540
rect 23632 12484 23636 12540
rect 23572 12480 23636 12484
rect 23652 12540 23716 12544
rect 23652 12484 23656 12540
rect 23656 12484 23712 12540
rect 23712 12484 23716 12540
rect 23652 12480 23716 12484
rect 23732 12540 23796 12544
rect 23732 12484 23736 12540
rect 23736 12484 23792 12540
rect 23792 12484 23796 12540
rect 23732 12480 23796 12484
rect 23812 12540 23876 12544
rect 23812 12484 23816 12540
rect 23816 12484 23872 12540
rect 23872 12484 23876 12540
rect 23812 12480 23876 12484
rect 28572 12540 28636 12544
rect 28572 12484 28576 12540
rect 28576 12484 28632 12540
rect 28632 12484 28636 12540
rect 28572 12480 28636 12484
rect 28652 12540 28716 12544
rect 28652 12484 28656 12540
rect 28656 12484 28712 12540
rect 28712 12484 28716 12540
rect 28652 12480 28716 12484
rect 28732 12540 28796 12544
rect 28732 12484 28736 12540
rect 28736 12484 28792 12540
rect 28792 12484 28796 12540
rect 28732 12480 28796 12484
rect 28812 12540 28876 12544
rect 28812 12484 28816 12540
rect 28816 12484 28872 12540
rect 28872 12484 28876 12540
rect 28812 12480 28876 12484
rect 33572 12540 33636 12544
rect 33572 12484 33576 12540
rect 33576 12484 33632 12540
rect 33632 12484 33636 12540
rect 33572 12480 33636 12484
rect 33652 12540 33716 12544
rect 33652 12484 33656 12540
rect 33656 12484 33712 12540
rect 33712 12484 33716 12540
rect 33652 12480 33716 12484
rect 33732 12540 33796 12544
rect 33732 12484 33736 12540
rect 33736 12484 33792 12540
rect 33792 12484 33796 12540
rect 33732 12480 33796 12484
rect 33812 12540 33876 12544
rect 33812 12484 33816 12540
rect 33816 12484 33872 12540
rect 33872 12484 33876 12540
rect 33812 12480 33876 12484
rect 38572 12540 38636 12544
rect 38572 12484 38576 12540
rect 38576 12484 38632 12540
rect 38632 12484 38636 12540
rect 38572 12480 38636 12484
rect 38652 12540 38716 12544
rect 38652 12484 38656 12540
rect 38656 12484 38712 12540
rect 38712 12484 38716 12540
rect 38652 12480 38716 12484
rect 38732 12540 38796 12544
rect 38732 12484 38736 12540
rect 38736 12484 38792 12540
rect 38792 12484 38796 12540
rect 38732 12480 38796 12484
rect 38812 12540 38876 12544
rect 38812 12484 38816 12540
rect 38816 12484 38872 12540
rect 38872 12484 38876 12540
rect 38812 12480 38876 12484
rect 43572 12540 43636 12544
rect 43572 12484 43576 12540
rect 43576 12484 43632 12540
rect 43632 12484 43636 12540
rect 43572 12480 43636 12484
rect 43652 12540 43716 12544
rect 43652 12484 43656 12540
rect 43656 12484 43712 12540
rect 43712 12484 43716 12540
rect 43652 12480 43716 12484
rect 43732 12540 43796 12544
rect 43732 12484 43736 12540
rect 43736 12484 43792 12540
rect 43792 12484 43796 12540
rect 43732 12480 43796 12484
rect 43812 12540 43876 12544
rect 43812 12484 43816 12540
rect 43816 12484 43872 12540
rect 43872 12484 43876 12540
rect 43812 12480 43876 12484
rect 30788 12276 30852 12340
rect 6072 11996 6136 12000
rect 6072 11940 6076 11996
rect 6076 11940 6132 11996
rect 6132 11940 6136 11996
rect 6072 11936 6136 11940
rect 6152 11996 6216 12000
rect 6152 11940 6156 11996
rect 6156 11940 6212 11996
rect 6212 11940 6216 11996
rect 6152 11936 6216 11940
rect 6232 11996 6296 12000
rect 6232 11940 6236 11996
rect 6236 11940 6292 11996
rect 6292 11940 6296 11996
rect 6232 11936 6296 11940
rect 6312 11996 6376 12000
rect 6312 11940 6316 11996
rect 6316 11940 6372 11996
rect 6372 11940 6376 11996
rect 6312 11936 6376 11940
rect 11072 11996 11136 12000
rect 11072 11940 11076 11996
rect 11076 11940 11132 11996
rect 11132 11940 11136 11996
rect 11072 11936 11136 11940
rect 11152 11996 11216 12000
rect 11152 11940 11156 11996
rect 11156 11940 11212 11996
rect 11212 11940 11216 11996
rect 11152 11936 11216 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 16072 11996 16136 12000
rect 16072 11940 16076 11996
rect 16076 11940 16132 11996
rect 16132 11940 16136 11996
rect 16072 11936 16136 11940
rect 16152 11996 16216 12000
rect 16152 11940 16156 11996
rect 16156 11940 16212 11996
rect 16212 11940 16216 11996
rect 16152 11936 16216 11940
rect 16232 11996 16296 12000
rect 16232 11940 16236 11996
rect 16236 11940 16292 11996
rect 16292 11940 16296 11996
rect 16232 11936 16296 11940
rect 16312 11996 16376 12000
rect 16312 11940 16316 11996
rect 16316 11940 16372 11996
rect 16372 11940 16376 11996
rect 16312 11936 16376 11940
rect 21072 11996 21136 12000
rect 21072 11940 21076 11996
rect 21076 11940 21132 11996
rect 21132 11940 21136 11996
rect 21072 11936 21136 11940
rect 21152 11996 21216 12000
rect 21152 11940 21156 11996
rect 21156 11940 21212 11996
rect 21212 11940 21216 11996
rect 21152 11936 21216 11940
rect 21232 11996 21296 12000
rect 21232 11940 21236 11996
rect 21236 11940 21292 11996
rect 21292 11940 21296 11996
rect 21232 11936 21296 11940
rect 21312 11996 21376 12000
rect 21312 11940 21316 11996
rect 21316 11940 21372 11996
rect 21372 11940 21376 11996
rect 21312 11936 21376 11940
rect 26072 11996 26136 12000
rect 26072 11940 26076 11996
rect 26076 11940 26132 11996
rect 26132 11940 26136 11996
rect 26072 11936 26136 11940
rect 26152 11996 26216 12000
rect 26152 11940 26156 11996
rect 26156 11940 26212 11996
rect 26212 11940 26216 11996
rect 26152 11936 26216 11940
rect 26232 11996 26296 12000
rect 26232 11940 26236 11996
rect 26236 11940 26292 11996
rect 26292 11940 26296 11996
rect 26232 11936 26296 11940
rect 26312 11996 26376 12000
rect 26312 11940 26316 11996
rect 26316 11940 26372 11996
rect 26372 11940 26376 11996
rect 26312 11936 26376 11940
rect 31072 11996 31136 12000
rect 31072 11940 31076 11996
rect 31076 11940 31132 11996
rect 31132 11940 31136 11996
rect 31072 11936 31136 11940
rect 31152 11996 31216 12000
rect 31152 11940 31156 11996
rect 31156 11940 31212 11996
rect 31212 11940 31216 11996
rect 31152 11936 31216 11940
rect 31232 11996 31296 12000
rect 31232 11940 31236 11996
rect 31236 11940 31292 11996
rect 31292 11940 31296 11996
rect 31232 11936 31296 11940
rect 31312 11996 31376 12000
rect 31312 11940 31316 11996
rect 31316 11940 31372 11996
rect 31372 11940 31376 11996
rect 31312 11936 31376 11940
rect 36072 11996 36136 12000
rect 36072 11940 36076 11996
rect 36076 11940 36132 11996
rect 36132 11940 36136 11996
rect 36072 11936 36136 11940
rect 36152 11996 36216 12000
rect 36152 11940 36156 11996
rect 36156 11940 36212 11996
rect 36212 11940 36216 11996
rect 36152 11936 36216 11940
rect 36232 11996 36296 12000
rect 36232 11940 36236 11996
rect 36236 11940 36292 11996
rect 36292 11940 36296 11996
rect 36232 11936 36296 11940
rect 36312 11996 36376 12000
rect 36312 11940 36316 11996
rect 36316 11940 36372 11996
rect 36372 11940 36376 11996
rect 36312 11936 36376 11940
rect 41072 11996 41136 12000
rect 41072 11940 41076 11996
rect 41076 11940 41132 11996
rect 41132 11940 41136 11996
rect 41072 11936 41136 11940
rect 41152 11996 41216 12000
rect 41152 11940 41156 11996
rect 41156 11940 41212 11996
rect 41212 11940 41216 11996
rect 41152 11936 41216 11940
rect 41232 11996 41296 12000
rect 41232 11940 41236 11996
rect 41236 11940 41292 11996
rect 41292 11940 41296 11996
rect 41232 11936 41296 11940
rect 41312 11996 41376 12000
rect 41312 11940 41316 11996
rect 41316 11940 41372 11996
rect 41372 11940 41376 11996
rect 41312 11936 41376 11940
rect 3572 11452 3636 11456
rect 3572 11396 3576 11452
rect 3576 11396 3632 11452
rect 3632 11396 3636 11452
rect 3572 11392 3636 11396
rect 3652 11452 3716 11456
rect 3652 11396 3656 11452
rect 3656 11396 3712 11452
rect 3712 11396 3716 11452
rect 3652 11392 3716 11396
rect 3732 11452 3796 11456
rect 3732 11396 3736 11452
rect 3736 11396 3792 11452
rect 3792 11396 3796 11452
rect 3732 11392 3796 11396
rect 3812 11452 3876 11456
rect 3812 11396 3816 11452
rect 3816 11396 3872 11452
rect 3872 11396 3876 11452
rect 3812 11392 3876 11396
rect 8572 11452 8636 11456
rect 8572 11396 8576 11452
rect 8576 11396 8632 11452
rect 8632 11396 8636 11452
rect 8572 11392 8636 11396
rect 8652 11452 8716 11456
rect 8652 11396 8656 11452
rect 8656 11396 8712 11452
rect 8712 11396 8716 11452
rect 8652 11392 8716 11396
rect 8732 11452 8796 11456
rect 8732 11396 8736 11452
rect 8736 11396 8792 11452
rect 8792 11396 8796 11452
rect 8732 11392 8796 11396
rect 8812 11452 8876 11456
rect 8812 11396 8816 11452
rect 8816 11396 8872 11452
rect 8872 11396 8876 11452
rect 8812 11392 8876 11396
rect 13572 11452 13636 11456
rect 13572 11396 13576 11452
rect 13576 11396 13632 11452
rect 13632 11396 13636 11452
rect 13572 11392 13636 11396
rect 13652 11452 13716 11456
rect 13652 11396 13656 11452
rect 13656 11396 13712 11452
rect 13712 11396 13716 11452
rect 13652 11392 13716 11396
rect 13732 11452 13796 11456
rect 13732 11396 13736 11452
rect 13736 11396 13792 11452
rect 13792 11396 13796 11452
rect 13732 11392 13796 11396
rect 13812 11452 13876 11456
rect 13812 11396 13816 11452
rect 13816 11396 13872 11452
rect 13872 11396 13876 11452
rect 13812 11392 13876 11396
rect 18572 11452 18636 11456
rect 18572 11396 18576 11452
rect 18576 11396 18632 11452
rect 18632 11396 18636 11452
rect 18572 11392 18636 11396
rect 18652 11452 18716 11456
rect 18652 11396 18656 11452
rect 18656 11396 18712 11452
rect 18712 11396 18716 11452
rect 18652 11392 18716 11396
rect 18732 11452 18796 11456
rect 18732 11396 18736 11452
rect 18736 11396 18792 11452
rect 18792 11396 18796 11452
rect 18732 11392 18796 11396
rect 18812 11452 18876 11456
rect 18812 11396 18816 11452
rect 18816 11396 18872 11452
rect 18872 11396 18876 11452
rect 18812 11392 18876 11396
rect 23572 11452 23636 11456
rect 23572 11396 23576 11452
rect 23576 11396 23632 11452
rect 23632 11396 23636 11452
rect 23572 11392 23636 11396
rect 23652 11452 23716 11456
rect 23652 11396 23656 11452
rect 23656 11396 23712 11452
rect 23712 11396 23716 11452
rect 23652 11392 23716 11396
rect 23732 11452 23796 11456
rect 23732 11396 23736 11452
rect 23736 11396 23792 11452
rect 23792 11396 23796 11452
rect 23732 11392 23796 11396
rect 23812 11452 23876 11456
rect 23812 11396 23816 11452
rect 23816 11396 23872 11452
rect 23872 11396 23876 11452
rect 23812 11392 23876 11396
rect 28572 11452 28636 11456
rect 28572 11396 28576 11452
rect 28576 11396 28632 11452
rect 28632 11396 28636 11452
rect 28572 11392 28636 11396
rect 28652 11452 28716 11456
rect 28652 11396 28656 11452
rect 28656 11396 28712 11452
rect 28712 11396 28716 11452
rect 28652 11392 28716 11396
rect 28732 11452 28796 11456
rect 28732 11396 28736 11452
rect 28736 11396 28792 11452
rect 28792 11396 28796 11452
rect 28732 11392 28796 11396
rect 28812 11452 28876 11456
rect 28812 11396 28816 11452
rect 28816 11396 28872 11452
rect 28872 11396 28876 11452
rect 28812 11392 28876 11396
rect 33572 11452 33636 11456
rect 33572 11396 33576 11452
rect 33576 11396 33632 11452
rect 33632 11396 33636 11452
rect 33572 11392 33636 11396
rect 33652 11452 33716 11456
rect 33652 11396 33656 11452
rect 33656 11396 33712 11452
rect 33712 11396 33716 11452
rect 33652 11392 33716 11396
rect 33732 11452 33796 11456
rect 33732 11396 33736 11452
rect 33736 11396 33792 11452
rect 33792 11396 33796 11452
rect 33732 11392 33796 11396
rect 33812 11452 33876 11456
rect 33812 11396 33816 11452
rect 33816 11396 33872 11452
rect 33872 11396 33876 11452
rect 33812 11392 33876 11396
rect 38572 11452 38636 11456
rect 38572 11396 38576 11452
rect 38576 11396 38632 11452
rect 38632 11396 38636 11452
rect 38572 11392 38636 11396
rect 38652 11452 38716 11456
rect 38652 11396 38656 11452
rect 38656 11396 38712 11452
rect 38712 11396 38716 11452
rect 38652 11392 38716 11396
rect 38732 11452 38796 11456
rect 38732 11396 38736 11452
rect 38736 11396 38792 11452
rect 38792 11396 38796 11452
rect 38732 11392 38796 11396
rect 38812 11452 38876 11456
rect 38812 11396 38816 11452
rect 38816 11396 38872 11452
rect 38872 11396 38876 11452
rect 38812 11392 38876 11396
rect 43572 11452 43636 11456
rect 43572 11396 43576 11452
rect 43576 11396 43632 11452
rect 43632 11396 43636 11452
rect 43572 11392 43636 11396
rect 43652 11452 43716 11456
rect 43652 11396 43656 11452
rect 43656 11396 43712 11452
rect 43712 11396 43716 11452
rect 43652 11392 43716 11396
rect 43732 11452 43796 11456
rect 43732 11396 43736 11452
rect 43736 11396 43792 11452
rect 43792 11396 43796 11452
rect 43732 11392 43796 11396
rect 43812 11452 43876 11456
rect 43812 11396 43816 11452
rect 43816 11396 43872 11452
rect 43872 11396 43876 11452
rect 43812 11392 43876 11396
rect 19012 11248 19076 11252
rect 19012 11192 19062 11248
rect 19062 11192 19076 11248
rect 19012 11188 19076 11192
rect 30788 11112 30852 11116
rect 30788 11056 30838 11112
rect 30838 11056 30852 11112
rect 30788 11052 30852 11056
rect 29316 10976 29380 10980
rect 29316 10920 29366 10976
rect 29366 10920 29380 10976
rect 29316 10916 29380 10920
rect 6072 10908 6136 10912
rect 6072 10852 6076 10908
rect 6076 10852 6132 10908
rect 6132 10852 6136 10908
rect 6072 10848 6136 10852
rect 6152 10908 6216 10912
rect 6152 10852 6156 10908
rect 6156 10852 6212 10908
rect 6212 10852 6216 10908
rect 6152 10848 6216 10852
rect 6232 10908 6296 10912
rect 6232 10852 6236 10908
rect 6236 10852 6292 10908
rect 6292 10852 6296 10908
rect 6232 10848 6296 10852
rect 6312 10908 6376 10912
rect 6312 10852 6316 10908
rect 6316 10852 6372 10908
rect 6372 10852 6376 10908
rect 6312 10848 6376 10852
rect 11072 10908 11136 10912
rect 11072 10852 11076 10908
rect 11076 10852 11132 10908
rect 11132 10852 11136 10908
rect 11072 10848 11136 10852
rect 11152 10908 11216 10912
rect 11152 10852 11156 10908
rect 11156 10852 11212 10908
rect 11212 10852 11216 10908
rect 11152 10848 11216 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 16072 10908 16136 10912
rect 16072 10852 16076 10908
rect 16076 10852 16132 10908
rect 16132 10852 16136 10908
rect 16072 10848 16136 10852
rect 16152 10908 16216 10912
rect 16152 10852 16156 10908
rect 16156 10852 16212 10908
rect 16212 10852 16216 10908
rect 16152 10848 16216 10852
rect 16232 10908 16296 10912
rect 16232 10852 16236 10908
rect 16236 10852 16292 10908
rect 16292 10852 16296 10908
rect 16232 10848 16296 10852
rect 16312 10908 16376 10912
rect 16312 10852 16316 10908
rect 16316 10852 16372 10908
rect 16372 10852 16376 10908
rect 16312 10848 16376 10852
rect 21072 10908 21136 10912
rect 21072 10852 21076 10908
rect 21076 10852 21132 10908
rect 21132 10852 21136 10908
rect 21072 10848 21136 10852
rect 21152 10908 21216 10912
rect 21152 10852 21156 10908
rect 21156 10852 21212 10908
rect 21212 10852 21216 10908
rect 21152 10848 21216 10852
rect 21232 10908 21296 10912
rect 21232 10852 21236 10908
rect 21236 10852 21292 10908
rect 21292 10852 21296 10908
rect 21232 10848 21296 10852
rect 21312 10908 21376 10912
rect 21312 10852 21316 10908
rect 21316 10852 21372 10908
rect 21372 10852 21376 10908
rect 21312 10848 21376 10852
rect 26072 10908 26136 10912
rect 26072 10852 26076 10908
rect 26076 10852 26132 10908
rect 26132 10852 26136 10908
rect 26072 10848 26136 10852
rect 26152 10908 26216 10912
rect 26152 10852 26156 10908
rect 26156 10852 26212 10908
rect 26212 10852 26216 10908
rect 26152 10848 26216 10852
rect 26232 10908 26296 10912
rect 26232 10852 26236 10908
rect 26236 10852 26292 10908
rect 26292 10852 26296 10908
rect 26232 10848 26296 10852
rect 26312 10908 26376 10912
rect 26312 10852 26316 10908
rect 26316 10852 26372 10908
rect 26372 10852 26376 10908
rect 26312 10848 26376 10852
rect 31072 10908 31136 10912
rect 31072 10852 31076 10908
rect 31076 10852 31132 10908
rect 31132 10852 31136 10908
rect 31072 10848 31136 10852
rect 31152 10908 31216 10912
rect 31152 10852 31156 10908
rect 31156 10852 31212 10908
rect 31212 10852 31216 10908
rect 31152 10848 31216 10852
rect 31232 10908 31296 10912
rect 31232 10852 31236 10908
rect 31236 10852 31292 10908
rect 31292 10852 31296 10908
rect 31232 10848 31296 10852
rect 31312 10908 31376 10912
rect 31312 10852 31316 10908
rect 31316 10852 31372 10908
rect 31372 10852 31376 10908
rect 31312 10848 31376 10852
rect 36072 10908 36136 10912
rect 36072 10852 36076 10908
rect 36076 10852 36132 10908
rect 36132 10852 36136 10908
rect 36072 10848 36136 10852
rect 36152 10908 36216 10912
rect 36152 10852 36156 10908
rect 36156 10852 36212 10908
rect 36212 10852 36216 10908
rect 36152 10848 36216 10852
rect 36232 10908 36296 10912
rect 36232 10852 36236 10908
rect 36236 10852 36292 10908
rect 36292 10852 36296 10908
rect 36232 10848 36296 10852
rect 36312 10908 36376 10912
rect 36312 10852 36316 10908
rect 36316 10852 36372 10908
rect 36372 10852 36376 10908
rect 36312 10848 36376 10852
rect 41072 10908 41136 10912
rect 41072 10852 41076 10908
rect 41076 10852 41132 10908
rect 41132 10852 41136 10908
rect 41072 10848 41136 10852
rect 41152 10908 41216 10912
rect 41152 10852 41156 10908
rect 41156 10852 41212 10908
rect 41212 10852 41216 10908
rect 41152 10848 41216 10852
rect 41232 10908 41296 10912
rect 41232 10852 41236 10908
rect 41236 10852 41292 10908
rect 41292 10852 41296 10908
rect 41232 10848 41296 10852
rect 41312 10908 41376 10912
rect 41312 10852 41316 10908
rect 41316 10852 41372 10908
rect 41372 10852 41376 10908
rect 41312 10848 41376 10852
rect 3572 10364 3636 10368
rect 3572 10308 3576 10364
rect 3576 10308 3632 10364
rect 3632 10308 3636 10364
rect 3572 10304 3636 10308
rect 3652 10364 3716 10368
rect 3652 10308 3656 10364
rect 3656 10308 3712 10364
rect 3712 10308 3716 10364
rect 3652 10304 3716 10308
rect 3732 10364 3796 10368
rect 3732 10308 3736 10364
rect 3736 10308 3792 10364
rect 3792 10308 3796 10364
rect 3732 10304 3796 10308
rect 3812 10364 3876 10368
rect 3812 10308 3816 10364
rect 3816 10308 3872 10364
rect 3872 10308 3876 10364
rect 3812 10304 3876 10308
rect 8572 10364 8636 10368
rect 8572 10308 8576 10364
rect 8576 10308 8632 10364
rect 8632 10308 8636 10364
rect 8572 10304 8636 10308
rect 8652 10364 8716 10368
rect 8652 10308 8656 10364
rect 8656 10308 8712 10364
rect 8712 10308 8716 10364
rect 8652 10304 8716 10308
rect 8732 10364 8796 10368
rect 8732 10308 8736 10364
rect 8736 10308 8792 10364
rect 8792 10308 8796 10364
rect 8732 10304 8796 10308
rect 8812 10364 8876 10368
rect 8812 10308 8816 10364
rect 8816 10308 8872 10364
rect 8872 10308 8876 10364
rect 8812 10304 8876 10308
rect 13572 10364 13636 10368
rect 13572 10308 13576 10364
rect 13576 10308 13632 10364
rect 13632 10308 13636 10364
rect 13572 10304 13636 10308
rect 13652 10364 13716 10368
rect 13652 10308 13656 10364
rect 13656 10308 13712 10364
rect 13712 10308 13716 10364
rect 13652 10304 13716 10308
rect 13732 10364 13796 10368
rect 13732 10308 13736 10364
rect 13736 10308 13792 10364
rect 13792 10308 13796 10364
rect 13732 10304 13796 10308
rect 13812 10364 13876 10368
rect 13812 10308 13816 10364
rect 13816 10308 13872 10364
rect 13872 10308 13876 10364
rect 13812 10304 13876 10308
rect 18572 10364 18636 10368
rect 18572 10308 18576 10364
rect 18576 10308 18632 10364
rect 18632 10308 18636 10364
rect 18572 10304 18636 10308
rect 18652 10364 18716 10368
rect 18652 10308 18656 10364
rect 18656 10308 18712 10364
rect 18712 10308 18716 10364
rect 18652 10304 18716 10308
rect 18732 10364 18796 10368
rect 18732 10308 18736 10364
rect 18736 10308 18792 10364
rect 18792 10308 18796 10364
rect 18732 10304 18796 10308
rect 18812 10364 18876 10368
rect 18812 10308 18816 10364
rect 18816 10308 18872 10364
rect 18872 10308 18876 10364
rect 18812 10304 18876 10308
rect 23572 10364 23636 10368
rect 23572 10308 23576 10364
rect 23576 10308 23632 10364
rect 23632 10308 23636 10364
rect 23572 10304 23636 10308
rect 23652 10364 23716 10368
rect 23652 10308 23656 10364
rect 23656 10308 23712 10364
rect 23712 10308 23716 10364
rect 23652 10304 23716 10308
rect 23732 10364 23796 10368
rect 23732 10308 23736 10364
rect 23736 10308 23792 10364
rect 23792 10308 23796 10364
rect 23732 10304 23796 10308
rect 23812 10364 23876 10368
rect 23812 10308 23816 10364
rect 23816 10308 23872 10364
rect 23872 10308 23876 10364
rect 23812 10304 23876 10308
rect 28572 10364 28636 10368
rect 28572 10308 28576 10364
rect 28576 10308 28632 10364
rect 28632 10308 28636 10364
rect 28572 10304 28636 10308
rect 28652 10364 28716 10368
rect 28652 10308 28656 10364
rect 28656 10308 28712 10364
rect 28712 10308 28716 10364
rect 28652 10304 28716 10308
rect 28732 10364 28796 10368
rect 28732 10308 28736 10364
rect 28736 10308 28792 10364
rect 28792 10308 28796 10364
rect 28732 10304 28796 10308
rect 28812 10364 28876 10368
rect 28812 10308 28816 10364
rect 28816 10308 28872 10364
rect 28872 10308 28876 10364
rect 28812 10304 28876 10308
rect 33572 10364 33636 10368
rect 33572 10308 33576 10364
rect 33576 10308 33632 10364
rect 33632 10308 33636 10364
rect 33572 10304 33636 10308
rect 33652 10364 33716 10368
rect 33652 10308 33656 10364
rect 33656 10308 33712 10364
rect 33712 10308 33716 10364
rect 33652 10304 33716 10308
rect 33732 10364 33796 10368
rect 33732 10308 33736 10364
rect 33736 10308 33792 10364
rect 33792 10308 33796 10364
rect 33732 10304 33796 10308
rect 33812 10364 33876 10368
rect 33812 10308 33816 10364
rect 33816 10308 33872 10364
rect 33872 10308 33876 10364
rect 33812 10304 33876 10308
rect 38572 10364 38636 10368
rect 38572 10308 38576 10364
rect 38576 10308 38632 10364
rect 38632 10308 38636 10364
rect 38572 10304 38636 10308
rect 38652 10364 38716 10368
rect 38652 10308 38656 10364
rect 38656 10308 38712 10364
rect 38712 10308 38716 10364
rect 38652 10304 38716 10308
rect 38732 10364 38796 10368
rect 38732 10308 38736 10364
rect 38736 10308 38792 10364
rect 38792 10308 38796 10364
rect 38732 10304 38796 10308
rect 38812 10364 38876 10368
rect 38812 10308 38816 10364
rect 38816 10308 38872 10364
rect 38872 10308 38876 10364
rect 38812 10304 38876 10308
rect 43572 10364 43636 10368
rect 43572 10308 43576 10364
rect 43576 10308 43632 10364
rect 43632 10308 43636 10364
rect 43572 10304 43636 10308
rect 43652 10364 43716 10368
rect 43652 10308 43656 10364
rect 43656 10308 43712 10364
rect 43712 10308 43716 10364
rect 43652 10304 43716 10308
rect 43732 10364 43796 10368
rect 43732 10308 43736 10364
rect 43736 10308 43792 10364
rect 43792 10308 43796 10364
rect 43732 10304 43796 10308
rect 43812 10364 43876 10368
rect 43812 10308 43816 10364
rect 43816 10308 43872 10364
rect 43872 10308 43876 10364
rect 43812 10304 43876 10308
rect 6072 9820 6136 9824
rect 6072 9764 6076 9820
rect 6076 9764 6132 9820
rect 6132 9764 6136 9820
rect 6072 9760 6136 9764
rect 6152 9820 6216 9824
rect 6152 9764 6156 9820
rect 6156 9764 6212 9820
rect 6212 9764 6216 9820
rect 6152 9760 6216 9764
rect 6232 9820 6296 9824
rect 6232 9764 6236 9820
rect 6236 9764 6292 9820
rect 6292 9764 6296 9820
rect 6232 9760 6296 9764
rect 6312 9820 6376 9824
rect 6312 9764 6316 9820
rect 6316 9764 6372 9820
rect 6372 9764 6376 9820
rect 6312 9760 6376 9764
rect 11072 9820 11136 9824
rect 11072 9764 11076 9820
rect 11076 9764 11132 9820
rect 11132 9764 11136 9820
rect 11072 9760 11136 9764
rect 11152 9820 11216 9824
rect 11152 9764 11156 9820
rect 11156 9764 11212 9820
rect 11212 9764 11216 9820
rect 11152 9760 11216 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 16072 9820 16136 9824
rect 16072 9764 16076 9820
rect 16076 9764 16132 9820
rect 16132 9764 16136 9820
rect 16072 9760 16136 9764
rect 16152 9820 16216 9824
rect 16152 9764 16156 9820
rect 16156 9764 16212 9820
rect 16212 9764 16216 9820
rect 16152 9760 16216 9764
rect 16232 9820 16296 9824
rect 16232 9764 16236 9820
rect 16236 9764 16292 9820
rect 16292 9764 16296 9820
rect 16232 9760 16296 9764
rect 16312 9820 16376 9824
rect 16312 9764 16316 9820
rect 16316 9764 16372 9820
rect 16372 9764 16376 9820
rect 16312 9760 16376 9764
rect 21072 9820 21136 9824
rect 21072 9764 21076 9820
rect 21076 9764 21132 9820
rect 21132 9764 21136 9820
rect 21072 9760 21136 9764
rect 21152 9820 21216 9824
rect 21152 9764 21156 9820
rect 21156 9764 21212 9820
rect 21212 9764 21216 9820
rect 21152 9760 21216 9764
rect 21232 9820 21296 9824
rect 21232 9764 21236 9820
rect 21236 9764 21292 9820
rect 21292 9764 21296 9820
rect 21232 9760 21296 9764
rect 21312 9820 21376 9824
rect 21312 9764 21316 9820
rect 21316 9764 21372 9820
rect 21372 9764 21376 9820
rect 21312 9760 21376 9764
rect 26072 9820 26136 9824
rect 26072 9764 26076 9820
rect 26076 9764 26132 9820
rect 26132 9764 26136 9820
rect 26072 9760 26136 9764
rect 26152 9820 26216 9824
rect 26152 9764 26156 9820
rect 26156 9764 26212 9820
rect 26212 9764 26216 9820
rect 26152 9760 26216 9764
rect 26232 9820 26296 9824
rect 26232 9764 26236 9820
rect 26236 9764 26292 9820
rect 26292 9764 26296 9820
rect 26232 9760 26296 9764
rect 26312 9820 26376 9824
rect 26312 9764 26316 9820
rect 26316 9764 26372 9820
rect 26372 9764 26376 9820
rect 26312 9760 26376 9764
rect 31072 9820 31136 9824
rect 31072 9764 31076 9820
rect 31076 9764 31132 9820
rect 31132 9764 31136 9820
rect 31072 9760 31136 9764
rect 31152 9820 31216 9824
rect 31152 9764 31156 9820
rect 31156 9764 31212 9820
rect 31212 9764 31216 9820
rect 31152 9760 31216 9764
rect 31232 9820 31296 9824
rect 31232 9764 31236 9820
rect 31236 9764 31292 9820
rect 31292 9764 31296 9820
rect 31232 9760 31296 9764
rect 31312 9820 31376 9824
rect 31312 9764 31316 9820
rect 31316 9764 31372 9820
rect 31372 9764 31376 9820
rect 31312 9760 31376 9764
rect 36072 9820 36136 9824
rect 36072 9764 36076 9820
rect 36076 9764 36132 9820
rect 36132 9764 36136 9820
rect 36072 9760 36136 9764
rect 36152 9820 36216 9824
rect 36152 9764 36156 9820
rect 36156 9764 36212 9820
rect 36212 9764 36216 9820
rect 36152 9760 36216 9764
rect 36232 9820 36296 9824
rect 36232 9764 36236 9820
rect 36236 9764 36292 9820
rect 36292 9764 36296 9820
rect 36232 9760 36296 9764
rect 36312 9820 36376 9824
rect 36312 9764 36316 9820
rect 36316 9764 36372 9820
rect 36372 9764 36376 9820
rect 36312 9760 36376 9764
rect 41072 9820 41136 9824
rect 41072 9764 41076 9820
rect 41076 9764 41132 9820
rect 41132 9764 41136 9820
rect 41072 9760 41136 9764
rect 41152 9820 41216 9824
rect 41152 9764 41156 9820
rect 41156 9764 41212 9820
rect 41212 9764 41216 9820
rect 41152 9760 41216 9764
rect 41232 9820 41296 9824
rect 41232 9764 41236 9820
rect 41236 9764 41292 9820
rect 41292 9764 41296 9820
rect 41232 9760 41296 9764
rect 41312 9820 41376 9824
rect 41312 9764 41316 9820
rect 41316 9764 41372 9820
rect 41372 9764 41376 9820
rect 41312 9760 41376 9764
rect 30236 9692 30300 9756
rect 28212 9616 28276 9620
rect 28212 9560 28226 9616
rect 28226 9560 28276 9616
rect 28212 9556 28276 9560
rect 32812 9556 32876 9620
rect 3572 9276 3636 9280
rect 3572 9220 3576 9276
rect 3576 9220 3632 9276
rect 3632 9220 3636 9276
rect 3572 9216 3636 9220
rect 3652 9276 3716 9280
rect 3652 9220 3656 9276
rect 3656 9220 3712 9276
rect 3712 9220 3716 9276
rect 3652 9216 3716 9220
rect 3732 9276 3796 9280
rect 3732 9220 3736 9276
rect 3736 9220 3792 9276
rect 3792 9220 3796 9276
rect 3732 9216 3796 9220
rect 3812 9276 3876 9280
rect 3812 9220 3816 9276
rect 3816 9220 3872 9276
rect 3872 9220 3876 9276
rect 3812 9216 3876 9220
rect 8572 9276 8636 9280
rect 8572 9220 8576 9276
rect 8576 9220 8632 9276
rect 8632 9220 8636 9276
rect 8572 9216 8636 9220
rect 8652 9276 8716 9280
rect 8652 9220 8656 9276
rect 8656 9220 8712 9276
rect 8712 9220 8716 9276
rect 8652 9216 8716 9220
rect 8732 9276 8796 9280
rect 8732 9220 8736 9276
rect 8736 9220 8792 9276
rect 8792 9220 8796 9276
rect 8732 9216 8796 9220
rect 8812 9276 8876 9280
rect 8812 9220 8816 9276
rect 8816 9220 8872 9276
rect 8872 9220 8876 9276
rect 8812 9216 8876 9220
rect 13572 9276 13636 9280
rect 13572 9220 13576 9276
rect 13576 9220 13632 9276
rect 13632 9220 13636 9276
rect 13572 9216 13636 9220
rect 13652 9276 13716 9280
rect 13652 9220 13656 9276
rect 13656 9220 13712 9276
rect 13712 9220 13716 9276
rect 13652 9216 13716 9220
rect 13732 9276 13796 9280
rect 13732 9220 13736 9276
rect 13736 9220 13792 9276
rect 13792 9220 13796 9276
rect 13732 9216 13796 9220
rect 13812 9276 13876 9280
rect 13812 9220 13816 9276
rect 13816 9220 13872 9276
rect 13872 9220 13876 9276
rect 13812 9216 13876 9220
rect 18572 9276 18636 9280
rect 18572 9220 18576 9276
rect 18576 9220 18632 9276
rect 18632 9220 18636 9276
rect 18572 9216 18636 9220
rect 18652 9276 18716 9280
rect 18652 9220 18656 9276
rect 18656 9220 18712 9276
rect 18712 9220 18716 9276
rect 18652 9216 18716 9220
rect 18732 9276 18796 9280
rect 18732 9220 18736 9276
rect 18736 9220 18792 9276
rect 18792 9220 18796 9276
rect 18732 9216 18796 9220
rect 18812 9276 18876 9280
rect 18812 9220 18816 9276
rect 18816 9220 18872 9276
rect 18872 9220 18876 9276
rect 18812 9216 18876 9220
rect 23572 9276 23636 9280
rect 23572 9220 23576 9276
rect 23576 9220 23632 9276
rect 23632 9220 23636 9276
rect 23572 9216 23636 9220
rect 23652 9276 23716 9280
rect 23652 9220 23656 9276
rect 23656 9220 23712 9276
rect 23712 9220 23716 9276
rect 23652 9216 23716 9220
rect 23732 9276 23796 9280
rect 23732 9220 23736 9276
rect 23736 9220 23792 9276
rect 23792 9220 23796 9276
rect 23732 9216 23796 9220
rect 23812 9276 23876 9280
rect 23812 9220 23816 9276
rect 23816 9220 23872 9276
rect 23872 9220 23876 9276
rect 23812 9216 23876 9220
rect 28572 9276 28636 9280
rect 28572 9220 28576 9276
rect 28576 9220 28632 9276
rect 28632 9220 28636 9276
rect 28572 9216 28636 9220
rect 28652 9276 28716 9280
rect 28652 9220 28656 9276
rect 28656 9220 28712 9276
rect 28712 9220 28716 9276
rect 28652 9216 28716 9220
rect 28732 9276 28796 9280
rect 28732 9220 28736 9276
rect 28736 9220 28792 9276
rect 28792 9220 28796 9276
rect 28732 9216 28796 9220
rect 28812 9276 28876 9280
rect 28812 9220 28816 9276
rect 28816 9220 28872 9276
rect 28872 9220 28876 9276
rect 28812 9216 28876 9220
rect 33572 9276 33636 9280
rect 33572 9220 33576 9276
rect 33576 9220 33632 9276
rect 33632 9220 33636 9276
rect 33572 9216 33636 9220
rect 33652 9276 33716 9280
rect 33652 9220 33656 9276
rect 33656 9220 33712 9276
rect 33712 9220 33716 9276
rect 33652 9216 33716 9220
rect 33732 9276 33796 9280
rect 33732 9220 33736 9276
rect 33736 9220 33792 9276
rect 33792 9220 33796 9276
rect 33732 9216 33796 9220
rect 33812 9276 33876 9280
rect 33812 9220 33816 9276
rect 33816 9220 33872 9276
rect 33872 9220 33876 9276
rect 33812 9216 33876 9220
rect 38572 9276 38636 9280
rect 38572 9220 38576 9276
rect 38576 9220 38632 9276
rect 38632 9220 38636 9276
rect 38572 9216 38636 9220
rect 38652 9276 38716 9280
rect 38652 9220 38656 9276
rect 38656 9220 38712 9276
rect 38712 9220 38716 9276
rect 38652 9216 38716 9220
rect 38732 9276 38796 9280
rect 38732 9220 38736 9276
rect 38736 9220 38792 9276
rect 38792 9220 38796 9276
rect 38732 9216 38796 9220
rect 38812 9276 38876 9280
rect 38812 9220 38816 9276
rect 38816 9220 38872 9276
rect 38872 9220 38876 9276
rect 38812 9216 38876 9220
rect 43572 9276 43636 9280
rect 43572 9220 43576 9276
rect 43576 9220 43632 9276
rect 43632 9220 43636 9276
rect 43572 9216 43636 9220
rect 43652 9276 43716 9280
rect 43652 9220 43656 9276
rect 43656 9220 43712 9276
rect 43712 9220 43716 9276
rect 43652 9216 43716 9220
rect 43732 9276 43796 9280
rect 43732 9220 43736 9276
rect 43736 9220 43792 9276
rect 43792 9220 43796 9276
rect 43732 9216 43796 9220
rect 43812 9276 43876 9280
rect 43812 9220 43816 9276
rect 43816 9220 43872 9276
rect 43872 9220 43876 9276
rect 43812 9216 43876 9220
rect 6072 8732 6136 8736
rect 6072 8676 6076 8732
rect 6076 8676 6132 8732
rect 6132 8676 6136 8732
rect 6072 8672 6136 8676
rect 6152 8732 6216 8736
rect 6152 8676 6156 8732
rect 6156 8676 6212 8732
rect 6212 8676 6216 8732
rect 6152 8672 6216 8676
rect 6232 8732 6296 8736
rect 6232 8676 6236 8732
rect 6236 8676 6292 8732
rect 6292 8676 6296 8732
rect 6232 8672 6296 8676
rect 6312 8732 6376 8736
rect 6312 8676 6316 8732
rect 6316 8676 6372 8732
rect 6372 8676 6376 8732
rect 6312 8672 6376 8676
rect 11072 8732 11136 8736
rect 11072 8676 11076 8732
rect 11076 8676 11132 8732
rect 11132 8676 11136 8732
rect 11072 8672 11136 8676
rect 11152 8732 11216 8736
rect 11152 8676 11156 8732
rect 11156 8676 11212 8732
rect 11212 8676 11216 8732
rect 11152 8672 11216 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 16072 8732 16136 8736
rect 16072 8676 16076 8732
rect 16076 8676 16132 8732
rect 16132 8676 16136 8732
rect 16072 8672 16136 8676
rect 16152 8732 16216 8736
rect 16152 8676 16156 8732
rect 16156 8676 16212 8732
rect 16212 8676 16216 8732
rect 16152 8672 16216 8676
rect 16232 8732 16296 8736
rect 16232 8676 16236 8732
rect 16236 8676 16292 8732
rect 16292 8676 16296 8732
rect 16232 8672 16296 8676
rect 16312 8732 16376 8736
rect 16312 8676 16316 8732
rect 16316 8676 16372 8732
rect 16372 8676 16376 8732
rect 16312 8672 16376 8676
rect 21072 8732 21136 8736
rect 21072 8676 21076 8732
rect 21076 8676 21132 8732
rect 21132 8676 21136 8732
rect 21072 8672 21136 8676
rect 21152 8732 21216 8736
rect 21152 8676 21156 8732
rect 21156 8676 21212 8732
rect 21212 8676 21216 8732
rect 21152 8672 21216 8676
rect 21232 8732 21296 8736
rect 21232 8676 21236 8732
rect 21236 8676 21292 8732
rect 21292 8676 21296 8732
rect 21232 8672 21296 8676
rect 21312 8732 21376 8736
rect 21312 8676 21316 8732
rect 21316 8676 21372 8732
rect 21372 8676 21376 8732
rect 21312 8672 21376 8676
rect 26072 8732 26136 8736
rect 26072 8676 26076 8732
rect 26076 8676 26132 8732
rect 26132 8676 26136 8732
rect 26072 8672 26136 8676
rect 26152 8732 26216 8736
rect 26152 8676 26156 8732
rect 26156 8676 26212 8732
rect 26212 8676 26216 8732
rect 26152 8672 26216 8676
rect 26232 8732 26296 8736
rect 26232 8676 26236 8732
rect 26236 8676 26292 8732
rect 26292 8676 26296 8732
rect 26232 8672 26296 8676
rect 26312 8732 26376 8736
rect 26312 8676 26316 8732
rect 26316 8676 26372 8732
rect 26372 8676 26376 8732
rect 26312 8672 26376 8676
rect 31072 8732 31136 8736
rect 31072 8676 31076 8732
rect 31076 8676 31132 8732
rect 31132 8676 31136 8732
rect 31072 8672 31136 8676
rect 31152 8732 31216 8736
rect 31152 8676 31156 8732
rect 31156 8676 31212 8732
rect 31212 8676 31216 8732
rect 31152 8672 31216 8676
rect 31232 8732 31296 8736
rect 31232 8676 31236 8732
rect 31236 8676 31292 8732
rect 31292 8676 31296 8732
rect 31232 8672 31296 8676
rect 31312 8732 31376 8736
rect 31312 8676 31316 8732
rect 31316 8676 31372 8732
rect 31372 8676 31376 8732
rect 31312 8672 31376 8676
rect 36072 8732 36136 8736
rect 36072 8676 36076 8732
rect 36076 8676 36132 8732
rect 36132 8676 36136 8732
rect 36072 8672 36136 8676
rect 36152 8732 36216 8736
rect 36152 8676 36156 8732
rect 36156 8676 36212 8732
rect 36212 8676 36216 8732
rect 36152 8672 36216 8676
rect 36232 8732 36296 8736
rect 36232 8676 36236 8732
rect 36236 8676 36292 8732
rect 36292 8676 36296 8732
rect 36232 8672 36296 8676
rect 36312 8732 36376 8736
rect 36312 8676 36316 8732
rect 36316 8676 36372 8732
rect 36372 8676 36376 8732
rect 36312 8672 36376 8676
rect 41072 8732 41136 8736
rect 41072 8676 41076 8732
rect 41076 8676 41132 8732
rect 41132 8676 41136 8732
rect 41072 8672 41136 8676
rect 41152 8732 41216 8736
rect 41152 8676 41156 8732
rect 41156 8676 41212 8732
rect 41212 8676 41216 8732
rect 41152 8672 41216 8676
rect 41232 8732 41296 8736
rect 41232 8676 41236 8732
rect 41236 8676 41292 8732
rect 41292 8676 41296 8732
rect 41232 8672 41296 8676
rect 41312 8732 41376 8736
rect 41312 8676 41316 8732
rect 41316 8676 41372 8732
rect 41372 8676 41376 8732
rect 41312 8672 41376 8676
rect 34284 8332 34348 8396
rect 34468 8392 34532 8396
rect 34468 8336 34482 8392
rect 34482 8336 34532 8392
rect 34468 8332 34532 8336
rect 3572 8188 3636 8192
rect 3572 8132 3576 8188
rect 3576 8132 3632 8188
rect 3632 8132 3636 8188
rect 3572 8128 3636 8132
rect 3652 8188 3716 8192
rect 3652 8132 3656 8188
rect 3656 8132 3712 8188
rect 3712 8132 3716 8188
rect 3652 8128 3716 8132
rect 3732 8188 3796 8192
rect 3732 8132 3736 8188
rect 3736 8132 3792 8188
rect 3792 8132 3796 8188
rect 3732 8128 3796 8132
rect 3812 8188 3876 8192
rect 3812 8132 3816 8188
rect 3816 8132 3872 8188
rect 3872 8132 3876 8188
rect 3812 8128 3876 8132
rect 8572 8188 8636 8192
rect 8572 8132 8576 8188
rect 8576 8132 8632 8188
rect 8632 8132 8636 8188
rect 8572 8128 8636 8132
rect 8652 8188 8716 8192
rect 8652 8132 8656 8188
rect 8656 8132 8712 8188
rect 8712 8132 8716 8188
rect 8652 8128 8716 8132
rect 8732 8188 8796 8192
rect 8732 8132 8736 8188
rect 8736 8132 8792 8188
rect 8792 8132 8796 8188
rect 8732 8128 8796 8132
rect 8812 8188 8876 8192
rect 8812 8132 8816 8188
rect 8816 8132 8872 8188
rect 8872 8132 8876 8188
rect 8812 8128 8876 8132
rect 13572 8188 13636 8192
rect 13572 8132 13576 8188
rect 13576 8132 13632 8188
rect 13632 8132 13636 8188
rect 13572 8128 13636 8132
rect 13652 8188 13716 8192
rect 13652 8132 13656 8188
rect 13656 8132 13712 8188
rect 13712 8132 13716 8188
rect 13652 8128 13716 8132
rect 13732 8188 13796 8192
rect 13732 8132 13736 8188
rect 13736 8132 13792 8188
rect 13792 8132 13796 8188
rect 13732 8128 13796 8132
rect 13812 8188 13876 8192
rect 13812 8132 13816 8188
rect 13816 8132 13872 8188
rect 13872 8132 13876 8188
rect 13812 8128 13876 8132
rect 18572 8188 18636 8192
rect 18572 8132 18576 8188
rect 18576 8132 18632 8188
rect 18632 8132 18636 8188
rect 18572 8128 18636 8132
rect 18652 8188 18716 8192
rect 18652 8132 18656 8188
rect 18656 8132 18712 8188
rect 18712 8132 18716 8188
rect 18652 8128 18716 8132
rect 18732 8188 18796 8192
rect 18732 8132 18736 8188
rect 18736 8132 18792 8188
rect 18792 8132 18796 8188
rect 18732 8128 18796 8132
rect 18812 8188 18876 8192
rect 18812 8132 18816 8188
rect 18816 8132 18872 8188
rect 18872 8132 18876 8188
rect 18812 8128 18876 8132
rect 23572 8188 23636 8192
rect 23572 8132 23576 8188
rect 23576 8132 23632 8188
rect 23632 8132 23636 8188
rect 23572 8128 23636 8132
rect 23652 8188 23716 8192
rect 23652 8132 23656 8188
rect 23656 8132 23712 8188
rect 23712 8132 23716 8188
rect 23652 8128 23716 8132
rect 23732 8188 23796 8192
rect 23732 8132 23736 8188
rect 23736 8132 23792 8188
rect 23792 8132 23796 8188
rect 23732 8128 23796 8132
rect 23812 8188 23876 8192
rect 23812 8132 23816 8188
rect 23816 8132 23872 8188
rect 23872 8132 23876 8188
rect 23812 8128 23876 8132
rect 28572 8188 28636 8192
rect 28572 8132 28576 8188
rect 28576 8132 28632 8188
rect 28632 8132 28636 8188
rect 28572 8128 28636 8132
rect 28652 8188 28716 8192
rect 28652 8132 28656 8188
rect 28656 8132 28712 8188
rect 28712 8132 28716 8188
rect 28652 8128 28716 8132
rect 28732 8188 28796 8192
rect 28732 8132 28736 8188
rect 28736 8132 28792 8188
rect 28792 8132 28796 8188
rect 28732 8128 28796 8132
rect 28812 8188 28876 8192
rect 28812 8132 28816 8188
rect 28816 8132 28872 8188
rect 28872 8132 28876 8188
rect 28812 8128 28876 8132
rect 33572 8188 33636 8192
rect 33572 8132 33576 8188
rect 33576 8132 33632 8188
rect 33632 8132 33636 8188
rect 33572 8128 33636 8132
rect 33652 8188 33716 8192
rect 33652 8132 33656 8188
rect 33656 8132 33712 8188
rect 33712 8132 33716 8188
rect 33652 8128 33716 8132
rect 33732 8188 33796 8192
rect 33732 8132 33736 8188
rect 33736 8132 33792 8188
rect 33792 8132 33796 8188
rect 33732 8128 33796 8132
rect 33812 8188 33876 8192
rect 33812 8132 33816 8188
rect 33816 8132 33872 8188
rect 33872 8132 33876 8188
rect 33812 8128 33876 8132
rect 38572 8188 38636 8192
rect 38572 8132 38576 8188
rect 38576 8132 38632 8188
rect 38632 8132 38636 8188
rect 38572 8128 38636 8132
rect 38652 8188 38716 8192
rect 38652 8132 38656 8188
rect 38656 8132 38712 8188
rect 38712 8132 38716 8188
rect 38652 8128 38716 8132
rect 38732 8188 38796 8192
rect 38732 8132 38736 8188
rect 38736 8132 38792 8188
rect 38792 8132 38796 8188
rect 38732 8128 38796 8132
rect 38812 8188 38876 8192
rect 38812 8132 38816 8188
rect 38816 8132 38872 8188
rect 38872 8132 38876 8188
rect 38812 8128 38876 8132
rect 43572 8188 43636 8192
rect 43572 8132 43576 8188
rect 43576 8132 43632 8188
rect 43632 8132 43636 8188
rect 43572 8128 43636 8132
rect 43652 8188 43716 8192
rect 43652 8132 43656 8188
rect 43656 8132 43712 8188
rect 43712 8132 43716 8188
rect 43652 8128 43716 8132
rect 43732 8188 43796 8192
rect 43732 8132 43736 8188
rect 43736 8132 43792 8188
rect 43792 8132 43796 8188
rect 43732 8128 43796 8132
rect 43812 8188 43876 8192
rect 43812 8132 43816 8188
rect 43816 8132 43872 8188
rect 43872 8132 43876 8188
rect 43812 8128 43876 8132
rect 25636 7788 25700 7852
rect 6072 7644 6136 7648
rect 6072 7588 6076 7644
rect 6076 7588 6132 7644
rect 6132 7588 6136 7644
rect 6072 7584 6136 7588
rect 6152 7644 6216 7648
rect 6152 7588 6156 7644
rect 6156 7588 6212 7644
rect 6212 7588 6216 7644
rect 6152 7584 6216 7588
rect 6232 7644 6296 7648
rect 6232 7588 6236 7644
rect 6236 7588 6292 7644
rect 6292 7588 6296 7644
rect 6232 7584 6296 7588
rect 6312 7644 6376 7648
rect 6312 7588 6316 7644
rect 6316 7588 6372 7644
rect 6372 7588 6376 7644
rect 6312 7584 6376 7588
rect 11072 7644 11136 7648
rect 11072 7588 11076 7644
rect 11076 7588 11132 7644
rect 11132 7588 11136 7644
rect 11072 7584 11136 7588
rect 11152 7644 11216 7648
rect 11152 7588 11156 7644
rect 11156 7588 11212 7644
rect 11212 7588 11216 7644
rect 11152 7584 11216 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 16072 7644 16136 7648
rect 16072 7588 16076 7644
rect 16076 7588 16132 7644
rect 16132 7588 16136 7644
rect 16072 7584 16136 7588
rect 16152 7644 16216 7648
rect 16152 7588 16156 7644
rect 16156 7588 16212 7644
rect 16212 7588 16216 7644
rect 16152 7584 16216 7588
rect 16232 7644 16296 7648
rect 16232 7588 16236 7644
rect 16236 7588 16292 7644
rect 16292 7588 16296 7644
rect 16232 7584 16296 7588
rect 16312 7644 16376 7648
rect 16312 7588 16316 7644
rect 16316 7588 16372 7644
rect 16372 7588 16376 7644
rect 16312 7584 16376 7588
rect 21072 7644 21136 7648
rect 21072 7588 21076 7644
rect 21076 7588 21132 7644
rect 21132 7588 21136 7644
rect 21072 7584 21136 7588
rect 21152 7644 21216 7648
rect 21152 7588 21156 7644
rect 21156 7588 21212 7644
rect 21212 7588 21216 7644
rect 21152 7584 21216 7588
rect 21232 7644 21296 7648
rect 21232 7588 21236 7644
rect 21236 7588 21292 7644
rect 21292 7588 21296 7644
rect 21232 7584 21296 7588
rect 21312 7644 21376 7648
rect 21312 7588 21316 7644
rect 21316 7588 21372 7644
rect 21372 7588 21376 7644
rect 21312 7584 21376 7588
rect 26072 7644 26136 7648
rect 26072 7588 26076 7644
rect 26076 7588 26132 7644
rect 26132 7588 26136 7644
rect 26072 7584 26136 7588
rect 26152 7644 26216 7648
rect 26152 7588 26156 7644
rect 26156 7588 26212 7644
rect 26212 7588 26216 7644
rect 26152 7584 26216 7588
rect 26232 7644 26296 7648
rect 26232 7588 26236 7644
rect 26236 7588 26292 7644
rect 26292 7588 26296 7644
rect 26232 7584 26296 7588
rect 26312 7644 26376 7648
rect 26312 7588 26316 7644
rect 26316 7588 26372 7644
rect 26372 7588 26376 7644
rect 26312 7584 26376 7588
rect 31072 7644 31136 7648
rect 31072 7588 31076 7644
rect 31076 7588 31132 7644
rect 31132 7588 31136 7644
rect 31072 7584 31136 7588
rect 31152 7644 31216 7648
rect 31152 7588 31156 7644
rect 31156 7588 31212 7644
rect 31212 7588 31216 7644
rect 31152 7584 31216 7588
rect 31232 7644 31296 7648
rect 31232 7588 31236 7644
rect 31236 7588 31292 7644
rect 31292 7588 31296 7644
rect 31232 7584 31296 7588
rect 31312 7644 31376 7648
rect 31312 7588 31316 7644
rect 31316 7588 31372 7644
rect 31372 7588 31376 7644
rect 31312 7584 31376 7588
rect 36072 7644 36136 7648
rect 36072 7588 36076 7644
rect 36076 7588 36132 7644
rect 36132 7588 36136 7644
rect 36072 7584 36136 7588
rect 36152 7644 36216 7648
rect 36152 7588 36156 7644
rect 36156 7588 36212 7644
rect 36212 7588 36216 7644
rect 36152 7584 36216 7588
rect 36232 7644 36296 7648
rect 36232 7588 36236 7644
rect 36236 7588 36292 7644
rect 36292 7588 36296 7644
rect 36232 7584 36296 7588
rect 36312 7644 36376 7648
rect 36312 7588 36316 7644
rect 36316 7588 36372 7644
rect 36372 7588 36376 7644
rect 36312 7584 36376 7588
rect 41072 7644 41136 7648
rect 41072 7588 41076 7644
rect 41076 7588 41132 7644
rect 41132 7588 41136 7644
rect 41072 7584 41136 7588
rect 41152 7644 41216 7648
rect 41152 7588 41156 7644
rect 41156 7588 41212 7644
rect 41212 7588 41216 7644
rect 41152 7584 41216 7588
rect 41232 7644 41296 7648
rect 41232 7588 41236 7644
rect 41236 7588 41292 7644
rect 41292 7588 41296 7644
rect 41232 7584 41296 7588
rect 41312 7644 41376 7648
rect 41312 7588 41316 7644
rect 41316 7588 41372 7644
rect 41372 7588 41376 7644
rect 41312 7584 41376 7588
rect 31892 7244 31956 7308
rect 3572 7100 3636 7104
rect 3572 7044 3576 7100
rect 3576 7044 3632 7100
rect 3632 7044 3636 7100
rect 3572 7040 3636 7044
rect 3652 7100 3716 7104
rect 3652 7044 3656 7100
rect 3656 7044 3712 7100
rect 3712 7044 3716 7100
rect 3652 7040 3716 7044
rect 3732 7100 3796 7104
rect 3732 7044 3736 7100
rect 3736 7044 3792 7100
rect 3792 7044 3796 7100
rect 3732 7040 3796 7044
rect 3812 7100 3876 7104
rect 3812 7044 3816 7100
rect 3816 7044 3872 7100
rect 3872 7044 3876 7100
rect 3812 7040 3876 7044
rect 8572 7100 8636 7104
rect 8572 7044 8576 7100
rect 8576 7044 8632 7100
rect 8632 7044 8636 7100
rect 8572 7040 8636 7044
rect 8652 7100 8716 7104
rect 8652 7044 8656 7100
rect 8656 7044 8712 7100
rect 8712 7044 8716 7100
rect 8652 7040 8716 7044
rect 8732 7100 8796 7104
rect 8732 7044 8736 7100
rect 8736 7044 8792 7100
rect 8792 7044 8796 7100
rect 8732 7040 8796 7044
rect 8812 7100 8876 7104
rect 8812 7044 8816 7100
rect 8816 7044 8872 7100
rect 8872 7044 8876 7100
rect 8812 7040 8876 7044
rect 13572 7100 13636 7104
rect 13572 7044 13576 7100
rect 13576 7044 13632 7100
rect 13632 7044 13636 7100
rect 13572 7040 13636 7044
rect 13652 7100 13716 7104
rect 13652 7044 13656 7100
rect 13656 7044 13712 7100
rect 13712 7044 13716 7100
rect 13652 7040 13716 7044
rect 13732 7100 13796 7104
rect 13732 7044 13736 7100
rect 13736 7044 13792 7100
rect 13792 7044 13796 7100
rect 13732 7040 13796 7044
rect 13812 7100 13876 7104
rect 13812 7044 13816 7100
rect 13816 7044 13872 7100
rect 13872 7044 13876 7100
rect 13812 7040 13876 7044
rect 18572 7100 18636 7104
rect 18572 7044 18576 7100
rect 18576 7044 18632 7100
rect 18632 7044 18636 7100
rect 18572 7040 18636 7044
rect 18652 7100 18716 7104
rect 18652 7044 18656 7100
rect 18656 7044 18712 7100
rect 18712 7044 18716 7100
rect 18652 7040 18716 7044
rect 18732 7100 18796 7104
rect 18732 7044 18736 7100
rect 18736 7044 18792 7100
rect 18792 7044 18796 7100
rect 18732 7040 18796 7044
rect 18812 7100 18876 7104
rect 18812 7044 18816 7100
rect 18816 7044 18872 7100
rect 18872 7044 18876 7100
rect 18812 7040 18876 7044
rect 23572 7100 23636 7104
rect 23572 7044 23576 7100
rect 23576 7044 23632 7100
rect 23632 7044 23636 7100
rect 23572 7040 23636 7044
rect 23652 7100 23716 7104
rect 23652 7044 23656 7100
rect 23656 7044 23712 7100
rect 23712 7044 23716 7100
rect 23652 7040 23716 7044
rect 23732 7100 23796 7104
rect 23732 7044 23736 7100
rect 23736 7044 23792 7100
rect 23792 7044 23796 7100
rect 23732 7040 23796 7044
rect 23812 7100 23876 7104
rect 23812 7044 23816 7100
rect 23816 7044 23872 7100
rect 23872 7044 23876 7100
rect 23812 7040 23876 7044
rect 28572 7100 28636 7104
rect 28572 7044 28576 7100
rect 28576 7044 28632 7100
rect 28632 7044 28636 7100
rect 28572 7040 28636 7044
rect 28652 7100 28716 7104
rect 28652 7044 28656 7100
rect 28656 7044 28712 7100
rect 28712 7044 28716 7100
rect 28652 7040 28716 7044
rect 28732 7100 28796 7104
rect 28732 7044 28736 7100
rect 28736 7044 28792 7100
rect 28792 7044 28796 7100
rect 28732 7040 28796 7044
rect 28812 7100 28876 7104
rect 28812 7044 28816 7100
rect 28816 7044 28872 7100
rect 28872 7044 28876 7100
rect 28812 7040 28876 7044
rect 33572 7100 33636 7104
rect 33572 7044 33576 7100
rect 33576 7044 33632 7100
rect 33632 7044 33636 7100
rect 33572 7040 33636 7044
rect 33652 7100 33716 7104
rect 33652 7044 33656 7100
rect 33656 7044 33712 7100
rect 33712 7044 33716 7100
rect 33652 7040 33716 7044
rect 33732 7100 33796 7104
rect 33732 7044 33736 7100
rect 33736 7044 33792 7100
rect 33792 7044 33796 7100
rect 33732 7040 33796 7044
rect 33812 7100 33876 7104
rect 33812 7044 33816 7100
rect 33816 7044 33872 7100
rect 33872 7044 33876 7100
rect 33812 7040 33876 7044
rect 38572 7100 38636 7104
rect 38572 7044 38576 7100
rect 38576 7044 38632 7100
rect 38632 7044 38636 7100
rect 38572 7040 38636 7044
rect 38652 7100 38716 7104
rect 38652 7044 38656 7100
rect 38656 7044 38712 7100
rect 38712 7044 38716 7100
rect 38652 7040 38716 7044
rect 38732 7100 38796 7104
rect 38732 7044 38736 7100
rect 38736 7044 38792 7100
rect 38792 7044 38796 7100
rect 38732 7040 38796 7044
rect 38812 7100 38876 7104
rect 38812 7044 38816 7100
rect 38816 7044 38872 7100
rect 38872 7044 38876 7100
rect 38812 7040 38876 7044
rect 43572 7100 43636 7104
rect 43572 7044 43576 7100
rect 43576 7044 43632 7100
rect 43632 7044 43636 7100
rect 43572 7040 43636 7044
rect 43652 7100 43716 7104
rect 43652 7044 43656 7100
rect 43656 7044 43712 7100
rect 43712 7044 43716 7100
rect 43652 7040 43716 7044
rect 43732 7100 43796 7104
rect 43732 7044 43736 7100
rect 43736 7044 43792 7100
rect 43792 7044 43796 7100
rect 43732 7040 43796 7044
rect 43812 7100 43876 7104
rect 43812 7044 43816 7100
rect 43816 7044 43872 7100
rect 43872 7044 43876 7100
rect 43812 7040 43876 7044
rect 23060 7032 23124 7036
rect 23060 6976 23074 7032
rect 23074 6976 23124 7032
rect 23060 6972 23124 6976
rect 9260 6896 9324 6900
rect 9260 6840 9274 6896
rect 9274 6840 9324 6896
rect 9260 6836 9324 6840
rect 17540 6836 17604 6900
rect 19748 6896 19812 6900
rect 19748 6840 19798 6896
rect 19798 6840 19812 6896
rect 19748 6836 19812 6840
rect 22876 6836 22940 6900
rect 24348 6896 24412 6900
rect 24348 6840 24362 6896
rect 24362 6840 24412 6896
rect 24348 6836 24412 6840
rect 25820 6836 25884 6900
rect 6072 6556 6136 6560
rect 6072 6500 6076 6556
rect 6076 6500 6132 6556
rect 6132 6500 6136 6556
rect 6072 6496 6136 6500
rect 6152 6556 6216 6560
rect 6152 6500 6156 6556
rect 6156 6500 6212 6556
rect 6212 6500 6216 6556
rect 6152 6496 6216 6500
rect 6232 6556 6296 6560
rect 6232 6500 6236 6556
rect 6236 6500 6292 6556
rect 6292 6500 6296 6556
rect 6232 6496 6296 6500
rect 6312 6556 6376 6560
rect 6312 6500 6316 6556
rect 6316 6500 6372 6556
rect 6372 6500 6376 6556
rect 6312 6496 6376 6500
rect 11072 6556 11136 6560
rect 11072 6500 11076 6556
rect 11076 6500 11132 6556
rect 11132 6500 11136 6556
rect 11072 6496 11136 6500
rect 11152 6556 11216 6560
rect 11152 6500 11156 6556
rect 11156 6500 11212 6556
rect 11212 6500 11216 6556
rect 11152 6496 11216 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 16072 6556 16136 6560
rect 16072 6500 16076 6556
rect 16076 6500 16132 6556
rect 16132 6500 16136 6556
rect 16072 6496 16136 6500
rect 16152 6556 16216 6560
rect 16152 6500 16156 6556
rect 16156 6500 16212 6556
rect 16212 6500 16216 6556
rect 16152 6496 16216 6500
rect 16232 6556 16296 6560
rect 16232 6500 16236 6556
rect 16236 6500 16292 6556
rect 16292 6500 16296 6556
rect 16232 6496 16296 6500
rect 16312 6556 16376 6560
rect 16312 6500 16316 6556
rect 16316 6500 16372 6556
rect 16372 6500 16376 6556
rect 16312 6496 16376 6500
rect 21072 6556 21136 6560
rect 21072 6500 21076 6556
rect 21076 6500 21132 6556
rect 21132 6500 21136 6556
rect 21072 6496 21136 6500
rect 21152 6556 21216 6560
rect 21152 6500 21156 6556
rect 21156 6500 21212 6556
rect 21212 6500 21216 6556
rect 21152 6496 21216 6500
rect 21232 6556 21296 6560
rect 21232 6500 21236 6556
rect 21236 6500 21292 6556
rect 21292 6500 21296 6556
rect 21232 6496 21296 6500
rect 21312 6556 21376 6560
rect 21312 6500 21316 6556
rect 21316 6500 21372 6556
rect 21372 6500 21376 6556
rect 21312 6496 21376 6500
rect 26072 6556 26136 6560
rect 26072 6500 26076 6556
rect 26076 6500 26132 6556
rect 26132 6500 26136 6556
rect 26072 6496 26136 6500
rect 26152 6556 26216 6560
rect 26152 6500 26156 6556
rect 26156 6500 26212 6556
rect 26212 6500 26216 6556
rect 26152 6496 26216 6500
rect 26232 6556 26296 6560
rect 26232 6500 26236 6556
rect 26236 6500 26292 6556
rect 26292 6500 26296 6556
rect 26232 6496 26296 6500
rect 26312 6556 26376 6560
rect 26312 6500 26316 6556
rect 26316 6500 26372 6556
rect 26372 6500 26376 6556
rect 26312 6496 26376 6500
rect 31072 6556 31136 6560
rect 31072 6500 31076 6556
rect 31076 6500 31132 6556
rect 31132 6500 31136 6556
rect 31072 6496 31136 6500
rect 31152 6556 31216 6560
rect 31152 6500 31156 6556
rect 31156 6500 31212 6556
rect 31212 6500 31216 6556
rect 31152 6496 31216 6500
rect 31232 6556 31296 6560
rect 31232 6500 31236 6556
rect 31236 6500 31292 6556
rect 31292 6500 31296 6556
rect 31232 6496 31296 6500
rect 31312 6556 31376 6560
rect 31312 6500 31316 6556
rect 31316 6500 31372 6556
rect 31372 6500 31376 6556
rect 31312 6496 31376 6500
rect 36072 6556 36136 6560
rect 36072 6500 36076 6556
rect 36076 6500 36132 6556
rect 36132 6500 36136 6556
rect 36072 6496 36136 6500
rect 36152 6556 36216 6560
rect 36152 6500 36156 6556
rect 36156 6500 36212 6556
rect 36212 6500 36216 6556
rect 36152 6496 36216 6500
rect 36232 6556 36296 6560
rect 36232 6500 36236 6556
rect 36236 6500 36292 6556
rect 36292 6500 36296 6556
rect 36232 6496 36296 6500
rect 36312 6556 36376 6560
rect 36312 6500 36316 6556
rect 36316 6500 36372 6556
rect 36372 6500 36376 6556
rect 36312 6496 36376 6500
rect 41072 6556 41136 6560
rect 41072 6500 41076 6556
rect 41076 6500 41132 6556
rect 41132 6500 41136 6556
rect 41072 6496 41136 6500
rect 41152 6556 41216 6560
rect 41152 6500 41156 6556
rect 41156 6500 41212 6556
rect 41212 6500 41216 6556
rect 41152 6496 41216 6500
rect 41232 6556 41296 6560
rect 41232 6500 41236 6556
rect 41236 6500 41292 6556
rect 41292 6500 41296 6556
rect 41232 6496 41296 6500
rect 41312 6556 41376 6560
rect 41312 6500 41316 6556
rect 41316 6500 41372 6556
rect 41372 6500 41376 6556
rect 41312 6496 41376 6500
rect 16988 6428 17052 6492
rect 26740 6020 26804 6084
rect 3572 6012 3636 6016
rect 3572 5956 3576 6012
rect 3576 5956 3632 6012
rect 3632 5956 3636 6012
rect 3572 5952 3636 5956
rect 3652 6012 3716 6016
rect 3652 5956 3656 6012
rect 3656 5956 3712 6012
rect 3712 5956 3716 6012
rect 3652 5952 3716 5956
rect 3732 6012 3796 6016
rect 3732 5956 3736 6012
rect 3736 5956 3792 6012
rect 3792 5956 3796 6012
rect 3732 5952 3796 5956
rect 3812 6012 3876 6016
rect 3812 5956 3816 6012
rect 3816 5956 3872 6012
rect 3872 5956 3876 6012
rect 3812 5952 3876 5956
rect 8572 6012 8636 6016
rect 8572 5956 8576 6012
rect 8576 5956 8632 6012
rect 8632 5956 8636 6012
rect 8572 5952 8636 5956
rect 8652 6012 8716 6016
rect 8652 5956 8656 6012
rect 8656 5956 8712 6012
rect 8712 5956 8716 6012
rect 8652 5952 8716 5956
rect 8732 6012 8796 6016
rect 8732 5956 8736 6012
rect 8736 5956 8792 6012
rect 8792 5956 8796 6012
rect 8732 5952 8796 5956
rect 8812 6012 8876 6016
rect 8812 5956 8816 6012
rect 8816 5956 8872 6012
rect 8872 5956 8876 6012
rect 8812 5952 8876 5956
rect 13572 6012 13636 6016
rect 13572 5956 13576 6012
rect 13576 5956 13632 6012
rect 13632 5956 13636 6012
rect 13572 5952 13636 5956
rect 13652 6012 13716 6016
rect 13652 5956 13656 6012
rect 13656 5956 13712 6012
rect 13712 5956 13716 6012
rect 13652 5952 13716 5956
rect 13732 6012 13796 6016
rect 13732 5956 13736 6012
rect 13736 5956 13792 6012
rect 13792 5956 13796 6012
rect 13732 5952 13796 5956
rect 13812 6012 13876 6016
rect 13812 5956 13816 6012
rect 13816 5956 13872 6012
rect 13872 5956 13876 6012
rect 13812 5952 13876 5956
rect 18572 6012 18636 6016
rect 18572 5956 18576 6012
rect 18576 5956 18632 6012
rect 18632 5956 18636 6012
rect 18572 5952 18636 5956
rect 18652 6012 18716 6016
rect 18652 5956 18656 6012
rect 18656 5956 18712 6012
rect 18712 5956 18716 6012
rect 18652 5952 18716 5956
rect 18732 6012 18796 6016
rect 18732 5956 18736 6012
rect 18736 5956 18792 6012
rect 18792 5956 18796 6012
rect 18732 5952 18796 5956
rect 18812 6012 18876 6016
rect 18812 5956 18816 6012
rect 18816 5956 18872 6012
rect 18872 5956 18876 6012
rect 18812 5952 18876 5956
rect 23572 6012 23636 6016
rect 23572 5956 23576 6012
rect 23576 5956 23632 6012
rect 23632 5956 23636 6012
rect 23572 5952 23636 5956
rect 23652 6012 23716 6016
rect 23652 5956 23656 6012
rect 23656 5956 23712 6012
rect 23712 5956 23716 6012
rect 23652 5952 23716 5956
rect 23732 6012 23796 6016
rect 23732 5956 23736 6012
rect 23736 5956 23792 6012
rect 23792 5956 23796 6012
rect 23732 5952 23796 5956
rect 23812 6012 23876 6016
rect 23812 5956 23816 6012
rect 23816 5956 23872 6012
rect 23872 5956 23876 6012
rect 23812 5952 23876 5956
rect 28572 6012 28636 6016
rect 28572 5956 28576 6012
rect 28576 5956 28632 6012
rect 28632 5956 28636 6012
rect 28572 5952 28636 5956
rect 28652 6012 28716 6016
rect 28652 5956 28656 6012
rect 28656 5956 28712 6012
rect 28712 5956 28716 6012
rect 28652 5952 28716 5956
rect 28732 6012 28796 6016
rect 28732 5956 28736 6012
rect 28736 5956 28792 6012
rect 28792 5956 28796 6012
rect 28732 5952 28796 5956
rect 28812 6012 28876 6016
rect 28812 5956 28816 6012
rect 28816 5956 28872 6012
rect 28872 5956 28876 6012
rect 28812 5952 28876 5956
rect 33572 6012 33636 6016
rect 33572 5956 33576 6012
rect 33576 5956 33632 6012
rect 33632 5956 33636 6012
rect 33572 5952 33636 5956
rect 33652 6012 33716 6016
rect 33652 5956 33656 6012
rect 33656 5956 33712 6012
rect 33712 5956 33716 6012
rect 33652 5952 33716 5956
rect 33732 6012 33796 6016
rect 33732 5956 33736 6012
rect 33736 5956 33792 6012
rect 33792 5956 33796 6012
rect 33732 5952 33796 5956
rect 33812 6012 33876 6016
rect 33812 5956 33816 6012
rect 33816 5956 33872 6012
rect 33872 5956 33876 6012
rect 33812 5952 33876 5956
rect 38572 6012 38636 6016
rect 38572 5956 38576 6012
rect 38576 5956 38632 6012
rect 38632 5956 38636 6012
rect 38572 5952 38636 5956
rect 38652 6012 38716 6016
rect 38652 5956 38656 6012
rect 38656 5956 38712 6012
rect 38712 5956 38716 6012
rect 38652 5952 38716 5956
rect 38732 6012 38796 6016
rect 38732 5956 38736 6012
rect 38736 5956 38792 6012
rect 38792 5956 38796 6012
rect 38732 5952 38796 5956
rect 38812 6012 38876 6016
rect 38812 5956 38816 6012
rect 38816 5956 38872 6012
rect 38872 5956 38876 6012
rect 38812 5952 38876 5956
rect 43572 6012 43636 6016
rect 43572 5956 43576 6012
rect 43576 5956 43632 6012
rect 43632 5956 43636 6012
rect 43572 5952 43636 5956
rect 43652 6012 43716 6016
rect 43652 5956 43656 6012
rect 43656 5956 43712 6012
rect 43712 5956 43716 6012
rect 43652 5952 43716 5956
rect 43732 6012 43796 6016
rect 43732 5956 43736 6012
rect 43736 5956 43792 6012
rect 43792 5956 43796 6012
rect 43732 5952 43796 5956
rect 43812 6012 43876 6016
rect 43812 5956 43816 6012
rect 43816 5956 43872 6012
rect 43872 5956 43876 6012
rect 43812 5952 43876 5956
rect 22692 5884 22756 5948
rect 25820 5748 25884 5812
rect 33180 5672 33244 5676
rect 33180 5616 33230 5672
rect 33230 5616 33244 5672
rect 33180 5612 33244 5616
rect 17540 5476 17604 5540
rect 19932 5536 19996 5540
rect 19932 5480 19946 5536
rect 19946 5480 19996 5536
rect 19932 5476 19996 5480
rect 21588 5476 21652 5540
rect 23244 5536 23308 5540
rect 23244 5480 23258 5536
rect 23258 5480 23308 5536
rect 6072 5468 6136 5472
rect 6072 5412 6076 5468
rect 6076 5412 6132 5468
rect 6132 5412 6136 5468
rect 6072 5408 6136 5412
rect 6152 5468 6216 5472
rect 6152 5412 6156 5468
rect 6156 5412 6212 5468
rect 6212 5412 6216 5468
rect 6152 5408 6216 5412
rect 6232 5468 6296 5472
rect 6232 5412 6236 5468
rect 6236 5412 6292 5468
rect 6292 5412 6296 5468
rect 6232 5408 6296 5412
rect 6312 5468 6376 5472
rect 6312 5412 6316 5468
rect 6316 5412 6372 5468
rect 6372 5412 6376 5468
rect 6312 5408 6376 5412
rect 11072 5468 11136 5472
rect 11072 5412 11076 5468
rect 11076 5412 11132 5468
rect 11132 5412 11136 5468
rect 11072 5408 11136 5412
rect 11152 5468 11216 5472
rect 11152 5412 11156 5468
rect 11156 5412 11212 5468
rect 11212 5412 11216 5468
rect 11152 5408 11216 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 16072 5468 16136 5472
rect 16072 5412 16076 5468
rect 16076 5412 16132 5468
rect 16132 5412 16136 5468
rect 16072 5408 16136 5412
rect 16152 5468 16216 5472
rect 16152 5412 16156 5468
rect 16156 5412 16212 5468
rect 16212 5412 16216 5468
rect 16152 5408 16216 5412
rect 16232 5468 16296 5472
rect 16232 5412 16236 5468
rect 16236 5412 16292 5468
rect 16292 5412 16296 5468
rect 16232 5408 16296 5412
rect 16312 5468 16376 5472
rect 16312 5412 16316 5468
rect 16316 5412 16372 5468
rect 16372 5412 16376 5468
rect 16312 5408 16376 5412
rect 21072 5468 21136 5472
rect 21072 5412 21076 5468
rect 21076 5412 21132 5468
rect 21132 5412 21136 5468
rect 21072 5408 21136 5412
rect 21152 5468 21216 5472
rect 21152 5412 21156 5468
rect 21156 5412 21212 5468
rect 21212 5412 21216 5468
rect 21152 5408 21216 5412
rect 21232 5468 21296 5472
rect 21232 5412 21236 5468
rect 21236 5412 21292 5468
rect 21292 5412 21296 5468
rect 21232 5408 21296 5412
rect 21312 5468 21376 5472
rect 21312 5412 21316 5468
rect 21316 5412 21372 5468
rect 21372 5412 21376 5468
rect 21312 5408 21376 5412
rect 21956 5400 22020 5404
rect 21956 5344 22006 5400
rect 22006 5344 22020 5400
rect 21956 5340 22020 5344
rect 23244 5476 23308 5480
rect 25452 5476 25516 5540
rect 26072 5468 26136 5472
rect 26072 5412 26076 5468
rect 26076 5412 26132 5468
rect 26132 5412 26136 5468
rect 26072 5408 26136 5412
rect 26152 5468 26216 5472
rect 26152 5412 26156 5468
rect 26156 5412 26212 5468
rect 26212 5412 26216 5468
rect 26152 5408 26216 5412
rect 26232 5468 26296 5472
rect 26232 5412 26236 5468
rect 26236 5412 26292 5468
rect 26292 5412 26296 5468
rect 26232 5408 26296 5412
rect 26312 5468 26376 5472
rect 26312 5412 26316 5468
rect 26316 5412 26372 5468
rect 26372 5412 26376 5468
rect 26312 5408 26376 5412
rect 31072 5468 31136 5472
rect 31072 5412 31076 5468
rect 31076 5412 31132 5468
rect 31132 5412 31136 5468
rect 31072 5408 31136 5412
rect 31152 5468 31216 5472
rect 31152 5412 31156 5468
rect 31156 5412 31212 5468
rect 31212 5412 31216 5468
rect 31152 5408 31216 5412
rect 31232 5468 31296 5472
rect 31232 5412 31236 5468
rect 31236 5412 31292 5468
rect 31292 5412 31296 5468
rect 31232 5408 31296 5412
rect 31312 5468 31376 5472
rect 31312 5412 31316 5468
rect 31316 5412 31372 5468
rect 31372 5412 31376 5468
rect 31312 5408 31376 5412
rect 36072 5468 36136 5472
rect 36072 5412 36076 5468
rect 36076 5412 36132 5468
rect 36132 5412 36136 5468
rect 36072 5408 36136 5412
rect 36152 5468 36216 5472
rect 36152 5412 36156 5468
rect 36156 5412 36212 5468
rect 36212 5412 36216 5468
rect 36152 5408 36216 5412
rect 36232 5468 36296 5472
rect 36232 5412 36236 5468
rect 36236 5412 36292 5468
rect 36292 5412 36296 5468
rect 36232 5408 36296 5412
rect 36312 5468 36376 5472
rect 36312 5412 36316 5468
rect 36316 5412 36372 5468
rect 36372 5412 36376 5468
rect 36312 5408 36376 5412
rect 41072 5468 41136 5472
rect 41072 5412 41076 5468
rect 41076 5412 41132 5468
rect 41132 5412 41136 5468
rect 41072 5408 41136 5412
rect 41152 5468 41216 5472
rect 41152 5412 41156 5468
rect 41156 5412 41212 5468
rect 41212 5412 41216 5468
rect 41152 5408 41216 5412
rect 41232 5468 41296 5472
rect 41232 5412 41236 5468
rect 41236 5412 41292 5468
rect 41292 5412 41296 5468
rect 41232 5408 41296 5412
rect 41312 5468 41376 5472
rect 41312 5412 41316 5468
rect 41316 5412 41372 5468
rect 41372 5412 41376 5468
rect 41312 5408 41376 5412
rect 19196 5204 19260 5268
rect 26556 5068 26620 5132
rect 3572 4924 3636 4928
rect 3572 4868 3576 4924
rect 3576 4868 3632 4924
rect 3632 4868 3636 4924
rect 3572 4864 3636 4868
rect 3652 4924 3716 4928
rect 3652 4868 3656 4924
rect 3656 4868 3712 4924
rect 3712 4868 3716 4924
rect 3652 4864 3716 4868
rect 3732 4924 3796 4928
rect 3732 4868 3736 4924
rect 3736 4868 3792 4924
rect 3792 4868 3796 4924
rect 3732 4864 3796 4868
rect 3812 4924 3876 4928
rect 3812 4868 3816 4924
rect 3816 4868 3872 4924
rect 3872 4868 3876 4924
rect 3812 4864 3876 4868
rect 8572 4924 8636 4928
rect 8572 4868 8576 4924
rect 8576 4868 8632 4924
rect 8632 4868 8636 4924
rect 8572 4864 8636 4868
rect 8652 4924 8716 4928
rect 8652 4868 8656 4924
rect 8656 4868 8712 4924
rect 8712 4868 8716 4924
rect 8652 4864 8716 4868
rect 8732 4924 8796 4928
rect 8732 4868 8736 4924
rect 8736 4868 8792 4924
rect 8792 4868 8796 4924
rect 8732 4864 8796 4868
rect 8812 4924 8876 4928
rect 8812 4868 8816 4924
rect 8816 4868 8872 4924
rect 8872 4868 8876 4924
rect 8812 4864 8876 4868
rect 13572 4924 13636 4928
rect 13572 4868 13576 4924
rect 13576 4868 13632 4924
rect 13632 4868 13636 4924
rect 13572 4864 13636 4868
rect 13652 4924 13716 4928
rect 13652 4868 13656 4924
rect 13656 4868 13712 4924
rect 13712 4868 13716 4924
rect 13652 4864 13716 4868
rect 13732 4924 13796 4928
rect 13732 4868 13736 4924
rect 13736 4868 13792 4924
rect 13792 4868 13796 4924
rect 13732 4864 13796 4868
rect 13812 4924 13876 4928
rect 13812 4868 13816 4924
rect 13816 4868 13872 4924
rect 13872 4868 13876 4924
rect 13812 4864 13876 4868
rect 18572 4924 18636 4928
rect 18572 4868 18576 4924
rect 18576 4868 18632 4924
rect 18632 4868 18636 4924
rect 18572 4864 18636 4868
rect 18652 4924 18716 4928
rect 18652 4868 18656 4924
rect 18656 4868 18712 4924
rect 18712 4868 18716 4924
rect 18652 4864 18716 4868
rect 18732 4924 18796 4928
rect 18732 4868 18736 4924
rect 18736 4868 18792 4924
rect 18792 4868 18796 4924
rect 18732 4864 18796 4868
rect 18812 4924 18876 4928
rect 18812 4868 18816 4924
rect 18816 4868 18872 4924
rect 18872 4868 18876 4924
rect 18812 4864 18876 4868
rect 23572 4924 23636 4928
rect 23572 4868 23576 4924
rect 23576 4868 23632 4924
rect 23632 4868 23636 4924
rect 23572 4864 23636 4868
rect 23652 4924 23716 4928
rect 23652 4868 23656 4924
rect 23656 4868 23712 4924
rect 23712 4868 23716 4924
rect 23652 4864 23716 4868
rect 23732 4924 23796 4928
rect 23732 4868 23736 4924
rect 23736 4868 23792 4924
rect 23792 4868 23796 4924
rect 23732 4864 23796 4868
rect 23812 4924 23876 4928
rect 23812 4868 23816 4924
rect 23816 4868 23872 4924
rect 23872 4868 23876 4924
rect 23812 4864 23876 4868
rect 28572 4924 28636 4928
rect 28572 4868 28576 4924
rect 28576 4868 28632 4924
rect 28632 4868 28636 4924
rect 28572 4864 28636 4868
rect 28652 4924 28716 4928
rect 28652 4868 28656 4924
rect 28656 4868 28712 4924
rect 28712 4868 28716 4924
rect 28652 4864 28716 4868
rect 28732 4924 28796 4928
rect 28732 4868 28736 4924
rect 28736 4868 28792 4924
rect 28792 4868 28796 4924
rect 28732 4864 28796 4868
rect 28812 4924 28876 4928
rect 28812 4868 28816 4924
rect 28816 4868 28872 4924
rect 28872 4868 28876 4924
rect 28812 4864 28876 4868
rect 33572 4924 33636 4928
rect 33572 4868 33576 4924
rect 33576 4868 33632 4924
rect 33632 4868 33636 4924
rect 33572 4864 33636 4868
rect 33652 4924 33716 4928
rect 33652 4868 33656 4924
rect 33656 4868 33712 4924
rect 33712 4868 33716 4924
rect 33652 4864 33716 4868
rect 33732 4924 33796 4928
rect 33732 4868 33736 4924
rect 33736 4868 33792 4924
rect 33792 4868 33796 4924
rect 33732 4864 33796 4868
rect 33812 4924 33876 4928
rect 33812 4868 33816 4924
rect 33816 4868 33872 4924
rect 33872 4868 33876 4924
rect 33812 4864 33876 4868
rect 38572 4924 38636 4928
rect 38572 4868 38576 4924
rect 38576 4868 38632 4924
rect 38632 4868 38636 4924
rect 38572 4864 38636 4868
rect 38652 4924 38716 4928
rect 38652 4868 38656 4924
rect 38656 4868 38712 4924
rect 38712 4868 38716 4924
rect 38652 4864 38716 4868
rect 38732 4924 38796 4928
rect 38732 4868 38736 4924
rect 38736 4868 38792 4924
rect 38792 4868 38796 4924
rect 38732 4864 38796 4868
rect 38812 4924 38876 4928
rect 38812 4868 38816 4924
rect 38816 4868 38872 4924
rect 38872 4868 38876 4924
rect 38812 4864 38876 4868
rect 43572 4924 43636 4928
rect 43572 4868 43576 4924
rect 43576 4868 43632 4924
rect 43632 4868 43636 4924
rect 43572 4864 43636 4868
rect 43652 4924 43716 4928
rect 43652 4868 43656 4924
rect 43656 4868 43712 4924
rect 43712 4868 43716 4924
rect 43652 4864 43716 4868
rect 43732 4924 43796 4928
rect 43732 4868 43736 4924
rect 43736 4868 43792 4924
rect 43792 4868 43796 4924
rect 43732 4864 43796 4868
rect 43812 4924 43876 4928
rect 43812 4868 43816 4924
rect 43816 4868 43872 4924
rect 43872 4868 43876 4924
rect 43812 4864 43876 4868
rect 22692 4660 22756 4724
rect 27660 4660 27724 4724
rect 6072 4380 6136 4384
rect 6072 4324 6076 4380
rect 6076 4324 6132 4380
rect 6132 4324 6136 4380
rect 6072 4320 6136 4324
rect 6152 4380 6216 4384
rect 6152 4324 6156 4380
rect 6156 4324 6212 4380
rect 6212 4324 6216 4380
rect 6152 4320 6216 4324
rect 6232 4380 6296 4384
rect 6232 4324 6236 4380
rect 6236 4324 6292 4380
rect 6292 4324 6296 4380
rect 6232 4320 6296 4324
rect 6312 4380 6376 4384
rect 6312 4324 6316 4380
rect 6316 4324 6372 4380
rect 6372 4324 6376 4380
rect 6312 4320 6376 4324
rect 11072 4380 11136 4384
rect 11072 4324 11076 4380
rect 11076 4324 11132 4380
rect 11132 4324 11136 4380
rect 11072 4320 11136 4324
rect 11152 4380 11216 4384
rect 11152 4324 11156 4380
rect 11156 4324 11212 4380
rect 11212 4324 11216 4380
rect 11152 4320 11216 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 16072 4380 16136 4384
rect 16072 4324 16076 4380
rect 16076 4324 16132 4380
rect 16132 4324 16136 4380
rect 16072 4320 16136 4324
rect 16152 4380 16216 4384
rect 16152 4324 16156 4380
rect 16156 4324 16212 4380
rect 16212 4324 16216 4380
rect 16152 4320 16216 4324
rect 16232 4380 16296 4384
rect 16232 4324 16236 4380
rect 16236 4324 16292 4380
rect 16292 4324 16296 4380
rect 16232 4320 16296 4324
rect 16312 4380 16376 4384
rect 16312 4324 16316 4380
rect 16316 4324 16372 4380
rect 16372 4324 16376 4380
rect 16312 4320 16376 4324
rect 21072 4380 21136 4384
rect 21072 4324 21076 4380
rect 21076 4324 21132 4380
rect 21132 4324 21136 4380
rect 21072 4320 21136 4324
rect 21152 4380 21216 4384
rect 21152 4324 21156 4380
rect 21156 4324 21212 4380
rect 21212 4324 21216 4380
rect 21152 4320 21216 4324
rect 21232 4380 21296 4384
rect 21232 4324 21236 4380
rect 21236 4324 21292 4380
rect 21292 4324 21296 4380
rect 21232 4320 21296 4324
rect 21312 4380 21376 4384
rect 21312 4324 21316 4380
rect 21316 4324 21372 4380
rect 21372 4324 21376 4380
rect 21312 4320 21376 4324
rect 26072 4380 26136 4384
rect 26072 4324 26076 4380
rect 26076 4324 26132 4380
rect 26132 4324 26136 4380
rect 26072 4320 26136 4324
rect 26152 4380 26216 4384
rect 26152 4324 26156 4380
rect 26156 4324 26212 4380
rect 26212 4324 26216 4380
rect 26152 4320 26216 4324
rect 26232 4380 26296 4384
rect 26232 4324 26236 4380
rect 26236 4324 26292 4380
rect 26292 4324 26296 4380
rect 26232 4320 26296 4324
rect 26312 4380 26376 4384
rect 26312 4324 26316 4380
rect 26316 4324 26372 4380
rect 26372 4324 26376 4380
rect 26312 4320 26376 4324
rect 31072 4380 31136 4384
rect 31072 4324 31076 4380
rect 31076 4324 31132 4380
rect 31132 4324 31136 4380
rect 31072 4320 31136 4324
rect 31152 4380 31216 4384
rect 31152 4324 31156 4380
rect 31156 4324 31212 4380
rect 31212 4324 31216 4380
rect 31152 4320 31216 4324
rect 31232 4380 31296 4384
rect 31232 4324 31236 4380
rect 31236 4324 31292 4380
rect 31292 4324 31296 4380
rect 31232 4320 31296 4324
rect 31312 4380 31376 4384
rect 31312 4324 31316 4380
rect 31316 4324 31372 4380
rect 31372 4324 31376 4380
rect 31312 4320 31376 4324
rect 36072 4380 36136 4384
rect 36072 4324 36076 4380
rect 36076 4324 36132 4380
rect 36132 4324 36136 4380
rect 36072 4320 36136 4324
rect 36152 4380 36216 4384
rect 36152 4324 36156 4380
rect 36156 4324 36212 4380
rect 36212 4324 36216 4380
rect 36152 4320 36216 4324
rect 36232 4380 36296 4384
rect 36232 4324 36236 4380
rect 36236 4324 36292 4380
rect 36292 4324 36296 4380
rect 36232 4320 36296 4324
rect 36312 4380 36376 4384
rect 36312 4324 36316 4380
rect 36316 4324 36372 4380
rect 36372 4324 36376 4380
rect 36312 4320 36376 4324
rect 41072 4380 41136 4384
rect 41072 4324 41076 4380
rect 41076 4324 41132 4380
rect 41132 4324 41136 4380
rect 41072 4320 41136 4324
rect 41152 4380 41216 4384
rect 41152 4324 41156 4380
rect 41156 4324 41212 4380
rect 41212 4324 41216 4380
rect 41152 4320 41216 4324
rect 41232 4380 41296 4384
rect 41232 4324 41236 4380
rect 41236 4324 41292 4380
rect 41292 4324 41296 4380
rect 41232 4320 41296 4324
rect 41312 4380 41376 4384
rect 41312 4324 41316 4380
rect 41316 4324 41372 4380
rect 41372 4324 41376 4380
rect 41312 4320 41376 4324
rect 19196 4040 19260 4044
rect 19196 3984 19210 4040
rect 19210 3984 19260 4040
rect 19196 3980 19260 3984
rect 25820 3980 25884 4044
rect 3572 3836 3636 3840
rect 3572 3780 3576 3836
rect 3576 3780 3632 3836
rect 3632 3780 3636 3836
rect 3572 3776 3636 3780
rect 3652 3836 3716 3840
rect 3652 3780 3656 3836
rect 3656 3780 3712 3836
rect 3712 3780 3716 3836
rect 3652 3776 3716 3780
rect 3732 3836 3796 3840
rect 3732 3780 3736 3836
rect 3736 3780 3792 3836
rect 3792 3780 3796 3836
rect 3732 3776 3796 3780
rect 3812 3836 3876 3840
rect 3812 3780 3816 3836
rect 3816 3780 3872 3836
rect 3872 3780 3876 3836
rect 3812 3776 3876 3780
rect 8572 3836 8636 3840
rect 8572 3780 8576 3836
rect 8576 3780 8632 3836
rect 8632 3780 8636 3836
rect 8572 3776 8636 3780
rect 8652 3836 8716 3840
rect 8652 3780 8656 3836
rect 8656 3780 8712 3836
rect 8712 3780 8716 3836
rect 8652 3776 8716 3780
rect 8732 3836 8796 3840
rect 8732 3780 8736 3836
rect 8736 3780 8792 3836
rect 8792 3780 8796 3836
rect 8732 3776 8796 3780
rect 8812 3836 8876 3840
rect 8812 3780 8816 3836
rect 8816 3780 8872 3836
rect 8872 3780 8876 3836
rect 8812 3776 8876 3780
rect 13572 3836 13636 3840
rect 13572 3780 13576 3836
rect 13576 3780 13632 3836
rect 13632 3780 13636 3836
rect 13572 3776 13636 3780
rect 13652 3836 13716 3840
rect 13652 3780 13656 3836
rect 13656 3780 13712 3836
rect 13712 3780 13716 3836
rect 13652 3776 13716 3780
rect 13732 3836 13796 3840
rect 13732 3780 13736 3836
rect 13736 3780 13792 3836
rect 13792 3780 13796 3836
rect 13732 3776 13796 3780
rect 13812 3836 13876 3840
rect 13812 3780 13816 3836
rect 13816 3780 13872 3836
rect 13872 3780 13876 3836
rect 13812 3776 13876 3780
rect 18572 3836 18636 3840
rect 18572 3780 18576 3836
rect 18576 3780 18632 3836
rect 18632 3780 18636 3836
rect 18572 3776 18636 3780
rect 18652 3836 18716 3840
rect 18652 3780 18656 3836
rect 18656 3780 18712 3836
rect 18712 3780 18716 3836
rect 18652 3776 18716 3780
rect 18732 3836 18796 3840
rect 18732 3780 18736 3836
rect 18736 3780 18792 3836
rect 18792 3780 18796 3836
rect 18732 3776 18796 3780
rect 18812 3836 18876 3840
rect 18812 3780 18816 3836
rect 18816 3780 18872 3836
rect 18872 3780 18876 3836
rect 18812 3776 18876 3780
rect 23572 3836 23636 3840
rect 23572 3780 23576 3836
rect 23576 3780 23632 3836
rect 23632 3780 23636 3836
rect 23572 3776 23636 3780
rect 23652 3836 23716 3840
rect 23652 3780 23656 3836
rect 23656 3780 23712 3836
rect 23712 3780 23716 3836
rect 23652 3776 23716 3780
rect 23732 3836 23796 3840
rect 23732 3780 23736 3836
rect 23736 3780 23792 3836
rect 23792 3780 23796 3836
rect 23732 3776 23796 3780
rect 23812 3836 23876 3840
rect 23812 3780 23816 3836
rect 23816 3780 23872 3836
rect 23872 3780 23876 3836
rect 23812 3776 23876 3780
rect 28572 3836 28636 3840
rect 28572 3780 28576 3836
rect 28576 3780 28632 3836
rect 28632 3780 28636 3836
rect 28572 3776 28636 3780
rect 28652 3836 28716 3840
rect 28652 3780 28656 3836
rect 28656 3780 28712 3836
rect 28712 3780 28716 3836
rect 28652 3776 28716 3780
rect 28732 3836 28796 3840
rect 28732 3780 28736 3836
rect 28736 3780 28792 3836
rect 28792 3780 28796 3836
rect 28732 3776 28796 3780
rect 28812 3836 28876 3840
rect 28812 3780 28816 3836
rect 28816 3780 28872 3836
rect 28872 3780 28876 3836
rect 28812 3776 28876 3780
rect 33572 3836 33636 3840
rect 33572 3780 33576 3836
rect 33576 3780 33632 3836
rect 33632 3780 33636 3836
rect 33572 3776 33636 3780
rect 33652 3836 33716 3840
rect 33652 3780 33656 3836
rect 33656 3780 33712 3836
rect 33712 3780 33716 3836
rect 33652 3776 33716 3780
rect 33732 3836 33796 3840
rect 33732 3780 33736 3836
rect 33736 3780 33792 3836
rect 33792 3780 33796 3836
rect 33732 3776 33796 3780
rect 33812 3836 33876 3840
rect 33812 3780 33816 3836
rect 33816 3780 33872 3836
rect 33872 3780 33876 3836
rect 33812 3776 33876 3780
rect 38572 3836 38636 3840
rect 38572 3780 38576 3836
rect 38576 3780 38632 3836
rect 38632 3780 38636 3836
rect 38572 3776 38636 3780
rect 38652 3836 38716 3840
rect 38652 3780 38656 3836
rect 38656 3780 38712 3836
rect 38712 3780 38716 3836
rect 38652 3776 38716 3780
rect 38732 3836 38796 3840
rect 38732 3780 38736 3836
rect 38736 3780 38792 3836
rect 38792 3780 38796 3836
rect 38732 3776 38796 3780
rect 38812 3836 38876 3840
rect 38812 3780 38816 3836
rect 38816 3780 38872 3836
rect 38872 3780 38876 3836
rect 38812 3776 38876 3780
rect 43572 3836 43636 3840
rect 43572 3780 43576 3836
rect 43576 3780 43632 3836
rect 43632 3780 43636 3836
rect 43572 3776 43636 3780
rect 43652 3836 43716 3840
rect 43652 3780 43656 3836
rect 43656 3780 43712 3836
rect 43712 3780 43716 3836
rect 43652 3776 43716 3780
rect 43732 3836 43796 3840
rect 43732 3780 43736 3836
rect 43736 3780 43792 3836
rect 43792 3780 43796 3836
rect 43732 3776 43796 3780
rect 43812 3836 43876 3840
rect 43812 3780 43816 3836
rect 43816 3780 43872 3836
rect 43872 3780 43876 3836
rect 43812 3776 43876 3780
rect 6072 3292 6136 3296
rect 6072 3236 6076 3292
rect 6076 3236 6132 3292
rect 6132 3236 6136 3292
rect 6072 3232 6136 3236
rect 6152 3292 6216 3296
rect 6152 3236 6156 3292
rect 6156 3236 6212 3292
rect 6212 3236 6216 3292
rect 6152 3232 6216 3236
rect 6232 3292 6296 3296
rect 6232 3236 6236 3292
rect 6236 3236 6292 3292
rect 6292 3236 6296 3292
rect 6232 3232 6296 3236
rect 6312 3292 6376 3296
rect 6312 3236 6316 3292
rect 6316 3236 6372 3292
rect 6372 3236 6376 3292
rect 6312 3232 6376 3236
rect 11072 3292 11136 3296
rect 11072 3236 11076 3292
rect 11076 3236 11132 3292
rect 11132 3236 11136 3292
rect 11072 3232 11136 3236
rect 11152 3292 11216 3296
rect 11152 3236 11156 3292
rect 11156 3236 11212 3292
rect 11212 3236 11216 3292
rect 11152 3232 11216 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 16072 3292 16136 3296
rect 16072 3236 16076 3292
rect 16076 3236 16132 3292
rect 16132 3236 16136 3292
rect 16072 3232 16136 3236
rect 16152 3292 16216 3296
rect 16152 3236 16156 3292
rect 16156 3236 16212 3292
rect 16212 3236 16216 3292
rect 16152 3232 16216 3236
rect 16232 3292 16296 3296
rect 16232 3236 16236 3292
rect 16236 3236 16292 3292
rect 16292 3236 16296 3292
rect 16232 3232 16296 3236
rect 16312 3292 16376 3296
rect 16312 3236 16316 3292
rect 16316 3236 16372 3292
rect 16372 3236 16376 3292
rect 16312 3232 16376 3236
rect 21072 3292 21136 3296
rect 21072 3236 21076 3292
rect 21076 3236 21132 3292
rect 21132 3236 21136 3292
rect 21072 3232 21136 3236
rect 21152 3292 21216 3296
rect 21152 3236 21156 3292
rect 21156 3236 21212 3292
rect 21212 3236 21216 3292
rect 21152 3232 21216 3236
rect 21232 3292 21296 3296
rect 21232 3236 21236 3292
rect 21236 3236 21292 3292
rect 21292 3236 21296 3292
rect 21232 3232 21296 3236
rect 21312 3292 21376 3296
rect 21312 3236 21316 3292
rect 21316 3236 21372 3292
rect 21372 3236 21376 3292
rect 21312 3232 21376 3236
rect 26072 3292 26136 3296
rect 26072 3236 26076 3292
rect 26076 3236 26132 3292
rect 26132 3236 26136 3292
rect 26072 3232 26136 3236
rect 26152 3292 26216 3296
rect 26152 3236 26156 3292
rect 26156 3236 26212 3292
rect 26212 3236 26216 3292
rect 26152 3232 26216 3236
rect 26232 3292 26296 3296
rect 26232 3236 26236 3292
rect 26236 3236 26292 3292
rect 26292 3236 26296 3292
rect 26232 3232 26296 3236
rect 26312 3292 26376 3296
rect 26312 3236 26316 3292
rect 26316 3236 26372 3292
rect 26372 3236 26376 3292
rect 26312 3232 26376 3236
rect 31072 3292 31136 3296
rect 31072 3236 31076 3292
rect 31076 3236 31132 3292
rect 31132 3236 31136 3292
rect 31072 3232 31136 3236
rect 31152 3292 31216 3296
rect 31152 3236 31156 3292
rect 31156 3236 31212 3292
rect 31212 3236 31216 3292
rect 31152 3232 31216 3236
rect 31232 3292 31296 3296
rect 31232 3236 31236 3292
rect 31236 3236 31292 3292
rect 31292 3236 31296 3292
rect 31232 3232 31296 3236
rect 31312 3292 31376 3296
rect 31312 3236 31316 3292
rect 31316 3236 31372 3292
rect 31372 3236 31376 3292
rect 31312 3232 31376 3236
rect 36072 3292 36136 3296
rect 36072 3236 36076 3292
rect 36076 3236 36132 3292
rect 36132 3236 36136 3292
rect 36072 3232 36136 3236
rect 36152 3292 36216 3296
rect 36152 3236 36156 3292
rect 36156 3236 36212 3292
rect 36212 3236 36216 3292
rect 36152 3232 36216 3236
rect 36232 3292 36296 3296
rect 36232 3236 36236 3292
rect 36236 3236 36292 3292
rect 36292 3236 36296 3292
rect 36232 3232 36296 3236
rect 36312 3292 36376 3296
rect 36312 3236 36316 3292
rect 36316 3236 36372 3292
rect 36372 3236 36376 3292
rect 36312 3232 36376 3236
rect 41072 3292 41136 3296
rect 41072 3236 41076 3292
rect 41076 3236 41132 3292
rect 41132 3236 41136 3292
rect 41072 3232 41136 3236
rect 41152 3292 41216 3296
rect 41152 3236 41156 3292
rect 41156 3236 41212 3292
rect 41212 3236 41216 3292
rect 41152 3232 41216 3236
rect 41232 3292 41296 3296
rect 41232 3236 41236 3292
rect 41236 3236 41292 3292
rect 41292 3236 41296 3292
rect 41232 3232 41296 3236
rect 41312 3292 41376 3296
rect 41312 3236 41316 3292
rect 41316 3236 41372 3292
rect 41372 3236 41376 3292
rect 41312 3232 41376 3236
rect 39988 3164 40052 3228
rect 28948 3028 29012 3092
rect 16988 2892 17052 2956
rect 3572 2748 3636 2752
rect 3572 2692 3576 2748
rect 3576 2692 3632 2748
rect 3632 2692 3636 2748
rect 3572 2688 3636 2692
rect 3652 2748 3716 2752
rect 3652 2692 3656 2748
rect 3656 2692 3712 2748
rect 3712 2692 3716 2748
rect 3652 2688 3716 2692
rect 3732 2748 3796 2752
rect 3732 2692 3736 2748
rect 3736 2692 3792 2748
rect 3792 2692 3796 2748
rect 3732 2688 3796 2692
rect 3812 2748 3876 2752
rect 3812 2692 3816 2748
rect 3816 2692 3872 2748
rect 3872 2692 3876 2748
rect 3812 2688 3876 2692
rect 8572 2748 8636 2752
rect 8572 2692 8576 2748
rect 8576 2692 8632 2748
rect 8632 2692 8636 2748
rect 8572 2688 8636 2692
rect 8652 2748 8716 2752
rect 8652 2692 8656 2748
rect 8656 2692 8712 2748
rect 8712 2692 8716 2748
rect 8652 2688 8716 2692
rect 8732 2748 8796 2752
rect 8732 2692 8736 2748
rect 8736 2692 8792 2748
rect 8792 2692 8796 2748
rect 8732 2688 8796 2692
rect 8812 2748 8876 2752
rect 8812 2692 8816 2748
rect 8816 2692 8872 2748
rect 8872 2692 8876 2748
rect 8812 2688 8876 2692
rect 13572 2748 13636 2752
rect 13572 2692 13576 2748
rect 13576 2692 13632 2748
rect 13632 2692 13636 2748
rect 13572 2688 13636 2692
rect 13652 2748 13716 2752
rect 13652 2692 13656 2748
rect 13656 2692 13712 2748
rect 13712 2692 13716 2748
rect 13652 2688 13716 2692
rect 13732 2748 13796 2752
rect 13732 2692 13736 2748
rect 13736 2692 13792 2748
rect 13792 2692 13796 2748
rect 13732 2688 13796 2692
rect 13812 2748 13876 2752
rect 13812 2692 13816 2748
rect 13816 2692 13872 2748
rect 13872 2692 13876 2748
rect 13812 2688 13876 2692
rect 18572 2748 18636 2752
rect 18572 2692 18576 2748
rect 18576 2692 18632 2748
rect 18632 2692 18636 2748
rect 18572 2688 18636 2692
rect 18652 2748 18716 2752
rect 18652 2692 18656 2748
rect 18656 2692 18712 2748
rect 18712 2692 18716 2748
rect 18652 2688 18716 2692
rect 18732 2748 18796 2752
rect 18732 2692 18736 2748
rect 18736 2692 18792 2748
rect 18792 2692 18796 2748
rect 18732 2688 18796 2692
rect 18812 2748 18876 2752
rect 18812 2692 18816 2748
rect 18816 2692 18872 2748
rect 18872 2692 18876 2748
rect 18812 2688 18876 2692
rect 23572 2748 23636 2752
rect 23572 2692 23576 2748
rect 23576 2692 23632 2748
rect 23632 2692 23636 2748
rect 23572 2688 23636 2692
rect 23652 2748 23716 2752
rect 23652 2692 23656 2748
rect 23656 2692 23712 2748
rect 23712 2692 23716 2748
rect 23652 2688 23716 2692
rect 23732 2748 23796 2752
rect 23732 2692 23736 2748
rect 23736 2692 23792 2748
rect 23792 2692 23796 2748
rect 23732 2688 23796 2692
rect 23812 2748 23876 2752
rect 23812 2692 23816 2748
rect 23816 2692 23872 2748
rect 23872 2692 23876 2748
rect 23812 2688 23876 2692
rect 28572 2748 28636 2752
rect 28572 2692 28576 2748
rect 28576 2692 28632 2748
rect 28632 2692 28636 2748
rect 28572 2688 28636 2692
rect 28652 2748 28716 2752
rect 28652 2692 28656 2748
rect 28656 2692 28712 2748
rect 28712 2692 28716 2748
rect 28652 2688 28716 2692
rect 28732 2748 28796 2752
rect 28732 2692 28736 2748
rect 28736 2692 28792 2748
rect 28792 2692 28796 2748
rect 28732 2688 28796 2692
rect 28812 2748 28876 2752
rect 28812 2692 28816 2748
rect 28816 2692 28872 2748
rect 28872 2692 28876 2748
rect 28812 2688 28876 2692
rect 33572 2748 33636 2752
rect 33572 2692 33576 2748
rect 33576 2692 33632 2748
rect 33632 2692 33636 2748
rect 33572 2688 33636 2692
rect 33652 2748 33716 2752
rect 33652 2692 33656 2748
rect 33656 2692 33712 2748
rect 33712 2692 33716 2748
rect 33652 2688 33716 2692
rect 33732 2748 33796 2752
rect 33732 2692 33736 2748
rect 33736 2692 33792 2748
rect 33792 2692 33796 2748
rect 33732 2688 33796 2692
rect 33812 2748 33876 2752
rect 33812 2692 33816 2748
rect 33816 2692 33872 2748
rect 33872 2692 33876 2748
rect 33812 2688 33876 2692
rect 38572 2748 38636 2752
rect 38572 2692 38576 2748
rect 38576 2692 38632 2748
rect 38632 2692 38636 2748
rect 38572 2688 38636 2692
rect 38652 2748 38716 2752
rect 38652 2692 38656 2748
rect 38656 2692 38712 2748
rect 38712 2692 38716 2748
rect 38652 2688 38716 2692
rect 38732 2748 38796 2752
rect 38732 2692 38736 2748
rect 38736 2692 38792 2748
rect 38792 2692 38796 2748
rect 38732 2688 38796 2692
rect 38812 2748 38876 2752
rect 38812 2692 38816 2748
rect 38816 2692 38872 2748
rect 38872 2692 38876 2748
rect 38812 2688 38876 2692
rect 43572 2748 43636 2752
rect 43572 2692 43576 2748
rect 43576 2692 43632 2748
rect 43632 2692 43636 2748
rect 43572 2688 43636 2692
rect 43652 2748 43716 2752
rect 43652 2692 43656 2748
rect 43656 2692 43712 2748
rect 43712 2692 43716 2748
rect 43652 2688 43716 2692
rect 43732 2748 43796 2752
rect 43732 2692 43736 2748
rect 43736 2692 43792 2748
rect 43792 2692 43796 2748
rect 43732 2688 43796 2692
rect 43812 2748 43876 2752
rect 43812 2692 43816 2748
rect 43816 2692 43872 2748
rect 43872 2692 43876 2748
rect 43812 2688 43876 2692
rect 22692 2348 22756 2412
rect 6072 2204 6136 2208
rect 6072 2148 6076 2204
rect 6076 2148 6132 2204
rect 6132 2148 6136 2204
rect 6072 2144 6136 2148
rect 6152 2204 6216 2208
rect 6152 2148 6156 2204
rect 6156 2148 6212 2204
rect 6212 2148 6216 2204
rect 6152 2144 6216 2148
rect 6232 2204 6296 2208
rect 6232 2148 6236 2204
rect 6236 2148 6292 2204
rect 6292 2148 6296 2204
rect 6232 2144 6296 2148
rect 6312 2204 6376 2208
rect 6312 2148 6316 2204
rect 6316 2148 6372 2204
rect 6372 2148 6376 2204
rect 6312 2144 6376 2148
rect 11072 2204 11136 2208
rect 11072 2148 11076 2204
rect 11076 2148 11132 2204
rect 11132 2148 11136 2204
rect 11072 2144 11136 2148
rect 11152 2204 11216 2208
rect 11152 2148 11156 2204
rect 11156 2148 11212 2204
rect 11212 2148 11216 2204
rect 11152 2144 11216 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 16072 2204 16136 2208
rect 16072 2148 16076 2204
rect 16076 2148 16132 2204
rect 16132 2148 16136 2204
rect 16072 2144 16136 2148
rect 16152 2204 16216 2208
rect 16152 2148 16156 2204
rect 16156 2148 16212 2204
rect 16212 2148 16216 2204
rect 16152 2144 16216 2148
rect 16232 2204 16296 2208
rect 16232 2148 16236 2204
rect 16236 2148 16292 2204
rect 16292 2148 16296 2204
rect 16232 2144 16296 2148
rect 16312 2204 16376 2208
rect 16312 2148 16316 2204
rect 16316 2148 16372 2204
rect 16372 2148 16376 2204
rect 16312 2144 16376 2148
rect 21072 2204 21136 2208
rect 21072 2148 21076 2204
rect 21076 2148 21132 2204
rect 21132 2148 21136 2204
rect 21072 2144 21136 2148
rect 21152 2204 21216 2208
rect 21152 2148 21156 2204
rect 21156 2148 21212 2204
rect 21212 2148 21216 2204
rect 21152 2144 21216 2148
rect 21232 2204 21296 2208
rect 21232 2148 21236 2204
rect 21236 2148 21292 2204
rect 21292 2148 21296 2204
rect 21232 2144 21296 2148
rect 21312 2204 21376 2208
rect 21312 2148 21316 2204
rect 21316 2148 21372 2204
rect 21372 2148 21376 2204
rect 21312 2144 21376 2148
rect 26072 2204 26136 2208
rect 26072 2148 26076 2204
rect 26076 2148 26132 2204
rect 26132 2148 26136 2204
rect 26072 2144 26136 2148
rect 26152 2204 26216 2208
rect 26152 2148 26156 2204
rect 26156 2148 26212 2204
rect 26212 2148 26216 2204
rect 26152 2144 26216 2148
rect 26232 2204 26296 2208
rect 26232 2148 26236 2204
rect 26236 2148 26292 2204
rect 26292 2148 26296 2204
rect 26232 2144 26296 2148
rect 26312 2204 26376 2208
rect 26312 2148 26316 2204
rect 26316 2148 26372 2204
rect 26372 2148 26376 2204
rect 26312 2144 26376 2148
rect 31072 2204 31136 2208
rect 31072 2148 31076 2204
rect 31076 2148 31132 2204
rect 31132 2148 31136 2204
rect 31072 2144 31136 2148
rect 31152 2204 31216 2208
rect 31152 2148 31156 2204
rect 31156 2148 31212 2204
rect 31212 2148 31216 2204
rect 31152 2144 31216 2148
rect 31232 2204 31296 2208
rect 31232 2148 31236 2204
rect 31236 2148 31292 2204
rect 31292 2148 31296 2204
rect 31232 2144 31296 2148
rect 31312 2204 31376 2208
rect 31312 2148 31316 2204
rect 31316 2148 31372 2204
rect 31372 2148 31376 2204
rect 31312 2144 31376 2148
rect 36072 2204 36136 2208
rect 36072 2148 36076 2204
rect 36076 2148 36132 2204
rect 36132 2148 36136 2204
rect 36072 2144 36136 2148
rect 36152 2204 36216 2208
rect 36152 2148 36156 2204
rect 36156 2148 36212 2204
rect 36212 2148 36216 2204
rect 36152 2144 36216 2148
rect 36232 2204 36296 2208
rect 36232 2148 36236 2204
rect 36236 2148 36292 2204
rect 36292 2148 36296 2204
rect 36232 2144 36296 2148
rect 36312 2204 36376 2208
rect 36312 2148 36316 2204
rect 36316 2148 36372 2204
rect 36372 2148 36376 2204
rect 36312 2144 36376 2148
rect 41072 2204 41136 2208
rect 41072 2148 41076 2204
rect 41076 2148 41132 2204
rect 41132 2148 41136 2204
rect 41072 2144 41136 2148
rect 41152 2204 41216 2208
rect 41152 2148 41156 2204
rect 41156 2148 41212 2204
rect 41212 2148 41216 2204
rect 41152 2144 41216 2148
rect 41232 2204 41296 2208
rect 41232 2148 41236 2204
rect 41236 2148 41292 2204
rect 41292 2148 41296 2204
rect 41232 2144 41296 2148
rect 41312 2204 41376 2208
rect 41312 2148 41316 2204
rect 41316 2148 41372 2204
rect 41372 2148 41376 2204
rect 41312 2144 41376 2148
rect 21588 2000 21652 2004
rect 21588 1944 21602 2000
rect 21602 1944 21652 2000
rect 21588 1940 21652 1944
rect 3572 1660 3636 1664
rect 3572 1604 3576 1660
rect 3576 1604 3632 1660
rect 3632 1604 3636 1660
rect 3572 1600 3636 1604
rect 3652 1660 3716 1664
rect 3652 1604 3656 1660
rect 3656 1604 3712 1660
rect 3712 1604 3716 1660
rect 3652 1600 3716 1604
rect 3732 1660 3796 1664
rect 3732 1604 3736 1660
rect 3736 1604 3792 1660
rect 3792 1604 3796 1660
rect 3732 1600 3796 1604
rect 3812 1660 3876 1664
rect 3812 1604 3816 1660
rect 3816 1604 3872 1660
rect 3872 1604 3876 1660
rect 3812 1600 3876 1604
rect 8572 1660 8636 1664
rect 8572 1604 8576 1660
rect 8576 1604 8632 1660
rect 8632 1604 8636 1660
rect 8572 1600 8636 1604
rect 8652 1660 8716 1664
rect 8652 1604 8656 1660
rect 8656 1604 8712 1660
rect 8712 1604 8716 1660
rect 8652 1600 8716 1604
rect 8732 1660 8796 1664
rect 8732 1604 8736 1660
rect 8736 1604 8792 1660
rect 8792 1604 8796 1660
rect 8732 1600 8796 1604
rect 8812 1660 8876 1664
rect 8812 1604 8816 1660
rect 8816 1604 8872 1660
rect 8872 1604 8876 1660
rect 8812 1600 8876 1604
rect 13572 1660 13636 1664
rect 13572 1604 13576 1660
rect 13576 1604 13632 1660
rect 13632 1604 13636 1660
rect 13572 1600 13636 1604
rect 13652 1660 13716 1664
rect 13652 1604 13656 1660
rect 13656 1604 13712 1660
rect 13712 1604 13716 1660
rect 13652 1600 13716 1604
rect 13732 1660 13796 1664
rect 13732 1604 13736 1660
rect 13736 1604 13792 1660
rect 13792 1604 13796 1660
rect 13732 1600 13796 1604
rect 13812 1660 13876 1664
rect 13812 1604 13816 1660
rect 13816 1604 13872 1660
rect 13872 1604 13876 1660
rect 13812 1600 13876 1604
rect 18572 1660 18636 1664
rect 18572 1604 18576 1660
rect 18576 1604 18632 1660
rect 18632 1604 18636 1660
rect 18572 1600 18636 1604
rect 18652 1660 18716 1664
rect 18652 1604 18656 1660
rect 18656 1604 18712 1660
rect 18712 1604 18716 1660
rect 18652 1600 18716 1604
rect 18732 1660 18796 1664
rect 18732 1604 18736 1660
rect 18736 1604 18792 1660
rect 18792 1604 18796 1660
rect 18732 1600 18796 1604
rect 18812 1660 18876 1664
rect 18812 1604 18816 1660
rect 18816 1604 18872 1660
rect 18872 1604 18876 1660
rect 18812 1600 18876 1604
rect 23572 1660 23636 1664
rect 23572 1604 23576 1660
rect 23576 1604 23632 1660
rect 23632 1604 23636 1660
rect 23572 1600 23636 1604
rect 23652 1660 23716 1664
rect 23652 1604 23656 1660
rect 23656 1604 23712 1660
rect 23712 1604 23716 1660
rect 23652 1600 23716 1604
rect 23732 1660 23796 1664
rect 23732 1604 23736 1660
rect 23736 1604 23792 1660
rect 23792 1604 23796 1660
rect 23732 1600 23796 1604
rect 23812 1660 23876 1664
rect 23812 1604 23816 1660
rect 23816 1604 23872 1660
rect 23872 1604 23876 1660
rect 23812 1600 23876 1604
rect 28572 1660 28636 1664
rect 28572 1604 28576 1660
rect 28576 1604 28632 1660
rect 28632 1604 28636 1660
rect 28572 1600 28636 1604
rect 28652 1660 28716 1664
rect 28652 1604 28656 1660
rect 28656 1604 28712 1660
rect 28712 1604 28716 1660
rect 28652 1600 28716 1604
rect 28732 1660 28796 1664
rect 28732 1604 28736 1660
rect 28736 1604 28792 1660
rect 28792 1604 28796 1660
rect 28732 1600 28796 1604
rect 28812 1660 28876 1664
rect 28812 1604 28816 1660
rect 28816 1604 28872 1660
rect 28872 1604 28876 1660
rect 28812 1600 28876 1604
rect 33572 1660 33636 1664
rect 33572 1604 33576 1660
rect 33576 1604 33632 1660
rect 33632 1604 33636 1660
rect 33572 1600 33636 1604
rect 33652 1660 33716 1664
rect 33652 1604 33656 1660
rect 33656 1604 33712 1660
rect 33712 1604 33716 1660
rect 33652 1600 33716 1604
rect 33732 1660 33796 1664
rect 33732 1604 33736 1660
rect 33736 1604 33792 1660
rect 33792 1604 33796 1660
rect 33732 1600 33796 1604
rect 33812 1660 33876 1664
rect 33812 1604 33816 1660
rect 33816 1604 33872 1660
rect 33872 1604 33876 1660
rect 33812 1600 33876 1604
rect 38572 1660 38636 1664
rect 38572 1604 38576 1660
rect 38576 1604 38632 1660
rect 38632 1604 38636 1660
rect 38572 1600 38636 1604
rect 38652 1660 38716 1664
rect 38652 1604 38656 1660
rect 38656 1604 38712 1660
rect 38712 1604 38716 1660
rect 38652 1600 38716 1604
rect 38732 1660 38796 1664
rect 38732 1604 38736 1660
rect 38736 1604 38792 1660
rect 38792 1604 38796 1660
rect 38732 1600 38796 1604
rect 38812 1660 38876 1664
rect 38812 1604 38816 1660
rect 38816 1604 38872 1660
rect 38872 1604 38876 1660
rect 38812 1600 38876 1604
rect 43572 1660 43636 1664
rect 43572 1604 43576 1660
rect 43576 1604 43632 1660
rect 43632 1604 43636 1660
rect 43572 1600 43636 1604
rect 43652 1660 43716 1664
rect 43652 1604 43656 1660
rect 43656 1604 43712 1660
rect 43712 1604 43716 1660
rect 43652 1600 43716 1604
rect 43732 1660 43796 1664
rect 43732 1604 43736 1660
rect 43736 1604 43792 1660
rect 43792 1604 43796 1660
rect 43732 1600 43796 1604
rect 43812 1660 43876 1664
rect 43812 1604 43816 1660
rect 43816 1604 43872 1660
rect 43872 1604 43876 1660
rect 43812 1600 43876 1604
rect 28948 1260 29012 1324
rect 34284 1260 34348 1324
rect 39988 1260 40052 1324
rect 34468 1124 34532 1188
rect 6072 1116 6136 1120
rect 6072 1060 6076 1116
rect 6076 1060 6132 1116
rect 6132 1060 6136 1116
rect 6072 1056 6136 1060
rect 6152 1116 6216 1120
rect 6152 1060 6156 1116
rect 6156 1060 6212 1116
rect 6212 1060 6216 1116
rect 6152 1056 6216 1060
rect 6232 1116 6296 1120
rect 6232 1060 6236 1116
rect 6236 1060 6292 1116
rect 6292 1060 6296 1116
rect 6232 1056 6296 1060
rect 6312 1116 6376 1120
rect 6312 1060 6316 1116
rect 6316 1060 6372 1116
rect 6372 1060 6376 1116
rect 6312 1056 6376 1060
rect 11072 1116 11136 1120
rect 11072 1060 11076 1116
rect 11076 1060 11132 1116
rect 11132 1060 11136 1116
rect 11072 1056 11136 1060
rect 11152 1116 11216 1120
rect 11152 1060 11156 1116
rect 11156 1060 11212 1116
rect 11212 1060 11216 1116
rect 11152 1056 11216 1060
rect 11232 1116 11296 1120
rect 11232 1060 11236 1116
rect 11236 1060 11292 1116
rect 11292 1060 11296 1116
rect 11232 1056 11296 1060
rect 11312 1116 11376 1120
rect 11312 1060 11316 1116
rect 11316 1060 11372 1116
rect 11372 1060 11376 1116
rect 11312 1056 11376 1060
rect 16072 1116 16136 1120
rect 16072 1060 16076 1116
rect 16076 1060 16132 1116
rect 16132 1060 16136 1116
rect 16072 1056 16136 1060
rect 16152 1116 16216 1120
rect 16152 1060 16156 1116
rect 16156 1060 16212 1116
rect 16212 1060 16216 1116
rect 16152 1056 16216 1060
rect 16232 1116 16296 1120
rect 16232 1060 16236 1116
rect 16236 1060 16292 1116
rect 16292 1060 16296 1116
rect 16232 1056 16296 1060
rect 16312 1116 16376 1120
rect 16312 1060 16316 1116
rect 16316 1060 16372 1116
rect 16372 1060 16376 1116
rect 16312 1056 16376 1060
rect 21072 1116 21136 1120
rect 21072 1060 21076 1116
rect 21076 1060 21132 1116
rect 21132 1060 21136 1116
rect 21072 1056 21136 1060
rect 21152 1116 21216 1120
rect 21152 1060 21156 1116
rect 21156 1060 21212 1116
rect 21212 1060 21216 1116
rect 21152 1056 21216 1060
rect 21232 1116 21296 1120
rect 21232 1060 21236 1116
rect 21236 1060 21292 1116
rect 21292 1060 21296 1116
rect 21232 1056 21296 1060
rect 21312 1116 21376 1120
rect 21312 1060 21316 1116
rect 21316 1060 21372 1116
rect 21372 1060 21376 1116
rect 21312 1056 21376 1060
rect 26072 1116 26136 1120
rect 26072 1060 26076 1116
rect 26076 1060 26132 1116
rect 26132 1060 26136 1116
rect 26072 1056 26136 1060
rect 26152 1116 26216 1120
rect 26152 1060 26156 1116
rect 26156 1060 26212 1116
rect 26212 1060 26216 1116
rect 26152 1056 26216 1060
rect 26232 1116 26296 1120
rect 26232 1060 26236 1116
rect 26236 1060 26292 1116
rect 26292 1060 26296 1116
rect 26232 1056 26296 1060
rect 26312 1116 26376 1120
rect 26312 1060 26316 1116
rect 26316 1060 26372 1116
rect 26372 1060 26376 1116
rect 26312 1056 26376 1060
rect 31072 1116 31136 1120
rect 31072 1060 31076 1116
rect 31076 1060 31132 1116
rect 31132 1060 31136 1116
rect 31072 1056 31136 1060
rect 31152 1116 31216 1120
rect 31152 1060 31156 1116
rect 31156 1060 31212 1116
rect 31212 1060 31216 1116
rect 31152 1056 31216 1060
rect 31232 1116 31296 1120
rect 31232 1060 31236 1116
rect 31236 1060 31292 1116
rect 31292 1060 31296 1116
rect 31232 1056 31296 1060
rect 31312 1116 31376 1120
rect 31312 1060 31316 1116
rect 31316 1060 31372 1116
rect 31372 1060 31376 1116
rect 31312 1056 31376 1060
rect 36072 1116 36136 1120
rect 36072 1060 36076 1116
rect 36076 1060 36132 1116
rect 36132 1060 36136 1116
rect 36072 1056 36136 1060
rect 36152 1116 36216 1120
rect 36152 1060 36156 1116
rect 36156 1060 36212 1116
rect 36212 1060 36216 1116
rect 36152 1056 36216 1060
rect 36232 1116 36296 1120
rect 36232 1060 36236 1116
rect 36236 1060 36292 1116
rect 36292 1060 36296 1116
rect 36232 1056 36296 1060
rect 36312 1116 36376 1120
rect 36312 1060 36316 1116
rect 36316 1060 36372 1116
rect 36372 1060 36376 1116
rect 36312 1056 36376 1060
rect 41072 1116 41136 1120
rect 41072 1060 41076 1116
rect 41076 1060 41132 1116
rect 41132 1060 41136 1116
rect 41072 1056 41136 1060
rect 41152 1116 41216 1120
rect 41152 1060 41156 1116
rect 41156 1060 41212 1116
rect 41212 1060 41216 1116
rect 41152 1056 41216 1060
rect 41232 1116 41296 1120
rect 41232 1060 41236 1116
rect 41236 1060 41292 1116
rect 41292 1060 41296 1116
rect 41232 1056 41296 1060
rect 41312 1116 41376 1120
rect 41312 1060 41316 1116
rect 41316 1060 41372 1116
rect 41372 1060 41376 1116
rect 41312 1056 41376 1060
<< metal4 >>
rect 3564 22336 3884 22896
rect 3564 22272 3572 22336
rect 3636 22272 3652 22336
rect 3716 22272 3732 22336
rect 3796 22272 3812 22336
rect 3876 22272 3884 22336
rect 3564 21248 3884 22272
rect 3564 21184 3572 21248
rect 3636 21184 3652 21248
rect 3716 21184 3732 21248
rect 3796 21184 3812 21248
rect 3876 21184 3884 21248
rect 3564 20160 3884 21184
rect 3564 20096 3572 20160
rect 3636 20096 3652 20160
rect 3716 20096 3732 20160
rect 3796 20096 3812 20160
rect 3876 20096 3884 20160
rect 3564 19072 3884 20096
rect 3564 19008 3572 19072
rect 3636 19008 3652 19072
rect 3716 19008 3732 19072
rect 3796 19008 3812 19072
rect 3876 19008 3884 19072
rect 3564 17984 3884 19008
rect 3564 17920 3572 17984
rect 3636 17920 3652 17984
rect 3716 17920 3732 17984
rect 3796 17920 3812 17984
rect 3876 17920 3884 17984
rect 3564 16896 3884 17920
rect 3564 16832 3572 16896
rect 3636 16832 3652 16896
rect 3716 16832 3732 16896
rect 3796 16832 3812 16896
rect 3876 16832 3884 16896
rect 3564 15808 3884 16832
rect 3564 15744 3572 15808
rect 3636 15744 3652 15808
rect 3716 15744 3732 15808
rect 3796 15744 3812 15808
rect 3876 15744 3884 15808
rect 3564 14720 3884 15744
rect 3564 14656 3572 14720
rect 3636 14656 3652 14720
rect 3716 14656 3732 14720
rect 3796 14656 3812 14720
rect 3876 14656 3884 14720
rect 3564 13632 3884 14656
rect 3564 13568 3572 13632
rect 3636 13568 3652 13632
rect 3716 13568 3732 13632
rect 3796 13568 3812 13632
rect 3876 13568 3884 13632
rect 3564 12544 3884 13568
rect 3564 12480 3572 12544
rect 3636 12480 3652 12544
rect 3716 12480 3732 12544
rect 3796 12480 3812 12544
rect 3876 12480 3884 12544
rect 3564 11456 3884 12480
rect 3564 11392 3572 11456
rect 3636 11392 3652 11456
rect 3716 11392 3732 11456
rect 3796 11392 3812 11456
rect 3876 11392 3884 11456
rect 3564 10368 3884 11392
rect 3564 10304 3572 10368
rect 3636 10304 3652 10368
rect 3716 10304 3732 10368
rect 3796 10304 3812 10368
rect 3876 10304 3884 10368
rect 3564 9280 3884 10304
rect 3564 9216 3572 9280
rect 3636 9216 3652 9280
rect 3716 9216 3732 9280
rect 3796 9216 3812 9280
rect 3876 9216 3884 9280
rect 3564 8192 3884 9216
rect 3564 8128 3572 8192
rect 3636 8128 3652 8192
rect 3716 8128 3732 8192
rect 3796 8128 3812 8192
rect 3876 8128 3884 8192
rect 3564 7104 3884 8128
rect 3564 7040 3572 7104
rect 3636 7040 3652 7104
rect 3716 7040 3732 7104
rect 3796 7040 3812 7104
rect 3876 7040 3884 7104
rect 3564 6016 3884 7040
rect 3564 5952 3572 6016
rect 3636 5952 3652 6016
rect 3716 5952 3732 6016
rect 3796 5952 3812 6016
rect 3876 5952 3884 6016
rect 3564 4928 3884 5952
rect 3564 4864 3572 4928
rect 3636 4864 3652 4928
rect 3716 4864 3732 4928
rect 3796 4864 3812 4928
rect 3876 4864 3884 4928
rect 3564 3840 3884 4864
rect 3564 3776 3572 3840
rect 3636 3776 3652 3840
rect 3716 3776 3732 3840
rect 3796 3776 3812 3840
rect 3876 3776 3884 3840
rect 3564 2752 3884 3776
rect 3564 2688 3572 2752
rect 3636 2688 3652 2752
rect 3716 2688 3732 2752
rect 3796 2688 3812 2752
rect 3876 2688 3884 2752
rect 3564 1664 3884 2688
rect 3564 1600 3572 1664
rect 3636 1600 3652 1664
rect 3716 1600 3732 1664
rect 3796 1600 3812 1664
rect 3876 1600 3884 1664
rect 3564 1040 3884 1600
rect 6064 22880 6384 22896
rect 6064 22816 6072 22880
rect 6136 22816 6152 22880
rect 6216 22816 6232 22880
rect 6296 22816 6312 22880
rect 6376 22816 6384 22880
rect 6064 21792 6384 22816
rect 6064 21728 6072 21792
rect 6136 21728 6152 21792
rect 6216 21728 6232 21792
rect 6296 21728 6312 21792
rect 6376 21728 6384 21792
rect 6064 20704 6384 21728
rect 6064 20640 6072 20704
rect 6136 20640 6152 20704
rect 6216 20640 6232 20704
rect 6296 20640 6312 20704
rect 6376 20640 6384 20704
rect 6064 19616 6384 20640
rect 6064 19552 6072 19616
rect 6136 19552 6152 19616
rect 6216 19552 6232 19616
rect 6296 19552 6312 19616
rect 6376 19552 6384 19616
rect 6064 18528 6384 19552
rect 6064 18464 6072 18528
rect 6136 18464 6152 18528
rect 6216 18464 6232 18528
rect 6296 18464 6312 18528
rect 6376 18464 6384 18528
rect 6064 17440 6384 18464
rect 6064 17376 6072 17440
rect 6136 17376 6152 17440
rect 6216 17376 6232 17440
rect 6296 17376 6312 17440
rect 6376 17376 6384 17440
rect 6064 16352 6384 17376
rect 6064 16288 6072 16352
rect 6136 16288 6152 16352
rect 6216 16288 6232 16352
rect 6296 16288 6312 16352
rect 6376 16288 6384 16352
rect 6064 15264 6384 16288
rect 6064 15200 6072 15264
rect 6136 15200 6152 15264
rect 6216 15200 6232 15264
rect 6296 15200 6312 15264
rect 6376 15200 6384 15264
rect 6064 14176 6384 15200
rect 6064 14112 6072 14176
rect 6136 14112 6152 14176
rect 6216 14112 6232 14176
rect 6296 14112 6312 14176
rect 6376 14112 6384 14176
rect 6064 13088 6384 14112
rect 6064 13024 6072 13088
rect 6136 13024 6152 13088
rect 6216 13024 6232 13088
rect 6296 13024 6312 13088
rect 6376 13024 6384 13088
rect 6064 12000 6384 13024
rect 6064 11936 6072 12000
rect 6136 11936 6152 12000
rect 6216 11936 6232 12000
rect 6296 11936 6312 12000
rect 6376 11936 6384 12000
rect 6064 10912 6384 11936
rect 6064 10848 6072 10912
rect 6136 10848 6152 10912
rect 6216 10848 6232 10912
rect 6296 10848 6312 10912
rect 6376 10848 6384 10912
rect 6064 9824 6384 10848
rect 6064 9760 6072 9824
rect 6136 9760 6152 9824
rect 6216 9760 6232 9824
rect 6296 9760 6312 9824
rect 6376 9760 6384 9824
rect 6064 8736 6384 9760
rect 6064 8672 6072 8736
rect 6136 8672 6152 8736
rect 6216 8672 6232 8736
rect 6296 8672 6312 8736
rect 6376 8672 6384 8736
rect 6064 7648 6384 8672
rect 6064 7584 6072 7648
rect 6136 7584 6152 7648
rect 6216 7584 6232 7648
rect 6296 7584 6312 7648
rect 6376 7584 6384 7648
rect 6064 6560 6384 7584
rect 6064 6496 6072 6560
rect 6136 6496 6152 6560
rect 6216 6496 6232 6560
rect 6296 6496 6312 6560
rect 6376 6496 6384 6560
rect 6064 5472 6384 6496
rect 6064 5408 6072 5472
rect 6136 5408 6152 5472
rect 6216 5408 6232 5472
rect 6296 5408 6312 5472
rect 6376 5408 6384 5472
rect 6064 4384 6384 5408
rect 6064 4320 6072 4384
rect 6136 4320 6152 4384
rect 6216 4320 6232 4384
rect 6296 4320 6312 4384
rect 6376 4320 6384 4384
rect 6064 3296 6384 4320
rect 6064 3232 6072 3296
rect 6136 3232 6152 3296
rect 6216 3232 6232 3296
rect 6296 3232 6312 3296
rect 6376 3232 6384 3296
rect 6064 2208 6384 3232
rect 6064 2144 6072 2208
rect 6136 2144 6152 2208
rect 6216 2144 6232 2208
rect 6296 2144 6312 2208
rect 6376 2144 6384 2208
rect 6064 1120 6384 2144
rect 6064 1056 6072 1120
rect 6136 1056 6152 1120
rect 6216 1056 6232 1120
rect 6296 1056 6312 1120
rect 6376 1056 6384 1120
rect 6064 1040 6384 1056
rect 8564 22336 8884 22896
rect 8564 22272 8572 22336
rect 8636 22272 8652 22336
rect 8716 22272 8732 22336
rect 8796 22272 8812 22336
rect 8876 22272 8884 22336
rect 8564 21248 8884 22272
rect 8564 21184 8572 21248
rect 8636 21184 8652 21248
rect 8716 21184 8732 21248
rect 8796 21184 8812 21248
rect 8876 21184 8884 21248
rect 8564 20160 8884 21184
rect 11064 22880 11384 22896
rect 11064 22816 11072 22880
rect 11136 22816 11152 22880
rect 11216 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11384 22880
rect 11064 21792 11384 22816
rect 11064 21728 11072 21792
rect 11136 21728 11152 21792
rect 11216 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11384 21792
rect 9259 20772 9325 20773
rect 9259 20708 9260 20772
rect 9324 20708 9325 20772
rect 9259 20707 9325 20708
rect 8564 20096 8572 20160
rect 8636 20096 8652 20160
rect 8716 20096 8732 20160
rect 8796 20096 8812 20160
rect 8876 20096 8884 20160
rect 8564 19072 8884 20096
rect 8564 19008 8572 19072
rect 8636 19008 8652 19072
rect 8716 19008 8732 19072
rect 8796 19008 8812 19072
rect 8876 19008 8884 19072
rect 8564 17984 8884 19008
rect 8564 17920 8572 17984
rect 8636 17920 8652 17984
rect 8716 17920 8732 17984
rect 8796 17920 8812 17984
rect 8876 17920 8884 17984
rect 8564 16896 8884 17920
rect 8564 16832 8572 16896
rect 8636 16832 8652 16896
rect 8716 16832 8732 16896
rect 8796 16832 8812 16896
rect 8876 16832 8884 16896
rect 8564 15808 8884 16832
rect 8564 15744 8572 15808
rect 8636 15744 8652 15808
rect 8716 15744 8732 15808
rect 8796 15744 8812 15808
rect 8876 15744 8884 15808
rect 8564 14720 8884 15744
rect 8564 14656 8572 14720
rect 8636 14656 8652 14720
rect 8716 14656 8732 14720
rect 8796 14656 8812 14720
rect 8876 14656 8884 14720
rect 8564 13632 8884 14656
rect 8564 13568 8572 13632
rect 8636 13568 8652 13632
rect 8716 13568 8732 13632
rect 8796 13568 8812 13632
rect 8876 13568 8884 13632
rect 8564 12544 8884 13568
rect 8564 12480 8572 12544
rect 8636 12480 8652 12544
rect 8716 12480 8732 12544
rect 8796 12480 8812 12544
rect 8876 12480 8884 12544
rect 8564 11456 8884 12480
rect 8564 11392 8572 11456
rect 8636 11392 8652 11456
rect 8716 11392 8732 11456
rect 8796 11392 8812 11456
rect 8876 11392 8884 11456
rect 8564 10368 8884 11392
rect 8564 10304 8572 10368
rect 8636 10304 8652 10368
rect 8716 10304 8732 10368
rect 8796 10304 8812 10368
rect 8876 10304 8884 10368
rect 8564 9280 8884 10304
rect 8564 9216 8572 9280
rect 8636 9216 8652 9280
rect 8716 9216 8732 9280
rect 8796 9216 8812 9280
rect 8876 9216 8884 9280
rect 8564 8192 8884 9216
rect 8564 8128 8572 8192
rect 8636 8128 8652 8192
rect 8716 8128 8732 8192
rect 8796 8128 8812 8192
rect 8876 8128 8884 8192
rect 8564 7104 8884 8128
rect 8564 7040 8572 7104
rect 8636 7040 8652 7104
rect 8716 7040 8732 7104
rect 8796 7040 8812 7104
rect 8876 7040 8884 7104
rect 8564 6016 8884 7040
rect 9262 6901 9322 20707
rect 11064 20704 11384 21728
rect 11064 20640 11072 20704
rect 11136 20640 11152 20704
rect 11216 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11384 20704
rect 11064 19616 11384 20640
rect 11064 19552 11072 19616
rect 11136 19552 11152 19616
rect 11216 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11384 19616
rect 11064 18528 11384 19552
rect 11064 18464 11072 18528
rect 11136 18464 11152 18528
rect 11216 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11384 18528
rect 11064 17440 11384 18464
rect 11064 17376 11072 17440
rect 11136 17376 11152 17440
rect 11216 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11384 17440
rect 11064 16352 11384 17376
rect 11064 16288 11072 16352
rect 11136 16288 11152 16352
rect 11216 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11384 16352
rect 11064 15264 11384 16288
rect 11064 15200 11072 15264
rect 11136 15200 11152 15264
rect 11216 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11384 15264
rect 11064 14176 11384 15200
rect 11064 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11384 14176
rect 11064 13088 11384 14112
rect 11064 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11384 13088
rect 11064 12000 11384 13024
rect 11064 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11384 12000
rect 11064 10912 11384 11936
rect 11064 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11384 10912
rect 11064 9824 11384 10848
rect 11064 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11384 9824
rect 11064 8736 11384 9760
rect 11064 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11384 8736
rect 11064 7648 11384 8672
rect 11064 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11384 7648
rect 9259 6900 9325 6901
rect 9259 6836 9260 6900
rect 9324 6836 9325 6900
rect 9259 6835 9325 6836
rect 8564 5952 8572 6016
rect 8636 5952 8652 6016
rect 8716 5952 8732 6016
rect 8796 5952 8812 6016
rect 8876 5952 8884 6016
rect 8564 4928 8884 5952
rect 8564 4864 8572 4928
rect 8636 4864 8652 4928
rect 8716 4864 8732 4928
rect 8796 4864 8812 4928
rect 8876 4864 8884 4928
rect 8564 3840 8884 4864
rect 8564 3776 8572 3840
rect 8636 3776 8652 3840
rect 8716 3776 8732 3840
rect 8796 3776 8812 3840
rect 8876 3776 8884 3840
rect 8564 2752 8884 3776
rect 8564 2688 8572 2752
rect 8636 2688 8652 2752
rect 8716 2688 8732 2752
rect 8796 2688 8812 2752
rect 8876 2688 8884 2752
rect 8564 1664 8884 2688
rect 8564 1600 8572 1664
rect 8636 1600 8652 1664
rect 8716 1600 8732 1664
rect 8796 1600 8812 1664
rect 8876 1600 8884 1664
rect 8564 1040 8884 1600
rect 11064 6560 11384 7584
rect 11064 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11384 6560
rect 11064 5472 11384 6496
rect 11064 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11384 5472
rect 11064 4384 11384 5408
rect 11064 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11384 4384
rect 11064 3296 11384 4320
rect 11064 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11384 3296
rect 11064 2208 11384 3232
rect 11064 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11384 2208
rect 11064 1120 11384 2144
rect 11064 1056 11072 1120
rect 11136 1056 11152 1120
rect 11216 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11384 1120
rect 11064 1040 11384 1056
rect 13564 22336 13884 22896
rect 13564 22272 13572 22336
rect 13636 22272 13652 22336
rect 13716 22272 13732 22336
rect 13796 22272 13812 22336
rect 13876 22272 13884 22336
rect 13564 21248 13884 22272
rect 13564 21184 13572 21248
rect 13636 21184 13652 21248
rect 13716 21184 13732 21248
rect 13796 21184 13812 21248
rect 13876 21184 13884 21248
rect 13564 20160 13884 21184
rect 13564 20096 13572 20160
rect 13636 20096 13652 20160
rect 13716 20096 13732 20160
rect 13796 20096 13812 20160
rect 13876 20096 13884 20160
rect 13564 19072 13884 20096
rect 13564 19008 13572 19072
rect 13636 19008 13652 19072
rect 13716 19008 13732 19072
rect 13796 19008 13812 19072
rect 13876 19008 13884 19072
rect 13564 17984 13884 19008
rect 13564 17920 13572 17984
rect 13636 17920 13652 17984
rect 13716 17920 13732 17984
rect 13796 17920 13812 17984
rect 13876 17920 13884 17984
rect 13564 16896 13884 17920
rect 13564 16832 13572 16896
rect 13636 16832 13652 16896
rect 13716 16832 13732 16896
rect 13796 16832 13812 16896
rect 13876 16832 13884 16896
rect 13564 15808 13884 16832
rect 13564 15744 13572 15808
rect 13636 15744 13652 15808
rect 13716 15744 13732 15808
rect 13796 15744 13812 15808
rect 13876 15744 13884 15808
rect 13564 14720 13884 15744
rect 13564 14656 13572 14720
rect 13636 14656 13652 14720
rect 13716 14656 13732 14720
rect 13796 14656 13812 14720
rect 13876 14656 13884 14720
rect 13564 13632 13884 14656
rect 13564 13568 13572 13632
rect 13636 13568 13652 13632
rect 13716 13568 13732 13632
rect 13796 13568 13812 13632
rect 13876 13568 13884 13632
rect 13564 12544 13884 13568
rect 13564 12480 13572 12544
rect 13636 12480 13652 12544
rect 13716 12480 13732 12544
rect 13796 12480 13812 12544
rect 13876 12480 13884 12544
rect 13564 11456 13884 12480
rect 13564 11392 13572 11456
rect 13636 11392 13652 11456
rect 13716 11392 13732 11456
rect 13796 11392 13812 11456
rect 13876 11392 13884 11456
rect 13564 10368 13884 11392
rect 13564 10304 13572 10368
rect 13636 10304 13652 10368
rect 13716 10304 13732 10368
rect 13796 10304 13812 10368
rect 13876 10304 13884 10368
rect 13564 9280 13884 10304
rect 13564 9216 13572 9280
rect 13636 9216 13652 9280
rect 13716 9216 13732 9280
rect 13796 9216 13812 9280
rect 13876 9216 13884 9280
rect 13564 8192 13884 9216
rect 13564 8128 13572 8192
rect 13636 8128 13652 8192
rect 13716 8128 13732 8192
rect 13796 8128 13812 8192
rect 13876 8128 13884 8192
rect 13564 7104 13884 8128
rect 13564 7040 13572 7104
rect 13636 7040 13652 7104
rect 13716 7040 13732 7104
rect 13796 7040 13812 7104
rect 13876 7040 13884 7104
rect 13564 6016 13884 7040
rect 13564 5952 13572 6016
rect 13636 5952 13652 6016
rect 13716 5952 13732 6016
rect 13796 5952 13812 6016
rect 13876 5952 13884 6016
rect 13564 4928 13884 5952
rect 13564 4864 13572 4928
rect 13636 4864 13652 4928
rect 13716 4864 13732 4928
rect 13796 4864 13812 4928
rect 13876 4864 13884 4928
rect 13564 3840 13884 4864
rect 13564 3776 13572 3840
rect 13636 3776 13652 3840
rect 13716 3776 13732 3840
rect 13796 3776 13812 3840
rect 13876 3776 13884 3840
rect 13564 2752 13884 3776
rect 13564 2688 13572 2752
rect 13636 2688 13652 2752
rect 13716 2688 13732 2752
rect 13796 2688 13812 2752
rect 13876 2688 13884 2752
rect 13564 1664 13884 2688
rect 13564 1600 13572 1664
rect 13636 1600 13652 1664
rect 13716 1600 13732 1664
rect 13796 1600 13812 1664
rect 13876 1600 13884 1664
rect 13564 1040 13884 1600
rect 16064 22880 16384 22896
rect 16064 22816 16072 22880
rect 16136 22816 16152 22880
rect 16216 22816 16232 22880
rect 16296 22816 16312 22880
rect 16376 22816 16384 22880
rect 16064 21792 16384 22816
rect 16064 21728 16072 21792
rect 16136 21728 16152 21792
rect 16216 21728 16232 21792
rect 16296 21728 16312 21792
rect 16376 21728 16384 21792
rect 16064 20704 16384 21728
rect 18564 22336 18884 22896
rect 21064 22880 21384 22896
rect 21064 22816 21072 22880
rect 21136 22816 21152 22880
rect 21216 22816 21232 22880
rect 21296 22816 21312 22880
rect 21376 22816 21384 22880
rect 19195 22540 19261 22541
rect 19195 22476 19196 22540
rect 19260 22476 19261 22540
rect 19195 22475 19261 22476
rect 18564 22272 18572 22336
rect 18636 22272 18652 22336
rect 18716 22272 18732 22336
rect 18796 22272 18812 22336
rect 18876 22272 18884 22336
rect 18564 21248 18884 22272
rect 18564 21184 18572 21248
rect 18636 21184 18652 21248
rect 18716 21184 18732 21248
rect 18796 21184 18812 21248
rect 18876 21184 18884 21248
rect 16987 20772 17053 20773
rect 16987 20708 16988 20772
rect 17052 20708 17053 20772
rect 16987 20707 17053 20708
rect 17539 20772 17605 20773
rect 17539 20708 17540 20772
rect 17604 20708 17605 20772
rect 17539 20707 17605 20708
rect 16064 20640 16072 20704
rect 16136 20640 16152 20704
rect 16216 20640 16232 20704
rect 16296 20640 16312 20704
rect 16376 20640 16384 20704
rect 16064 19616 16384 20640
rect 16064 19552 16072 19616
rect 16136 19552 16152 19616
rect 16216 19552 16232 19616
rect 16296 19552 16312 19616
rect 16376 19552 16384 19616
rect 16064 18528 16384 19552
rect 16064 18464 16072 18528
rect 16136 18464 16152 18528
rect 16216 18464 16232 18528
rect 16296 18464 16312 18528
rect 16376 18464 16384 18528
rect 16064 17440 16384 18464
rect 16064 17376 16072 17440
rect 16136 17376 16152 17440
rect 16216 17376 16232 17440
rect 16296 17376 16312 17440
rect 16376 17376 16384 17440
rect 16064 16352 16384 17376
rect 16064 16288 16072 16352
rect 16136 16288 16152 16352
rect 16216 16288 16232 16352
rect 16296 16288 16312 16352
rect 16376 16288 16384 16352
rect 16064 15264 16384 16288
rect 16064 15200 16072 15264
rect 16136 15200 16152 15264
rect 16216 15200 16232 15264
rect 16296 15200 16312 15264
rect 16376 15200 16384 15264
rect 16064 14176 16384 15200
rect 16064 14112 16072 14176
rect 16136 14112 16152 14176
rect 16216 14112 16232 14176
rect 16296 14112 16312 14176
rect 16376 14112 16384 14176
rect 16064 13088 16384 14112
rect 16064 13024 16072 13088
rect 16136 13024 16152 13088
rect 16216 13024 16232 13088
rect 16296 13024 16312 13088
rect 16376 13024 16384 13088
rect 16064 12000 16384 13024
rect 16064 11936 16072 12000
rect 16136 11936 16152 12000
rect 16216 11936 16232 12000
rect 16296 11936 16312 12000
rect 16376 11936 16384 12000
rect 16064 10912 16384 11936
rect 16064 10848 16072 10912
rect 16136 10848 16152 10912
rect 16216 10848 16232 10912
rect 16296 10848 16312 10912
rect 16376 10848 16384 10912
rect 16064 9824 16384 10848
rect 16064 9760 16072 9824
rect 16136 9760 16152 9824
rect 16216 9760 16232 9824
rect 16296 9760 16312 9824
rect 16376 9760 16384 9824
rect 16064 8736 16384 9760
rect 16064 8672 16072 8736
rect 16136 8672 16152 8736
rect 16216 8672 16232 8736
rect 16296 8672 16312 8736
rect 16376 8672 16384 8736
rect 16064 7648 16384 8672
rect 16064 7584 16072 7648
rect 16136 7584 16152 7648
rect 16216 7584 16232 7648
rect 16296 7584 16312 7648
rect 16376 7584 16384 7648
rect 16064 6560 16384 7584
rect 16064 6496 16072 6560
rect 16136 6496 16152 6560
rect 16216 6496 16232 6560
rect 16296 6496 16312 6560
rect 16376 6496 16384 6560
rect 16064 5472 16384 6496
rect 16990 6493 17050 20707
rect 17542 6901 17602 20707
rect 18564 20160 18884 21184
rect 18564 20096 18572 20160
rect 18636 20096 18652 20160
rect 18716 20096 18732 20160
rect 18796 20096 18812 20160
rect 18876 20096 18884 20160
rect 18564 19072 18884 20096
rect 18564 19008 18572 19072
rect 18636 19008 18652 19072
rect 18716 19008 18732 19072
rect 18796 19008 18812 19072
rect 18876 19008 18884 19072
rect 18564 17984 18884 19008
rect 18564 17920 18572 17984
rect 18636 17920 18652 17984
rect 18716 17920 18732 17984
rect 18796 17920 18812 17984
rect 18876 17920 18884 17984
rect 18564 16896 18884 17920
rect 18564 16832 18572 16896
rect 18636 16832 18652 16896
rect 18716 16832 18732 16896
rect 18796 16832 18812 16896
rect 18876 16832 18884 16896
rect 18564 15808 18884 16832
rect 18564 15744 18572 15808
rect 18636 15744 18652 15808
rect 18716 15744 18732 15808
rect 18796 15744 18812 15808
rect 18876 15744 18884 15808
rect 18564 14720 18884 15744
rect 18564 14656 18572 14720
rect 18636 14656 18652 14720
rect 18716 14656 18732 14720
rect 18796 14656 18812 14720
rect 18876 14656 18884 14720
rect 18564 13632 18884 14656
rect 19011 14516 19077 14517
rect 19011 14452 19012 14516
rect 19076 14452 19077 14516
rect 19011 14451 19077 14452
rect 18564 13568 18572 13632
rect 18636 13568 18652 13632
rect 18716 13568 18732 13632
rect 18796 13568 18812 13632
rect 18876 13568 18884 13632
rect 18564 12544 18884 13568
rect 18564 12480 18572 12544
rect 18636 12480 18652 12544
rect 18716 12480 18732 12544
rect 18796 12480 18812 12544
rect 18876 12480 18884 12544
rect 18564 11456 18884 12480
rect 18564 11392 18572 11456
rect 18636 11392 18652 11456
rect 18716 11392 18732 11456
rect 18796 11392 18812 11456
rect 18876 11392 18884 11456
rect 18564 10368 18884 11392
rect 19014 11253 19074 14451
rect 19011 11252 19077 11253
rect 19011 11188 19012 11252
rect 19076 11188 19077 11252
rect 19011 11187 19077 11188
rect 18564 10304 18572 10368
rect 18636 10304 18652 10368
rect 18716 10304 18732 10368
rect 18796 10304 18812 10368
rect 18876 10304 18884 10368
rect 18564 9280 18884 10304
rect 18564 9216 18572 9280
rect 18636 9216 18652 9280
rect 18716 9216 18732 9280
rect 18796 9216 18812 9280
rect 18876 9216 18884 9280
rect 18564 8192 18884 9216
rect 18564 8128 18572 8192
rect 18636 8128 18652 8192
rect 18716 8128 18732 8192
rect 18796 8128 18812 8192
rect 18876 8128 18884 8192
rect 18564 7104 18884 8128
rect 18564 7040 18572 7104
rect 18636 7040 18652 7104
rect 18716 7040 18732 7104
rect 18796 7040 18812 7104
rect 18876 7040 18884 7104
rect 17539 6900 17605 6901
rect 17539 6836 17540 6900
rect 17604 6836 17605 6900
rect 17539 6835 17605 6836
rect 16987 6492 17053 6493
rect 16987 6428 16988 6492
rect 17052 6428 17053 6492
rect 16987 6427 17053 6428
rect 16064 5408 16072 5472
rect 16136 5408 16152 5472
rect 16216 5408 16232 5472
rect 16296 5408 16312 5472
rect 16376 5408 16384 5472
rect 16064 4384 16384 5408
rect 16064 4320 16072 4384
rect 16136 4320 16152 4384
rect 16216 4320 16232 4384
rect 16296 4320 16312 4384
rect 16376 4320 16384 4384
rect 16064 3296 16384 4320
rect 16064 3232 16072 3296
rect 16136 3232 16152 3296
rect 16216 3232 16232 3296
rect 16296 3232 16312 3296
rect 16376 3232 16384 3296
rect 16064 2208 16384 3232
rect 16990 2957 17050 6427
rect 17542 5541 17602 6835
rect 18564 6016 18884 7040
rect 18564 5952 18572 6016
rect 18636 5952 18652 6016
rect 18716 5952 18732 6016
rect 18796 5952 18812 6016
rect 18876 5952 18884 6016
rect 17539 5540 17605 5541
rect 17539 5476 17540 5540
rect 17604 5476 17605 5540
rect 17539 5475 17605 5476
rect 18564 4928 18884 5952
rect 19198 5269 19258 22475
rect 21064 21792 21384 22816
rect 21064 21728 21072 21792
rect 21136 21728 21152 21792
rect 21216 21728 21232 21792
rect 21296 21728 21312 21792
rect 21376 21728 21384 21792
rect 19931 21724 19997 21725
rect 19931 21660 19932 21724
rect 19996 21660 19997 21724
rect 19931 21659 19997 21660
rect 19747 20772 19813 20773
rect 19747 20708 19748 20772
rect 19812 20708 19813 20772
rect 19747 20707 19813 20708
rect 19750 6901 19810 20707
rect 19747 6900 19813 6901
rect 19747 6836 19748 6900
rect 19812 6836 19813 6900
rect 19747 6835 19813 6836
rect 19934 5541 19994 21659
rect 21064 20704 21384 21728
rect 23564 22336 23884 22896
rect 23564 22272 23572 22336
rect 23636 22272 23652 22336
rect 23716 22272 23732 22336
rect 23796 22272 23812 22336
rect 23876 22272 23884 22336
rect 23564 21248 23884 22272
rect 26064 22880 26384 22896
rect 26064 22816 26072 22880
rect 26136 22816 26152 22880
rect 26216 22816 26232 22880
rect 26296 22816 26312 22880
rect 26376 22816 26384 22880
rect 25819 22132 25885 22133
rect 25819 22068 25820 22132
rect 25884 22068 25885 22132
rect 25819 22067 25885 22068
rect 23564 21184 23572 21248
rect 23636 21184 23652 21248
rect 23716 21184 23732 21248
rect 23796 21184 23812 21248
rect 23876 21184 23884 21248
rect 21587 20772 21653 20773
rect 21587 20708 21588 20772
rect 21652 20708 21653 20772
rect 21587 20707 21653 20708
rect 23243 20772 23309 20773
rect 23243 20708 23244 20772
rect 23308 20708 23309 20772
rect 23243 20707 23309 20708
rect 21064 20640 21072 20704
rect 21136 20640 21152 20704
rect 21216 20640 21232 20704
rect 21296 20640 21312 20704
rect 21376 20640 21384 20704
rect 21064 19616 21384 20640
rect 21064 19552 21072 19616
rect 21136 19552 21152 19616
rect 21216 19552 21232 19616
rect 21296 19552 21312 19616
rect 21376 19552 21384 19616
rect 21064 18528 21384 19552
rect 21064 18464 21072 18528
rect 21136 18464 21152 18528
rect 21216 18464 21232 18528
rect 21296 18464 21312 18528
rect 21376 18464 21384 18528
rect 21064 17440 21384 18464
rect 21064 17376 21072 17440
rect 21136 17376 21152 17440
rect 21216 17376 21232 17440
rect 21296 17376 21312 17440
rect 21376 17376 21384 17440
rect 21064 16352 21384 17376
rect 21064 16288 21072 16352
rect 21136 16288 21152 16352
rect 21216 16288 21232 16352
rect 21296 16288 21312 16352
rect 21376 16288 21384 16352
rect 21064 15264 21384 16288
rect 21064 15200 21072 15264
rect 21136 15200 21152 15264
rect 21216 15200 21232 15264
rect 21296 15200 21312 15264
rect 21376 15200 21384 15264
rect 21064 14176 21384 15200
rect 21064 14112 21072 14176
rect 21136 14112 21152 14176
rect 21216 14112 21232 14176
rect 21296 14112 21312 14176
rect 21376 14112 21384 14176
rect 21064 13088 21384 14112
rect 21064 13024 21072 13088
rect 21136 13024 21152 13088
rect 21216 13024 21232 13088
rect 21296 13024 21312 13088
rect 21376 13024 21384 13088
rect 21064 12000 21384 13024
rect 21064 11936 21072 12000
rect 21136 11936 21152 12000
rect 21216 11936 21232 12000
rect 21296 11936 21312 12000
rect 21376 11936 21384 12000
rect 21064 10912 21384 11936
rect 21064 10848 21072 10912
rect 21136 10848 21152 10912
rect 21216 10848 21232 10912
rect 21296 10848 21312 10912
rect 21376 10848 21384 10912
rect 21064 9824 21384 10848
rect 21064 9760 21072 9824
rect 21136 9760 21152 9824
rect 21216 9760 21232 9824
rect 21296 9760 21312 9824
rect 21376 9760 21384 9824
rect 21064 8736 21384 9760
rect 21064 8672 21072 8736
rect 21136 8672 21152 8736
rect 21216 8672 21232 8736
rect 21296 8672 21312 8736
rect 21376 8672 21384 8736
rect 21064 7648 21384 8672
rect 21064 7584 21072 7648
rect 21136 7584 21152 7648
rect 21216 7584 21232 7648
rect 21296 7584 21312 7648
rect 21376 7584 21384 7648
rect 21064 6560 21384 7584
rect 21064 6496 21072 6560
rect 21136 6496 21152 6560
rect 21216 6496 21232 6560
rect 21296 6496 21312 6560
rect 21376 6496 21384 6560
rect 19931 5540 19997 5541
rect 19931 5476 19932 5540
rect 19996 5476 19997 5540
rect 19931 5475 19997 5476
rect 21064 5472 21384 6496
rect 21590 5541 21650 20707
rect 23059 19820 23125 19821
rect 23059 19756 23060 19820
rect 23124 19756 23125 19820
rect 23059 19755 23125 19756
rect 21955 18732 22021 18733
rect 21955 18668 21956 18732
rect 22020 18668 22021 18732
rect 21955 18667 22021 18668
rect 21587 5540 21653 5541
rect 21587 5476 21588 5540
rect 21652 5476 21653 5540
rect 21587 5475 21653 5476
rect 21064 5408 21072 5472
rect 21136 5408 21152 5472
rect 21216 5408 21232 5472
rect 21296 5408 21312 5472
rect 21376 5408 21384 5472
rect 19195 5268 19261 5269
rect 19195 5204 19196 5268
rect 19260 5204 19261 5268
rect 19195 5203 19261 5204
rect 18564 4864 18572 4928
rect 18636 4864 18652 4928
rect 18716 4864 18732 4928
rect 18796 4864 18812 4928
rect 18876 4864 18884 4928
rect 18564 3840 18884 4864
rect 19198 4045 19258 5203
rect 21064 4384 21384 5408
rect 21064 4320 21072 4384
rect 21136 4320 21152 4384
rect 21216 4320 21232 4384
rect 21296 4320 21312 4384
rect 21376 4320 21384 4384
rect 19195 4044 19261 4045
rect 19195 3980 19196 4044
rect 19260 3980 19261 4044
rect 19195 3979 19261 3980
rect 18564 3776 18572 3840
rect 18636 3776 18652 3840
rect 18716 3776 18732 3840
rect 18796 3776 18812 3840
rect 18876 3776 18884 3840
rect 16987 2956 17053 2957
rect 16987 2892 16988 2956
rect 17052 2892 17053 2956
rect 16987 2891 17053 2892
rect 16064 2144 16072 2208
rect 16136 2144 16152 2208
rect 16216 2144 16232 2208
rect 16296 2144 16312 2208
rect 16376 2144 16384 2208
rect 16064 1120 16384 2144
rect 16064 1056 16072 1120
rect 16136 1056 16152 1120
rect 16216 1056 16232 1120
rect 16296 1056 16312 1120
rect 16376 1056 16384 1120
rect 16064 1040 16384 1056
rect 18564 2752 18884 3776
rect 18564 2688 18572 2752
rect 18636 2688 18652 2752
rect 18716 2688 18732 2752
rect 18796 2688 18812 2752
rect 18876 2688 18884 2752
rect 18564 1664 18884 2688
rect 18564 1600 18572 1664
rect 18636 1600 18652 1664
rect 18716 1600 18732 1664
rect 18796 1600 18812 1664
rect 18876 1600 18884 1664
rect 18564 1040 18884 1600
rect 21064 3296 21384 4320
rect 21064 3232 21072 3296
rect 21136 3232 21152 3296
rect 21216 3232 21232 3296
rect 21296 3232 21312 3296
rect 21376 3232 21384 3296
rect 21064 2208 21384 3232
rect 21064 2144 21072 2208
rect 21136 2144 21152 2208
rect 21216 2144 21232 2208
rect 21296 2144 21312 2208
rect 21376 2144 21384 2208
rect 21064 1120 21384 2144
rect 21590 2005 21650 5475
rect 21958 5405 22018 18667
rect 22875 17236 22941 17237
rect 22875 17172 22876 17236
rect 22940 17172 22941 17236
rect 22875 17171 22941 17172
rect 22691 14924 22757 14925
rect 22691 14860 22692 14924
rect 22756 14860 22757 14924
rect 22691 14859 22757 14860
rect 22694 5949 22754 14859
rect 22878 6901 22938 17171
rect 23062 7037 23122 19755
rect 23059 7036 23125 7037
rect 23059 6972 23060 7036
rect 23124 6972 23125 7036
rect 23059 6971 23125 6972
rect 22875 6900 22941 6901
rect 22875 6836 22876 6900
rect 22940 6836 22941 6900
rect 22875 6835 22941 6836
rect 22691 5948 22757 5949
rect 22691 5884 22692 5948
rect 22756 5884 22757 5948
rect 22691 5883 22757 5884
rect 23246 5541 23306 20707
rect 23564 20160 23884 21184
rect 25451 20772 25517 20773
rect 25451 20708 25452 20772
rect 25516 20708 25517 20772
rect 25451 20707 25517 20708
rect 23564 20096 23572 20160
rect 23636 20096 23652 20160
rect 23716 20096 23732 20160
rect 23796 20096 23812 20160
rect 23876 20096 23884 20160
rect 23564 19072 23884 20096
rect 24347 19412 24413 19413
rect 24347 19348 24348 19412
rect 24412 19348 24413 19412
rect 24347 19347 24413 19348
rect 23564 19008 23572 19072
rect 23636 19008 23652 19072
rect 23716 19008 23732 19072
rect 23796 19008 23812 19072
rect 23876 19008 23884 19072
rect 23564 17984 23884 19008
rect 23564 17920 23572 17984
rect 23636 17920 23652 17984
rect 23716 17920 23732 17984
rect 23796 17920 23812 17984
rect 23876 17920 23884 17984
rect 23564 16896 23884 17920
rect 23564 16832 23572 16896
rect 23636 16832 23652 16896
rect 23716 16832 23732 16896
rect 23796 16832 23812 16896
rect 23876 16832 23884 16896
rect 23564 15808 23884 16832
rect 23564 15744 23572 15808
rect 23636 15744 23652 15808
rect 23716 15744 23732 15808
rect 23796 15744 23812 15808
rect 23876 15744 23884 15808
rect 23564 14720 23884 15744
rect 23564 14656 23572 14720
rect 23636 14656 23652 14720
rect 23716 14656 23732 14720
rect 23796 14656 23812 14720
rect 23876 14656 23884 14720
rect 23564 13632 23884 14656
rect 23564 13568 23572 13632
rect 23636 13568 23652 13632
rect 23716 13568 23732 13632
rect 23796 13568 23812 13632
rect 23876 13568 23884 13632
rect 23564 12544 23884 13568
rect 23564 12480 23572 12544
rect 23636 12480 23652 12544
rect 23716 12480 23732 12544
rect 23796 12480 23812 12544
rect 23876 12480 23884 12544
rect 23564 11456 23884 12480
rect 23564 11392 23572 11456
rect 23636 11392 23652 11456
rect 23716 11392 23732 11456
rect 23796 11392 23812 11456
rect 23876 11392 23884 11456
rect 23564 10368 23884 11392
rect 23564 10304 23572 10368
rect 23636 10304 23652 10368
rect 23716 10304 23732 10368
rect 23796 10304 23812 10368
rect 23876 10304 23884 10368
rect 23564 9280 23884 10304
rect 23564 9216 23572 9280
rect 23636 9216 23652 9280
rect 23716 9216 23732 9280
rect 23796 9216 23812 9280
rect 23876 9216 23884 9280
rect 23564 8192 23884 9216
rect 23564 8128 23572 8192
rect 23636 8128 23652 8192
rect 23716 8128 23732 8192
rect 23796 8128 23812 8192
rect 23876 8128 23884 8192
rect 23564 7104 23884 8128
rect 23564 7040 23572 7104
rect 23636 7040 23652 7104
rect 23716 7040 23732 7104
rect 23796 7040 23812 7104
rect 23876 7040 23884 7104
rect 23564 6016 23884 7040
rect 24350 6901 24410 19347
rect 24347 6900 24413 6901
rect 24347 6836 24348 6900
rect 24412 6836 24413 6900
rect 24347 6835 24413 6836
rect 23564 5952 23572 6016
rect 23636 5952 23652 6016
rect 23716 5952 23732 6016
rect 23796 5952 23812 6016
rect 23876 5952 23884 6016
rect 23243 5540 23309 5541
rect 23243 5476 23244 5540
rect 23308 5476 23309 5540
rect 23243 5475 23309 5476
rect 21955 5404 22021 5405
rect 21955 5340 21956 5404
rect 22020 5340 22021 5404
rect 21955 5339 22021 5340
rect 23564 4928 23884 5952
rect 25454 5541 25514 20707
rect 25635 19820 25701 19821
rect 25635 19756 25636 19820
rect 25700 19756 25701 19820
rect 25635 19755 25701 19756
rect 25638 7853 25698 19755
rect 25635 7852 25701 7853
rect 25635 7788 25636 7852
rect 25700 7788 25701 7852
rect 25635 7787 25701 7788
rect 25822 6901 25882 22067
rect 26064 21792 26384 22816
rect 28564 22336 28884 22896
rect 28564 22272 28572 22336
rect 28636 22272 28652 22336
rect 28716 22272 28732 22336
rect 28796 22272 28812 22336
rect 28876 22272 28884 22336
rect 28211 22132 28277 22133
rect 28211 22068 28212 22132
rect 28276 22068 28277 22132
rect 28211 22067 28277 22068
rect 26064 21728 26072 21792
rect 26136 21728 26152 21792
rect 26216 21728 26232 21792
rect 26296 21728 26312 21792
rect 26376 21728 26384 21792
rect 26064 20704 26384 21728
rect 26739 21724 26805 21725
rect 26739 21660 26740 21724
rect 26804 21660 26805 21724
rect 26739 21659 26805 21660
rect 26742 20909 26802 21659
rect 27659 21180 27725 21181
rect 27659 21116 27660 21180
rect 27724 21116 27725 21180
rect 27659 21115 27725 21116
rect 26739 20908 26805 20909
rect 26739 20844 26740 20908
rect 26804 20844 26805 20908
rect 26739 20843 26805 20844
rect 26064 20640 26072 20704
rect 26136 20640 26152 20704
rect 26216 20640 26232 20704
rect 26296 20640 26312 20704
rect 26376 20640 26384 20704
rect 26064 19616 26384 20640
rect 26555 20364 26621 20365
rect 26555 20300 26556 20364
rect 26620 20300 26621 20364
rect 26555 20299 26621 20300
rect 26064 19552 26072 19616
rect 26136 19552 26152 19616
rect 26216 19552 26232 19616
rect 26296 19552 26312 19616
rect 26376 19552 26384 19616
rect 26064 18528 26384 19552
rect 26064 18464 26072 18528
rect 26136 18464 26152 18528
rect 26216 18464 26232 18528
rect 26296 18464 26312 18528
rect 26376 18464 26384 18528
rect 26064 17440 26384 18464
rect 26064 17376 26072 17440
rect 26136 17376 26152 17440
rect 26216 17376 26232 17440
rect 26296 17376 26312 17440
rect 26376 17376 26384 17440
rect 26064 16352 26384 17376
rect 26064 16288 26072 16352
rect 26136 16288 26152 16352
rect 26216 16288 26232 16352
rect 26296 16288 26312 16352
rect 26376 16288 26384 16352
rect 26064 15264 26384 16288
rect 26064 15200 26072 15264
rect 26136 15200 26152 15264
rect 26216 15200 26232 15264
rect 26296 15200 26312 15264
rect 26376 15200 26384 15264
rect 26064 14176 26384 15200
rect 26064 14112 26072 14176
rect 26136 14112 26152 14176
rect 26216 14112 26232 14176
rect 26296 14112 26312 14176
rect 26376 14112 26384 14176
rect 26064 13088 26384 14112
rect 26064 13024 26072 13088
rect 26136 13024 26152 13088
rect 26216 13024 26232 13088
rect 26296 13024 26312 13088
rect 26376 13024 26384 13088
rect 26064 12000 26384 13024
rect 26064 11936 26072 12000
rect 26136 11936 26152 12000
rect 26216 11936 26232 12000
rect 26296 11936 26312 12000
rect 26376 11936 26384 12000
rect 26064 10912 26384 11936
rect 26064 10848 26072 10912
rect 26136 10848 26152 10912
rect 26216 10848 26232 10912
rect 26296 10848 26312 10912
rect 26376 10848 26384 10912
rect 26064 9824 26384 10848
rect 26064 9760 26072 9824
rect 26136 9760 26152 9824
rect 26216 9760 26232 9824
rect 26296 9760 26312 9824
rect 26376 9760 26384 9824
rect 26064 8736 26384 9760
rect 26064 8672 26072 8736
rect 26136 8672 26152 8736
rect 26216 8672 26232 8736
rect 26296 8672 26312 8736
rect 26376 8672 26384 8736
rect 26064 7648 26384 8672
rect 26064 7584 26072 7648
rect 26136 7584 26152 7648
rect 26216 7584 26232 7648
rect 26296 7584 26312 7648
rect 26376 7584 26384 7648
rect 25819 6900 25885 6901
rect 25819 6836 25820 6900
rect 25884 6836 25885 6900
rect 25819 6835 25885 6836
rect 26064 6560 26384 7584
rect 26064 6496 26072 6560
rect 26136 6496 26152 6560
rect 26216 6496 26232 6560
rect 26296 6496 26312 6560
rect 26376 6496 26384 6560
rect 25819 5812 25885 5813
rect 25819 5748 25820 5812
rect 25884 5748 25885 5812
rect 25819 5747 25885 5748
rect 25451 5540 25517 5541
rect 25451 5476 25452 5540
rect 25516 5476 25517 5540
rect 25451 5475 25517 5476
rect 23564 4864 23572 4928
rect 23636 4864 23652 4928
rect 23716 4864 23732 4928
rect 23796 4864 23812 4928
rect 23876 4864 23884 4928
rect 22691 4724 22757 4725
rect 22691 4660 22692 4724
rect 22756 4660 22757 4724
rect 22691 4659 22757 4660
rect 22694 2413 22754 4659
rect 23564 3840 23884 4864
rect 25822 4045 25882 5747
rect 26064 5472 26384 6496
rect 26064 5408 26072 5472
rect 26136 5408 26152 5472
rect 26216 5408 26232 5472
rect 26296 5408 26312 5472
rect 26376 5408 26384 5472
rect 26064 4384 26384 5408
rect 26558 5133 26618 20299
rect 26742 6085 26802 20843
rect 27662 20773 27722 21115
rect 27659 20772 27725 20773
rect 27659 20708 27660 20772
rect 27724 20708 27725 20772
rect 27659 20707 27725 20708
rect 26923 16012 26989 16013
rect 26923 15948 26924 16012
rect 26988 15948 26989 16012
rect 26923 15947 26989 15948
rect 26926 14109 26986 15947
rect 26923 14108 26989 14109
rect 26923 14044 26924 14108
rect 26988 14044 26989 14108
rect 26923 14043 26989 14044
rect 26739 6084 26805 6085
rect 26739 6020 26740 6084
rect 26804 6020 26805 6084
rect 26739 6019 26805 6020
rect 26555 5132 26621 5133
rect 26555 5068 26556 5132
rect 26620 5068 26621 5132
rect 26555 5067 26621 5068
rect 27662 4725 27722 20707
rect 28214 9621 28274 22067
rect 28564 21248 28884 22272
rect 28564 21184 28572 21248
rect 28636 21184 28652 21248
rect 28716 21184 28732 21248
rect 28796 21184 28812 21248
rect 28876 21184 28884 21248
rect 28564 20160 28884 21184
rect 28564 20096 28572 20160
rect 28636 20096 28652 20160
rect 28716 20096 28732 20160
rect 28796 20096 28812 20160
rect 28876 20096 28884 20160
rect 28564 19072 28884 20096
rect 28564 19008 28572 19072
rect 28636 19008 28652 19072
rect 28716 19008 28732 19072
rect 28796 19008 28812 19072
rect 28876 19008 28884 19072
rect 28564 17984 28884 19008
rect 28564 17920 28572 17984
rect 28636 17920 28652 17984
rect 28716 17920 28732 17984
rect 28796 17920 28812 17984
rect 28876 17920 28884 17984
rect 28564 16896 28884 17920
rect 31064 22880 31384 22896
rect 31064 22816 31072 22880
rect 31136 22816 31152 22880
rect 31216 22816 31232 22880
rect 31296 22816 31312 22880
rect 31376 22816 31384 22880
rect 31064 21792 31384 22816
rect 31064 21728 31072 21792
rect 31136 21728 31152 21792
rect 31216 21728 31232 21792
rect 31296 21728 31312 21792
rect 31376 21728 31384 21792
rect 31064 20704 31384 21728
rect 33564 22336 33884 22896
rect 33564 22272 33572 22336
rect 33636 22272 33652 22336
rect 33716 22272 33732 22336
rect 33796 22272 33812 22336
rect 33876 22272 33884 22336
rect 33564 21248 33884 22272
rect 33564 21184 33572 21248
rect 33636 21184 33652 21248
rect 33716 21184 33732 21248
rect 33796 21184 33812 21248
rect 33876 21184 33884 21248
rect 31891 20772 31957 20773
rect 31891 20708 31892 20772
rect 31956 20708 31957 20772
rect 31891 20707 31957 20708
rect 31064 20640 31072 20704
rect 31136 20640 31152 20704
rect 31216 20640 31232 20704
rect 31296 20640 31312 20704
rect 31376 20640 31384 20704
rect 31064 19616 31384 20640
rect 31064 19552 31072 19616
rect 31136 19552 31152 19616
rect 31216 19552 31232 19616
rect 31296 19552 31312 19616
rect 31376 19552 31384 19616
rect 31064 18528 31384 19552
rect 31064 18464 31072 18528
rect 31136 18464 31152 18528
rect 31216 18464 31232 18528
rect 31296 18464 31312 18528
rect 31376 18464 31384 18528
rect 30419 17508 30485 17509
rect 30419 17444 30420 17508
rect 30484 17444 30485 17508
rect 30419 17443 30485 17444
rect 28564 16832 28572 16896
rect 28636 16832 28652 16896
rect 28716 16832 28732 16896
rect 28796 16832 28812 16896
rect 28876 16832 28884 16896
rect 28564 15808 28884 16832
rect 30235 16012 30301 16013
rect 30235 15948 30236 16012
rect 30300 15948 30301 16012
rect 30235 15947 30301 15948
rect 28564 15744 28572 15808
rect 28636 15744 28652 15808
rect 28716 15744 28732 15808
rect 28796 15744 28812 15808
rect 28876 15744 28884 15808
rect 28564 14720 28884 15744
rect 29315 14924 29381 14925
rect 29315 14860 29316 14924
rect 29380 14860 29381 14924
rect 29315 14859 29381 14860
rect 28564 14656 28572 14720
rect 28636 14656 28652 14720
rect 28716 14656 28732 14720
rect 28796 14656 28812 14720
rect 28876 14656 28884 14720
rect 28564 13632 28884 14656
rect 28564 13568 28572 13632
rect 28636 13568 28652 13632
rect 28716 13568 28732 13632
rect 28796 13568 28812 13632
rect 28876 13568 28884 13632
rect 28564 12544 28884 13568
rect 28564 12480 28572 12544
rect 28636 12480 28652 12544
rect 28716 12480 28732 12544
rect 28796 12480 28812 12544
rect 28876 12480 28884 12544
rect 28564 11456 28884 12480
rect 28564 11392 28572 11456
rect 28636 11392 28652 11456
rect 28716 11392 28732 11456
rect 28796 11392 28812 11456
rect 28876 11392 28884 11456
rect 28564 10368 28884 11392
rect 29318 10981 29378 14859
rect 29315 10980 29381 10981
rect 29315 10916 29316 10980
rect 29380 10916 29381 10980
rect 29315 10915 29381 10916
rect 28564 10304 28572 10368
rect 28636 10304 28652 10368
rect 28716 10304 28732 10368
rect 28796 10304 28812 10368
rect 28876 10304 28884 10368
rect 28211 9620 28277 9621
rect 28211 9556 28212 9620
rect 28276 9556 28277 9620
rect 28211 9555 28277 9556
rect 28564 9280 28884 10304
rect 30238 9757 30298 15947
rect 30422 12749 30482 17443
rect 31064 17440 31384 18464
rect 31064 17376 31072 17440
rect 31136 17376 31152 17440
rect 31216 17376 31232 17440
rect 31296 17376 31312 17440
rect 31376 17376 31384 17440
rect 31064 16352 31384 17376
rect 31064 16288 31072 16352
rect 31136 16288 31152 16352
rect 31216 16288 31232 16352
rect 31296 16288 31312 16352
rect 31376 16288 31384 16352
rect 31064 15264 31384 16288
rect 31064 15200 31072 15264
rect 31136 15200 31152 15264
rect 31216 15200 31232 15264
rect 31296 15200 31312 15264
rect 31376 15200 31384 15264
rect 30787 14380 30853 14381
rect 30787 14316 30788 14380
rect 30852 14316 30853 14380
rect 30787 14315 30853 14316
rect 30419 12748 30485 12749
rect 30419 12684 30420 12748
rect 30484 12684 30485 12748
rect 30419 12683 30485 12684
rect 30790 12341 30850 14315
rect 31064 14176 31384 15200
rect 31064 14112 31072 14176
rect 31136 14112 31152 14176
rect 31216 14112 31232 14176
rect 31296 14112 31312 14176
rect 31376 14112 31384 14176
rect 31064 13088 31384 14112
rect 31064 13024 31072 13088
rect 31136 13024 31152 13088
rect 31216 13024 31232 13088
rect 31296 13024 31312 13088
rect 31376 13024 31384 13088
rect 30787 12340 30853 12341
rect 30787 12276 30788 12340
rect 30852 12276 30853 12340
rect 30787 12275 30853 12276
rect 30790 11117 30850 12275
rect 31064 12000 31384 13024
rect 31064 11936 31072 12000
rect 31136 11936 31152 12000
rect 31216 11936 31232 12000
rect 31296 11936 31312 12000
rect 31376 11936 31384 12000
rect 30787 11116 30853 11117
rect 30787 11052 30788 11116
rect 30852 11052 30853 11116
rect 30787 11051 30853 11052
rect 31064 10912 31384 11936
rect 31064 10848 31072 10912
rect 31136 10848 31152 10912
rect 31216 10848 31232 10912
rect 31296 10848 31312 10912
rect 31376 10848 31384 10912
rect 31064 9824 31384 10848
rect 31064 9760 31072 9824
rect 31136 9760 31152 9824
rect 31216 9760 31232 9824
rect 31296 9760 31312 9824
rect 31376 9760 31384 9824
rect 30235 9756 30301 9757
rect 30235 9692 30236 9756
rect 30300 9692 30301 9756
rect 30235 9691 30301 9692
rect 28564 9216 28572 9280
rect 28636 9216 28652 9280
rect 28716 9216 28732 9280
rect 28796 9216 28812 9280
rect 28876 9216 28884 9280
rect 28564 8192 28884 9216
rect 28564 8128 28572 8192
rect 28636 8128 28652 8192
rect 28716 8128 28732 8192
rect 28796 8128 28812 8192
rect 28876 8128 28884 8192
rect 28564 7104 28884 8128
rect 28564 7040 28572 7104
rect 28636 7040 28652 7104
rect 28716 7040 28732 7104
rect 28796 7040 28812 7104
rect 28876 7040 28884 7104
rect 28564 6016 28884 7040
rect 28564 5952 28572 6016
rect 28636 5952 28652 6016
rect 28716 5952 28732 6016
rect 28796 5952 28812 6016
rect 28876 5952 28884 6016
rect 28564 4928 28884 5952
rect 28564 4864 28572 4928
rect 28636 4864 28652 4928
rect 28716 4864 28732 4928
rect 28796 4864 28812 4928
rect 28876 4864 28884 4928
rect 27659 4724 27725 4725
rect 27659 4660 27660 4724
rect 27724 4660 27725 4724
rect 27659 4659 27725 4660
rect 26064 4320 26072 4384
rect 26136 4320 26152 4384
rect 26216 4320 26232 4384
rect 26296 4320 26312 4384
rect 26376 4320 26384 4384
rect 25819 4044 25885 4045
rect 25819 3980 25820 4044
rect 25884 3980 25885 4044
rect 25819 3979 25885 3980
rect 23564 3776 23572 3840
rect 23636 3776 23652 3840
rect 23716 3776 23732 3840
rect 23796 3776 23812 3840
rect 23876 3776 23884 3840
rect 23564 2752 23884 3776
rect 23564 2688 23572 2752
rect 23636 2688 23652 2752
rect 23716 2688 23732 2752
rect 23796 2688 23812 2752
rect 23876 2688 23884 2752
rect 22691 2412 22757 2413
rect 22691 2348 22692 2412
rect 22756 2348 22757 2412
rect 22691 2347 22757 2348
rect 21587 2004 21653 2005
rect 21587 1940 21588 2004
rect 21652 1940 21653 2004
rect 21587 1939 21653 1940
rect 21064 1056 21072 1120
rect 21136 1056 21152 1120
rect 21216 1056 21232 1120
rect 21296 1056 21312 1120
rect 21376 1056 21384 1120
rect 21064 1040 21384 1056
rect 23564 1664 23884 2688
rect 23564 1600 23572 1664
rect 23636 1600 23652 1664
rect 23716 1600 23732 1664
rect 23796 1600 23812 1664
rect 23876 1600 23884 1664
rect 23564 1040 23884 1600
rect 26064 3296 26384 4320
rect 26064 3232 26072 3296
rect 26136 3232 26152 3296
rect 26216 3232 26232 3296
rect 26296 3232 26312 3296
rect 26376 3232 26384 3296
rect 26064 2208 26384 3232
rect 26064 2144 26072 2208
rect 26136 2144 26152 2208
rect 26216 2144 26232 2208
rect 26296 2144 26312 2208
rect 26376 2144 26384 2208
rect 26064 1120 26384 2144
rect 26064 1056 26072 1120
rect 26136 1056 26152 1120
rect 26216 1056 26232 1120
rect 26296 1056 26312 1120
rect 26376 1056 26384 1120
rect 26064 1040 26384 1056
rect 28564 3840 28884 4864
rect 28564 3776 28572 3840
rect 28636 3776 28652 3840
rect 28716 3776 28732 3840
rect 28796 3776 28812 3840
rect 28876 3776 28884 3840
rect 28564 2752 28884 3776
rect 31064 8736 31384 9760
rect 31064 8672 31072 8736
rect 31136 8672 31152 8736
rect 31216 8672 31232 8736
rect 31296 8672 31312 8736
rect 31376 8672 31384 8736
rect 31064 7648 31384 8672
rect 31064 7584 31072 7648
rect 31136 7584 31152 7648
rect 31216 7584 31232 7648
rect 31296 7584 31312 7648
rect 31376 7584 31384 7648
rect 31064 6560 31384 7584
rect 31894 7309 31954 20707
rect 33564 20160 33884 21184
rect 33564 20096 33572 20160
rect 33636 20096 33652 20160
rect 33716 20096 33732 20160
rect 33796 20096 33812 20160
rect 33876 20096 33884 20160
rect 33564 19072 33884 20096
rect 33564 19008 33572 19072
rect 33636 19008 33652 19072
rect 33716 19008 33732 19072
rect 33796 19008 33812 19072
rect 33876 19008 33884 19072
rect 33564 17984 33884 19008
rect 33564 17920 33572 17984
rect 33636 17920 33652 17984
rect 33716 17920 33732 17984
rect 33796 17920 33812 17984
rect 33876 17920 33884 17984
rect 32811 17236 32877 17237
rect 32811 17172 32812 17236
rect 32876 17172 32877 17236
rect 32811 17171 32877 17172
rect 32814 9621 32874 17171
rect 33564 16896 33884 17920
rect 33564 16832 33572 16896
rect 33636 16832 33652 16896
rect 33716 16832 33732 16896
rect 33796 16832 33812 16896
rect 33876 16832 33884 16896
rect 33179 16556 33245 16557
rect 33179 16492 33180 16556
rect 33244 16492 33245 16556
rect 33179 16491 33245 16492
rect 32811 9620 32877 9621
rect 32811 9556 32812 9620
rect 32876 9556 32877 9620
rect 32811 9555 32877 9556
rect 31891 7308 31957 7309
rect 31891 7244 31892 7308
rect 31956 7244 31957 7308
rect 31891 7243 31957 7244
rect 31064 6496 31072 6560
rect 31136 6496 31152 6560
rect 31216 6496 31232 6560
rect 31296 6496 31312 6560
rect 31376 6496 31384 6560
rect 31064 5472 31384 6496
rect 33182 5677 33242 16491
rect 33564 15808 33884 16832
rect 33564 15744 33572 15808
rect 33636 15744 33652 15808
rect 33716 15744 33732 15808
rect 33796 15744 33812 15808
rect 33876 15744 33884 15808
rect 33564 14720 33884 15744
rect 33564 14656 33572 14720
rect 33636 14656 33652 14720
rect 33716 14656 33732 14720
rect 33796 14656 33812 14720
rect 33876 14656 33884 14720
rect 33564 13632 33884 14656
rect 33564 13568 33572 13632
rect 33636 13568 33652 13632
rect 33716 13568 33732 13632
rect 33796 13568 33812 13632
rect 33876 13568 33884 13632
rect 33564 12544 33884 13568
rect 33564 12480 33572 12544
rect 33636 12480 33652 12544
rect 33716 12480 33732 12544
rect 33796 12480 33812 12544
rect 33876 12480 33884 12544
rect 33564 11456 33884 12480
rect 33564 11392 33572 11456
rect 33636 11392 33652 11456
rect 33716 11392 33732 11456
rect 33796 11392 33812 11456
rect 33876 11392 33884 11456
rect 33564 10368 33884 11392
rect 33564 10304 33572 10368
rect 33636 10304 33652 10368
rect 33716 10304 33732 10368
rect 33796 10304 33812 10368
rect 33876 10304 33884 10368
rect 33564 9280 33884 10304
rect 33564 9216 33572 9280
rect 33636 9216 33652 9280
rect 33716 9216 33732 9280
rect 33796 9216 33812 9280
rect 33876 9216 33884 9280
rect 33564 8192 33884 9216
rect 36064 22880 36384 22896
rect 36064 22816 36072 22880
rect 36136 22816 36152 22880
rect 36216 22816 36232 22880
rect 36296 22816 36312 22880
rect 36376 22816 36384 22880
rect 36064 21792 36384 22816
rect 36064 21728 36072 21792
rect 36136 21728 36152 21792
rect 36216 21728 36232 21792
rect 36296 21728 36312 21792
rect 36376 21728 36384 21792
rect 36064 20704 36384 21728
rect 36064 20640 36072 20704
rect 36136 20640 36152 20704
rect 36216 20640 36232 20704
rect 36296 20640 36312 20704
rect 36376 20640 36384 20704
rect 36064 19616 36384 20640
rect 36064 19552 36072 19616
rect 36136 19552 36152 19616
rect 36216 19552 36232 19616
rect 36296 19552 36312 19616
rect 36376 19552 36384 19616
rect 36064 18528 36384 19552
rect 36064 18464 36072 18528
rect 36136 18464 36152 18528
rect 36216 18464 36232 18528
rect 36296 18464 36312 18528
rect 36376 18464 36384 18528
rect 36064 17440 36384 18464
rect 36064 17376 36072 17440
rect 36136 17376 36152 17440
rect 36216 17376 36232 17440
rect 36296 17376 36312 17440
rect 36376 17376 36384 17440
rect 36064 16352 36384 17376
rect 36064 16288 36072 16352
rect 36136 16288 36152 16352
rect 36216 16288 36232 16352
rect 36296 16288 36312 16352
rect 36376 16288 36384 16352
rect 36064 15264 36384 16288
rect 36064 15200 36072 15264
rect 36136 15200 36152 15264
rect 36216 15200 36232 15264
rect 36296 15200 36312 15264
rect 36376 15200 36384 15264
rect 36064 14176 36384 15200
rect 36064 14112 36072 14176
rect 36136 14112 36152 14176
rect 36216 14112 36232 14176
rect 36296 14112 36312 14176
rect 36376 14112 36384 14176
rect 36064 13088 36384 14112
rect 36064 13024 36072 13088
rect 36136 13024 36152 13088
rect 36216 13024 36232 13088
rect 36296 13024 36312 13088
rect 36376 13024 36384 13088
rect 36064 12000 36384 13024
rect 36064 11936 36072 12000
rect 36136 11936 36152 12000
rect 36216 11936 36232 12000
rect 36296 11936 36312 12000
rect 36376 11936 36384 12000
rect 36064 10912 36384 11936
rect 36064 10848 36072 10912
rect 36136 10848 36152 10912
rect 36216 10848 36232 10912
rect 36296 10848 36312 10912
rect 36376 10848 36384 10912
rect 36064 9824 36384 10848
rect 36064 9760 36072 9824
rect 36136 9760 36152 9824
rect 36216 9760 36232 9824
rect 36296 9760 36312 9824
rect 36376 9760 36384 9824
rect 36064 8736 36384 9760
rect 36064 8672 36072 8736
rect 36136 8672 36152 8736
rect 36216 8672 36232 8736
rect 36296 8672 36312 8736
rect 36376 8672 36384 8736
rect 34283 8396 34349 8397
rect 34283 8332 34284 8396
rect 34348 8332 34349 8396
rect 34283 8331 34349 8332
rect 34467 8396 34533 8397
rect 34467 8332 34468 8396
rect 34532 8332 34533 8396
rect 34467 8331 34533 8332
rect 33564 8128 33572 8192
rect 33636 8128 33652 8192
rect 33716 8128 33732 8192
rect 33796 8128 33812 8192
rect 33876 8128 33884 8192
rect 33564 7104 33884 8128
rect 33564 7040 33572 7104
rect 33636 7040 33652 7104
rect 33716 7040 33732 7104
rect 33796 7040 33812 7104
rect 33876 7040 33884 7104
rect 33564 6016 33884 7040
rect 33564 5952 33572 6016
rect 33636 5952 33652 6016
rect 33716 5952 33732 6016
rect 33796 5952 33812 6016
rect 33876 5952 33884 6016
rect 33179 5676 33245 5677
rect 33179 5612 33180 5676
rect 33244 5612 33245 5676
rect 33179 5611 33245 5612
rect 31064 5408 31072 5472
rect 31136 5408 31152 5472
rect 31216 5408 31232 5472
rect 31296 5408 31312 5472
rect 31376 5408 31384 5472
rect 31064 4384 31384 5408
rect 31064 4320 31072 4384
rect 31136 4320 31152 4384
rect 31216 4320 31232 4384
rect 31296 4320 31312 4384
rect 31376 4320 31384 4384
rect 31064 3296 31384 4320
rect 31064 3232 31072 3296
rect 31136 3232 31152 3296
rect 31216 3232 31232 3296
rect 31296 3232 31312 3296
rect 31376 3232 31384 3296
rect 28947 3092 29013 3093
rect 28947 3028 28948 3092
rect 29012 3028 29013 3092
rect 28947 3027 29013 3028
rect 28564 2688 28572 2752
rect 28636 2688 28652 2752
rect 28716 2688 28732 2752
rect 28796 2688 28812 2752
rect 28876 2688 28884 2752
rect 28564 1664 28884 2688
rect 28564 1600 28572 1664
rect 28636 1600 28652 1664
rect 28716 1600 28732 1664
rect 28796 1600 28812 1664
rect 28876 1600 28884 1664
rect 28564 1040 28884 1600
rect 28950 1325 29010 3027
rect 31064 2208 31384 3232
rect 31064 2144 31072 2208
rect 31136 2144 31152 2208
rect 31216 2144 31232 2208
rect 31296 2144 31312 2208
rect 31376 2144 31384 2208
rect 28947 1324 29013 1325
rect 28947 1260 28948 1324
rect 29012 1260 29013 1324
rect 28947 1259 29013 1260
rect 31064 1120 31384 2144
rect 31064 1056 31072 1120
rect 31136 1056 31152 1120
rect 31216 1056 31232 1120
rect 31296 1056 31312 1120
rect 31376 1056 31384 1120
rect 31064 1040 31384 1056
rect 33564 4928 33884 5952
rect 33564 4864 33572 4928
rect 33636 4864 33652 4928
rect 33716 4864 33732 4928
rect 33796 4864 33812 4928
rect 33876 4864 33884 4928
rect 33564 3840 33884 4864
rect 33564 3776 33572 3840
rect 33636 3776 33652 3840
rect 33716 3776 33732 3840
rect 33796 3776 33812 3840
rect 33876 3776 33884 3840
rect 33564 2752 33884 3776
rect 33564 2688 33572 2752
rect 33636 2688 33652 2752
rect 33716 2688 33732 2752
rect 33796 2688 33812 2752
rect 33876 2688 33884 2752
rect 33564 1664 33884 2688
rect 33564 1600 33572 1664
rect 33636 1600 33652 1664
rect 33716 1600 33732 1664
rect 33796 1600 33812 1664
rect 33876 1600 33884 1664
rect 33564 1040 33884 1600
rect 34286 1325 34346 8331
rect 34283 1324 34349 1325
rect 34283 1260 34284 1324
rect 34348 1260 34349 1324
rect 34283 1259 34349 1260
rect 34470 1189 34530 8331
rect 36064 7648 36384 8672
rect 36064 7584 36072 7648
rect 36136 7584 36152 7648
rect 36216 7584 36232 7648
rect 36296 7584 36312 7648
rect 36376 7584 36384 7648
rect 36064 6560 36384 7584
rect 36064 6496 36072 6560
rect 36136 6496 36152 6560
rect 36216 6496 36232 6560
rect 36296 6496 36312 6560
rect 36376 6496 36384 6560
rect 36064 5472 36384 6496
rect 36064 5408 36072 5472
rect 36136 5408 36152 5472
rect 36216 5408 36232 5472
rect 36296 5408 36312 5472
rect 36376 5408 36384 5472
rect 36064 4384 36384 5408
rect 36064 4320 36072 4384
rect 36136 4320 36152 4384
rect 36216 4320 36232 4384
rect 36296 4320 36312 4384
rect 36376 4320 36384 4384
rect 36064 3296 36384 4320
rect 36064 3232 36072 3296
rect 36136 3232 36152 3296
rect 36216 3232 36232 3296
rect 36296 3232 36312 3296
rect 36376 3232 36384 3296
rect 36064 2208 36384 3232
rect 36064 2144 36072 2208
rect 36136 2144 36152 2208
rect 36216 2144 36232 2208
rect 36296 2144 36312 2208
rect 36376 2144 36384 2208
rect 34467 1188 34533 1189
rect 34467 1124 34468 1188
rect 34532 1124 34533 1188
rect 34467 1123 34533 1124
rect 36064 1120 36384 2144
rect 36064 1056 36072 1120
rect 36136 1056 36152 1120
rect 36216 1056 36232 1120
rect 36296 1056 36312 1120
rect 36376 1056 36384 1120
rect 36064 1040 36384 1056
rect 38564 22336 38884 22896
rect 38564 22272 38572 22336
rect 38636 22272 38652 22336
rect 38716 22272 38732 22336
rect 38796 22272 38812 22336
rect 38876 22272 38884 22336
rect 38564 21248 38884 22272
rect 38564 21184 38572 21248
rect 38636 21184 38652 21248
rect 38716 21184 38732 21248
rect 38796 21184 38812 21248
rect 38876 21184 38884 21248
rect 38564 20160 38884 21184
rect 38564 20096 38572 20160
rect 38636 20096 38652 20160
rect 38716 20096 38732 20160
rect 38796 20096 38812 20160
rect 38876 20096 38884 20160
rect 38564 19072 38884 20096
rect 38564 19008 38572 19072
rect 38636 19008 38652 19072
rect 38716 19008 38732 19072
rect 38796 19008 38812 19072
rect 38876 19008 38884 19072
rect 38564 17984 38884 19008
rect 38564 17920 38572 17984
rect 38636 17920 38652 17984
rect 38716 17920 38732 17984
rect 38796 17920 38812 17984
rect 38876 17920 38884 17984
rect 38564 16896 38884 17920
rect 38564 16832 38572 16896
rect 38636 16832 38652 16896
rect 38716 16832 38732 16896
rect 38796 16832 38812 16896
rect 38876 16832 38884 16896
rect 38564 15808 38884 16832
rect 38564 15744 38572 15808
rect 38636 15744 38652 15808
rect 38716 15744 38732 15808
rect 38796 15744 38812 15808
rect 38876 15744 38884 15808
rect 38564 14720 38884 15744
rect 38564 14656 38572 14720
rect 38636 14656 38652 14720
rect 38716 14656 38732 14720
rect 38796 14656 38812 14720
rect 38876 14656 38884 14720
rect 38564 13632 38884 14656
rect 38564 13568 38572 13632
rect 38636 13568 38652 13632
rect 38716 13568 38732 13632
rect 38796 13568 38812 13632
rect 38876 13568 38884 13632
rect 38564 12544 38884 13568
rect 38564 12480 38572 12544
rect 38636 12480 38652 12544
rect 38716 12480 38732 12544
rect 38796 12480 38812 12544
rect 38876 12480 38884 12544
rect 38564 11456 38884 12480
rect 38564 11392 38572 11456
rect 38636 11392 38652 11456
rect 38716 11392 38732 11456
rect 38796 11392 38812 11456
rect 38876 11392 38884 11456
rect 38564 10368 38884 11392
rect 38564 10304 38572 10368
rect 38636 10304 38652 10368
rect 38716 10304 38732 10368
rect 38796 10304 38812 10368
rect 38876 10304 38884 10368
rect 38564 9280 38884 10304
rect 38564 9216 38572 9280
rect 38636 9216 38652 9280
rect 38716 9216 38732 9280
rect 38796 9216 38812 9280
rect 38876 9216 38884 9280
rect 38564 8192 38884 9216
rect 38564 8128 38572 8192
rect 38636 8128 38652 8192
rect 38716 8128 38732 8192
rect 38796 8128 38812 8192
rect 38876 8128 38884 8192
rect 38564 7104 38884 8128
rect 38564 7040 38572 7104
rect 38636 7040 38652 7104
rect 38716 7040 38732 7104
rect 38796 7040 38812 7104
rect 38876 7040 38884 7104
rect 38564 6016 38884 7040
rect 38564 5952 38572 6016
rect 38636 5952 38652 6016
rect 38716 5952 38732 6016
rect 38796 5952 38812 6016
rect 38876 5952 38884 6016
rect 38564 4928 38884 5952
rect 38564 4864 38572 4928
rect 38636 4864 38652 4928
rect 38716 4864 38732 4928
rect 38796 4864 38812 4928
rect 38876 4864 38884 4928
rect 38564 3840 38884 4864
rect 38564 3776 38572 3840
rect 38636 3776 38652 3840
rect 38716 3776 38732 3840
rect 38796 3776 38812 3840
rect 38876 3776 38884 3840
rect 38564 2752 38884 3776
rect 41064 22880 41384 22896
rect 41064 22816 41072 22880
rect 41136 22816 41152 22880
rect 41216 22816 41232 22880
rect 41296 22816 41312 22880
rect 41376 22816 41384 22880
rect 41064 21792 41384 22816
rect 41064 21728 41072 21792
rect 41136 21728 41152 21792
rect 41216 21728 41232 21792
rect 41296 21728 41312 21792
rect 41376 21728 41384 21792
rect 41064 20704 41384 21728
rect 41064 20640 41072 20704
rect 41136 20640 41152 20704
rect 41216 20640 41232 20704
rect 41296 20640 41312 20704
rect 41376 20640 41384 20704
rect 41064 19616 41384 20640
rect 41064 19552 41072 19616
rect 41136 19552 41152 19616
rect 41216 19552 41232 19616
rect 41296 19552 41312 19616
rect 41376 19552 41384 19616
rect 41064 18528 41384 19552
rect 41064 18464 41072 18528
rect 41136 18464 41152 18528
rect 41216 18464 41232 18528
rect 41296 18464 41312 18528
rect 41376 18464 41384 18528
rect 41064 17440 41384 18464
rect 41064 17376 41072 17440
rect 41136 17376 41152 17440
rect 41216 17376 41232 17440
rect 41296 17376 41312 17440
rect 41376 17376 41384 17440
rect 41064 16352 41384 17376
rect 41064 16288 41072 16352
rect 41136 16288 41152 16352
rect 41216 16288 41232 16352
rect 41296 16288 41312 16352
rect 41376 16288 41384 16352
rect 41064 15264 41384 16288
rect 41064 15200 41072 15264
rect 41136 15200 41152 15264
rect 41216 15200 41232 15264
rect 41296 15200 41312 15264
rect 41376 15200 41384 15264
rect 41064 14176 41384 15200
rect 41064 14112 41072 14176
rect 41136 14112 41152 14176
rect 41216 14112 41232 14176
rect 41296 14112 41312 14176
rect 41376 14112 41384 14176
rect 41064 13088 41384 14112
rect 41064 13024 41072 13088
rect 41136 13024 41152 13088
rect 41216 13024 41232 13088
rect 41296 13024 41312 13088
rect 41376 13024 41384 13088
rect 41064 12000 41384 13024
rect 41064 11936 41072 12000
rect 41136 11936 41152 12000
rect 41216 11936 41232 12000
rect 41296 11936 41312 12000
rect 41376 11936 41384 12000
rect 41064 10912 41384 11936
rect 41064 10848 41072 10912
rect 41136 10848 41152 10912
rect 41216 10848 41232 10912
rect 41296 10848 41312 10912
rect 41376 10848 41384 10912
rect 41064 9824 41384 10848
rect 41064 9760 41072 9824
rect 41136 9760 41152 9824
rect 41216 9760 41232 9824
rect 41296 9760 41312 9824
rect 41376 9760 41384 9824
rect 41064 8736 41384 9760
rect 41064 8672 41072 8736
rect 41136 8672 41152 8736
rect 41216 8672 41232 8736
rect 41296 8672 41312 8736
rect 41376 8672 41384 8736
rect 41064 7648 41384 8672
rect 41064 7584 41072 7648
rect 41136 7584 41152 7648
rect 41216 7584 41232 7648
rect 41296 7584 41312 7648
rect 41376 7584 41384 7648
rect 41064 6560 41384 7584
rect 41064 6496 41072 6560
rect 41136 6496 41152 6560
rect 41216 6496 41232 6560
rect 41296 6496 41312 6560
rect 41376 6496 41384 6560
rect 41064 5472 41384 6496
rect 41064 5408 41072 5472
rect 41136 5408 41152 5472
rect 41216 5408 41232 5472
rect 41296 5408 41312 5472
rect 41376 5408 41384 5472
rect 41064 4384 41384 5408
rect 41064 4320 41072 4384
rect 41136 4320 41152 4384
rect 41216 4320 41232 4384
rect 41296 4320 41312 4384
rect 41376 4320 41384 4384
rect 41064 3296 41384 4320
rect 41064 3232 41072 3296
rect 41136 3232 41152 3296
rect 41216 3232 41232 3296
rect 41296 3232 41312 3296
rect 41376 3232 41384 3296
rect 39987 3228 40053 3229
rect 39987 3164 39988 3228
rect 40052 3164 40053 3228
rect 39987 3163 40053 3164
rect 38564 2688 38572 2752
rect 38636 2688 38652 2752
rect 38716 2688 38732 2752
rect 38796 2688 38812 2752
rect 38876 2688 38884 2752
rect 38564 1664 38884 2688
rect 38564 1600 38572 1664
rect 38636 1600 38652 1664
rect 38716 1600 38732 1664
rect 38796 1600 38812 1664
rect 38876 1600 38884 1664
rect 38564 1040 38884 1600
rect 39990 1325 40050 3163
rect 41064 2208 41384 3232
rect 41064 2144 41072 2208
rect 41136 2144 41152 2208
rect 41216 2144 41232 2208
rect 41296 2144 41312 2208
rect 41376 2144 41384 2208
rect 39987 1324 40053 1325
rect 39987 1260 39988 1324
rect 40052 1260 40053 1324
rect 39987 1259 40053 1260
rect 41064 1120 41384 2144
rect 41064 1056 41072 1120
rect 41136 1056 41152 1120
rect 41216 1056 41232 1120
rect 41296 1056 41312 1120
rect 41376 1056 41384 1120
rect 41064 1040 41384 1056
rect 43564 22336 43884 22896
rect 43564 22272 43572 22336
rect 43636 22272 43652 22336
rect 43716 22272 43732 22336
rect 43796 22272 43812 22336
rect 43876 22272 43884 22336
rect 43564 21248 43884 22272
rect 43564 21184 43572 21248
rect 43636 21184 43652 21248
rect 43716 21184 43732 21248
rect 43796 21184 43812 21248
rect 43876 21184 43884 21248
rect 43564 20160 43884 21184
rect 43564 20096 43572 20160
rect 43636 20096 43652 20160
rect 43716 20096 43732 20160
rect 43796 20096 43812 20160
rect 43876 20096 43884 20160
rect 43564 19072 43884 20096
rect 43564 19008 43572 19072
rect 43636 19008 43652 19072
rect 43716 19008 43732 19072
rect 43796 19008 43812 19072
rect 43876 19008 43884 19072
rect 43564 17984 43884 19008
rect 43564 17920 43572 17984
rect 43636 17920 43652 17984
rect 43716 17920 43732 17984
rect 43796 17920 43812 17984
rect 43876 17920 43884 17984
rect 43564 16896 43884 17920
rect 43564 16832 43572 16896
rect 43636 16832 43652 16896
rect 43716 16832 43732 16896
rect 43796 16832 43812 16896
rect 43876 16832 43884 16896
rect 43564 15808 43884 16832
rect 43564 15744 43572 15808
rect 43636 15744 43652 15808
rect 43716 15744 43732 15808
rect 43796 15744 43812 15808
rect 43876 15744 43884 15808
rect 43564 14720 43884 15744
rect 43564 14656 43572 14720
rect 43636 14656 43652 14720
rect 43716 14656 43732 14720
rect 43796 14656 43812 14720
rect 43876 14656 43884 14720
rect 43564 13632 43884 14656
rect 43564 13568 43572 13632
rect 43636 13568 43652 13632
rect 43716 13568 43732 13632
rect 43796 13568 43812 13632
rect 43876 13568 43884 13632
rect 43564 12544 43884 13568
rect 43564 12480 43572 12544
rect 43636 12480 43652 12544
rect 43716 12480 43732 12544
rect 43796 12480 43812 12544
rect 43876 12480 43884 12544
rect 43564 11456 43884 12480
rect 43564 11392 43572 11456
rect 43636 11392 43652 11456
rect 43716 11392 43732 11456
rect 43796 11392 43812 11456
rect 43876 11392 43884 11456
rect 43564 10368 43884 11392
rect 43564 10304 43572 10368
rect 43636 10304 43652 10368
rect 43716 10304 43732 10368
rect 43796 10304 43812 10368
rect 43876 10304 43884 10368
rect 43564 9280 43884 10304
rect 43564 9216 43572 9280
rect 43636 9216 43652 9280
rect 43716 9216 43732 9280
rect 43796 9216 43812 9280
rect 43876 9216 43884 9280
rect 43564 8192 43884 9216
rect 43564 8128 43572 8192
rect 43636 8128 43652 8192
rect 43716 8128 43732 8192
rect 43796 8128 43812 8192
rect 43876 8128 43884 8192
rect 43564 7104 43884 8128
rect 43564 7040 43572 7104
rect 43636 7040 43652 7104
rect 43716 7040 43732 7104
rect 43796 7040 43812 7104
rect 43876 7040 43884 7104
rect 43564 6016 43884 7040
rect 43564 5952 43572 6016
rect 43636 5952 43652 6016
rect 43716 5952 43732 6016
rect 43796 5952 43812 6016
rect 43876 5952 43884 6016
rect 43564 4928 43884 5952
rect 43564 4864 43572 4928
rect 43636 4864 43652 4928
rect 43716 4864 43732 4928
rect 43796 4864 43812 4928
rect 43876 4864 43884 4928
rect 43564 3840 43884 4864
rect 43564 3776 43572 3840
rect 43636 3776 43652 3840
rect 43716 3776 43732 3840
rect 43796 3776 43812 3840
rect 43876 3776 43884 3840
rect 43564 2752 43884 3776
rect 43564 2688 43572 2752
rect 43636 2688 43652 2752
rect 43716 2688 43732 2752
rect 43796 2688 43812 2752
rect 43876 2688 43884 2752
rect 43564 1664 43884 2688
rect 43564 1600 43572 1664
rect 43636 1600 43652 1664
rect 43716 1600 43732 1664
rect 43796 1600 43812 1664
rect 43876 1600 43884 1664
rect 43564 1040 43884 1600
use sky130_fd_sc_hd__clkbuf_4  _073_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _074_
timestamp 1688980957
transform 1 0 27968 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _075_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _077_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _079_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 1688980957
transform 1 0 27968 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _081_
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 1688980957
transform 1 0 32568 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _084_
timestamp 1688980957
transform 1 0 28704 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1688980957
transform 1 0 28152 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp 1688980957
transform 1 0 34040 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _087_
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1688980957
transform 1 0 28428 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp 1688980957
transform 1 0 34500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1688980957
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1688980957
transform 1 0 28888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 1688980957
transform 1 0 35144 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1688980957
transform 1 0 28704 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp 1688980957
transform 1 0 36616 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 1688980957
transform 1 0 30360 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1688980957
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1688980957
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 1688980957
transform 1 0 39192 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1688980957
transform 1 0 30912 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _104_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41768 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp 1688980957
transform 1 0 38732 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _106_
timestamp 1688980957
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1688980957
transform 1 0 32936 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1688980957
transform 1 0 34040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp 1688980957
transform 1 0 40296 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1688980957
transform 1 0 32568 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1688980957
transform 1 0 41860 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _113_
timestamp 1688980957
transform 1 0 31464 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1688980957
transform 1 0 31464 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _115_
timestamp 1688980957
transform 1 0 42596 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1688980957
transform 1 0 32660 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1688980957
transform 1 0 32292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1688980957
transform 1 0 42504 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _119_
timestamp 1688980957
transform 1 0 31832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _121_
timestamp 1688980957
transform 1 0 42872 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1688980957
transform 1 0 33488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1688980957
transform 1 0 42136 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 1688980957
transform 1 0 31832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1688980957
transform 1 0 31464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 1688980957
transform 1 0 32936 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1688980957
transform 1 0 32108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1688980957
transform 1 0 34040 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _131_
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 1688980957
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1688980957
transform 1 0 31280 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1688980957
transform 1 0 30176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _136_
timestamp 1688980957
transform 1 0 37536 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _138_
timestamp 1688980957
transform 1 0 33488 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 1688980957
transform 1 0 28520 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1688980957
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _141_
timestamp 1688980957
transform 1 0 35880 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1688980957
transform 1 0 29072 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _144_
timestamp 1688980957
transform 1 0 35880 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1688980957
transform 1 0 29900 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1688980957
transform 1 0 28704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 1688980957
transform 1 0 35696 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _148_
timestamp 1688980957
transform 1 0 30084 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1688980957
transform 1 0 29716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _150_
timestamp 1688980957
transform 1 0 37628 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp 1688980957
transform 1 0 30912 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1688980957
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _153_
timestamp 1688980957
transform 1 0 40848 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 1688980957
transform 1 0 32384 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1688980957
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp 1688980957
transform 1 0 40296 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1688980957
transform 1 0 33304 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1688980957
transform 1 0 33672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp 1688980957
transform 1 0 40756 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1688980957
transform 1 0 32844 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _161_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1688980957
transform 1 0 40388 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _163_
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp 1688980957
transform 1 0 25944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp 1688980957
transform 1 0 38088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1688980957
transform 1 0 32660 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 1688980957
transform 1 0 42872 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp 1688980957
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _171_
timestamp 1688980957
transform 1 0 42596 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _173_
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1688980957
transform 1 0 42320 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _175_
timestamp 1688980957
transform 1 0 33672 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _176_
timestamp 1688980957
transform 1 0 34040 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _177_
timestamp 1688980957
transform 1 0 15824 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1688980957
transform 1 0 26128 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _180_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _181_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1688980957
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1688980957
transform 1 0 2760 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1688980957
transform 1 0 3864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1688980957
transform 1 0 6440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1688980957
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _189_
timestamp 1688980957
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _191_
timestamp 1688980957
transform 1 0 10120 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1688980957
transform 1 0 12788 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1688980957
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1688980957
transform 1 0 17204 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1688980957
transform 1 0 19688 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1688980957
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1688980957
transform 1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1688980957
transform 1 0 22724 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1688980957
transform 1 0 24932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1688980957
transform 1 0 25392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1688980957
transform 1 0 27048 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1688980957
transform 1 0 25944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 1688980957
transform 1 0 32844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1688980957
transform 1 0 29992 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1688980957
transform 1 0 5152 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1688980957
transform 1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1688980957
transform 1 0 11132 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1688980957
transform 1 0 11960 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1688980957
transform 1 0 12236 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1688980957
transform 1 0 16192 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1688980957
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _233__113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _233_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1688980957
transform 1 0 18676 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _235_
timestamp 1688980957
transform 1 0 19688 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1688980957
transform 1 0 20792 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1688980957
transform 1 0 21528 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1688980957
transform 1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1688980957
transform 1 0 25852 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1688980957
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1688980957
transform 1 0 31096 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1688980957
transform 1 0 33672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1688980957
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1688980957
transform 1 0 35604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1688980957
transform 1 0 38732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1688980957
transform 1 0 44068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__S
timestamp 1688980957
transform 1 0 44528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1688980957
transform 1 0 44528 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__S
timestamp 1688980957
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__S
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__S
timestamp 1688980957
transform 1 0 6532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__S
timestamp 1688980957
transform 1 0 6624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__S
timestamp 1688980957
transform 1 0 44528 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__S
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__S
timestamp 1688980957
transform 1 0 43240 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__S
timestamp 1688980957
transform 1 0 44068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__S
timestamp 1688980957
transform 1 0 44528 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1688980957
transform 1 0 44160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1688980957
transform 1 0 44712 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__S
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__S
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__S
timestamp 1688980957
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__S
timestamp 1688980957
transform 1 0 44988 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__S
timestamp 1688980957
transform 1 0 8372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__S
timestamp 1688980957
transform 1 0 44068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__S
timestamp 1688980957
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__S
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1688980957
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1688980957
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1688980957
transform 1 0 4324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1688980957
transform 1 0 5060 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1688980957
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1688980957
transform 1 0 6256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1688980957
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1688980957
transform 1 0 9936 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1688980957
transform 1 0 10672 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1688980957
transform 1 0 11592 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1688980957
transform 1 0 12144 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1688980957
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1688980957
transform 1 0 12604 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1688980957
transform 1 0 12696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1688980957
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1688980957
transform 1 0 13616 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1688980957
transform 1 0 40940 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1688980957
transform 1 0 43148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1688980957
transform 1 0 43792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._121__A
timestamp 1688980957
transform 1 0 41400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._121__C
timestamp 1688980957
transform 1 0 41952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._122__A
timestamp 1688980957
transform 1 0 42504 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._124__A
timestamp 1688980957
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._124__B
timestamp 1688980957
transform 1 0 37720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._124__C_N
timestamp 1688980957
transform 1 0 37536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._124__D_N
timestamp 1688980957
transform 1 0 12788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._125__A
timestamp 1688980957
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._125__B
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._125__C
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._125__D_N
timestamp 1688980957
transform 1 0 34224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._126__A
timestamp 1688980957
transform 1 0 37904 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._126__B
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._126__D_N
timestamp 1688980957
transform 1 0 38640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._127__B
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._127__C
timestamp 1688980957
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._127__D
timestamp 1688980957
transform 1 0 36156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._129__A
timestamp 1688980957
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._129__B
timestamp 1688980957
transform 1 0 20884 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._129__C_N
timestamp 1688980957
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._129__D_N
timestamp 1688980957
transform 1 0 19136 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._130__A
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._130__B
timestamp 1688980957
transform 1 0 33672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._130__C_N
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._130__D_N
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._131__A
timestamp 1688980957
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._131__B
timestamp 1688980957
transform 1 0 19964 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._131__C_N
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._131__D_N
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._132__A
timestamp 1688980957
transform 1 0 23460 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._132__B
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._132__C
timestamp 1688980957
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._132__D
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._141__A
timestamp 1688980957
transform 1 0 41952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._143__B1
timestamp 1688980957
transform 1 0 41400 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._181__A0
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._181__S
timestamp 1688980957
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._183__A0
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._183__S
timestamp 1688980957
transform 1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._185__A0
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._185__S
timestamp 1688980957
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._187__A0
timestamp 1688980957
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._187__S
timestamp 1688980957
transform 1 0 1288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._189__A0
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._189__S
timestamp 1688980957
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._191__A0
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._191__S
timestamp 1688980957
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._193__A0
timestamp 1688980957
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._193__S
timestamp 1688980957
transform 1 0 6900 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._195__A0
timestamp 1688980957
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._195__S
timestamp 1688980957
transform 1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._197__A0
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._197__S
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._200__A0
timestamp 1688980957
transform 1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._202__A0
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._204__A0
timestamp 1688980957
transform 1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._206__A0
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._208__A0
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._210__A0
timestamp 1688980957
transform 1 0 10580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._212__A0
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._214__A0
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._216__A0
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._218__A0
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._221__A0
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._223__A0
timestamp 1688980957
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._225__A0
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._227__A0
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._229__A0
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._231__A0
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._233__A0
timestamp 1688980957
transform 1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._237__A0
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._241__A0
timestamp 1688980957
transform 1 0 14168 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._243__A0
timestamp 1688980957
transform 1 0 41216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._245__CLK
timestamp 1688980957
transform 1 0 42964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._245__RESET_B
timestamp 1688980957
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._246__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._246__RESET_B
timestamp 1688980957
transform 1 0 43792 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._247__CLK
timestamp 1688980957
transform 1 0 42688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._247__RESET_B
timestamp 1688980957
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._248__CLK
timestamp 1688980957
transform 1 0 41584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._248__RESET_B
timestamp 1688980957
transform 1 0 41952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._249__CLK
timestamp 1688980957
transform 1 0 43056 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._249__RESET_B
timestamp 1688980957
transform 1 0 42596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._250__CLK
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._250__SET_B
timestamp 1688980957
transform 1 0 42688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._251__CLK
timestamp 1688980957
transform 1 0 41952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._251__RESET_B
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._252__CLK
timestamp 1688980957
transform 1 0 41768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._252__RESET_B
timestamp 1688980957
transform 1 0 42136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._253__CLK
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._253__RESET_B
timestamp 1688980957
transform 1 0 42688 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._254__CLK
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._254__RESET_B
timestamp 1688980957
transform 1 0 42964 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._255__CLK
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._255__RESET_B
timestamp 1688980957
transform 1 0 1012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._256__CLK
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._256__RESET_B
timestamp 1688980957
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._257__CLK
timestamp 1688980957
transform 1 0 1472 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._257__RESET_B
timestamp 1688980957
transform 1 0 1012 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._258__CLK
timestamp 1688980957
transform 1 0 1012 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._258__RESET_B
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._259__CLK
timestamp 1688980957
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._259__RESET_B
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._260__CLK
timestamp 1688980957
transform 1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._260__RESET_B
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._261__CLK
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._261__RESET_B
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._262__CLK
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._262__RESET_B
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._263__CLK
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._263__RESET_B
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._264__CLK
timestamp 1688980957
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._264__RESET_B
timestamp 1688980957
transform 1 0 7636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._265__CLK
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._265__RESET_B
timestamp 1688980957
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._266__CLK
timestamp 1688980957
transform 1 0 8004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._266__RESET_B
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._267__CLK
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._267__RESET_B
timestamp 1688980957
transform 1 0 6440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._268__CLK
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._268__RESET_B
timestamp 1688980957
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._269__CLK
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._269__RESET_B
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._270__CLK
timestamp 1688980957
transform 1 0 6808 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._270__RESET_B
timestamp 1688980957
transform 1 0 7176 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._271__CLK
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._271__RESET_B
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._272__CLK
timestamp 1688980957
transform 1 0 8372 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._272__RESET_B
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._273__CLK
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._273__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._274__CLK
timestamp 1688980957
transform 1 0 8740 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._274__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._275__CLK
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._275__RESET_B
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._276__CLK
timestamp 1688980957
transform 1 0 10120 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._276__RESET_B
timestamp 1688980957
transform 1 0 11776 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._277__CLK
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._277__RESET_B
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._278__CLK
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._278__RESET_B
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._279__CLK
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._279__RESET_B
timestamp 1688980957
transform 1 0 17572 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._280__CLK
timestamp 1688980957
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._280__RESET_B
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._281__CLK
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._281__RESET_B
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._282__CLK
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._282__RESET_B
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._283__CLK
timestamp 1688980957
transform 1 0 12512 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._283__RESET_B
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._284__CLK
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._284__RESET_B
timestamp 1688980957
transform 1 0 41308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._285__CLK
timestamp 1688980957
transform 1 0 42228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._285__RESET_B
timestamp 1688980957
transform 1 0 41952 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._286__CLK
timestamp 1688980957
transform 1 0 11684 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._286__RESET_B
timestamp 1688980957
transform 1 0 41860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._287__CLK
timestamp 1688980957
transform 1 0 41400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ConfigFSM_inst._287__RESET_B
timestamp 1688980957
transform 1 0 41032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._186__A
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._187__A
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._191__A
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._193__A
timestamp 1688980957
transform 1 0 10672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._194__S
timestamp 1688980957
transform 1 0 35604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._196__S
timestamp 1688980957
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._198__S
timestamp 1688980957
transform 1 0 41952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._200__S
timestamp 1688980957
transform 1 0 42044 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._202__S
timestamp 1688980957
transform 1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._204__S
timestamp 1688980957
transform 1 0 44712 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._206__S
timestamp 1688980957
transform 1 0 43240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._208__S
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._210__A
timestamp 1688980957
transform 1 0 44528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._231__A
timestamp 1688980957
transform 1 0 43056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._252__S
timestamp 1688980957
transform 1 0 44896 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._254__S
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._256__S
timestamp 1688980957
transform 1 0 9476 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._258__S
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._261__A
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._282__A
timestamp 1688980957
transform 1 0 44896 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._303__A
timestamp 1688980957
transform 1 0 44528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._324__S
timestamp 1688980957
transform 1 0 44804 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._326__S
timestamp 1688980957
transform 1 0 43792 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._362__CLK
timestamp 1688980957
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._362__RESET_B
timestamp 1688980957
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._363__CLK
timestamp 1688980957
transform 1 0 14168 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._363__RESET_B
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._364__CLK
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._364__RESET_B
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._365__CLK
timestamp 1688980957
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._365__RESET_B
timestamp 1688980957
transform 1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._366__CLK
timestamp 1688980957
transform 1 0 17296 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._366__RESET_B
timestamp 1688980957
transform 1 0 36156 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._367__CLK
timestamp 1688980957
transform 1 0 41308 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._367__RESET_B
timestamp 1688980957
transform 1 0 41952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._368__CLK
timestamp 1688980957
transform 1 0 42412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._368__RESET_B
timestamp 1688980957
transform 1 0 42780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._369__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._369__RESET_B
timestamp 1688980957
transform 1 0 43516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._370__CLK
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._370__RESET_B
timestamp 1688980957
transform 1 0 44804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._371__CLK
timestamp 1688980957
transform 1 0 44896 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._371__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._372__CLK
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._372__RESET_B
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._373__CLK
timestamp 1688980957
transform 1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._373__RESET_B
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._374__CLK
timestamp 1688980957
transform 1 0 8004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._374__RESET_B
timestamp 1688980957
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._375__CLK
timestamp 1688980957
transform 1 0 44528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._375__RESET_B
timestamp 1688980957
transform 1 0 43700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._376__CLK
timestamp 1688980957
transform 1 0 6164 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._376__RESET_B
timestamp 1688980957
transform 1 0 5796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._377__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._377__RESET_B
timestamp 1688980957
transform 1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._378__CLK
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._378__RESET_B
timestamp 1688980957
transform 1 0 4692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._379__CLK
timestamp 1688980957
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._379__RESET_B
timestamp 1688980957
transform 1 0 6164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._380__CLK
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._380__RESET_B
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._381__CLK
timestamp 1688980957
transform 1 0 44528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._381__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._382__CLK
timestamp 1688980957
transform 1 0 44528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._382__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._383__CLK
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._383__RESET_B
timestamp 1688980957
transform 1 0 44804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._384__CLK
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._384__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._385__CLK
timestamp 1688980957
transform 1 0 45080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._385__RESET_B
timestamp 1688980957
transform 1 0 43608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._386__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._386__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._387__CLK
timestamp 1688980957
transform 1 0 44896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._387__RESET_B
timestamp 1688980957
transform 1 0 43792 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._388__CLK
timestamp 1688980957
transform 1 0 4968 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._388__RESET_B
timestamp 1688980957
transform 1 0 4232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._389__CLK
timestamp 1688980957
transform 1 0 3128 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._389__RESET_B
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._390__CLK
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._390__RESET_B
timestamp 1688980957
transform 1 0 1564 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._391__CLK
timestamp 1688980957
transform 1 0 1196 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._391__RESET_B
timestamp 1688980957
transform 1 0 1012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._392__CLK
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._392__RESET_B
timestamp 1688980957
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._393__CLK
timestamp 1688980957
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._393__RESET_B
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._394__CLK
timestamp 1688980957
transform 1 0 44896 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._394__RESET_B
timestamp 1688980957
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._395__CLK
timestamp 1688980957
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._395__RESET_B
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._396__CLK
timestamp 1688980957
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._396__RESET_B
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._397__CLK
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._397__RESET_B
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._398__CLK
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._398__RESET_B
timestamp 1688980957
transform 1 0 22816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._399__CLK
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._399__RESET_B
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._400__CLK
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._400__RESET_B
timestamp 1688980957
transform 1 0 41308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._401__CLK
timestamp 1688980957
transform 1 0 42688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._401__RESET_B
timestamp 1688980957
transform 1 0 43056 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._402__CLK
timestamp 1688980957
transform 1 0 43608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._402__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._403__CLK
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._403__RESET_B
timestamp 1688980957
transform 1 0 45080 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._404__CLK
timestamp 1688980957
transform 1 0 43976 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._404__RESET_B
timestamp 1688980957
transform 1 0 44160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._405__CLK
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._405__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._406__CLK
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._406__RESET_B
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._407__CLK
timestamp 1688980957
transform 1 0 44896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._407__RESET_B
timestamp 1688980957
transform 1 0 44528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._408__CLK
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._408__RESET_B
timestamp 1688980957
transform 1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._409__CLK
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._409__RESET_B
timestamp 1688980957
transform 1 0 7268 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._410__CLK
timestamp 1688980957
transform 1 0 5428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._410__RESET_B
timestamp 1688980957
transform 1 0 5060 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._411__CLK
timestamp 1688980957
transform 1 0 6900 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._411__RESET_B
timestamp 1688980957
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._412__CLK
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._412__RESET_B
timestamp 1688980957
transform 1 0 3956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._413__CLK
timestamp 1688980957
transform 1 0 44528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._413__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._414__CLK
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._414__RESET_B
timestamp 1688980957
transform 1 0 44160 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._415__CLK
timestamp 1688980957
transform 1 0 43056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._415__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._416__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._416__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._417__CLK
timestamp 1688980957
transform 1 0 44528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._417__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._418__CLK
timestamp 1688980957
transform 1 0 43056 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._418__RESET_B
timestamp 1688980957
transform 1 0 43424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._419__CLK
timestamp 1688980957
transform 1 0 42688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._419__RESET_B
timestamp 1688980957
transform 1 0 44160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._420__CLK
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._420__RESET_B
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._421__CLK
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._421__RESET_B
timestamp 1688980957
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._422__CLK
timestamp 1688980957
transform 1 0 5060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._422__RESET_B
timestamp 1688980957
transform 1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._423__CLK
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._423__RESET_B
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._424__CLK
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._424__RESET_B
timestamp 1688980957
transform 1 0 6256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._425__CLK
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._425__RESET_B
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._426__CLK
timestamp 1688980957
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._426__RESET_B
timestamp 1688980957
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._427__CLK
timestamp 1688980957
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._427__RESET_B
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._428__CLK
timestamp 1688980957
transform 1 0 8004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._428__RESET_B
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._429__CLK
timestamp 1688980957
transform 1 0 920 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._429__RESET_B
timestamp 1688980957
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._430__CLK
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._430__RESET_B
timestamp 1688980957
transform 1 0 3864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._431__CLK
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._431__RESET_B
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._432__CLK
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._432__RESET_B
timestamp 1688980957
transform 1 0 8372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._433__CLK
timestamp 1688980957
transform 1 0 9292 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._433__RESET_B
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._434__CLK
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._434__RESET_B
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._435__CLK
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._435__RESET_B
timestamp 1688980957
transform 1 0 4692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._436__CLK
timestamp 1688980957
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._436__RESET_B
timestamp 1688980957
transform 1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._437__CLK
timestamp 1688980957
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._437__RESET_B
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._438__CLK
timestamp 1688980957
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._438__RESET_B
timestamp 1688980957
transform 1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._439__CLK
timestamp 1688980957
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._439__RESET_B
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._440__CLK
timestamp 1688980957
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._440__RESET_B
timestamp 1688980957
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._441__CLK
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._441__RESET_B
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._442__CLK
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._442__RESET_B
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._443__CLK
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._443__RESET_B
timestamp 1688980957
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._444__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._444__RESET_B
timestamp 1688980957
transform 1 0 6992 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._445__CLK
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._445__RESET_B
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._446__CLK
timestamp 1688980957
transform 1 0 6440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._446__RESET_B
timestamp 1688980957
transform 1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._447__CLK
timestamp 1688980957
transform 1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._447__RESET_B
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._448__CLK
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._448__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._449__CLK
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._449__RESET_B
timestamp 1688980957
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._450__CLK
timestamp 1688980957
transform 1 0 9016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._450__RESET_B
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._451__CLK
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._451__RESET_B
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._452__CLK
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._452__RESET_B
timestamp 1688980957
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._453__CLK
timestamp 1688980957
transform 1 0 9384 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Inst_bitbang._453__RESET_B
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0597__A_N
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0612__A
timestamp 1688980957
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0623__B
timestamp 1688980957
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0623__C_N
timestamp 1688980957
transform 1 0 28336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0623__D_N
timestamp 1688980957
transform 1 0 25300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0624__A
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0629__A
timestamp 1688980957
transform 1 0 25852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0629__C_N
timestamp 1688980957
transform 1 0 26496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0632__B
timestamp 1688980957
transform 1 0 25300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0633__B_N
timestamp 1688980957
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0636__A1
timestamp 1688980957
transform 1 0 26496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0636__A2
timestamp 1688980957
transform 1 0 26404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0655__B1
timestamp 1688980957
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0656__A
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0662__A
timestamp 1688980957
transform 1 0 30636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0759__A1
timestamp 1688980957
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0763__A0
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0763__A1
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0829__A1
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0829__B2
timestamp 1688980957
transform 1 0 26772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0833__A1
timestamp 1688980957
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0840__A1
timestamp 1688980957
transform 1 0 43608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0842__A1
timestamp 1688980957
transform 1 0 43516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0844__A1
timestamp 1688980957
transform 1 0 43240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0846__A1
timestamp 1688980957
transform 1 0 43700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0848__A1
timestamp 1688980957
transform 1 0 42504 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0855__A1
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0855__B2
timestamp 1688980957
transform 1 0 24656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0859__A1
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0859__B2
timestamp 1688980957
transform 1 0 26036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0863__A1
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0870__A1
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0872__A1
timestamp 1688980957
transform 1 0 43424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0874__A1
timestamp 1688980957
transform 1 0 44988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0876__A1
timestamp 1688980957
transform 1 0 43792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0878__A1
timestamp 1688980957
transform 1 0 42780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0892__B1
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0911__S
timestamp 1688980957
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0976__A
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0978__A1
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0978__B2
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._0999__B1
timestamp 1688980957
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1013__A0
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1018__A0
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1027__A0
timestamp 1688980957
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1034__A0
timestamp 1688980957
transform 1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1040__A0
timestamp 1688980957
transform 1 0 23460 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1107__A1
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1107__B2
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1114__A1
timestamp 1688980957
transform 1 0 44528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1116__A1
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1118__A1
timestamp 1688980957
transform 1 0 44528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1120__A1
timestamp 1688980957
transform 1 0 44160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1122__A1
timestamp 1688980957
transform 1 0 44528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1132__A1
timestamp 1688980957
transform 1 0 41952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1134__A1
timestamp 1688980957
transform 1 0 42136 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1136__A1
timestamp 1688980957
transform 1 0 41308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1138__A1
timestamp 1688980957
transform 1 0 41216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1140__A1
timestamp 1688980957
transform 1 0 42688 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1144__A
timestamp 1688980957
transform 1 0 30084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1144__B
timestamp 1688980957
transform 1 0 32568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1150__A1
timestamp 1688980957
transform 1 0 33304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1152__A1
timestamp 1688980957
transform 1 0 31832 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1154__A1
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1156__A1
timestamp 1688980957
transform 1 0 33672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1158__A1
timestamp 1688980957
transform 1 0 36708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1178__CLK
timestamp 1688980957
transform 1 0 40204 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1178__RESET_B
timestamp 1688980957
transform 1 0 39376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1179__CLK
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1179__SET_B
timestamp 1688980957
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1180__CLK
timestamp 1688980957
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1180__RESET_B
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1181__CLK
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1181__RESET_B
timestamp 1688980957
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1182__CLK
timestamp 1688980957
transform 1 0 32384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1182__RESET_B
timestamp 1688980957
transform 1 0 31832 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1183__CLK
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1183__RESET_B
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1184__CLK
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1184__RESET_B
timestamp 1688980957
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1185__CLK
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1185__RESET_B
timestamp 1688980957
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1186__CLK
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1186__RESET_B
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1187__CLK
timestamp 1688980957
transform 1 0 38824 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1187__RESET_B
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1188__CLK
timestamp 1688980957
transform 1 0 40020 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1188__RESET_B
timestamp 1688980957
transform 1 0 40572 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1189__CLK
timestamp 1688980957
transform 1 0 43056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1189__RESET_B
timestamp 1688980957
transform 1 0 42872 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1190__CLK
timestamp 1688980957
transform 1 0 41676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1190__RESET_B
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1191__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1191__RESET_B
timestamp 1688980957
transform 1 0 43608 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1192__CLK
timestamp 1688980957
transform 1 0 43516 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1192__RESET_B
timestamp 1688980957
transform 1 0 42780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1193__CLK
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1193__RESET_B
timestamp 1688980957
transform 1 0 43792 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1194__CLK
timestamp 1688980957
transform 1 0 41216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1194__RESET_B
timestamp 1688980957
transform 1 0 43792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1195__CLK
timestamp 1688980957
transform 1 0 42504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1195__RESET_B
timestamp 1688980957
transform 1 0 42228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1196__CLK
timestamp 1688980957
transform 1 0 42596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1196__RESET_B
timestamp 1688980957
transform 1 0 42964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1197__CLK
timestamp 1688980957
transform 1 0 42872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1197__RESET_B
timestamp 1688980957
transform 1 0 43700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1198__CLK
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1198__RESET_B
timestamp 1688980957
transform 1 0 43884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1199__CLK
timestamp 1688980957
transform 1 0 43884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1199__RESET_B
timestamp 1688980957
transform 1 0 43608 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1200__CLK
timestamp 1688980957
transform 1 0 43056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1200__RESET_B
timestamp 1688980957
transform 1 0 43424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1201__CLK
timestamp 1688980957
transform 1 0 43976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1201__RESET_B
timestamp 1688980957
transform 1 0 44344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1202__CLK
timestamp 1688980957
transform 1 0 43056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1202__RESET_B
timestamp 1688980957
transform 1 0 43792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1203__CLK
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1203__RESET_B
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1204__CLK
timestamp 1688980957
transform 1 0 44160 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1204__RESET_B
timestamp 1688980957
transform 1 0 44528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1205__CLK
timestamp 1688980957
transform 1 0 43976 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1205__RESET_B
timestamp 1688980957
transform 1 0 44344 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1206__CLK
timestamp 1688980957
transform 1 0 43516 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1206__RESET_B
timestamp 1688980957
transform 1 0 43884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1207__CLK
timestamp 1688980957
transform 1 0 43884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1207__RESET_B
timestamp 1688980957
transform 1 0 43884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1208__CLK
timestamp 1688980957
transform 1 0 43148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1208__RESET_B
timestamp 1688980957
transform 1 0 43884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1209__CLK
timestamp 1688980957
transform 1 0 44160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1209__RESET_B
timestamp 1688980957
transform 1 0 44528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1210__CLK
timestamp 1688980957
transform 1 0 43424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1210__RESET_B
timestamp 1688980957
transform 1 0 43792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1211__CLK
timestamp 1688980957
transform 1 0 40756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1211__SET_B
timestamp 1688980957
transform 1 0 42504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1212__CLK
timestamp 1688980957
transform 1 0 41032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1212__RESET_B
timestamp 1688980957
transform 1 0 41400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1213__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1213__RESET_B
timestamp 1688980957
transform 1 0 43332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1214__CLK
timestamp 1688980957
transform 1 0 40572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1214__RESET_B
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1215__CLK
timestamp 1688980957
transform 1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1215__RESET_B
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1216__CLK
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1216__SET_B
timestamp 1688980957
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1217__CLK
timestamp 1688980957
transform 1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1217__RESET_B
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1218__CLK
timestamp 1688980957
transform 1 0 20700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1218__RESET_B
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1219__CLK
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1219__RESET_B
timestamp 1688980957
transform 1 0 43884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1220__CLK
timestamp 1688980957
transform 1 0 42688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1220__RESET_B
timestamp 1688980957
transform 1 0 43056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1221__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1221__RESET_B
timestamp 1688980957
transform 1 0 43976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1222__CLK
timestamp 1688980957
transform 1 0 43976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1222__RESET_B
timestamp 1688980957
transform 1 0 43424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1223__CLK
timestamp 1688980957
transform 1 0 44068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1223__RESET_B
timestamp 1688980957
transform 1 0 44436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1224__CLK
timestamp 1688980957
transform 1 0 44528 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1224__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1225__CLK
timestamp 1688980957
transform 1 0 42872 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1225__RESET_B
timestamp 1688980957
transform 1 0 42688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1226__CLK
timestamp 1688980957
transform 1 0 43608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1226__RESET_B
timestamp 1688980957
transform 1 0 43976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1227__CLK
timestamp 1688980957
transform 1 0 25576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1227__RESET_B
timestamp 1688980957
transform 1 0 25024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1228__CLK
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1228__RESET_B
timestamp 1688980957
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1229__CLK
timestamp 1688980957
transform 1 0 25576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1229__RESET_B
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1230__CLK
timestamp 1688980957
transform 1 0 43516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1230__RESET_B
timestamp 1688980957
transform 1 0 44896 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1231__CLK
timestamp 1688980957
transform 1 0 43056 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1231__RESET_B
timestamp 1688980957
transform 1 0 43792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1232__CLK
timestamp 1688980957
transform 1 0 43148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1232__RESET_B
timestamp 1688980957
transform 1 0 43516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1233__CLK
timestamp 1688980957
transform 1 0 43424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1233__RESET_B
timestamp 1688980957
transform 1 0 43792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1234__CLK
timestamp 1688980957
transform 1 0 44528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1234__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1235__CLK
timestamp 1688980957
transform 1 0 44252 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1235__RESET_B
timestamp 1688980957
transform 1 0 44620 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1236__CLK
timestamp 1688980957
transform 1 0 42412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1236__RESET_B
timestamp 1688980957
transform 1 0 42780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1237__CLK
timestamp 1688980957
transform 1 0 43056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1237__RESET_B
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1238__CLK
timestamp 1688980957
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1238__SET_B
timestamp 1688980957
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1239__CLK
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1239__RESET_B
timestamp 1688980957
transform 1 0 22356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1240__CLK
timestamp 1688980957
transform 1 0 21896 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1240__RESET_B
timestamp 1688980957
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1241__CLK
timestamp 1688980957
transform 1 0 25852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1241__RESET_B
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1242__CLK
timestamp 1688980957
transform 1 0 26036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1242__RESET_B
timestamp 1688980957
transform 1 0 26496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1243__CLK
timestamp 1688980957
transform 1 0 35512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1243__RESET_B
timestamp 1688980957
transform 1 0 36432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1244__CLK
timestamp 1688980957
transform 1 0 13156 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1245__CLK
timestamp 1688980957
transform 1 0 33120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1245__RESET_B
timestamp 1688980957
transform 1 0 32752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1246__CLK
timestamp 1688980957
transform 1 0 26772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1246__RESET_B
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1247__CLK
timestamp 1688980957
transform 1 0 30360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1247__RESET_B
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1248__CLK
timestamp 1688980957
transform 1 0 29072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1248__RESET_B
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1249__CLK
timestamp 1688980957
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1249__RESET_B
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1250__CLK
timestamp 1688980957
transform 1 0 36800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1250__RESET_B
timestamp 1688980957
transform 1 0 39376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1251__CLK
timestamp 1688980957
transform 1 0 24472 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1251__RESET_B
timestamp 1688980957
transform 1 0 35512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1252__CLK
timestamp 1688980957
transform 1 0 32200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1252__RESET_B
timestamp 1688980957
transform 1 0 32936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1253__CLK
timestamp 1688980957
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1253__RESET_B
timestamp 1688980957
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1254__CLK
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1254__RESET_B
timestamp 1688980957
transform 1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1255__CLK
timestamp 1688980957
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1255__RESET_B
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1256__CLK
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1256__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1257__CLK
timestamp 1688980957
transform 1 0 9844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1257__RESET_B
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1258__CLK
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1258__RESET_B
timestamp 1688980957
transform 1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1259__CLK
timestamp 1688980957
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1259__RESET_B
timestamp 1688980957
transform 1 0 10948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1260__CLK
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1260__RESET_B
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1261__CLK
timestamp 1688980957
transform 1 0 7636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1261__RESET_B
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1262__CLK
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1262__RESET_B
timestamp 1688980957
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1263__CLK
timestamp 1688980957
transform 1 0 11684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1263__RESET_B
timestamp 1688980957
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1264__CLK
timestamp 1688980957
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1264__RESET_B
timestamp 1688980957
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1265__CLK
timestamp 1688980957
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1265__RESET_B
timestamp 1688980957
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1266__CLK
timestamp 1688980957
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1266__RESET_B
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1267__CLK
timestamp 1688980957
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1267__RESET_B
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1268__CLK
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1268__RESET_B
timestamp 1688980957
transform 1 0 31556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1269__CLK
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1269__RESET_B
timestamp 1688980957
transform 1 0 36800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1270__CLK
timestamp 1688980957
transform 1 0 38640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1270__RESET_B
timestamp 1688980957
transform 1 0 40204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1271__CLK
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1272__CLK
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1272__RESET_B
timestamp 1688980957
transform 1 0 42872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1273__CLK
timestamp 1688980957
transform 1 0 42688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1273__RESET_B
timestamp 1688980957
transform 1 0 43240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1274__CLK
timestamp 1688980957
transform 1 0 43424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1274__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1275__CLK
timestamp 1688980957
transform 1 0 42780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1275__RESET_B
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1276__CLK
timestamp 1688980957
transform 1 0 44252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1276__RESET_B
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1277__CLK
timestamp 1688980957
transform 1 0 38732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1277__RESET_B
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1278__CLK
timestamp 1688980957
transform 1 0 43700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1278__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1279__CLK
timestamp 1688980957
transform 1 0 44160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1279__RESET_B
timestamp 1688980957
transform 1 0 44528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1280__CLK
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1280__RESET_B
timestamp 1688980957
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1281__CLK
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1281__RESET_B
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1282__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1282__RESET_B
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1283__CLK
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1283__RESET_B
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1284__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1284__RESET_B
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1285__CLK
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1285__RESET_B
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1286__CLK
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1286__RESET_B
timestamp 1688980957
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1287__CLK
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1287__RESET_B
timestamp 1688980957
transform 1 0 4140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1288__CLK
timestamp 1688980957
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1288__RESET_B
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1289__CLK
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1289__RESET_B
timestamp 1688980957
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1290__CLK
timestamp 1688980957
transform 1 0 4232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1290__RESET_B
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1291__CLK
timestamp 1688980957
transform 1 0 3864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1291__RESET_B
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1292__CLK
timestamp 1688980957
transform 1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1292__RESET_B
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1293__CLK
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1293__RESET_B
timestamp 1688980957
transform 1 0 6348 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1294__CLK
timestamp 1688980957
transform 1 0 7360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1294__RESET_B
timestamp 1688980957
transform 1 0 8004 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1295__CLK
timestamp 1688980957
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1295__RESET_B
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1296__CLK
timestamp 1688980957
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1296__RESET_B
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1297__CLK
timestamp 1688980957
transform 1 0 9476 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1297__RESET_B
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1298__CLK
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1298__RESET_B
timestamp 1688980957
transform 1 0 8004 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1299__CLK
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1299__RESET_B
timestamp 1688980957
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1300__CLK
timestamp 1688980957
transform 1 0 10948 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1300__RESET_B
timestamp 1688980957
transform 1 0 10580 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1301__CLK
timestamp 1688980957
transform 1 0 11316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1301__RESET_B
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1302__CLK
timestamp 1688980957
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1302__RESET_B
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1303__CLK
timestamp 1688980957
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1303__RESET_B
timestamp 1688980957
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1304__CLK
timestamp 1688980957
transform 1 0 21252 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1304__RESET_B
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1305__CLK
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1305__RESET_B
timestamp 1688980957
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1306__CLK
timestamp 1688980957
transform 1 0 22264 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1306__RESET_B
timestamp 1688980957
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1307__CLK
timestamp 1688980957
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1307__RESET_B
timestamp 1688980957
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1308__CLK
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1308__RESET_B
timestamp 1688980957
transform 1 0 20056 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1309__CLK
timestamp 1688980957
transform 1 0 13156 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1309__RESET_B
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1310__CLK
timestamp 1688980957
transform 1 0 12788 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1310__RESET_B
timestamp 1688980957
transform 1 0 13892 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1311__CLK
timestamp 1688980957
transform 1 0 11776 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1311__SET_B
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1312__CLK
timestamp 1688980957
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1312__SET_B
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1313__CLK
timestamp 1688980957
transform 1 0 12052 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1313__RESET_B
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1314__CLK
timestamp 1688980957
transform 1 0 12420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1314__SET_B
timestamp 1688980957
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1315__CLK
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1315__SET_B
timestamp 1688980957
transform 1 0 12052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1316__CLK
timestamp 1688980957
transform 1 0 12420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1316__SET_B
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1317__CLK
timestamp 1688980957
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1317__SET_B
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1318__CLK
timestamp 1688980957
transform 1 0 10580 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1318__SET_B
timestamp 1688980957
transform 1 0 13156 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1319__CLK
timestamp 1688980957
transform 1 0 13156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1319__RESET_B
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1320__CLK
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1320__RESET_B
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1321__CLK
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1321__SET_B
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1322__CLK
timestamp 1688980957
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1322__RESET_B
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1323__CLK
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1323__RESET_B
timestamp 1688980957
transform 1 0 26404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1324__CLK
timestamp 1688980957
transform 1 0 44528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1324__RESET_B
timestamp 1688980957
transform 1 0 43884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1325__CLK
timestamp 1688980957
transform 1 0 44528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1325__RESET_B
timestamp 1688980957
transform 1 0 44160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1326__CLK
timestamp 1688980957
transform 1 0 44528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1326__RESET_B
timestamp 1688980957
transform 1 0 43884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1327__CLK
timestamp 1688980957
transform 1 0 43792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1327__RESET_B
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1328__CLK
timestamp 1688980957
transform 1 0 44160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1328__RESET_B
timestamp 1688980957
transform 1 0 44896 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1329__CLK
timestamp 1688980957
transform 1 0 43700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1329__RESET_B
timestamp 1688980957
transform 1 0 44068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1330__CLK
timestamp 1688980957
transform 1 0 44620 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1330__RESET_B
timestamp 1688980957
transform 1 0 44988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1331__CLK
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1331__RESET_B
timestamp 1688980957
transform 1 0 44252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1332__CLK
timestamp 1688980957
transform 1 0 40848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1332__RESET_B
timestamp 1688980957
transform 1 0 41216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1333__CLK
timestamp 1688980957
transform 1 0 38732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1333__RESET_B
timestamp 1688980957
transform 1 0 40480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1334__CLK
timestamp 1688980957
transform 1 0 43332 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1334__RESET_B
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1335__CLK
timestamp 1688980957
transform 1 0 42872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1335__RESET_B
timestamp 1688980957
transform 1 0 43240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1336__CLK
timestamp 1688980957
transform 1 0 41584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1336__RESET_B
timestamp 1688980957
transform 1 0 41952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1337__CLK
timestamp 1688980957
transform 1 0 42320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1337__RESET_B
timestamp 1688980957
transform 1 0 42688 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1338__CLK
timestamp 1688980957
transform 1 0 41952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1338__RESET_B
timestamp 1688980957
transform 1 0 41676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1339__CLK
timestamp 1688980957
transform 1 0 26036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1339__RESET_B
timestamp 1688980957
transform 1 0 25944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1340__CLK
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1340__RESET_B
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1341__CLK
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1341__RESET_B
timestamp 1688980957
transform 1 0 17940 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1342__CLK
timestamp 1688980957
transform 1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1342__RESET_B
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1343__CLK
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1343__RESET_B
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1344__CLK
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1344__RESET_B
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1345__CLK
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1345__RESET_B
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1346__CLK
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1346__RESET_B
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1347__CLK
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1347__RESET_B
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1348__CLK
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1348__RESET_B
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1349__CLK
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1349__RESET_B
timestamp 1688980957
transform 1 0 12420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1350__CLK
timestamp 1688980957
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1350__RESET_B
timestamp 1688980957
transform 1 0 13156 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1351__CLK
timestamp 1688980957
transform 1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1351__RESET_B
timestamp 1688980957
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1352__CLK
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1352__RESET_B
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1353__CLK
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1353__SET_B
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1354__CLK
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1355__CLK
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1356__CLK
timestamp 1688980957
transform 1 0 34040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1357__CLK
timestamp 1688980957
transform 1 0 36524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1358__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1359__CLK
timestamp 1688980957
transform 1 0 37076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1360__CLK
timestamp 1688980957
transform 1 0 35512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1361__CLK
timestamp 1688980957
transform 1 0 37628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1362__CLK
timestamp 1688980957
transform 1 0 20884 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1362__RESET_B
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1363__CLK
timestamp 1688980957
transform 1 0 14260 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1363__RESET_B
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1364__CLK
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1364__RESET_B
timestamp 1688980957
transform 1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1365__CLK
timestamp 1688980957
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1365__RESET_B
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1366__CLK
timestamp 1688980957
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1366__RESET_B
timestamp 1688980957
transform 1 0 24748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1367__CLK
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1367__RESET_B
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1368__CLK
timestamp 1688980957
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1368__RESET_B
timestamp 1688980957
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1369__CLK
timestamp 1688980957
transform 1 0 14628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1369__RESET_B
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1370__CLK
timestamp 1688980957
transform 1 0 20976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_INST_config_UART._1370__RESET_B
timestamp 1688980957
transform 1 0 21344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew111_A
timestamp 1688980957
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew112_A
timestamp 1688980957
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1688980957
transform 1 0 5428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1688980957
transform 1 0 42780 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__and2b_1  ConfigFSM_inst._120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27048 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  ConfigFSM_inst._121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27876 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  ConfigFSM_inst._122_
timestamp 1688980957
transform 1 0 29164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  ConfigFSM_inst._123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  ConfigFSM_inst._124_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  ConfigFSM_inst._125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  ConfigFSM_inst._126_
timestamp 1688980957
transform 1 0 24932 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  ConfigFSM_inst._127_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25300 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  ConfigFSM_inst._128_
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  ConfigFSM_inst._129_
timestamp 1688980957
transform 1 0 22724 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  ConfigFSM_inst._130_
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  ConfigFSM_inst._131_
timestamp 1688980957
transform 1 0 23552 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  ConfigFSM_inst._132_
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  ConfigFSM_inst._133_
timestamp 1688980957
transform 1 0 24564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  ConfigFSM_inst._134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26404 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  ConfigFSM_inst._135_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._136_
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  ConfigFSM_inst._137_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  ConfigFSM_inst._138_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  ConfigFSM_inst._139_
timestamp 1688980957
transform 1 0 30176 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  ConfigFSM_inst._140_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28796 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_4  ConfigFSM_inst._141_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  ConfigFSM_inst._142_
timestamp 1688980957
transform 1 0 26680 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  ConfigFSM_inst._143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  ConfigFSM_inst._144_
timestamp 1688980957
transform 1 0 25944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  ConfigFSM_inst._145_
timestamp 1688980957
transform 1 0 27692 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  ConfigFSM_inst._146_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  ConfigFSM_inst._147_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  ConfigFSM_inst._148_
timestamp 1688980957
transform 1 0 25392 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._149_
timestamp 1688980957
transform 1 0 28520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  ConfigFSM_inst._150_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28888 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._151_
timestamp 1688980957
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  ConfigFSM_inst._152_
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._153_
timestamp 1688980957
transform 1 0 31096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  ConfigFSM_inst._154_
timestamp 1688980957
transform 1 0 30544 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._155_
timestamp 1688980957
transform 1 0 34040 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  ConfigFSM_inst._156_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  ConfigFSM_inst._157_
timestamp 1688980957
transform 1 0 32108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  ConfigFSM_inst._158_
timestamp 1688980957
transform 1 0 29992 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._159_
timestamp 1688980957
transform 1 0 35880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  ConfigFSM_inst._160_
timestamp 1688980957
transform 1 0 27232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._161_
timestamp 1688980957
transform 1 0 25116 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  ConfigFSM_inst._162_
timestamp 1688980957
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ConfigFSM_inst._163_
timestamp 1688980957
transform 1 0 28796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  ConfigFSM_inst._164_
timestamp 1688980957
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  ConfigFSM_inst._165_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._166_
timestamp 1688980957
transform 1 0 30728 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._167_
timestamp 1688980957
transform 1 0 33212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  ConfigFSM_inst._168_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  ConfigFSM_inst._169_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  ConfigFSM_inst._170_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  ConfigFSM_inst._171_
timestamp 1688980957
transform 1 0 33304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  ConfigFSM_inst._172_
timestamp 1688980957
transform 1 0 33488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  ConfigFSM_inst._173_
timestamp 1688980957
transform 1 0 31464 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  ConfigFSM_inst._174_
timestamp 1688980957
transform 1 0 31096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  ConfigFSM_inst._175_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  ConfigFSM_inst._176_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  ConfigFSM_inst._177_
timestamp 1688980957
transform 1 0 29716 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  ConfigFSM_inst._178_
timestamp 1688980957
transform 1 0 28520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  ConfigFSM_inst._179_
timestamp 1688980957
transform 1 0 29072 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  ConfigFSM_inst._180_
timestamp 1688980957
transform 1 0 28244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._181_
timestamp 1688980957
transform 1 0 3128 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._182_
timestamp 1688980957
transform 1 0 920 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._183_
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._184_
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._185_
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._186_
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._187_
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._188_
timestamp 1688980957
transform 1 0 3312 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._189_
timestamp 1688980957
transform 1 0 4140 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._190_
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._191_
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._192_
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._193_
timestamp 1688980957
transform 1 0 5888 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._194_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._195_
timestamp 1688980957
transform 1 0 6716 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._196_
timestamp 1688980957
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._197_
timestamp 1688980957
transform 1 0 8280 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._198_
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ConfigFSM_inst._199_
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._200_
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._201_
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._202_
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._203_
timestamp 1688980957
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._204_
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._205_
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._206_
timestamp 1688980957
transform 1 0 10948 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._207_
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._208_
timestamp 1688980957
transform 1 0 11684 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._209_
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._210_
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._211_
timestamp 1688980957
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._212_
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._213_
timestamp 1688980957
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._214_
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._215_
timestamp 1688980957
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._216_
timestamp 1688980957
transform 1 0 16008 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._217_
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._218_
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._219_
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ConfigFSM_inst._220_
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._221_
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._222_
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._223_
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._224_
timestamp 1688980957
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._225_
timestamp 1688980957
transform 1 0 19780 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._226_
timestamp 1688980957
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._227_
timestamp 1688980957
transform 1 0 21160 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._228_
timestamp 1688980957
transform 1 0 20424 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._229_
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._230_
timestamp 1688980957
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._231_
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._232_
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._233_
timestamp 1688980957
transform 1 0 23092 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._234_
timestamp 1688980957
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._235_
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._236_
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._237_
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._238_
timestamp 1688980957
transform 1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._239_
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._240_
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._241_
timestamp 1688980957
transform 1 0 25024 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._242_
timestamp 1688980957
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ConfigFSM_inst._243_
timestamp 1688980957
transform 1 0 25852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ConfigFSM_inst._244_
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  ConfigFSM_inst._245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  ConfigFSM_inst._246_
timestamp 1688980957
transform 1 0 31924 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._247_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31648 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  ConfigFSM_inst._248_
timestamp 1688980957
transform 1 0 29164 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._249_
timestamp 1688980957
transform 1 0 28152 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  ConfigFSM_inst._250_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  ConfigFSM_inst._251_
timestamp 1688980957
transform 1 0 26588 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._252_
timestamp 1688980957
transform 1 0 25760 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._253_
timestamp 1688980957
transform 1 0 26312 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._254_
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._255_
timestamp 1688980957
transform 1 0 1196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._256_
timestamp 1688980957
transform 1 0 1196 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._257_
timestamp 1688980957
transform 1 0 1472 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._258_
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._259_
timestamp 1688980957
transform 1 0 3312 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._260_
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._261_
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._262_
timestamp 1688980957
transform 1 0 5888 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._263_
timestamp 1688980957
transform 1 0 6532 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._264_
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._265_
timestamp 1688980957
transform 1 0 8648 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._266_
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._267_
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._268_
timestamp 1688980957
transform 1 0 11316 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._269_
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._270_
timestamp 1688980957
transform 1 0 12512 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._271_
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._272_
timestamp 1688980957
transform 1 0 14260 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._273_
timestamp 1688980957
transform 1 0 14996 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._274_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._275_
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._276_
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._277_
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._278_
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._279_
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._280_
timestamp 1688980957
transform 1 0 21252 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._281_
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._282_
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._283_
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._284_
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._285_
timestamp 1688980957
transform 1 0 25576 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._286_
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  ConfigFSM_inst._287_
timestamp 1688980957
transform 1 0 25392 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_20
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_24
timestamp 1688980957
transform 1 0 2668 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_47
timestamp 1688980957
transform 1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65
timestamp 1688980957
transform 1 0 6440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_74
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_92
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_101
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 10580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_119
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_128
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_146
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_155
timestamp 1688980957
transform 1 0 14720 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_164
timestamp 1688980957
transform 1 0 15548 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_173
timestamp 1688980957
transform 1 0 16376 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_182 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_188
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_192
timestamp 1688980957
transform 1 0 18124 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_201
timestamp 1688980957
transform 1 0 18952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_209
timestamp 1688980957
transform 1 0 19688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_218
timestamp 1688980957
transform 1 0 20516 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_236
timestamp 1688980957
transform 1 0 22172 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23000 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_256
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_278
timestamp 1688980957
transform 1 0 26036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_293
timestamp 1688980957
transform 1 0 27416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_321
timestamp 1688980957
transform 1 0 29992 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_371
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 36432 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_455
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_460
timestamp 1688980957
transform 1 0 42780 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_464
timestamp 1688980957
transform 1 0 43148 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_469
timestamp 1688980957
transform 1 0 43608 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 43976 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_480
timestamp 1688980957
transform 1 0 44620 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_3
timestamp 1688980957
transform 1 0 736 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_7
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_10
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_14
timestamp 1688980957
transform 1 0 1748 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_21
timestamp 1688980957
transform 1 0 2392 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_27
timestamp 1688980957
transform 1 0 2944 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_34
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4048 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_47
timestamp 1688980957
transform 1 0 4784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 5428 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1688980957
transform 1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_65
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_71
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_75
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_82
timestamp 1688980957
transform 1 0 8004 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_88
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_95
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_103
timestamp 1688980957
transform 1 0 9936 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 10580 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_119
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_154
timestamp 1688980957
transform 1 0 14628 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_158
timestamp 1688980957
transform 1 0 14996 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1688980957
transform 1 0 15640 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_174
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_180
timestamp 1688980957
transform 1 0 17020 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_197
timestamp 1688980957
transform 1 0 18584 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_201
timestamp 1688980957
transform 1 0 18952 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19320 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_212
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_220
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_234
timestamp 1688980957
transform 1 0 21988 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26128 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1688980957
transform 1 0 31832 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_416
timestamp 1688980957
transform 1 0 38732 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_443
timestamp 1688980957
transform 1 0 41216 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 41584 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_449
timestamp 1688980957
transform 1 0 41768 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_453
timestamp 1688980957
transform 1 0 42136 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_457
timestamp 1688980957
transform 1 0 42504 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_461
timestamp 1688980957
transform 1 0 42872 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_465
timestamp 1688980957
transform 1 0 43240 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_469
timestamp 1688980957
transform 1 0 43608 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_473
timestamp 1688980957
transform 1 0 43976 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_477
timestamp 1688980957
transform 1 0 44344 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_481
timestamp 1688980957
transform 1 0 44712 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_485
timestamp 1688980957
transform 1 0 45080 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3
timestamp 1688980957
transform 1 0 736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_8
timestamp 1688980957
transform 1 0 1196 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_15
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_49
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_55
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_59
timestamp 1688980957
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_63
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_67
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_74
timestamp 1688980957
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_80
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_90
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_103
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_124
timestamp 1688980957
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_132
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_136
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_147
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_170
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1688980957
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_231
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_300
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_309
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_448
timestamp 1688980957
transform 1 0 41676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_452
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_456
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_460
timestamp 1688980957
transform 1 0 42780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_464
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_468
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_472
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_477
timestamp 1688980957
transform 1 0 44344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_481
timestamp 1688980957
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_485
timestamp 1688980957
transform 1 0 45080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_6
timestamp 1688980957
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_31
timestamp 1688980957
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_46
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_52
timestamp 1688980957
transform 1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_79
timestamp 1688980957
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_83
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1688980957
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_123
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_127
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_153
timestamp 1688980957
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_159
timestamp 1688980957
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_164
timestamp 1688980957
transform 1 0 15548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_178
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_220
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_326
timestamp 1688980957
transform 1 0 30452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 1688980957
transform 1 0 31188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_337
timestamp 1688980957
transform 1 0 31464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_362
timestamp 1688980957
transform 1 0 33764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_387
timestamp 1688980957
transform 1 0 36064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_442
timestamp 1688980957
transform 1 0 41124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_446
timestamp 1688980957
transform 1 0 41492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_449
timestamp 1688980957
transform 1 0 41768 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_453
timestamp 1688980957
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_457
timestamp 1688980957
transform 1 0 42504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_461
timestamp 1688980957
transform 1 0 42872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_465
timestamp 1688980957
transform 1 0 43240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1688980957
transform 1 0 736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_8
timestamp 1688980957
transform 1 0 1196 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_12
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_16
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_20
timestamp 1688980957
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_24
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_51
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_56
timestamp 1688980957
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_60
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_67
timestamp 1688980957
transform 1 0 6624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_77
timestamp 1688980957
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_81
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_114
timestamp 1688980957
transform 1 0 10948 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 13432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_151
timestamp 1688980957
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 18584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_248
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_262
timestamp 1688980957
transform 1 0 24564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_266
timestamp 1688980957
transform 1 0 24932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_296
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_336
timestamp 1688980957
transform 1 0 31372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_359
timestamp 1688980957
transform 1 0 33488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 33856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_375
timestamp 1688980957
transform 1 0 34960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_394
timestamp 1688980957
transform 1 0 36708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_416
timestamp 1688980957
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_441
timestamp 1688980957
transform 1 0 41032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_445
timestamp 1688980957
transform 1 0 41400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_449
timestamp 1688980957
transform 1 0 41768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_453
timestamp 1688980957
transform 1 0 42136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_457
timestamp 1688980957
transform 1 0 42504 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_461
timestamp 1688980957
transform 1 0 42872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_465
timestamp 1688980957
transform 1 0 43240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_469
timestamp 1688980957
transform 1 0 43608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_473
timestamp 1688980957
transform 1 0 43976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_481
timestamp 1688980957
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_485
timestamp 1688980957
transform 1 0 45080 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 1688980957
transform 1 0 736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_28
timestamp 1688980957
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_32
timestamp 1688980957
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_60
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_86
timestamp 1688980957
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_143
timestamp 1688980957
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_153
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_160
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_164
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_199
timestamp 1688980957
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_209
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_219
timestamp 1688980957
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21160 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_255
timestamp 1688980957
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_260
timestamp 1688980957
transform 1 0 24380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_287
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_301
timestamp 1688980957
transform 1 0 28152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_337
timestamp 1688980957
transform 1 0 31464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_365
timestamp 1688980957
transform 1 0 34040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_386
timestamp 1688980957
transform 1 0 35972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1688980957
transform 1 0 36340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_393
timestamp 1688980957
transform 1 0 36616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_397
timestamp 1688980957
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_401
timestamp 1688980957
transform 1 0 37352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 1688980957
transform 1 0 37720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 41584 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_449
timestamp 1688980957
transform 1 0 41768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_453
timestamp 1688980957
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_457
timestamp 1688980957
transform 1 0 42504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_461
timestamp 1688980957
transform 1 0 42872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_465
timestamp 1688980957
transform 1 0 43240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_469
timestamp 1688980957
transform 1 0 43608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_473
timestamp 1688980957
transform 1 0 43976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_477
timestamp 1688980957
transform 1 0 44344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_481
timestamp 1688980957
transform 1 0 44712 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_485
timestamp 1688980957
transform 1 0 45080 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_38
timestamp 1688980957
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_69
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_75
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_80
timestamp 1688980957
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_94
timestamp 1688980957
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_102
timestamp 1688980957
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_113
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_118
timestamp 1688980957
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_145
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_172
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1688980957
transform 1 0 18584 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_204
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_214
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_218
timestamp 1688980957
transform 1 0 20516 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_221
timestamp 1688980957
transform 1 0 20792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_262
timestamp 1688980957
transform 1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 28704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_316
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_340
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_403
timestamp 1688980957
transform 1 0 37536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_407
timestamp 1688980957
transform 1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_413
timestamp 1688980957
transform 1 0 38456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_439
timestamp 1688980957
transform 1 0 40848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_443
timestamp 1688980957
transform 1 0 41216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_447
timestamp 1688980957
transform 1 0 41584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_451
timestamp 1688980957
transform 1 0 41952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_455
timestamp 1688980957
transform 1 0 42320 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_459
timestamp 1688980957
transform 1 0 42688 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_463
timestamp 1688980957
transform 1 0 43056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_467
timestamp 1688980957
transform 1 0 43424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_471
timestamp 1688980957
transform 1 0 43792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44160 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_481
timestamp 1688980957
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_485
timestamp 1688980957
transform 1 0 45080 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 1688980957
transform 1 0 736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_8
timestamp 1688980957
transform 1 0 1196 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_25
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_29
timestamp 1688980957
transform 1 0 3128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_33
timestamp 1688980957
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_38
timestamp 1688980957
transform 1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_45
timestamp 1688980957
transform 1 0 4600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_72
timestamp 1688980957
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_76
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_80
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_88
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_92
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_96
timestamp 1688980957
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_100
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_104
timestamp 1688980957
transform 1 0 10028 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_108
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_118
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_122
timestamp 1688980957
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_129
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_133
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_136
timestamp 1688980957
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_140
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_144
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_232
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_236
timestamp 1688980957
transform 1 0 22172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_240
timestamp 1688980957
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_260
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_276
timestamp 1688980957
transform 1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_366
timestamp 1688980957
transform 1 0 34132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_396
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_400
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_404
timestamp 1688980957
transform 1 0 37628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_443
timestamp 1688980957
transform 1 0 41216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 41584 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_449
timestamp 1688980957
transform 1 0 41768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_453
timestamp 1688980957
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_457
timestamp 1688980957
transform 1 0 42504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_461
timestamp 1688980957
transform 1 0 42872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_465
timestamp 1688980957
transform 1 0 43240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_469
timestamp 1688980957
transform 1 0 43608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_473
timestamp 1688980957
transform 1 0 43976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_477
timestamp 1688980957
transform 1 0 44344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_481
timestamp 1688980957
transform 1 0 44712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_485
timestamp 1688980957
transform 1 0 45080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1688980957
transform 1 0 736 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_10
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_33
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1688980957
transform 1 0 3864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_40
timestamp 1688980957
transform 1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_45
timestamp 1688980957
transform 1 0 4600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_51
timestamp 1688980957
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_55
timestamp 1688980957
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_59
timestamp 1688980957
transform 1 0 5888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_65
timestamp 1688980957
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_69
timestamp 1688980957
transform 1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_73
timestamp 1688980957
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_77
timestamp 1688980957
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_81
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_89
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_92
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_96
timestamp 1688980957
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_100
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_104
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_108
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_112
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_116
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_120
timestamp 1688980957
transform 1 0 11500 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_124
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_128
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_132
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_136
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_145
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_149
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_170
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1688980957
transform 1 0 18308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_232
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_236
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_242
timestamp 1688980957
transform 1 0 22724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_262
timestamp 1688980957
transform 1 0 24564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_303
timestamp 1688980957
transform 1 0 28336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 33856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_372
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_407
timestamp 1688980957
transform 1 0 37904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_418
timestamp 1688980957
transform 1 0 38916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_461
timestamp 1688980957
transform 1 0 42872 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_465
timestamp 1688980957
transform 1 0 43240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_469
timestamp 1688980957
transform 1 0 43608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1688980957
transform 1 0 43976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44344 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_481
timestamp 1688980957
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_485
timestamp 1688980957
transform 1 0 45080 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 736 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 1840 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 2944 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 1688980957
transform 1 0 6440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_68
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_76
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_80
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_88
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_92
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_96
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_100
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_104
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_108
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_120
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_124
timestamp 1688980957
transform 1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_132
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_140
timestamp 1688980957
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_144
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_186
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_190
timestamp 1688980957
transform 1 0 17940 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_232
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_258
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_262
timestamp 1688980957
transform 1 0 24564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_266
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp 1688980957
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_295
timestamp 1688980957
transform 1 0 27600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_314
timestamp 1688980957
transform 1 0 29348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_337
timestamp 1688980957
transform 1 0 31464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_365
timestamp 1688980957
transform 1 0 34040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 36432 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_393
timestamp 1688980957
transform 1 0 36616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 41584 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_467
timestamp 1688980957
transform 1 0 43424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_471
timestamp 1688980957
transform 1 0 43792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_475
timestamp 1688980957
transform 1 0 44160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_479
timestamp 1688980957
transform 1 0 44528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_483
timestamp 1688980957
transform 1 0 44896 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 736 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3128 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5336 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_65
timestamp 1688980957
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_69
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_72
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_76
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_80
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_89
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_92
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_96
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_100
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_108
timestamp 1688980957
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_112
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_116
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_120
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_124
timestamp 1688980957
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_128
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_132
timestamp 1688980957
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_136
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_148
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_152
timestamp 1688980957
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_188
timestamp 1688980957
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_192
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_197
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_201
timestamp 1688980957
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_216
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_222
timestamp 1688980957
transform 1 0 20884 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_257
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_261
timestamp 1688980957
transform 1 0 24472 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_265
timestamp 1688980957
transform 1 0 24840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_269
timestamp 1688980957
transform 1 0 25208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_280
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_284
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_288
timestamp 1688980957
transform 1 0 26956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_292
timestamp 1688980957
transform 1 0 27324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_296
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_336
timestamp 1688980957
transform 1 0 31372 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_370
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_399
timestamp 1688980957
transform 1 0 37168 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_418
timestamp 1688980957
transform 1 0 38916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_470
timestamp 1688980957
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_474
timestamp 1688980957
transform 1 0 44068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_481
timestamp 1688980957
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_485
timestamp 1688980957
transform 1 0 45080 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 736 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 5520 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_69
timestamp 1688980957
transform 1 0 6808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_77
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_80
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_84
timestamp 1688980957
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_88
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_120
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_124
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_128
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_132
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_136
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_144
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_148
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_152
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_197
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_267
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_271
timestamp 1688980957
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_275
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_337
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_358
timestamp 1688980957
transform 1 0 33396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_379
timestamp 1688980957
transform 1 0 35328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_390
timestamp 1688980957
transform 1 0 36340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_393
timestamp 1688980957
transform 1 0 36616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_404
timestamp 1688980957
transform 1 0 37628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_440
timestamp 1688980957
transform 1 0 40940 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 41584 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_458
timestamp 1688980957
transform 1 0 42596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_462
timestamp 1688980957
transform 1 0 42964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_466
timestamp 1688980957
transform 1 0 43332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_470
timestamp 1688980957
transform 1 0 43700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_474
timestamp 1688980957
transform 1 0 44068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_478
timestamp 1688980957
transform 1 0 44436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_482
timestamp 1688980957
transform 1 0 44804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_486
timestamp 1688980957
transform 1 0 45172 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 736 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3128 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_77
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_80
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_124
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_129
timestamp 1688980957
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_161
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_190
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_256
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 28704 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_334
timestamp 1688980957
transform 1 0 31188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_375
timestamp 1688980957
transform 1 0 34960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_406
timestamp 1688980957
transform 1 0 37812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_410
timestamp 1688980957
transform 1 0 38180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_414
timestamp 1688980957
transform 1 0 38548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_418
timestamp 1688980957
transform 1 0 38916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_464
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_468
timestamp 1688980957
transform 1 0 43516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_472
timestamp 1688980957
transform 1 0 43884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_481
timestamp 1688980957
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_485
timestamp 1688980957
transform 1 0 45080 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 736 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_61
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_66
timestamp 1688980957
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_70
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_76
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_80
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_84
timestamp 1688980957
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_88
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_120
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_160
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_164
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_175
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_180
timestamp 1688980957
transform 1 0 17020 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_319
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_334
timestamp 1688980957
transform 1 0 31188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 36432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_433
timestamp 1688980957
transform 1 0 40296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 1688980957
transform 1 0 41492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_469
timestamp 1688980957
transform 1 0 43608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_473
timestamp 1688980957
transform 1 0 43976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_477
timestamp 1688980957
transform 1 0 44344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_481
timestamp 1688980957
transform 1 0 44712 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_485
timestamp 1688980957
transform 1 0 45080 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_7
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1688980957
transform 1 0 2208 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_62
timestamp 1688980957
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_68
timestamp 1688980957
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_72
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_76
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_80
timestamp 1688980957
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_100
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_107
timestamp 1688980957
transform 1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_112
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_150
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_155
timestamp 1688980957
transform 1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_159
timestamp 1688980957
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_163
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_197
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_238
timestamp 1688980957
transform 1 0 22356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_274
timestamp 1688980957
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_278
timestamp 1688980957
transform 1 0 26036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_355
timestamp 1688980957
transform 1 0 33120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_393
timestamp 1688980957
transform 1 0 36616 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_468
timestamp 1688980957
transform 1 0 43516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_472
timestamp 1688980957
transform 1 0 43884 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_477
timestamp 1688980957
transform 1 0 44344 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_481
timestamp 1688980957
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_485
timestamp 1688980957
transform 1 0 45080 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 736 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_27
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_35
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_64
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_68
timestamp 1688980957
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_72
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_76
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1688980957
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_124
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 1688980957
transform 1 0 12696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_157
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_214
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_233
timestamp 1688980957
transform 1 0 21896 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_271
timestamp 1688980957
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_275
timestamp 1688980957
transform 1 0 25760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_342
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_352
timestamp 1688980957
transform 1 0 32844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_367
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_436
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_440
timestamp 1688980957
transform 1 0 40940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_455
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_459
timestamp 1688980957
transform 1 0 42688 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_463
timestamp 1688980957
transform 1 0 43056 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 736 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 2944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_134
timestamp 1688980957
transform 1 0 12788 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_156
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_186
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_302
timestamp 1688980957
transform 1 0 28244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 33856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_412
timestamp 1688980957
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_430
timestamp 1688980957
transform 1 0 40020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_434
timestamp 1688980957
transform 1 0 40388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_455
timestamp 1688980957
transform 1 0 42320 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_459
timestamp 1688980957
transform 1 0 42688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_463
timestamp 1688980957
transform 1 0 43056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_467
timestamp 1688980957
transform 1 0 43424 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_471
timestamp 1688980957
transform 1 0 43792 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 1688980957
transform 1 0 44160 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_477
timestamp 1688980957
transform 1 0 44344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_481
timestamp 1688980957
transform 1 0 44712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_485
timestamp 1688980957
transform 1 0 45080 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 736 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1688980957
transform 1 0 2944 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_49
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_63
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_67
timestamp 1688980957
transform 1 0 6624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_70
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_74
timestamp 1688980957
transform 1 0 7268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_78
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_165
timestamp 1688980957
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_178
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_242
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_268
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_272
timestamp 1688980957
transform 1 0 25484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_276
timestamp 1688980957
transform 1 0 25852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_310
timestamp 1688980957
transform 1 0 28980 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_327
timestamp 1688980957
transform 1 0 30544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_396
timestamp 1688980957
transform 1 0 36892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_400
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_446
timestamp 1688980957
transform 1 0 41492 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_452
timestamp 1688980957
transform 1 0 42044 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_456
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_460
timestamp 1688980957
transform 1 0 42780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_464
timestamp 1688980957
transform 1 0 43148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_468
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_472
timestamp 1688980957
transform 1 0 43884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_476
timestamp 1688980957
transform 1 0 44252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_480
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_484
timestamp 1688980957
transform 1 0 44988 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 736 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 2944 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3128 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_51
timestamp 1688980957
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_55
timestamp 1688980957
transform 1 0 5520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_59
timestamp 1688980957
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_64
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_68
timestamp 1688980957
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_72
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_76
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_80
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_100
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_113
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_132
timestamp 1688980957
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_136
timestamp 1688980957
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_156
timestamp 1688980957
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 1688980957
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_183
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1688980957
transform 1 0 18584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_201
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_205
timestamp 1688980957
transform 1 0 19320 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_208
timestamp 1688980957
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_215
timestamp 1688980957
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_219
timestamp 1688980957
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_241
timestamp 1688980957
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_253
timestamp 1688980957
transform 1 0 23736 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_268
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_272
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_276
timestamp 1688980957
transform 1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_302
timestamp 1688980957
transform 1 0 28244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_321
timestamp 1688980957
transform 1 0 29992 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_368
timestamp 1688980957
transform 1 0 34316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_393
timestamp 1688980957
transform 1 0 36616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_397
timestamp 1688980957
transform 1 0 36984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_441
timestamp 1688980957
transform 1 0 41032 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_451
timestamp 1688980957
transform 1 0 41952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_455
timestamp 1688980957
transform 1 0 42320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_459
timestamp 1688980957
transform 1 0 42688 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_463
timestamp 1688980957
transform 1 0 43056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_467
timestamp 1688980957
transform 1 0 43424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_471
timestamp 1688980957
transform 1 0 43792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44160 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44344 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_481
timestamp 1688980957
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_485
timestamp 1688980957
transform 1 0 45080 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 736 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_47
timestamp 1688980957
transform 1 0 4784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_77
timestamp 1688980957
transform 1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_82
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_86
timestamp 1688980957
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_90
timestamp 1688980957
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_94
timestamp 1688980957
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_107
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_123
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_216
timestamp 1688980957
transform 1 0 20332 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_228
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_333
timestamp 1688980957
transform 1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_345
timestamp 1688980957
transform 1 0 32200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_349
timestamp 1688980957
transform 1 0 32568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_353
timestamp 1688980957
transform 1 0 32936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_379
timestamp 1688980957
transform 1 0 35328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_383
timestamp 1688980957
transform 1 0 35696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 36432 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_439
timestamp 1688980957
transform 1 0 40848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_443
timestamp 1688980957
transform 1 0 41216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1688980957
transform 1 0 41584 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_449
timestamp 1688980957
transform 1 0 41768 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_453
timestamp 1688980957
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_457
timestamp 1688980957
transform 1 0 42504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_461
timestamp 1688980957
transform 1 0 42872 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 736 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 1840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 2944 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3128 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_79
timestamp 1688980957
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_91
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_95
timestamp 1688980957
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_119
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_124
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_133
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13064 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_141
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_158
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_179
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_185
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_221
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_244
timestamp 1688980957
transform 1 0 22908 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27232 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_305
timestamp 1688980957
transform 1 0 28520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_309
timestamp 1688980957
transform 1 0 28888 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_339
timestamp 1688980957
transform 1 0 31648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_343
timestamp 1688980957
transform 1 0 32016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_353
timestamp 1688980957
transform 1 0 32936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_418
timestamp 1688980957
transform 1 0 38916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_430
timestamp 1688980957
transform 1 0 40020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_434
timestamp 1688980957
transform 1 0 40388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_438
timestamp 1688980957
transform 1 0 40756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_442
timestamp 1688980957
transform 1 0 41124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_446
timestamp 1688980957
transform 1 0 41492 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_450
timestamp 1688980957
transform 1 0 41860 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_454
timestamp 1688980957
transform 1 0 42228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_458
timestamp 1688980957
transform 1 0 42596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_462
timestamp 1688980957
transform 1 0 42964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_466
timestamp 1688980957
transform 1 0 43332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_470
timestamp 1688980957
transform 1 0 43700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_474
timestamp 1688980957
transform 1 0 44068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44344 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_481
timestamp 1688980957
transform 1 0 44712 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_485
timestamp 1688980957
transform 1 0 45080 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 736 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4048 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_45
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_77
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_82
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_86
timestamp 1688980957
transform 1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_132
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1688980957
transform 1 0 23000 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26128 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_286
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_296
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_314
timestamp 1688980957
transform 1 0 29348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_326
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_330
timestamp 1688980957
transform 1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_377
timestamp 1688980957
transform 1 0 35144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_390
timestamp 1688980957
transform 1 0 36340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_413
timestamp 1688980957
transform 1 0 38456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_433
timestamp 1688980957
transform 1 0 40296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_437
timestamp 1688980957
transform 1 0 40664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41032 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_445
timestamp 1688980957
transform 1 0 41400 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_449
timestamp 1688980957
transform 1 0 41768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_453
timestamp 1688980957
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_457
timestamp 1688980957
transform 1 0 42504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_461
timestamp 1688980957
transform 1 0 42872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_465
timestamp 1688980957
transform 1 0 43240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_469
timestamp 1688980957
transform 1 0 43608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_473
timestamp 1688980957
transform 1 0 43976 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_477
timestamp 1688980957
transform 1 0 44344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_481
timestamp 1688980957
transform 1 0 44712 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_485
timestamp 1688980957
transform 1 0 45080 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 736 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 2944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_34
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_38
timestamp 1688980957
transform 1 0 3956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_44
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_48
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_52
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_60
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_172
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_210
timestamp 1688980957
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_263
timestamp 1688980957
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_290
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_320
timestamp 1688980957
transform 1 0 29900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_324
timestamp 1688980957
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_362
timestamp 1688980957
transform 1 0 33764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_408
timestamp 1688980957
transform 1 0 37996 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_418
timestamp 1688980957
transform 1 0 38916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_441
timestamp 1688980957
transform 1 0 41032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_445
timestamp 1688980957
transform 1 0 41400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_449
timestamp 1688980957
transform 1 0 41768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_453
timestamp 1688980957
transform 1 0 42136 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_457
timestamp 1688980957
transform 1 0 42504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_461
timestamp 1688980957
transform 1 0 42872 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_465
timestamp 1688980957
transform 1 0 43240 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_469
timestamp 1688980957
transform 1 0 43608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_473
timestamp 1688980957
transform 1 0 43976 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44344 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_481
timestamp 1688980957
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_485
timestamp 1688980957
transform 1 0 45080 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1688980957
transform 1 0 736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_11
timestamp 1688980957
transform 1 0 1472 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_34
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1688980957
transform 1 0 5704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_67
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_71
timestamp 1688980957
transform 1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 15824 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_182
timestamp 1688980957
transform 1 0 17204 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_232
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_262
timestamp 1688980957
transform 1 0 24564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_315
timestamp 1688980957
transform 1 0 29440 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_337
timestamp 1688980957
transform 1 0 31464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_347
timestamp 1688980957
transform 1 0 32384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_351
timestamp 1688980957
transform 1 0 32752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_381
timestamp 1688980957
transform 1 0 35512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_393
timestamp 1688980957
transform 1 0 36616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_445
timestamp 1688980957
transform 1 0 41400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_458
timestamp 1688980957
transform 1 0 42596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_462
timestamp 1688980957
transform 1 0 42964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_466
timestamp 1688980957
transform 1 0 43332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_470
timestamp 1688980957
transform 1 0 43700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_474
timestamp 1688980957
transform 1 0 44068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_478
timestamp 1688980957
transform 1 0 44436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_482
timestamp 1688980957
transform 1 0 44804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_486
timestamp 1688980957
transform 1 0 45172 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 736 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 2944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_35
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_38
timestamp 1688980957
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_69
timestamp 1688980957
transform 1 0 6808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_74
timestamp 1688980957
transform 1 0 7268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1688980957
transform 1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_179
timestamp 1688980957
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_183
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_186
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_204
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_260
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 28704 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_325
timestamp 1688980957
transform 1 0 30360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_339
timestamp 1688980957
transform 1 0 31648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_343
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_347
timestamp 1688980957
transform 1 0 32384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_351
timestamp 1688980957
transform 1 0 32752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_355
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 33856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_378
timestamp 1688980957
transform 1 0 35236 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_390
timestamp 1688980957
transform 1 0 36340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_394
timestamp 1688980957
transform 1 0 36708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_404
timestamp 1688980957
transform 1 0 37628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_409
timestamp 1688980957
transform 1 0 38088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_441
timestamp 1688980957
transform 1 0 41032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_445
timestamp 1688980957
transform 1 0 41400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_457
timestamp 1688980957
transform 1 0 42504 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_461
timestamp 1688980957
transform 1 0 42872 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_465
timestamp 1688980957
transform 1 0 43240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_469
timestamp 1688980957
transform 1 0 43608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_473
timestamp 1688980957
transform 1 0 43976 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_481
timestamp 1688980957
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_485
timestamp 1688980957
transform 1 0 45080 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_6
timestamp 1688980957
transform 1 0 1012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_18
timestamp 1688980957
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_30
timestamp 1688980957
transform 1 0 3220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_36
timestamp 1688980957
transform 1 0 3772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_77
timestamp 1688980957
transform 1 0 7544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_108
timestamp 1688980957
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_128
timestamp 1688980957
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_147
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_151
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_155
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_187
timestamp 1688980957
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_191
timestamp 1688980957
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_194
timestamp 1688980957
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_198
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_202
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_206
timestamp 1688980957
transform 1 0 19412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_217
timestamp 1688980957
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_243
timestamp 1688980957
transform 1 0 22816 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_262
timestamp 1688980957
transform 1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_329
timestamp 1688980957
transform 1 0 30728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_357
timestamp 1688980957
transform 1 0 33304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_361
timestamp 1688980957
transform 1 0 33672 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_386
timestamp 1688980957
transform 1 0 35972 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_402
timestamp 1688980957
transform 1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_406
timestamp 1688980957
transform 1 0 37812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_410
timestamp 1688980957
transform 1 0 38180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_414
timestamp 1688980957
transform 1 0 38548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_427
timestamp 1688980957
transform 1 0 39744 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_469
timestamp 1688980957
transform 1 0 43608 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_473
timestamp 1688980957
transform 1 0 43976 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_477
timestamp 1688980957
transform 1 0 44344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_481
timestamp 1688980957
transform 1 0 44712 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 736 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 2944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_35
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_39
timestamp 1688980957
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_70
timestamp 1688980957
transform 1 0 6900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_130
timestamp 1688980957
transform 1 0 12420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13248 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_151
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_191
timestamp 1688980957
transform 1 0 18032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 18400 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_197
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_202
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_211
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_231
timestamp 1688980957
transform 1 0 21712 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_241
timestamp 1688980957
transform 1 0 22632 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_293
timestamp 1688980957
transform 1 0 27416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_324
timestamp 1688980957
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_410
timestamp 1688980957
transform 1 0 38180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_465
timestamp 1688980957
transform 1 0 43240 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_469
timestamp 1688980957
transform 1 0 43608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_473
timestamp 1688980957
transform 1 0 43976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_477
timestamp 1688980957
transform 1 0 44344 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_481
timestamp 1688980957
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_485
timestamp 1688980957
transform 1 0 45080 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 736 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_27
timestamp 1688980957
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_32
timestamp 1688980957
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_36
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_40
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_44
timestamp 1688980957
transform 1 0 4508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_48
timestamp 1688980957
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 5520 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_67
timestamp 1688980957
transform 1 0 6624 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_73
timestamp 1688980957
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_77
timestamp 1688980957
transform 1 0 7544 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_101
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_133
timestamp 1688980957
transform 1 0 12696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_158
timestamp 1688980957
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16008 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_212
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_220
timestamp 1688980957
transform 1 0 20700 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21160 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1688980957
transform 1 0 26036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_285
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_314
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_357
timestamp 1688980957
transform 1 0 33304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 36432 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_469
timestamp 1688980957
transform 1 0 43608 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_473
timestamp 1688980957
transform 1 0 43976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_477
timestamp 1688980957
transform 1 0 44344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_481
timestamp 1688980957
transform 1 0 44712 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_485
timestamp 1688980957
transform 1 0 45080 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 736 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 1840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 2944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_35
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_39
timestamp 1688980957
transform 1 0 4048 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_43
timestamp 1688980957
transform 1 0 4416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_67
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_72
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_76
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_80
timestamp 1688980957
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_146
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_150
timestamp 1688980957
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 18400 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_280
timestamp 1688980957
transform 1 0 26220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_284
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_288
timestamp 1688980957
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_323
timestamp 1688980957
transform 1 0 30176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_327
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 33856 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_403
timestamp 1688980957
transform 1 0 37536 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_470
timestamp 1688980957
transform 1 0 43700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_474
timestamp 1688980957
transform 1 0 44068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_481
timestamp 1688980957
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_485
timestamp 1688980957
transform 1 0 45080 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 736 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_27
timestamp 1688980957
transform 1 0 2944 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_33
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_64
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_73
timestamp 1688980957
transform 1 0 7176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_79
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_85
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_98
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_108
timestamp 1688980957
transform 1 0 10396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_153
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_188
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_220
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_229
timestamp 1688980957
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_232
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_236
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_276
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_355
timestamp 1688980957
transform 1 0 33120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_359
timestamp 1688980957
transform 1 0 33488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_363
timestamp 1688980957
transform 1 0 33856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_367
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_389
timestamp 1688980957
transform 1 0 36248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_396
timestamp 1688980957
transform 1 0 36892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_400
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_404
timestamp 1688980957
transform 1 0 37628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_434
timestamp 1688980957
transform 1 0 40388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_458
timestamp 1688980957
transform 1 0 42596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_462
timestamp 1688980957
transform 1 0 42964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_466
timestamp 1688980957
transform 1 0 43332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_470
timestamp 1688980957
transform 1 0 43700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_474
timestamp 1688980957
transform 1 0 44068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_478
timestamp 1688980957
transform 1 0 44436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_482
timestamp 1688980957
transform 1 0 44804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_486
timestamp 1688980957
transform 1 0 45172 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 736 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 1840 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_92
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_103
timestamp 1688980957
transform 1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_109
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_122
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_135
timestamp 1688980957
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16192 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_177
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_191
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_205
timestamp 1688980957
transform 1 0 19320 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_209
timestamp 1688980957
transform 1 0 19688 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_227
timestamp 1688980957
transform 1 0 21344 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_231
timestamp 1688980957
transform 1 0 21712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_236
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_262
timestamp 1688980957
transform 1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_329
timestamp 1688980957
transform 1 0 30728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_369
timestamp 1688980957
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_379
timestamp 1688980957
transform 1 0 35328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_392
timestamp 1688980957
transform 1 0 36524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_396
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_418
timestamp 1688980957
transform 1 0 38916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_430
timestamp 1688980957
transform 1 0 40020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_466
timestamp 1688980957
transform 1 0 43332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_470
timestamp 1688980957
transform 1 0 43700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_474
timestamp 1688980957
transform 1 0 44068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_477
timestamp 1688980957
transform 1 0 44344 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_481
timestamp 1688980957
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_485
timestamp 1688980957
transform 1 0 45080 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 736 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 1688980957
transform 1 0 2944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_35
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_108
timestamp 1688980957
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp 1688980957
transform 1 0 10856 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11224 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_132
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_138
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18216 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1688980957
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_234
timestamp 1688980957
transform 1 0 21988 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_275
timestamp 1688980957
transform 1 0 25760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26128 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26312 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_344
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_371
timestamp 1688980957
transform 1 0 34592 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_393
timestamp 1688980957
transform 1 0 36616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_434
timestamp 1688980957
transform 1 0 40388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_469
timestamp 1688980957
transform 1 0 43608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_473
timestamp 1688980957
transform 1 0 43976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_477
timestamp 1688980957
transform 1 0 44344 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_481
timestamp 1688980957
transform 1 0 44712 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_485
timestamp 1688980957
transform 1 0 45080 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 736 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 2944 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3128 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_49
timestamp 1688980957
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_58
timestamp 1688980957
transform 1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_76
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_135
timestamp 1688980957
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_177
timestamp 1688980957
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_200
timestamp 1688980957
transform 1 0 18860 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_239
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 28704 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_309
timestamp 1688980957
transform 1 0 28888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_313
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_324
timestamp 1688980957
transform 1 0 30268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_418
timestamp 1688980957
transform 1 0 38916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_462
timestamp 1688980957
transform 1 0 42964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_466
timestamp 1688980957
transform 1 0 43332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_470
timestamp 1688980957
transform 1 0 43700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_474
timestamp 1688980957
transform 1 0 44068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_477
timestamp 1688980957
transform 1 0 44344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_481
timestamp 1688980957
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_485
timestamp 1688980957
transform 1 0 45080 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 736 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 1840 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 2944 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4048 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1688980957
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_61
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_65
timestamp 1688980957
transform 1 0 6440 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_69
timestamp 1688980957
transform 1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_73
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_80
timestamp 1688980957
transform 1 0 7820 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_84
timestamp 1688980957
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 10672 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_133
timestamp 1688980957
transform 1 0 12696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_155
timestamp 1688980957
transform 1 0 14720 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_195
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_231
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_235
timestamp 1688980957
transform 1 0 22080 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_239
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_263
timestamp 1688980957
transform 1 0 24656 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_276
timestamp 1688980957
transform 1 0 25852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_285
timestamp 1688980957
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_289
timestamp 1688980957
transform 1 0 27048 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_305
timestamp 1688980957
transform 1 0 28520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_311
timestamp 1688980957
transform 1 0 29072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_328
timestamp 1688980957
transform 1 0 30636 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_368
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 36432 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_393
timestamp 1688980957
transform 1 0 36616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_420
timestamp 1688980957
transform 1 0 39100 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 41584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_467
timestamp 1688980957
transform 1 0 43424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_471
timestamp 1688980957
transform 1 0 43792 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_475
timestamp 1688980957
transform 1 0 44160 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_479
timestamp 1688980957
transform 1 0 44528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_483
timestamp 1688980957
transform 1 0 44896 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 736 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 2944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3128 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_39
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_45
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_48
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_52
timestamp 1688980957
transform 1 0 5244 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_56
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_60
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_64
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_68
timestamp 1688980957
transform 1 0 6716 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_72
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_76
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_80
timestamp 1688980957
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_89
timestamp 1688980957
transform 1 0 8648 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_92
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_99
timestamp 1688980957
transform 1 0 9568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_127
timestamp 1688980957
transform 1 0 12144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_132
timestamp 1688980957
transform 1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_136
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1688980957
transform 1 0 13432 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_147
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_158
timestamp 1688980957
transform 1 0 14996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_180
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_208
timestamp 1688980957
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_224
timestamp 1688980957
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_228
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_236
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_240
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_244
timestamp 1688980957
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_248
timestamp 1688980957
transform 1 0 23276 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_262
timestamp 1688980957
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_274
timestamp 1688980957
transform 1 0 25668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_278
timestamp 1688980957
transform 1 0 26036 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 28704 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_336
timestamp 1688980957
transform 1 0 31372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_359
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 33856 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_371
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_375
timestamp 1688980957
transform 1 0 34960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_386
timestamp 1688980957
transform 1 0 35972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_390
timestamp 1688980957
transform 1 0 36340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_414
timestamp 1688980957
transform 1 0 38548 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_418
timestamp 1688980957
transform 1 0 38916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_474
timestamp 1688980957
transform 1 0 44068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44344 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_481
timestamp 1688980957
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_485
timestamp 1688980957
transform 1 0 45080 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 736 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_35
timestamp 1688980957
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_61
timestamp 1688980957
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_65
timestamp 1688980957
transform 1 0 6440 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_69
timestamp 1688980957
transform 1 0 6808 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_72
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_76
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_80
timestamp 1688980957
transform 1 0 7820 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_84
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_88
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_92
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_96
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_100
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_104
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_108
timestamp 1688980957
transform 1 0 10396 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_113
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_117
timestamp 1688980957
transform 1 0 11224 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_120
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_124
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_128
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_132
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_136
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_140
timestamp 1688980957
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_144
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_213
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_243
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_247
timestamp 1688980957
transform 1 0 23184 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_259
timestamp 1688980957
transform 1 0 24288 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_272
timestamp 1688980957
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_276
timestamp 1688980957
transform 1 0 25852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_348
timestamp 1688980957
transform 1 0 32476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_379
timestamp 1688980957
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_402
timestamp 1688980957
transform 1 0 37444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_423
timestamp 1688980957
transform 1 0 39376 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_446
timestamp 1688980957
transform 1 0 41492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_461
timestamp 1688980957
transform 1 0 42872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_465
timestamp 1688980957
transform 1 0 43240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_469
timestamp 1688980957
transform 1 0 43608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_473
timestamp 1688980957
transform 1 0 43976 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_477
timestamp 1688980957
transform 1 0 44344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_481
timestamp 1688980957
transform 1 0 44712 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_485
timestamp 1688980957
transform 1 0 45080 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_6
timestamp 1688980957
transform 1 0 1012 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_18
timestamp 1688980957
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_37
timestamp 1688980957
transform 1 0 3864 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_49
timestamp 1688980957
transform 1 0 4968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5336 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_56
timestamp 1688980957
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_60
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 8648 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_112
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_116
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_120
timestamp 1688980957
transform 1 0 11500 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_124
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_128
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_132
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_136
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1688980957
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_145
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_149
timestamp 1688980957
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 23460 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_273
timestamp 1688980957
transform 1 0 25576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_338
timestamp 1688980957
transform 1 0 31556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_459
timestamp 1688980957
transform 1 0 42688 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_463
timestamp 1688980957
transform 1 0 43056 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_467
timestamp 1688980957
transform 1 0 43424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_471
timestamp 1688980957
transform 1 0 43792 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_475
timestamp 1688980957
transform 1 0 44160 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_477
timestamp 1688980957
transform 1 0 44344 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 736 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 1840 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 2944 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 5520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_57
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_62
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_66
timestamp 1688980957
transform 1 0 6532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_70
timestamp 1688980957
transform 1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_74
timestamp 1688980957
transform 1 0 7268 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_78
timestamp 1688980957
transform 1 0 7636 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_82
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_86
timestamp 1688980957
transform 1 0 8372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_90
timestamp 1688980957
transform 1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_94
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_98
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_102
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_106
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_117
timestamp 1688980957
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_121
timestamp 1688980957
transform 1 0 11592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_125
timestamp 1688980957
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_129
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_133
timestamp 1688980957
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_141
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 15732 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_186
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_207
timestamp 1688980957
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_229
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_305
timestamp 1688980957
transform 1 0 28520 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1688980957
transform 1 0 31188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_442
timestamp 1688980957
transform 1 0 41124 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_446
timestamp 1688980957
transform 1 0 41492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_449
timestamp 1688980957
transform 1 0 41768 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_453
timestamp 1688980957
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_457
timestamp 1688980957
transform 1 0 42504 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_461
timestamp 1688980957
transform 1 0 42872 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_465
timestamp 1688980957
transform 1 0 43240 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_469
timestamp 1688980957
transform 1 0 43608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_473
timestamp 1688980957
transform 1 0 43976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_477
timestamp 1688980957
transform 1 0 44344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_481
timestamp 1688980957
transform 1 0 44712 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_485
timestamp 1688980957
transform 1 0 45080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_3
timestamp 1688980957
transform 1 0 736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_13
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_20
timestamp 1688980957
transform 1 0 2300 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_24
timestamp 1688980957
transform 1 0 2668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_33
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_40
timestamp 1688980957
transform 1 0 4140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_44
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_48
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_52
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1688980957
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_61
timestamp 1688980957
transform 1 0 6072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_68
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_77
timestamp 1688980957
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_81
timestamp 1688980957
transform 1 0 7912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_88
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9016 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_100
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_108
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_116
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_120
timestamp 1688980957
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_126
timestamp 1688980957
transform 1 0 12052 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_130
timestamp 1688980957
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_141
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_145
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_185
timestamp 1688980957
transform 1 0 17480 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_189
timestamp 1688980957
transform 1 0 17848 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_207
timestamp 1688980957
transform 1 0 19504 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_238
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_253
timestamp 1688980957
transform 1 0 23736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_269
timestamp 1688980957
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_313
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_327
timestamp 1688980957
transform 1 0 30544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_385
timestamp 1688980957
transform 1 0 35880 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_415
timestamp 1688980957
transform 1 0 38640 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 1688980957
transform 1 0 39008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_430
timestamp 1688980957
transform 1 0 40020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_434
timestamp 1688980957
transform 1 0 40388 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_438
timestamp 1688980957
transform 1 0 40756 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_442
timestamp 1688980957
transform 1 0 41124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_446
timestamp 1688980957
transform 1 0 41492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_450
timestamp 1688980957
transform 1 0 41860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_454
timestamp 1688980957
transform 1 0 42228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_458
timestamp 1688980957
transform 1 0 42596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_462
timestamp 1688980957
transform 1 0 42964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_466
timestamp 1688980957
transform 1 0 43332 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_470
timestamp 1688980957
transform 1 0 43700 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_474
timestamp 1688980957
transform 1 0 44068 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_477
timestamp 1688980957
transform 1 0 44344 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_481
timestamp 1688980957
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_485
timestamp 1688980957
transform 1 0 45080 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_3
timestamp 1688980957
transform 1 0 736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_9
timestamp 1688980957
transform 1 0 1288 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_19
timestamp 1688980957
transform 1 0 2208 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_27
timestamp 1688980957
transform 1 0 2944 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4048 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_49
timestamp 1688980957
transform 1 0 4968 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 5520 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_63
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_69
timestamp 1688980957
transform 1 0 6808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_79
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_91
timestamp 1688980957
transform 1 0 8832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_99
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1688980957
transform 1 0 10488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_113
timestamp 1688980957
transform 1 0 10856 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_121
timestamp 1688980957
transform 1 0 11592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_129
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_139
timestamp 1688980957
transform 1 0 13248 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_141
timestamp 1688980957
transform 1 0 13432 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_151
timestamp 1688980957
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_159
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_179
timestamp 1688980957
transform 1 0 16928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_189
timestamp 1688980957
transform 1 0 17848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18216 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_201
timestamp 1688980957
transform 1 0 18952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_209
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_219
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_232
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_241
timestamp 1688980957
transform 1 0 22632 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_249
timestamp 1688980957
transform 1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_253
timestamp 1688980957
transform 1 0 23736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_259
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_269
timestamp 1688980957
transform 1 0 25208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_274
timestamp 1688980957
transform 1 0 25668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26128 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_284
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_292
timestamp 1688980957
transform 1 0 27324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_303
timestamp 1688980957
transform 1 0 28336 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31280 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_380
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1688980957
transform 1 0 36340 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_424
timestamp 1688980957
transform 1 0 39468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_428
timestamp 1688980957
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_432
timestamp 1688980957
transform 1 0 40204 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_438
timestamp 1688980957
transform 1 0 40756 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_442
timestamp 1688980957
transform 1 0 41124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_449
timestamp 1688980957
transform 1 0 41768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_453
timestamp 1688980957
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_458
timestamp 1688980957
transform 1 0 42596 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_462
timestamp 1688980957
transform 1 0 42964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_468
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_472
timestamp 1688980957
transform 1 0 43884 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_480
timestamp 1688980957
transform 1 0 44620 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43424 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 44988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 33396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 40480 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 41400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 43240 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 44344 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 44988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 36156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 36616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 36892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 38456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 33672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 38548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 40664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 40572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 40848 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 41124 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 41400 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 41768 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 42504 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 43332 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 33396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 44344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 35144 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 35788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 37720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 39192 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 39560 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  input36
timestamp 1688980957
transform 1 0 43424 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 736 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 736 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  Inst_bitbang._181_
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  Inst_bitbang._182_
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  Inst_bitbang._183_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  Inst_bitbang._184_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_4  Inst_bitbang._185_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_4  Inst_bitbang._186_
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  Inst_bitbang._187_
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  Inst_bitbang._188_
timestamp 1688980957
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._189_
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  Inst_bitbang._190_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  Inst_bitbang._191_
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  Inst_bitbang._192_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  Inst_bitbang._193_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._194_
timestamp 1688980957
transform 1 0 25392 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._195_
timestamp 1688980957
transform 1 0 23368 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._196_
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._197_
timestamp 1688980957
transform 1 0 26312 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._198_
timestamp 1688980957
transform 1 0 31464 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._199_
timestamp 1688980957
transform 1 0 33120 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._200_
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._201_
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._202_
timestamp 1688980957
transform 1 0 35144 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._203_
timestamp 1688980957
transform 1 0 33672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._204_
timestamp 1688980957
transform 1 0 35328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._205_
timestamp 1688980957
transform 1 0 35052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._206_
timestamp 1688980957
transform 1 0 35696 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._207_
timestamp 1688980957
transform 1 0 35972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._208_
timestamp 1688980957
transform 1 0 37720 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._209_
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  Inst_bitbang._210_
timestamp 1688980957
transform 1 0 41124 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._211_
timestamp 1688980957
transform 1 0 37996 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._212_
timestamp 1688980957
transform 1 0 38548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._213_
timestamp 1688980957
transform 1 0 38088 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._214_
timestamp 1688980957
transform 1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._215_
timestamp 1688980957
transform 1 0 41032 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._216_
timestamp 1688980957
transform 1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._217_
timestamp 1688980957
transform 1 0 41768 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._218_
timestamp 1688980957
transform 1 0 40112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._219_
timestamp 1688980957
transform 1 0 41768 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._220_
timestamp 1688980957
transform 1 0 42596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._221_
timestamp 1688980957
transform 1 0 41860 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._222_
timestamp 1688980957
transform 1 0 42688 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._223_
timestamp 1688980957
transform 1 0 41768 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._224_
timestamp 1688980957
transform 1 0 41400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._225_
timestamp 1688980957
transform 1 0 41676 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._226_
timestamp 1688980957
transform 1 0 42964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._227_
timestamp 1688980957
transform 1 0 38916 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._228_
timestamp 1688980957
transform 1 0 37260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._229_
timestamp 1688980957
transform 1 0 37536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._230_
timestamp 1688980957
transform 1 0 36984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  Inst_bitbang._231_
timestamp 1688980957
transform 1 0 37904 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._232_
timestamp 1688980957
transform 1 0 35512 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._233_
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._234_
timestamp 1688980957
transform 1 0 35512 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._235_
timestamp 1688980957
transform 1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._236_
timestamp 1688980957
transform 1 0 37076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._237_
timestamp 1688980957
transform 1 0 36616 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._238_
timestamp 1688980957
transform 1 0 35052 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._239_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._240_
timestamp 1688980957
transform 1 0 34776 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._241_
timestamp 1688980957
transform 1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._242_
timestamp 1688980957
transform 1 0 37720 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._243_
timestamp 1688980957
transform 1 0 40020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._244_
timestamp 1688980957
transform 1 0 40020 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._245_
timestamp 1688980957
transform 1 0 40296 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._246_
timestamp 1688980957
transform 1 0 39192 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._247_
timestamp 1688980957
transform 1 0 40940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._248_
timestamp 1688980957
transform 1 0 40020 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._249_
timestamp 1688980957
transform 1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._250_
timestamp 1688980957
transform 1 0 39192 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._251_
timestamp 1688980957
transform 1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._252_
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._253_
timestamp 1688980957
transform 1 0 37260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._254_
timestamp 1688980957
transform 1 0 41768 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._255_
timestamp 1688980957
transform 1 0 41308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._256_
timestamp 1688980957
transform 1 0 41768 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._257_
timestamp 1688980957
transform 1 0 41032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._258_
timestamp 1688980957
transform 1 0 41492 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._259_
timestamp 1688980957
transform 1 0 41216 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  Inst_bitbang._260_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  Inst_bitbang._261_
timestamp 1688980957
transform 1 0 37812 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._262_
timestamp 1688980957
transform 1 0 23460 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._263_
timestamp 1688980957
transform 1 0 23184 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._264_
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._265_
timestamp 1688980957
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._266_
timestamp 1688980957
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._267_
timestamp 1688980957
transform 1 0 25576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._268_
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._269_
timestamp 1688980957
transform 1 0 32568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._270_
timestamp 1688980957
transform 1 0 33672 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._271_
timestamp 1688980957
transform 1 0 33396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._272_
timestamp 1688980957
transform 1 0 34500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._273_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._274_
timestamp 1688980957
transform 1 0 35696 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._275_
timestamp 1688980957
transform 1 0 36156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._276_
timestamp 1688980957
transform 1 0 36616 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._277_
timestamp 1688980957
transform 1 0 36248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._278_
timestamp 1688980957
transform 1 0 36616 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._279_
timestamp 1688980957
transform 1 0 37444 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._280_
timestamp 1688980957
transform 1 0 37444 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._281_
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  Inst_bitbang._282_
timestamp 1688980957
transform 1 0 40112 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._283_
timestamp 1688980957
transform 1 0 39560 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._284_
timestamp 1688980957
transform 1 0 38364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._285_
timestamp 1688980957
transform 1 0 39560 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._286_
timestamp 1688980957
transform 1 0 41032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._287_
timestamp 1688980957
transform 1 0 41032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._288_
timestamp 1688980957
transform 1 0 41308 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._289_
timestamp 1688980957
transform 1 0 40848 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._290_
timestamp 1688980957
transform 1 0 40572 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._291_
timestamp 1688980957
transform 1 0 40848 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._292_
timestamp 1688980957
transform 1 0 40572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._293_
timestamp 1688980957
transform 1 0 41308 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._294_
timestamp 1688980957
transform 1 0 41032 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._295_
timestamp 1688980957
transform 1 0 41124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._296_
timestamp 1688980957
transform 1 0 41768 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._297_
timestamp 1688980957
transform 1 0 39744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._298_
timestamp 1688980957
transform 1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._299_
timestamp 1688980957
transform 1 0 36800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._300_
timestamp 1688980957
transform 1 0 38548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._301_
timestamp 1688980957
transform 1 0 36984 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._302_
timestamp 1688980957
transform 1 0 36708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  Inst_bitbang._303_
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._304_
timestamp 1688980957
transform 1 0 36340 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._305_
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._306_
timestamp 1688980957
transform 1 0 36708 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._307_
timestamp 1688980957
transform 1 0 34408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._308_
timestamp 1688980957
transform 1 0 34960 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._309_
timestamp 1688980957
transform 1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._310_
timestamp 1688980957
transform 1 0 34132 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._311_
timestamp 1688980957
transform 1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._312_
timestamp 1688980957
transform 1 0 36800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._313_
timestamp 1688980957
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._314_
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._315_
timestamp 1688980957
transform 1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._316_
timestamp 1688980957
transform 1 0 39928 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._317_
timestamp 1688980957
transform 1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._318_
timestamp 1688980957
transform 1 0 39560 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._319_
timestamp 1688980957
transform 1 0 38180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._320_
timestamp 1688980957
transform 1 0 40756 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._321_
timestamp 1688980957
transform 1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._322_
timestamp 1688980957
transform 1 0 39008 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._323_
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._324_
timestamp 1688980957
transform 1 0 40112 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._325_
timestamp 1688980957
transform 1 0 39376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._326_
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._327_
timestamp 1688980957
transform 1 0 39560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  Inst_bitbang._328_
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  Inst_bitbang._329_
timestamp 1688980957
transform 1 0 10120 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._330_
timestamp 1688980957
transform 1 0 10856 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._331_
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._332_
timestamp 1688980957
transform 1 0 12328 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._333_
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._334_
timestamp 1688980957
transform 1 0 11500 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._335_
timestamp 1688980957
transform 1 0 10304 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._336_
timestamp 1688980957
transform 1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._337_
timestamp 1688980957
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._338_
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._339_
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._340_
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._341_
timestamp 1688980957
transform 1 0 8280 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._342_
timestamp 1688980957
transform 1 0 7360 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._343_
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._344_
timestamp 1688980957
transform 1 0 9568 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._345_
timestamp 1688980957
transform 1 0 7636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._346_
timestamp 1688980957
transform 1 0 7360 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._347_
timestamp 1688980957
transform 1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._348_
timestamp 1688980957
transform 1 0 9476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._349_
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._350_
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._351_
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._352_
timestamp 1688980957
transform 1 0 10672 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._353_
timestamp 1688980957
transform 1 0 10488 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._354_
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._355_
timestamp 1688980957
transform 1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._356_
timestamp 1688980957
transform 1 0 12512 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._357_
timestamp 1688980957
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._358_
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._359_
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  Inst_bitbang._360_
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Inst_bitbang._361_
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._362_
timestamp 1688980957
transform 1 0 15088 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  Inst_bitbang._363_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._364_
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._365_
timestamp 1688980957
transform 1 0 15088 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._366_
timestamp 1688980957
transform 1 0 23736 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._367_
timestamp 1688980957
transform 1 0 26312 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._368_
timestamp 1688980957
transform 1 0 30728 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._369_
timestamp 1688980957
transform 1 0 33304 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._370_
timestamp 1688980957
transform 1 0 34040 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._371_
timestamp 1688980957
transform 1 0 34684 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._372_
timestamp 1688980957
transform 1 0 36616 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._373_
timestamp 1688980957
transform 1 0 35880 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._374_
timestamp 1688980957
transform 1 0 37536 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._375_
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._376_
timestamp 1688980957
transform 1 0 39192 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._377_
timestamp 1688980957
transform 1 0 39652 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._378_
timestamp 1688980957
transform 1 0 42228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._379_
timestamp 1688980957
transform 1 0 41768 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._380_
timestamp 1688980957
transform 1 0 41768 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._381_
timestamp 1688980957
transform 1 0 41768 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._382_
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._383_
timestamp 1688980957
transform 1 0 36708 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._384_
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._385_
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._386_
timestamp 1688980957
transform 1 0 34684 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._387_
timestamp 1688980957
transform 1 0 34132 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._388_
timestamp 1688980957
transform 1 0 33856 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._389_
timestamp 1688980957
transform 1 0 36616 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._390_
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._391_
timestamp 1688980957
transform 1 0 38824 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._392_
timestamp 1688980957
transform 1 0 39192 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._393_
timestamp 1688980957
transform 1 0 39192 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._394_
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._395_
timestamp 1688980957
transform 1 0 41032 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._396_
timestamp 1688980957
transform 1 0 41032 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._397_
timestamp 1688980957
transform 1 0 41768 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._398_
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._399_
timestamp 1688980957
transform 1 0 23552 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._400_
timestamp 1688980957
transform 1 0 25300 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._401_
timestamp 1688980957
transform 1 0 31464 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._402_
timestamp 1688980957
transform 1 0 34040 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._403_
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._404_
timestamp 1688980957
transform 1 0 36248 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._405_
timestamp 1688980957
transform 1 0 35972 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._406_
timestamp 1688980957
transform 1 0 38456 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._407_
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._408_
timestamp 1688980957
transform 1 0 39192 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._409_
timestamp 1688980957
transform 1 0 39192 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._410_
timestamp 1688980957
transform 1 0 40388 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._411_
timestamp 1688980957
transform 1 0 40664 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._412_
timestamp 1688980957
transform 1 0 41032 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._413_
timestamp 1688980957
transform 1 0 39836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._414_
timestamp 1688980957
transform 1 0 40480 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._415_
timestamp 1688980957
transform 1 0 38456 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._416_
timestamp 1688980957
transform 1 0 36616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._417_
timestamp 1688980957
transform 1 0 35144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._418_
timestamp 1688980957
transform 1 0 35236 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._419_
timestamp 1688980957
transform 1 0 34040 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._420_
timestamp 1688980957
transform 1 0 34040 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._421_
timestamp 1688980957
transform 1 0 35880 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._422_
timestamp 1688980957
transform 1 0 36616 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._423_
timestamp 1688980957
transform 1 0 38456 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._424_
timestamp 1688980957
transform 1 0 38088 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._425_
timestamp 1688980957
transform 1 0 37720 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._426_
timestamp 1688980957
transform 1 0 38916 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._427_
timestamp 1688980957
transform 1 0 39192 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._428_
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._429_
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._430_
timestamp 1688980957
transform 1 0 1840 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._431_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._432_
timestamp 1688980957
transform 1 0 6348 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._433_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._434_
timestamp 1688980957
transform 1 0 1748 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._435_
timestamp 1688980957
transform 1 0 3772 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  Inst_bitbang._436_
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._437_
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._438_
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._439_
timestamp 1688980957
transform 1 0 10580 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._440_
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._441_
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._442_
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._443_
timestamp 1688980957
transform 1 0 7728 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._444_
timestamp 1688980957
transform 1 0 8280 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._445_
timestamp 1688980957
transform 1 0 8280 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._446_
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._447_
timestamp 1688980957
transform 1 0 8740 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._448_
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._449_
timestamp 1688980957
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._450_
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._451_
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._452_
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  Inst_bitbang._453_
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0589_
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0590_
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._0591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0592_
timestamp 1688980957
transform 1 0 20516 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0593_
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0594_
timestamp 1688980957
transform 1 0 19320 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0595_
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0596_
timestamp 1688980957
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  INST_config_UART._0597_
timestamp 1688980957
transform 1 0 21896 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._0598_
timestamp 1688980957
transform 1 0 17940 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0599_
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0600_
timestamp 1688980957
transform 1 0 32292 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0601_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35972 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0602_
timestamp 1688980957
transform 1 0 34868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  INST_config_UART._0603_
timestamp 1688980957
transform 1 0 35328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  INST_config_UART._0604_
timestamp 1688980957
transform 1 0 39100 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  INST_config_UART._0605_
timestamp 1688980957
transform 1 0 39744 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0606_
timestamp 1688980957
transform 1 0 37720 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0607_
timestamp 1688980957
transform 1 0 40296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  INST_config_UART._0608_
timestamp 1688980957
transform 1 0 36708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0609_
timestamp 1688980957
transform 1 0 37720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  INST_config_UART._0610_
timestamp 1688980957
transform 1 0 36984 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  INST_config_UART._0611_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33304 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0612_
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  INST_config_UART._0613_
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  INST_config_UART._0614_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18584 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0615_
timestamp 1688980957
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  INST_config_UART._0616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0617_
timestamp 1688980957
transform 1 0 29716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._0618_
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0619_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0620_
timestamp 1688980957
transform 1 0 18584 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0621_
timestamp 1688980957
transform 1 0 17664 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  INST_config_UART._0622_
timestamp 1688980957
transform 1 0 24012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  INST_config_UART._0623_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0624_
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0625_
timestamp 1688980957
transform 1 0 23552 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0626_
timestamp 1688980957
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0627_
timestamp 1688980957
transform 1 0 24564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0628_
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  INST_config_UART._0629_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0630_
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  INST_config_UART._0631_
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  INST_config_UART._0632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._0633_
timestamp 1688980957
transform 1 0 23092 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0634_
timestamp 1688980957
transform 1 0 23736 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  INST_config_UART._0635_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o311ai_4  INST_config_UART._0636_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_2  INST_config_UART._0637_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21988 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  INST_config_UART._0638_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  INST_config_UART._0639_
timestamp 1688980957
transform 1 0 28888 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._0640_
timestamp 1688980957
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0641_
timestamp 1688980957
transform 1 0 29716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  INST_config_UART._0642_
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._0643_
timestamp 1688980957
transform 1 0 30544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0644_
timestamp 1688980957
transform 1 0 30084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0645_
timestamp 1688980957
transform 1 0 28520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._0646_
timestamp 1688980957
transform 1 0 29624 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0647_
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  INST_config_UART._0648_
timestamp 1688980957
transform 1 0 28152 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0649_
timestamp 1688980957
transform 1 0 28428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0650_
timestamp 1688980957
transform 1 0 17848 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0651_
timestamp 1688980957
transform 1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0652_
timestamp 1688980957
transform 1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0653_
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0654_
timestamp 1688980957
transform 1 0 19320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  INST_config_UART._0655_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0656_
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0657_
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0658_
timestamp 1688980957
transform 1 0 22816 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0659_
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0660_
timestamp 1688980957
transform 1 0 27324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0661_
timestamp 1688980957
transform 1 0 27968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0662_
timestamp 1688980957
transform 1 0 26312 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0663_
timestamp 1688980957
transform 1 0 26956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  INST_config_UART._0664_
timestamp 1688980957
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0665_
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0666_
timestamp 1688980957
transform 1 0 21344 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0667_
timestamp 1688980957
transform 1 0 18676 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0668_
timestamp 1688980957
transform 1 0 17480 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0669_
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0670_
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0671_
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0672_
timestamp 1688980957
transform 1 0 17296 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0673_
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0674_
timestamp 1688980957
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0675_
timestamp 1688980957
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0676_
timestamp 1688980957
transform 1 0 20424 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0677_
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  INST_config_UART._0678_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0679_
timestamp 1688980957
transform 1 0 18584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0680_
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0681_
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._0682_
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0683_
timestamp 1688980957
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0684_
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0685_
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0686_
timestamp 1688980957
transform 1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0687_
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0688_
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0689_
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._0690_
timestamp 1688980957
transform 1 0 16928 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0691_
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0692_
timestamp 1688980957
transform 1 0 14904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0693_
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0694_
timestamp 1688980957
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0695_
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0696_
timestamp 1688980957
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0697_
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0698_
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0699_
timestamp 1688980957
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0700_
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0701_
timestamp 1688980957
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0702_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0703_
timestamp 1688980957
transform 1 0 16744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0704_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0705_
timestamp 1688980957
transform 1 0 19320 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0706_
timestamp 1688980957
transform 1 0 20148 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0707_
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0708_
timestamp 1688980957
transform 1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0709_
timestamp 1688980957
transform 1 0 3864 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0710_
timestamp 1688980957
transform 1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0711_
timestamp 1688980957
transform 1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0712_
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0713_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0714_
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0715_
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0716_
timestamp 1688980957
transform 1 0 4784 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0717_
timestamp 1688980957
transform 1 0 5336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0718_
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0719_
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0720_
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0721_
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0722_
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0723_
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  INST_config_UART._0724_
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0725_
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0726_
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0727_
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  INST_config_UART._0728_
timestamp 1688980957
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0729_
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0730_
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0731_
timestamp 1688980957
transform 1 0 4048 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0732_
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0733_
timestamp 1688980957
transform 1 0 3496 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0734_
timestamp 1688980957
transform 1 0 4324 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0735_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  INST_config_UART._0736_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0737_
timestamp 1688980957
transform 1 0 5520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0738_
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0739_
timestamp 1688980957
transform 1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0740_
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0741_
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0742_
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0743_
timestamp 1688980957
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0744_
timestamp 1688980957
transform 1 0 7544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0745_
timestamp 1688980957
transform 1 0 7544 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0746_
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0747_
timestamp 1688980957
transform 1 0 9108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0748_
timestamp 1688980957
transform 1 0 9292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0749_
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0750_
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0751_
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0752_
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0753_
timestamp 1688980957
transform 1 0 11868 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0754_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0755_
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._0756_
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0757_
timestamp 1688980957
transform 1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0758_
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0759_
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0760_
timestamp 1688980957
transform 1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0761_
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0762_
timestamp 1688980957
transform 1 0 20332 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0763_
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0764_
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0765_
timestamp 1688980957
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0766_
timestamp 1688980957
transform 1 0 28612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0767_
timestamp 1688980957
transform 1 0 28888 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0768_
timestamp 1688980957
transform 1 0 27324 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0769_
timestamp 1688980957
transform 1 0 27140 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0770_
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0771_
timestamp 1688980957
transform 1 0 28060 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0772_
timestamp 1688980957
transform 1 0 27324 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  INST_config_UART._0773_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28612 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0774_
timestamp 1688980957
transform 1 0 28152 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0775_
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0776_
timestamp 1688980957
transform 1 0 27600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0777_
timestamp 1688980957
transform 1 0 31464 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0778_
timestamp 1688980957
transform 1 0 29716 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0779_
timestamp 1688980957
transform 1 0 30176 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0780_
timestamp 1688980957
transform 1 0 30728 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0781_
timestamp 1688980957
transform 1 0 28336 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0782_
timestamp 1688980957
transform 1 0 27784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0783_
timestamp 1688980957
transform 1 0 29992 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0784_
timestamp 1688980957
transform 1 0 28612 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0785_
timestamp 1688980957
transform 1 0 29440 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0786_
timestamp 1688980957
transform 1 0 29348 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0787_
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._0788_
timestamp 1688980957
transform 1 0 28888 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._0789_
timestamp 1688980957
transform 1 0 29624 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0790_
timestamp 1688980957
transform 1 0 33764 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0791_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0792_
timestamp 1688980957
transform 1 0 31464 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0793_
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0794_
timestamp 1688980957
transform 1 0 30360 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0795_
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0796_
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0797_
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0798_
timestamp 1688980957
transform 1 0 30820 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0799_
timestamp 1688980957
transform 1 0 28152 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0800_
timestamp 1688980957
transform 1 0 30084 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0801_
timestamp 1688980957
transform 1 0 30728 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  INST_config_UART._0802_
timestamp 1688980957
transform 1 0 31832 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0803_
timestamp 1688980957
transform 1 0 36616 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0804_
timestamp 1688980957
transform 1 0 30728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0805_
timestamp 1688980957
transform 1 0 35696 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0806_
timestamp 1688980957
transform 1 0 30544 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0807_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0808_
timestamp 1688980957
transform 1 0 30544 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0809_
timestamp 1688980957
transform 1 0 33396 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0810_
timestamp 1688980957
transform 1 0 30820 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0811_
timestamp 1688980957
transform 1 0 32292 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0812_
timestamp 1688980957
transform 1 0 34132 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0813_
timestamp 1688980957
transform 1 0 33672 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0814_
timestamp 1688980957
transform 1 0 30912 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0815_
timestamp 1688980957
transform 1 0 31464 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0816_
timestamp 1688980957
transform 1 0 32660 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0817_
timestamp 1688980957
transform 1 0 30728 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0818_
timestamp 1688980957
transform 1 0 30912 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0819_
timestamp 1688980957
transform 1 0 31280 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0820_
timestamp 1688980957
transform 1 0 30452 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0821_
timestamp 1688980957
transform 1 0 32660 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0822_
timestamp 1688980957
transform 1 0 30912 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0823_
timestamp 1688980957
transform 1 0 32752 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  INST_config_UART._0824_
timestamp 1688980957
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0825_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0826_
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._0827_
timestamp 1688980957
transform 1 0 24840 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0828_
timestamp 1688980957
transform 1 0 21252 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0829_
timestamp 1688980957
transform 1 0 25024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0830_
timestamp 1688980957
transform 1 0 20424 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0831_
timestamp 1688980957
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0832_
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0833_
timestamp 1688980957
transform 1 0 20424 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0834_
timestamp 1688980957
transform 1 0 19596 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0835_
timestamp 1688980957
transform 1 0 34684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0836_
timestamp 1688980957
transform 1 0 38088 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0837_
timestamp 1688980957
transform 1 0 35880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0838_
timestamp 1688980957
transform 1 0 37260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0839_
timestamp 1688980957
transform 1 0 36156 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0840_
timestamp 1688980957
transform 1 0 38272 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0841_
timestamp 1688980957
transform 1 0 37168 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0842_
timestamp 1688980957
transform 1 0 39192 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0843_
timestamp 1688980957
transform 1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0844_
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0845_
timestamp 1688980957
transform 1 0 37536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0846_
timestamp 1688980957
transform 1 0 39192 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0847_
timestamp 1688980957
transform 1 0 38548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0848_
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0849_
timestamp 1688980957
transform 1 0 36616 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0850_
timestamp 1688980957
transform 1 0 35880 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0851_
timestamp 1688980957
transform 1 0 35052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0852_
timestamp 1688980957
transform 1 0 22816 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0853_
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0854_
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0855_
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0856_
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0857_
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0858_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0859_
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0860_
timestamp 1688980957
transform 1 0 21252 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0861_
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._0862_
timestamp 1688980957
transform 1 0 21252 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0863_
timestamp 1688980957
transform 1 0 21988 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0864_
timestamp 1688980957
transform 1 0 19596 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0865_
timestamp 1688980957
transform 1 0 34868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0866_
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0867_
timestamp 1688980957
transform 1 0 33672 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0868_
timestamp 1688980957
transform 1 0 35144 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0869_
timestamp 1688980957
transform 1 0 33396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0870_
timestamp 1688980957
transform 1 0 38088 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0871_
timestamp 1688980957
transform 1 0 37812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0872_
timestamp 1688980957
transform 1 0 38272 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0873_
timestamp 1688980957
transform 1 0 40020 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0874_
timestamp 1688980957
transform 1 0 41768 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0875_
timestamp 1688980957
transform 1 0 41124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0876_
timestamp 1688980957
transform 1 0 38916 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0877_
timestamp 1688980957
transform 1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0878_
timestamp 1688980957
transform 1 0 35696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0879_
timestamp 1688980957
transform 1 0 36064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0880_
timestamp 1688980957
transform 1 0 35512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0881_
timestamp 1688980957
transform 1 0 35236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0882_
timestamp 1688980957
transform 1 0 22908 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0883_
timestamp 1688980957
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  INST_config_UART._0884_
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  INST_config_UART._0885_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0886_
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  INST_config_UART._0887_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0888_
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0889_
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0890_
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0891_
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  INST_config_UART._0892_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22816 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0893_
timestamp 1688980957
transform 1 0 22816 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0894_
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  INST_config_UART._0895_
timestamp 1688980957
transform 1 0 24656 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0896_
timestamp 1688980957
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0897_
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0898_
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0899_
timestamp 1688980957
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0900_
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  INST_config_UART._0901_
timestamp 1688980957
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0902_
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  INST_config_UART._0903_
timestamp 1688980957
transform 1 0 10856 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  INST_config_UART._0904_
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0905_
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0906_
timestamp 1688980957
transform 1 0 14720 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0907_
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._0908_
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  INST_config_UART._0909_
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0910_
timestamp 1688980957
transform 1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0911_
timestamp 1688980957
transform 1 0 16008 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0912_
timestamp 1688980957
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0913_
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0914_
timestamp 1688980957
transform 1 0 25944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0915_
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0916_
timestamp 1688980957
transform 1 0 26312 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0917_
timestamp 1688980957
transform 1 0 24564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0918_
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0919_
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0920_
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0921_
timestamp 1688980957
transform 1 0 25024 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0922_
timestamp 1688980957
transform 1 0 24748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0923_
timestamp 1688980957
transform 1 0 24840 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0924_
timestamp 1688980957
transform 1 0 25576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0925_
timestamp 1688980957
transform 1 0 24748 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0926_
timestamp 1688980957
transform 1 0 25484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0927_
timestamp 1688980957
transform 1 0 25392 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._0928_
timestamp 1688980957
transform 1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._0929_
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._0930_
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0931_
timestamp 1688980957
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0932_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0933_
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0934_
timestamp 1688980957
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0935_
timestamp 1688980957
transform 1 0 9200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0936_
timestamp 1688980957
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0937_
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0938_
timestamp 1688980957
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._0939_
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  INST_config_UART._0940_
timestamp 1688980957
transform 1 0 10212 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0941_
timestamp 1688980957
transform 1 0 9108 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0942_
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0943_
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0944_
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0945_
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0946_
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0947_
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0948_
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0949_
timestamp 1688980957
transform 1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._0950_
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  INST_config_UART._0951_
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0952_
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  INST_config_UART._0953_
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  INST_config_UART._0954_
timestamp 1688980957
transform 1 0 11684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0955_
timestamp 1688980957
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0956_
timestamp 1688980957
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0957_
timestamp 1688980957
transform 1 0 12420 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0958_
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0959_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  INST_config_UART._0960_
timestamp 1688980957
transform 1 0 12972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0961_
timestamp 1688980957
transform 1 0 13432 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0962_
timestamp 1688980957
transform 1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0963_
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0964_
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0965_
timestamp 1688980957
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._0966_
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._0967_
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0968_
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0969_
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0970_
timestamp 1688980957
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._0971_
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  INST_config_UART._0972_
timestamp 1688980957
transform 1 0 18584 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  INST_config_UART._0973_
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  INST_config_UART._0974_
timestamp 1688980957
transform 1 0 16376 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  INST_config_UART._0975_
timestamp 1688980957
transform 1 0 16836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._0976_
timestamp 1688980957
transform 1 0 16376 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0977_
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._0978_
timestamp 1688980957
transform 1 0 16928 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0979_
timestamp 1688980957
transform 1 0 32200 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0980_
timestamp 1688980957
transform 1 0 32568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0981_
timestamp 1688980957
transform 1 0 33396 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0982_
timestamp 1688980957
transform 1 0 34040 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0983_
timestamp 1688980957
transform 1 0 33488 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0984_
timestamp 1688980957
transform 1 0 33212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0985_
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0986_
timestamp 1688980957
transform 1 0 28888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0987_
timestamp 1688980957
transform 1 0 34040 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0988_
timestamp 1688980957
transform 1 0 31464 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0989_
timestamp 1688980957
transform 1 0 30728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0990_
timestamp 1688980957
transform 1 0 28060 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0991_
timestamp 1688980957
transform 1 0 32660 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0992_
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._0993_
timestamp 1688980957
transform 1 0 36156 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._0994_
timestamp 1688980957
transform 1 0 32476 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._0995_
timestamp 1688980957
transform 1 0 21804 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._0996_
timestamp 1688980957
transform 1 0 19412 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._0997_
timestamp 1688980957
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._0998_
timestamp 1688980957
transform 1 0 20056 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  INST_config_UART._0999_
timestamp 1688980957
transform 1 0 20608 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._1000_
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._1001_
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._1002_
timestamp 1688980957
transform 1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._1003_
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  INST_config_UART._1004_
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1005_
timestamp 1688980957
transform 1 0 18768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1006_
timestamp 1688980957
transform 1 0 21252 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  INST_config_UART._1007_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._1008_
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  INST_config_UART._1009_
timestamp 1688980957
transform 1 0 20424 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  INST_config_UART._1010_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1011_
timestamp 1688980957
transform 1 0 20056 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1012_
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1013_
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._1014_
timestamp 1688980957
transform 1 0 20148 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._1015_
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  INST_config_UART._1016_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1017_
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1018_
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._1019_
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1020_
timestamp 1688980957
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._1021_
timestamp 1688980957
transform 1 0 20332 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1022_
timestamp 1688980957
transform 1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1023_
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._1024_
timestamp 1688980957
transform 1 0 19320 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1025_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._1026_
timestamp 1688980957
transform 1 0 20424 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1027_
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1028_
timestamp 1688980957
transform 1 0 22356 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1029_
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1030_
timestamp 1688980957
transform 1 0 22908 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1031_
timestamp 1688980957
transform 1 0 20148 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1032_
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1033_
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1034_
timestamp 1688980957
transform 1 0 23736 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._1035_
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1036_
timestamp 1688980957
transform 1 0 21160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  INST_config_UART._1037_
timestamp 1688980957
transform 1 0 18308 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._1038_
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  INST_config_UART._1039_
timestamp 1688980957
transform 1 0 20332 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1040_
timestamp 1688980957
transform 1 0 22816 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1041_
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1042_
timestamp 1688980957
transform 1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1043_
timestamp 1688980957
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  INST_config_UART._1044_
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1045_
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1046_
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  INST_config_UART._1047_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1048_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  INST_config_UART._1049_
timestamp 1688980957
transform 1 0 18952 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1050_
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._1051_
timestamp 1688980957
transform 1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1052_
timestamp 1688980957
transform 1 0 23736 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  INST_config_UART._1053_
timestamp 1688980957
transform 1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1054_
timestamp 1688980957
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  INST_config_UART._1055_
timestamp 1688980957
transform 1 0 18584 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1056_
timestamp 1688980957
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._1057_
timestamp 1688980957
transform 1 0 19320 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  INST_config_UART._1058_
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._1059_
timestamp 1688980957
transform 1 0 19596 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_2  INST_config_UART._1060_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  INST_config_UART._1061_
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  INST_config_UART._1062_
timestamp 1688980957
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  INST_config_UART._1063_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  INST_config_UART._1064_
timestamp 1688980957
transform 1 0 15456 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1065_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1066_
timestamp 1688980957
transform 1 0 16008 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._1067_
timestamp 1688980957
transform 1 0 16744 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1068_
timestamp 1688980957
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1069_
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1070_
timestamp 1688980957
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1071_
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  INST_config_UART._1072_
timestamp 1688980957
transform 1 0 15640 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  INST_config_UART._1073_
timestamp 1688980957
transform 1 0 16744 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  INST_config_UART._1074_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  INST_config_UART._1075_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._1076_
timestamp 1688980957
transform 1 0 17756 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1077_
timestamp 1688980957
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  INST_config_UART._1078_
timestamp 1688980957
transform 1 0 16008 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  INST_config_UART._1079_
timestamp 1688980957
transform 1 0 15456 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1080_
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._1081_
timestamp 1688980957
transform 1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  INST_config_UART._1082_
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  INST_config_UART._1083_
timestamp 1688980957
transform 1 0 14352 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  INST_config_UART._1084_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  INST_config_UART._1085_
timestamp 1688980957
transform 1 0 15364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1086_
timestamp 1688980957
transform 1 0 16008 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1087_
timestamp 1688980957
transform 1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1088_
timestamp 1688980957
transform 1 0 15364 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1089_
timestamp 1688980957
transform 1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  INST_config_UART._1090_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__a31oi_2  INST_config_UART._1091_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._1092_
timestamp 1688980957
transform 1 0 16836 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._1093_
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1094_
timestamp 1688980957
transform 1 0 16928 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1095_
timestamp 1688980957
transform 1 0 15088 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1096_
timestamp 1688980957
transform 1 0 14628 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  INST_config_UART._1097_
timestamp 1688980957
transform 1 0 17664 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  INST_config_UART._1098_
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  INST_config_UART._1099_
timestamp 1688980957
transform 1 0 17112 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  INST_config_UART._1100_
timestamp 1688980957
transform 1 0 16836 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._1101_
timestamp 1688980957
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  INST_config_UART._1102_
timestamp 1688980957
transform 1 0 16100 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  INST_config_UART._1103_
timestamp 1688980957
transform 1 0 15272 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1104_
timestamp 1688980957
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  INST_config_UART._1105_
timestamp 1688980957
transform 1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  INST_config_UART._1106_
timestamp 1688980957
transform 1 0 23736 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  INST_config_UART._1107_
timestamp 1688980957
transform 1 0 22356 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1108_
timestamp 1688980957
transform 1 0 20608 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._1109_
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1110_
timestamp 1688980957
transform 1 0 36708 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1111_
timestamp 1688980957
transform 1 0 36616 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1112_
timestamp 1688980957
transform 1 0 36616 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1113_
timestamp 1688980957
transform 1 0 36248 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1114_
timestamp 1688980957
transform 1 0 38272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1115_
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1116_
timestamp 1688980957
transform 1 0 38272 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1117_
timestamp 1688980957
transform 1 0 37996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1118_
timestamp 1688980957
transform 1 0 40296 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1119_
timestamp 1688980957
transform 1 0 41124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1120_
timestamp 1688980957
transform 1 0 39192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1121_
timestamp 1688980957
transform 1 0 38640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1122_
timestamp 1688980957
transform 1 0 35880 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1123_
timestamp 1688980957
transform 1 0 34776 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1124_
timestamp 1688980957
transform 1 0 35328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1125_
timestamp 1688980957
transform 1 0 36156 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1126_
timestamp 1688980957
transform 1 0 20148 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._1127_
timestamp 1688980957
transform 1 0 21252 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1128_
timestamp 1688980957
transform 1 0 32660 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1129_
timestamp 1688980957
transform 1 0 31096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1130_
timestamp 1688980957
transform 1 0 31556 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1131_
timestamp 1688980957
transform 1 0 30544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1132_
timestamp 1688980957
transform 1 0 33856 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1133_
timestamp 1688980957
transform 1 0 34040 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1134_
timestamp 1688980957
transform 1 0 33120 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1135_
timestamp 1688980957
transform 1 0 33120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1136_
timestamp 1688980957
transform 1 0 34040 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1137_
timestamp 1688980957
transform 1 0 33304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1138_
timestamp 1688980957
transform 1 0 34684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1139_
timestamp 1688980957
transform 1 0 33580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1140_
timestamp 1688980957
transform 1 0 34040 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1141_
timestamp 1688980957
transform 1 0 33488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1142_
timestamp 1688980957
transform 1 0 23460 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1143_
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  INST_config_UART._1144_
timestamp 1688980957
transform 1 0 26680 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  INST_config_UART._1145_
timestamp 1688980957
transform 1 0 25668 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1146_
timestamp 1688980957
transform 1 0 27784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1147_
timestamp 1688980957
transform 1 0 28060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1148_
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1149_
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1150_
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1151_
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1152_
timestamp 1688980957
transform 1 0 27784 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1153_
timestamp 1688980957
transform 1 0 29624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1154_
timestamp 1688980957
transform 1 0 28888 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1155_
timestamp 1688980957
transform 1 0 28520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1156_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1157_
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1158_
timestamp 1688980957
transform 1 0 27784 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1159_
timestamp 1688980957
transform 1 0 26404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1160_
timestamp 1688980957
transform 1 0 28612 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1161_
timestamp 1688980957
transform 1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1162_
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1163_
timestamp 1688980957
transform 1 0 22724 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1164_
timestamp 1688980957
transform 1 0 18676 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1165_
timestamp 1688980957
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1166_
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1167_
timestamp 1688980957
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  INST_config_UART._1168_
timestamp 1688980957
transform 1 0 21620 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1169_
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1170_
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1171_
timestamp 1688980957
transform 1 0 18676 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1172_
timestamp 1688980957
transform 1 0 17664 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1173_
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1174_
timestamp 1688980957
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  INST_config_UART._1175_
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  INST_config_UART._1176_
timestamp 1688980957
transform 1 0 21896 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  INST_config_UART._1177_
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1178_
timestamp 1688980957
transform 1 0 26128 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1179_
timestamp 1688980957
transform 1 0 16008 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1180_
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1181_
timestamp 1688980957
transform 1 0 16652 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1182_
timestamp 1688980957
transform 1 0 24104 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1183_
timestamp 1688980957
transform 1 0 17480 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1184_
timestamp 1688980957
transform 1 0 19872 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1185_
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1186_
timestamp 1688980957
transform 1 0 21068 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1187_
timestamp 1688980957
transform 1 0 26220 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1188_
timestamp 1688980957
transform 1 0 26312 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1189_
timestamp 1688980957
transform 1 0 28152 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1190_
timestamp 1688980957
transform 1 0 28888 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1191_
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1192_
timestamp 1688980957
transform 1 0 28888 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1193_
timestamp 1688980957
transform 1 0 29072 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1194_
timestamp 1688980957
transform 1 0 29440 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1195_
timestamp 1688980957
transform 1 0 30728 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1196_
timestamp 1688980957
transform 1 0 31464 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1197_
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1198_
timestamp 1688980957
transform 1 0 28428 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1199_
timestamp 1688980957
transform 1 0 28888 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1200_
timestamp 1688980957
transform 1 0 28888 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1201_
timestamp 1688980957
transform 1 0 29532 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1202_
timestamp 1688980957
transform 1 0 30728 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1203_
timestamp 1688980957
transform 1 0 29532 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1204_
timestamp 1688980957
transform 1 0 32292 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1205_
timestamp 1688980957
transform 1 0 31832 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1206_
timestamp 1688980957
transform 1 0 30452 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1207_
timestamp 1688980957
transform 1 0 31924 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1208_
timestamp 1688980957
transform 1 0 30820 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1209_
timestamp 1688980957
transform 1 0 31464 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1210_
timestamp 1688980957
transform 1 0 30912 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  INST_config_UART._1211_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27600 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1212_
timestamp 1688980957
transform 1 0 30084 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1213_
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1214_
timestamp 1688980957
transform 1 0 28980 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1215_
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_2  INST_config_UART._1216_
timestamp 1688980957
transform 1 0 19136 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1217_
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1218_
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1219_
timestamp 1688980957
transform 1 0 36616 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1220_
timestamp 1688980957
transform 1 0 36616 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1221_
timestamp 1688980957
transform 1 0 38456 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1222_
timestamp 1688980957
transform 1 0 39652 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1223_
timestamp 1688980957
transform 1 0 37812 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1224_
timestamp 1688980957
transform 1 0 39192 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1225_
timestamp 1688980957
transform 1 0 34408 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1226_
timestamp 1688980957
transform 1 0 34500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  INST_config_UART._1227_
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1228_
timestamp 1688980957
transform 1 0 24104 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1229_
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1230_
timestamp 1688980957
transform 1 0 33488 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1231_
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1232_
timestamp 1688980957
transform 1 0 37444 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1233_
timestamp 1688980957
transform 1 0 39192 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1234_
timestamp 1688980957
transform 1 0 39192 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1235_
timestamp 1688980957
transform 1 0 39284 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1236_
timestamp 1688980957
transform 1 0 35420 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1237_
timestamp 1688980957
transform 1 0 35880 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1238_
timestamp 1688980957
transform 1 0 19872 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1239_
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1240_
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1241_
timestamp 1688980957
transform 1 0 22816 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1242_
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1243_
timestamp 1688980957
transform 1 0 26312 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1244_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1245_
timestamp 1688980957
transform 1 0 25116 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1246_
timestamp 1688980957
transform 1 0 24840 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1247_
timestamp 1688980957
transform 1 0 24196 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1248_
timestamp 1688980957
transform 1 0 25576 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1249_
timestamp 1688980957
transform 1 0 25024 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1250_
timestamp 1688980957
transform 1 0 26404 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1251_
timestamp 1688980957
transform 1 0 24564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1252_
timestamp 1688980957
transform 1 0 25392 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1253_
timestamp 1688980957
transform 1 0 6348 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1254_
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1255_
timestamp 1688980957
transform 1 0 8280 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1256_
timestamp 1688980957
transform 1 0 8648 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1257_
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1258_
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1259_
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1260_
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1261_
timestamp 1688980957
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1262_
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1263_
timestamp 1688980957
transform 1 0 13432 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1264_
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1265_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1266_
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1267_
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1268_
timestamp 1688980957
transform 1 0 26312 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1269_
timestamp 1688980957
transform 1 0 26128 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1270_
timestamp 1688980957
transform 1 0 28152 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1271_
timestamp 1688980957
transform 1 0 16008 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1272_
timestamp 1688980957
transform 1 0 31464 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1273_
timestamp 1688980957
transform 1 0 32016 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1274_
timestamp 1688980957
transform 1 0 31648 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1275_
timestamp 1688980957
transform 1 0 26588 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1276_
timestamp 1688980957
transform 1 0 31556 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1277_
timestamp 1688980957
transform 1 0 26220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1278_
timestamp 1688980957
transform 1 0 32108 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1279_
timestamp 1688980957
transform 1 0 32476 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  INST_config_UART._1280_
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1281_
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1282_
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1283_
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1284_
timestamp 1688980957
transform 1 0 5704 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1285_
timestamp 1688980957
transform 1 0 5244 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1286_
timestamp 1688980957
transform 1 0 5704 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1287_
timestamp 1688980957
transform 1 0 4968 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1288_
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1289_
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1290_
timestamp 1688980957
transform 1 0 4784 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1291_
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1292_
timestamp 1688980957
transform 1 0 3772 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1293_
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1294_
timestamp 1688980957
transform 1 0 6348 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1295_
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1296_
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1297_
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1298_
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1299_
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1300_
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1301_
timestamp 1688980957
transform 1 0 11040 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1302_
timestamp 1688980957
transform 1 0 12696 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1303_
timestamp 1688980957
transform 1 0 18124 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1304_
timestamp 1688980957
transform 1 0 18584 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1305_
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1306_
timestamp 1688980957
transform 1 0 20608 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1307_
timestamp 1688980957
transform 1 0 20240 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1308_
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1309_
timestamp 1688980957
transform 1 0 17664 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1310_
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1311_
timestamp 1688980957
transform 1 0 14352 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1312_
timestamp 1688980957
transform 1 0 13800 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1313_
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1314_
timestamp 1688980957
transform 1 0 15088 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1315_
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1316_
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1317_
timestamp 1688980957
transform 1 0 13432 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1318_
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  INST_config_UART._1319_
timestamp 1688980957
transform 1 0 14904 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1320_
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  INST_config_UART._1321_
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1322_
timestamp 1688980957
transform 1 0 14628 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1323_
timestamp 1688980957
transform 1 0 24012 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1324_
timestamp 1688980957
transform 1 0 36616 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1325_
timestamp 1688980957
transform 1 0 35880 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1326_
timestamp 1688980957
transform 1 0 37904 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1327_
timestamp 1688980957
transform 1 0 38456 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1328_
timestamp 1688980957
transform 1 0 39192 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1329_
timestamp 1688980957
transform 1 0 39192 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1330_
timestamp 1688980957
transform 1 0 34408 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1331_
timestamp 1688980957
transform 1 0 34040 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1332_
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1333_
timestamp 1688980957
transform 1 0 30820 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1334_
timestamp 1688980957
transform 1 0 33304 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1335_
timestamp 1688980957
transform 1 0 34040 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1336_
timestamp 1688980957
transform 1 0 32844 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1337_
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1338_
timestamp 1688980957
transform 1 0 33304 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1339_
timestamp 1688980957
transform 1 0 22356 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1340_
timestamp 1688980957
transform 1 0 19504 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1341_
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1342_
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1343_
timestamp 1688980957
transform 1 0 16836 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1344_
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1345_
timestamp 1688980957
transform 1 0 16376 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1346_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1347_
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1348_
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1349_
timestamp 1688980957
transform 1 0 14812 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1350_
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1351_
timestamp 1688980957
transform 1 0 16100 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  INST_config_UART._1352_
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_4  INST_config_UART._1353_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43056 0 -1 11968
box -38 -48 2246 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1354_
timestamp 1688980957
transform 1 0 27324 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1355_
timestamp 1688980957
transform 1 0 26312 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1356_
timestamp 1688980957
transform 1 0 27140 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1357_
timestamp 1688980957
transform 1 0 28336 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1358_
timestamp 1688980957
transform 1 0 27968 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1359_
timestamp 1688980957
transform 1 0 26864 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1360_
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  INST_config_UART._1361_
timestamp 1688980957
transform 1 0 28888 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1362_
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1363_
timestamp 1688980957
transform 1 0 16652 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1364_
timestamp 1688980957
transform 1 0 20700 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1365_
timestamp 1688980957
transform 1 0 19780 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1366_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  INST_config_UART._1367_
timestamp 1688980957
transform 1 0 17204 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1368_
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1369_
timestamp 1688980957
transform 1 0 19044 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  INST_config_UART._1370_
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  load_slew111
timestamp 1688980957
transform 1 0 26956 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  load_slew112
timestamp 1688980957
transform 1 0 41676 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform 1 0 44712 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1688980957
transform 1 0 920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1688980957
transform 1 0 10120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output42
timestamp 1688980957
transform 1 0 11040 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1688980957
transform 1 0 17480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1688980957
transform 1 0 18584 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1688980957
transform 1 0 1840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 1688980957
transform 1 0 19136 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1688980957
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1688980957
transform 1 0 21160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output55
timestamp 1688980957
transform 1 0 22080 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1688980957
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1688980957
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output58
timestamp 1688980957
transform 1 0 24656 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1688980957
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1688980957
transform 1 0 26680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 28888 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 3128 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 29440 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform 1 0 30360 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1688980957
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1688980957
transform 1 0 4600 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1688980957
transform 1 0 6440 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1688980957
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1688980957
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 32292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1688980957
transform 1 0 9384 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform 1 0 10212 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 16008 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1688980957
transform 1 0 16836 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 1932 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform 1 0 20148 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 24564 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 26312 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 28152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform 1 0 5244 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 6072 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 6716 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 27600 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform 1 0 736 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 30728 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 30176 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 31464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 32752 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45540 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 45540 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 45540 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 45540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 45540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 45540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 45540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 45540 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 45540 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 45540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 45540 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 45540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 45540 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 45540 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 45540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 45540 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 45540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 45540 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 460 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 45540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 45540 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 45540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 45540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 45540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 45540 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 45540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 45540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 460 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 45540 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 13340 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 15916 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 18492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21068 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 23644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 26220 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 28796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 31372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 33948 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 36524 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39100 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 41676 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 44252 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 26220 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 31372 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 36524 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 41676 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 39100 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 5612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 39100 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 44252 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 5612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 36524 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 39100 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 44252 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 41676 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 39100 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 44252 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 36524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 41676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 39100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 41676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 39100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 44252 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 5612 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 44252 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 5612 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 36524 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 41676 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 5612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 41676 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3036 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 39100 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 44252 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 5612 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 41676 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 39100 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 44252 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 5612 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 41676 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 3036 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 39100 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 44252 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 5612 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 41676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 39100 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 41676 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 3036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 39100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 44252 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 5612 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 13340 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 28796 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 33948 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 39100 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 41676 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 44252 0 -1 22848
box -38 -48 130 592
<< labels >>
flabel metal3 s 45840 2728 46300 2848 0 FreeSans 480 0 0 0 CLK
port 0 nsew signal input
flabel metal3 s 45840 20680 46300 20800 0 FreeSans 480 0 0 0 ComActive
port 1 nsew signal tristate
flabel metal2 s 846 23840 902 24300 0 FreeSans 224 90 0 0 ConfigWriteData[0]
port 2 nsew signal tristate
flabel metal2 s 10046 23840 10102 24300 0 FreeSans 224 90 0 0 ConfigWriteData[10]
port 3 nsew signal tristate
flabel metal2 s 10966 23840 11022 24300 0 FreeSans 224 90 0 0 ConfigWriteData[11]
port 4 nsew signal tristate
flabel metal2 s 11886 23840 11942 24300 0 FreeSans 224 90 0 0 ConfigWriteData[12]
port 5 nsew signal tristate
flabel metal2 s 12806 23840 12862 24300 0 FreeSans 224 90 0 0 ConfigWriteData[13]
port 6 nsew signal tristate
flabel metal2 s 13726 23840 13782 24300 0 FreeSans 224 90 0 0 ConfigWriteData[14]
port 7 nsew signal tristate
flabel metal2 s 14646 23840 14702 24300 0 FreeSans 224 90 0 0 ConfigWriteData[15]
port 8 nsew signal tristate
flabel metal2 s 15566 23840 15622 24300 0 FreeSans 224 90 0 0 ConfigWriteData[16]
port 9 nsew signal tristate
flabel metal2 s 16486 23840 16542 24300 0 FreeSans 224 90 0 0 ConfigWriteData[17]
port 10 nsew signal tristate
flabel metal2 s 17406 23840 17462 24300 0 FreeSans 224 90 0 0 ConfigWriteData[18]
port 11 nsew signal tristate
flabel metal2 s 18326 23840 18382 24300 0 FreeSans 224 90 0 0 ConfigWriteData[19]
port 12 nsew signal tristate
flabel metal2 s 1766 23840 1822 24300 0 FreeSans 224 90 0 0 ConfigWriteData[1]
port 13 nsew signal tristate
flabel metal2 s 19246 23840 19302 24300 0 FreeSans 224 90 0 0 ConfigWriteData[20]
port 14 nsew signal tristate
flabel metal2 s 20166 23840 20222 24300 0 FreeSans 224 90 0 0 ConfigWriteData[21]
port 15 nsew signal tristate
flabel metal2 s 21086 23840 21142 24300 0 FreeSans 224 90 0 0 ConfigWriteData[22]
port 16 nsew signal tristate
flabel metal2 s 22006 23840 22062 24300 0 FreeSans 224 90 0 0 ConfigWriteData[23]
port 17 nsew signal tristate
flabel metal2 s 22926 23840 22982 24300 0 FreeSans 224 90 0 0 ConfigWriteData[24]
port 18 nsew signal tristate
flabel metal2 s 23846 23840 23902 24300 0 FreeSans 224 90 0 0 ConfigWriteData[25]
port 19 nsew signal tristate
flabel metal2 s 24766 23840 24822 24300 0 FreeSans 224 90 0 0 ConfigWriteData[26]
port 20 nsew signal tristate
flabel metal2 s 25686 23840 25742 24300 0 FreeSans 224 90 0 0 ConfigWriteData[27]
port 21 nsew signal tristate
flabel metal2 s 26606 23840 26662 24300 0 FreeSans 224 90 0 0 ConfigWriteData[28]
port 22 nsew signal tristate
flabel metal2 s 27526 23840 27582 24300 0 FreeSans 224 90 0 0 ConfigWriteData[29]
port 23 nsew signal tristate
flabel metal2 s 2686 23840 2742 24300 0 FreeSans 224 90 0 0 ConfigWriteData[2]
port 24 nsew signal tristate
flabel metal2 s 28446 23840 28502 24300 0 FreeSans 224 90 0 0 ConfigWriteData[30]
port 25 nsew signal tristate
flabel metal2 s 29366 23840 29422 24300 0 FreeSans 224 90 0 0 ConfigWriteData[31]
port 26 nsew signal tristate
flabel metal2 s 3606 23840 3662 24300 0 FreeSans 224 90 0 0 ConfigWriteData[3]
port 27 nsew signal tristate
flabel metal2 s 4526 23840 4582 24300 0 FreeSans 224 90 0 0 ConfigWriteData[4]
port 28 nsew signal tristate
flabel metal2 s 5446 23840 5502 24300 0 FreeSans 224 90 0 0 ConfigWriteData[5]
port 29 nsew signal tristate
flabel metal2 s 6366 23840 6422 24300 0 FreeSans 224 90 0 0 ConfigWriteData[6]
port 30 nsew signal tristate
flabel metal2 s 7286 23840 7342 24300 0 FreeSans 224 90 0 0 ConfigWriteData[7]
port 31 nsew signal tristate
flabel metal2 s 8206 23840 8262 24300 0 FreeSans 224 90 0 0 ConfigWriteData[8]
port 32 nsew signal tristate
flabel metal2 s 9126 23840 9182 24300 0 FreeSans 224 90 0 0 ConfigWriteData[9]
port 33 nsew signal tristate
flabel metal2 s 30286 23840 30342 24300 0 FreeSans 224 90 0 0 ConfigWriteStrobe
port 34 nsew signal tristate
flabel metal2 s 1030 -300 1086 160 0 FreeSans 224 90 0 0 FrameAddressRegister[0]
port 35 nsew signal tristate
flabel metal2 s 9310 -300 9366 160 0 FreeSans 224 90 0 0 FrameAddressRegister[10]
port 36 nsew signal tristate
flabel metal2 s 10138 -300 10194 160 0 FreeSans 224 90 0 0 FrameAddressRegister[11]
port 37 nsew signal tristate
flabel metal2 s 10966 -300 11022 160 0 FreeSans 224 90 0 0 FrameAddressRegister[12]
port 38 nsew signal tristate
flabel metal2 s 11794 -300 11850 160 0 FreeSans 224 90 0 0 FrameAddressRegister[13]
port 39 nsew signal tristate
flabel metal2 s 12622 -300 12678 160 0 FreeSans 224 90 0 0 FrameAddressRegister[14]
port 40 nsew signal tristate
flabel metal2 s 13450 -300 13506 160 0 FreeSans 224 90 0 0 FrameAddressRegister[15]
port 41 nsew signal tristate
flabel metal2 s 14278 -300 14334 160 0 FreeSans 224 90 0 0 FrameAddressRegister[16]
port 42 nsew signal tristate
flabel metal2 s 15106 -300 15162 160 0 FreeSans 224 90 0 0 FrameAddressRegister[17]
port 43 nsew signal tristate
flabel metal2 s 15934 -300 15990 160 0 FreeSans 224 90 0 0 FrameAddressRegister[18]
port 44 nsew signal tristate
flabel metal2 s 16762 -300 16818 160 0 FreeSans 224 90 0 0 FrameAddressRegister[19]
port 45 nsew signal tristate
flabel metal2 s 1858 -300 1914 160 0 FreeSans 224 90 0 0 FrameAddressRegister[1]
port 46 nsew signal tristate
flabel metal2 s 17590 -300 17646 160 0 FreeSans 224 90 0 0 FrameAddressRegister[20]
port 47 nsew signal tristate
flabel metal2 s 18418 -300 18474 160 0 FreeSans 224 90 0 0 FrameAddressRegister[21]
port 48 nsew signal tristate
flabel metal2 s 19246 -300 19302 160 0 FreeSans 224 90 0 0 FrameAddressRegister[22]
port 49 nsew signal tristate
flabel metal2 s 20074 -300 20130 160 0 FreeSans 224 90 0 0 FrameAddressRegister[23]
port 50 nsew signal tristate
flabel metal2 s 20902 -300 20958 160 0 FreeSans 224 90 0 0 FrameAddressRegister[24]
port 51 nsew signal tristate
flabel metal2 s 21730 -300 21786 160 0 FreeSans 224 90 0 0 FrameAddressRegister[25]
port 52 nsew signal tristate
flabel metal2 s 22558 -300 22614 160 0 FreeSans 224 90 0 0 FrameAddressRegister[26]
port 53 nsew signal tristate
flabel metal2 s 23386 -300 23442 160 0 FreeSans 224 90 0 0 FrameAddressRegister[27]
port 54 nsew signal tristate
flabel metal2 s 24214 -300 24270 160 0 FreeSans 224 90 0 0 FrameAddressRegister[28]
port 55 nsew signal tristate
flabel metal2 s 25042 -300 25098 160 0 FreeSans 224 90 0 0 FrameAddressRegister[29]
port 56 nsew signal tristate
flabel metal2 s 2686 -300 2742 160 0 FreeSans 224 90 0 0 FrameAddressRegister[2]
port 57 nsew signal tristate
flabel metal2 s 25870 -300 25926 160 0 FreeSans 224 90 0 0 FrameAddressRegister[30]
port 58 nsew signal tristate
flabel metal2 s 26698 -300 26754 160 0 FreeSans 224 90 0 0 FrameAddressRegister[31]
port 59 nsew signal tristate
flabel metal2 s 3514 -300 3570 160 0 FreeSans 224 90 0 0 FrameAddressRegister[3]
port 60 nsew signal tristate
flabel metal2 s 4342 -300 4398 160 0 FreeSans 224 90 0 0 FrameAddressRegister[4]
port 61 nsew signal tristate
flabel metal2 s 5170 -300 5226 160 0 FreeSans 224 90 0 0 FrameAddressRegister[5]
port 62 nsew signal tristate
flabel metal2 s 5998 -300 6054 160 0 FreeSans 224 90 0 0 FrameAddressRegister[6]
port 63 nsew signal tristate
flabel metal2 s 6826 -300 6882 160 0 FreeSans 224 90 0 0 FrameAddressRegister[7]
port 64 nsew signal tristate
flabel metal2 s 7654 -300 7710 160 0 FreeSans 224 90 0 0 FrameAddressRegister[8]
port 65 nsew signal tristate
flabel metal2 s 8482 -300 8538 160 0 FreeSans 224 90 0 0 FrameAddressRegister[9]
port 66 nsew signal tristate
flabel metal2 s 27526 -300 27582 160 0 FreeSans 224 90 0 0 LongFrameStrobe
port 67 nsew signal tristate
flabel metal3 s -300 8712 160 8832 0 FreeSans 480 0 0 0 ReceiveLED
port 68 nsew signal tristate
flabel metal2 s 28354 -300 28410 160 0 FreeSans 224 90 0 0 RowSelect[0]
port 69 nsew signal tristate
flabel metal2 s 29182 -300 29238 160 0 FreeSans 224 90 0 0 RowSelect[1]
port 70 nsew signal tristate
flabel metal2 s 30010 -300 30066 160 0 FreeSans 224 90 0 0 RowSelect[2]
port 71 nsew signal tristate
flabel metal2 s 30838 -300 30894 160 0 FreeSans 224 90 0 0 RowSelect[3]
port 72 nsew signal tristate
flabel metal2 s 31666 -300 31722 160 0 FreeSans 224 90 0 0 RowSelect[4]
port 73 nsew signal tristate
flabel metal3 s 45840 14696 46300 14816 0 FreeSans 480 0 0 0 Rx
port 74 nsew signal input
flabel metal2 s 31206 23840 31262 24300 0 FreeSans 224 90 0 0 SelfWriteData[0]
port 75 nsew signal input
flabel metal2 s 40406 23840 40462 24300 0 FreeSans 224 90 0 0 SelfWriteData[10]
port 76 nsew signal input
flabel metal2 s 41326 23840 41382 24300 0 FreeSans 224 90 0 0 SelfWriteData[11]
port 77 nsew signal input
flabel metal2 s 42246 23840 42302 24300 0 FreeSans 224 90 0 0 SelfWriteData[12]
port 78 nsew signal input
flabel metal2 s 43166 23840 43222 24300 0 FreeSans 224 90 0 0 SelfWriteData[13]
port 79 nsew signal input
flabel metal2 s 44086 23840 44142 24300 0 FreeSans 224 90 0 0 SelfWriteData[14]
port 80 nsew signal input
flabel metal2 s 45006 23840 45062 24300 0 FreeSans 224 90 0 0 SelfWriteData[15]
port 81 nsew signal input
flabel metal2 s 32494 -300 32550 160 0 FreeSans 224 90 0 0 SelfWriteData[16]
port 82 nsew signal input
flabel metal2 s 33322 -300 33378 160 0 FreeSans 224 90 0 0 SelfWriteData[17]
port 83 nsew signal input
flabel metal2 s 34150 -300 34206 160 0 FreeSans 224 90 0 0 SelfWriteData[18]
port 84 nsew signal input
flabel metal2 s 34978 -300 35034 160 0 FreeSans 224 90 0 0 SelfWriteData[19]
port 85 nsew signal input
flabel metal2 s 32126 23840 32182 24300 0 FreeSans 224 90 0 0 SelfWriteData[1]
port 86 nsew signal input
flabel metal2 s 35806 -300 35862 160 0 FreeSans 224 90 0 0 SelfWriteData[20]
port 87 nsew signal input
flabel metal2 s 36634 -300 36690 160 0 FreeSans 224 90 0 0 SelfWriteData[21]
port 88 nsew signal input
flabel metal2 s 37462 -300 37518 160 0 FreeSans 224 90 0 0 SelfWriteData[22]
port 89 nsew signal input
flabel metal2 s 38290 -300 38346 160 0 FreeSans 224 90 0 0 SelfWriteData[23]
port 90 nsew signal input
flabel metal2 s 39118 -300 39174 160 0 FreeSans 224 90 0 0 SelfWriteData[24]
port 91 nsew signal input
flabel metal2 s 39946 -300 40002 160 0 FreeSans 224 90 0 0 SelfWriteData[25]
port 92 nsew signal input
flabel metal2 s 40774 -300 40830 160 0 FreeSans 224 90 0 0 SelfWriteData[26]
port 93 nsew signal input
flabel metal2 s 41602 -300 41658 160 0 FreeSans 224 90 0 0 SelfWriteData[27]
port 94 nsew signal input
flabel metal2 s 42430 -300 42486 160 0 FreeSans 224 90 0 0 SelfWriteData[28]
port 95 nsew signal input
flabel metal2 s 43258 -300 43314 160 0 FreeSans 224 90 0 0 SelfWriteData[29]
port 96 nsew signal input
flabel metal2 s 33046 23840 33102 24300 0 FreeSans 224 90 0 0 SelfWriteData[2]
port 97 nsew signal input
flabel metal2 s 44086 -300 44142 160 0 FreeSans 224 90 0 0 SelfWriteData[30]
port 98 nsew signal input
flabel metal2 s 44914 -300 44970 160 0 FreeSans 224 90 0 0 SelfWriteData[31]
port 99 nsew signal input
flabel metal2 s 33966 23840 34022 24300 0 FreeSans 224 90 0 0 SelfWriteData[3]
port 100 nsew signal input
flabel metal2 s 34886 23840 34942 24300 0 FreeSans 224 90 0 0 SelfWriteData[4]
port 101 nsew signal input
flabel metal2 s 35806 23840 35862 24300 0 FreeSans 224 90 0 0 SelfWriteData[5]
port 102 nsew signal input
flabel metal2 s 36726 23840 36782 24300 0 FreeSans 224 90 0 0 SelfWriteData[6]
port 103 nsew signal input
flabel metal2 s 37646 23840 37702 24300 0 FreeSans 224 90 0 0 SelfWriteData[7]
port 104 nsew signal input
flabel metal2 s 38566 23840 38622 24300 0 FreeSans 224 90 0 0 SelfWriteData[8]
port 105 nsew signal input
flabel metal2 s 39486 23840 39542 24300 0 FreeSans 224 90 0 0 SelfWriteData[9]
port 106 nsew signal input
flabel metal3 s -300 2728 160 2848 0 FreeSans 480 0 0 0 SelfWriteStrobe
port 107 nsew signal input
flabel metal3 s 45840 8712 46300 8832 0 FreeSans 480 0 0 0 resetn
port 108 nsew signal input
flabel metal3 s -300 14696 160 14816 0 FreeSans 480 0 0 0 s_clk
port 109 nsew signal input
flabel metal3 s -300 20680 160 20800 0 FreeSans 480 0 0 0 s_data
port 110 nsew signal input
flabel metal4 s 3564 1040 3884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 8564 1040 8884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 13564 1040 13884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 18564 1040 18884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 23564 1040 23884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 28564 1040 28884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 33564 1040 33884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 38564 1040 38884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 43564 1040 43884 22896 0 FreeSans 1920 90 0 0 vccd1
port 111 nsew power bidirectional
flabel metal4 s 6064 1040 6384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 11064 1040 11384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 16064 1040 16384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 21064 1040 21384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 26064 1040 26384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 31064 1040 31384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 36064 1040 36384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
flabel metal4 s 41064 1040 41384 22896 0 FreeSans 1920 90 0 0 vssd1
port 112 nsew ground bidirectional
rlabel metal1 23000 22304 23000 22304 0 vccd1
rlabel metal1 23000 22848 23000 22848 0 vssd1
rlabel metal3 45272 2788 45272 2788 0 CLK
rlabel metal3 45548 20740 45548 20740 0 ComActive
rlabel metal1 27646 5610 27646 5610 0 ConfigFSM_inst.FSM_Reset
rlabel metal1 1794 2482 1794 2482 0 ConfigFSM_inst.FrameAddressRegister\[0\]
rlabel metal1 10166 1938 10166 1938 0 ConfigFSM_inst.FrameAddressRegister\[10\]
rlabel metal2 10534 2349 10534 2349 0 ConfigFSM_inst.FrameAddressRegister\[11\]
rlabel metal1 11592 1938 11592 1938 0 ConfigFSM_inst.FrameAddressRegister\[12\]
rlabel metal2 12190 4080 12190 4080 0 ConfigFSM_inst.FrameAddressRegister\[13\]
rlabel metal2 12512 1938 12512 1938 0 ConfigFSM_inst.FrameAddressRegister\[14\]
rlabel metal1 14122 2414 14122 2414 0 ConfigFSM_inst.FrameAddressRegister\[15\]
rlabel metal2 14536 1938 14536 1938 0 ConfigFSM_inst.FrameAddressRegister\[16\]
rlabel metal1 16284 2618 16284 2618 0 ConfigFSM_inst.FrameAddressRegister\[17\]
rlabel metal1 16514 1938 16514 1938 0 ConfigFSM_inst.FrameAddressRegister\[18\]
rlabel metal1 18768 2482 18768 2482 0 ConfigFSM_inst.FrameAddressRegister\[19\]
rlabel metal2 2346 3196 2346 3196 0 ConfigFSM_inst.FrameAddressRegister\[1\]
rlabel metal1 18906 2890 18906 2890 0 ConfigFSM_inst.FrameAddressRegister\[21\]
rlabel metal1 20562 2958 20562 2958 0 ConfigFSM_inst.FrameAddressRegister\[22\]
rlabel metal2 21666 2176 21666 2176 0 ConfigFSM_inst.FrameAddressRegister\[23\]
rlabel metal1 20516 3366 20516 3366 0 ConfigFSM_inst.FrameAddressRegister\[24\]
rlabel metal2 22034 2873 22034 2873 0 ConfigFSM_inst.FrameAddressRegister\[25\]
rlabel metal1 22448 2618 22448 2618 0 ConfigFSM_inst.FrameAddressRegister\[26\]
rlabel metal1 23920 2618 23920 2618 0 ConfigFSM_inst.FrameAddressRegister\[27\]
rlabel metal2 22540 1326 22540 1326 0 ConfigFSM_inst.FrameAddressRegister\[28\]
rlabel metal1 24426 1734 24426 1734 0 ConfigFSM_inst.FrameAddressRegister\[29\]
rlabel metal1 2944 1938 2944 1938 0 ConfigFSM_inst.FrameAddressRegister\[2\]
rlabel metal1 26404 2618 26404 2618 0 ConfigFSM_inst.FrameAddressRegister\[30\]
rlabel metal1 27324 2618 27324 2618 0 ConfigFSM_inst.FrameAddressRegister\[31\]
rlabel metal1 4048 1938 4048 1938 0 ConfigFSM_inst.FrameAddressRegister\[3\]
rlabel metal2 4692 1938 4692 1938 0 ConfigFSM_inst.FrameAddressRegister\[4\]
rlabel metal1 5474 4046 5474 4046 0 ConfigFSM_inst.FrameAddressRegister\[5\]
rlabel metal1 6578 1938 6578 1938 0 ConfigFSM_inst.FrameAddressRegister\[6\]
rlabel metal1 7452 3162 7452 3162 0 ConfigFSM_inst.FrameAddressRegister\[7\]
rlabel metal1 8142 1938 8142 1938 0 ConfigFSM_inst.FrameAddressRegister\[8\]
rlabel metal1 9752 2414 9752 2414 0 ConfigFSM_inst.FrameAddressRegister\[9\]
rlabel metal1 33304 1326 33304 1326 0 ConfigFSM_inst.FrameShiftState\[0\]
rlabel metal1 30222 2822 30222 2822 0 ConfigFSM_inst.FrameShiftState\[1\]
rlabel metal1 33810 1394 33810 1394 0 ConfigFSM_inst.FrameShiftState\[2\]
rlabel metal1 29394 2414 29394 2414 0 ConfigFSM_inst.FrameShiftState\[3\]
rlabel metal1 30130 2482 30130 2482 0 ConfigFSM_inst.FrameShiftState\[4\]
rlabel metal1 25438 1904 25438 1904 0 ConfigFSM_inst.FrameStrobe
rlabel via2 33902 1309 33902 1309 0 ConfigFSM_inst.RowSelect\[0\]
rlabel metal1 31050 2074 31050 2074 0 ConfigFSM_inst.RowSelect\[1\]
rlabel metal1 34546 1292 34546 1292 0 ConfigFSM_inst.RowSelect\[2\]
rlabel metal1 33442 2414 33442 2414 0 ConfigFSM_inst.RowSelect\[3\]
rlabel metal1 35880 1326 35880 1326 0 ConfigFSM_inst.RowSelect\[4\]
rlabel metal2 1978 22338 1978 22338 0 ConfigFSM_inst.WriteData\[0\]
rlabel metal2 20102 1088 20102 1088 0 ConfigFSM_inst.WriteData\[10\]
rlabel metal2 22310 22583 22310 22583 0 ConfigFSM_inst.WriteData\[11\]
rlabel metal2 32522 19737 32522 19737 0 ConfigFSM_inst.WriteData\[12\]
rlabel metal2 13110 19363 13110 19363 0 ConfigFSM_inst.WriteData\[13\]
rlabel metal1 33718 16592 33718 16592 0 ConfigFSM_inst.WriteData\[14\]
rlabel metal2 14168 15572 14168 15572 0 ConfigFSM_inst.WriteData\[15\]
rlabel metal2 32890 5933 32890 5933 0 ConfigFSM_inst.WriteData\[16\]
rlabel metal1 17158 21998 17158 21998 0 ConfigFSM_inst.WriteData\[17\]
rlabel metal1 17480 21998 17480 21998 0 ConfigFSM_inst.WriteData\[18\]
rlabel metal2 12650 21165 12650 21165 0 ConfigFSM_inst.WriteData\[19\]
rlabel metal1 2254 21964 2254 21964 0 ConfigFSM_inst.WriteData\[1\]
rlabel metal1 19872 21998 19872 21998 0 ConfigFSM_inst.WriteData\[20\]
rlabel metal1 13110 21862 13110 21862 0 ConfigFSM_inst.WriteData\[21\]
rlabel metal1 14582 2618 14582 2618 0 ConfigFSM_inst.WriteData\[22\]
rlabel metal2 21574 1394 21574 1394 0 ConfigFSM_inst.WriteData\[23\]
rlabel metal3 19757 21692 19757 21692 0 ConfigFSM_inst.WriteData\[24\]
rlabel metal1 20930 1768 20930 1768 0 ConfigFSM_inst.WriteData\[25\]
rlabel metal2 14858 3927 14858 3927 0 ConfigFSM_inst.WriteData\[26\]
rlabel metal3 25737 22100 25737 22100 0 ConfigFSM_inst.WriteData\[27\]
rlabel metal1 27370 22610 27370 22610 0 ConfigFSM_inst.WriteData\[28\]
rlabel metal3 25921 19788 25921 19788 0 ConfigFSM_inst.WriteData\[29\]
rlabel metal1 2576 2414 2576 2414 0 ConfigFSM_inst.WriteData\[2\]
rlabel metal1 14214 952 14214 952 0 ConfigFSM_inst.WriteData\[30\]
rlabel via2 43838 20315 43838 20315 0 ConfigFSM_inst.WriteData\[31\]
rlabel metal1 28152 22406 28152 22406 0 ConfigFSM_inst.WriteData\[3\]
rlabel metal2 19274 2227 19274 2227 0 ConfigFSM_inst.WriteData\[4\]
rlabel metal2 6026 22610 6026 22610 0 ConfigFSM_inst.WriteData\[5\]
rlabel metal1 29210 22474 29210 22474 0 ConfigFSM_inst.WriteData\[6\]
rlabel metal1 18354 1224 18354 1224 0 ConfigFSM_inst.WriteData\[7\]
rlabel metal1 8234 22610 8234 22610 0 ConfigFSM_inst.WriteData\[8\]
rlabel metal1 9384 22406 9384 22406 0 ConfigFSM_inst.WriteData\[9\]
rlabel metal1 24610 2074 24610 2074 0 ConfigFSM_inst._000_
rlabel metal1 27278 1870 27278 1870 0 ConfigFSM_inst._001_
rlabel metal1 26588 5202 26588 5202 0 ConfigFSM_inst._002_
rlabel metal1 27646 2346 27646 2346 0 ConfigFSM_inst._003_
rlabel metal1 26174 4046 26174 4046 0 ConfigFSM_inst._004_
rlabel metal1 32384 2482 32384 2482 0 ConfigFSM_inst._005_
rlabel metal1 32476 1530 32476 1530 0 ConfigFSM_inst._006_
rlabel metal1 31970 3128 31970 3128 0 ConfigFSM_inst._007_
rlabel metal1 29532 3570 29532 3570 0 ConfigFSM_inst._008_
rlabel metal1 28520 1870 28520 1870 0 ConfigFSM_inst._009_
rlabel metal1 1426 4046 1426 4046 0 ConfigFSM_inst._010_
rlabel metal1 1564 4658 1564 4658 0 ConfigFSM_inst._011_
rlabel metal1 1886 2618 1886 2618 0 ConfigFSM_inst._012_
rlabel metal1 3404 2074 3404 2074 0 ConfigFSM_inst._013_
rlabel metal2 4462 3264 4462 3264 0 ConfigFSM_inst._014_
rlabel metal1 4232 4182 4232 4182 0 ConfigFSM_inst._015_
rlabel metal1 5658 4250 5658 4250 0 ConfigFSM_inst._016_
rlabel metal1 6348 3094 6348 3094 0 ConfigFSM_inst._017_
rlabel metal1 6900 4046 6900 4046 0 ConfigFSM_inst._018_
rlabel metal1 8510 3162 8510 3162 0 ConfigFSM_inst._019_
rlabel metal2 8970 3434 8970 3434 0 ConfigFSM_inst._020_
rlabel metal1 9430 4182 9430 4182 0 ConfigFSM_inst._021_
rlabel metal1 10626 2074 10626 2074 0 ConfigFSM_inst._022_
rlabel metal1 11454 3570 11454 3570 0 ConfigFSM_inst._023_
rlabel metal1 11960 4182 11960 4182 0 ConfigFSM_inst._024_
rlabel metal1 12650 2074 12650 2074 0 ConfigFSM_inst._025_
rlabel metal1 13202 2958 13202 2958 0 ConfigFSM_inst._026_
rlabel metal2 14628 2346 14628 2346 0 ConfigFSM_inst._027_
rlabel metal1 15502 3162 15502 3162 0 ConfigFSM_inst._028_
rlabel metal1 17388 2074 17388 2074 0 ConfigFSM_inst._029_
rlabel metal1 17342 3128 17342 3128 0 ConfigFSM_inst._030_
rlabel metal1 19320 3094 19320 3094 0 ConfigFSM_inst._031_
rlabel metal1 20332 2074 20332 2074 0 ConfigFSM_inst._032_
rlabel metal1 20746 3162 20746 3162 0 ConfigFSM_inst._033_
rlabel metal1 21482 3128 21482 3128 0 ConfigFSM_inst._034_
rlabel metal2 21574 4250 21574 4250 0 ConfigFSM_inst._035_
rlabel metal1 22310 2074 22310 2074 0 ConfigFSM_inst._036_
rlabel metal2 22126 4828 22126 4828 0 ConfigFSM_inst._037_
rlabel metal2 23046 2414 23046 2414 0 ConfigFSM_inst._038_
rlabel metal1 24426 3128 24426 3128 0 ConfigFSM_inst._039_
rlabel metal1 26128 2482 26128 2482 0 ConfigFSM_inst._040_
rlabel metal2 28382 5644 28382 5644 0 ConfigFSM_inst._041_
rlabel metal2 28290 5270 28290 5270 0 ConfigFSM_inst._042_
rlabel metal1 30038 1972 30038 1972 0 ConfigFSM_inst._043_
rlabel metal1 27488 4216 27488 4216 0 ConfigFSM_inst._044_
rlabel metal2 25806 4556 25806 4556 0 ConfigFSM_inst._045_
rlabel metal1 25392 5542 25392 5542 0 ConfigFSM_inst._046_
rlabel metal2 25714 4284 25714 4284 0 ConfigFSM_inst._047_
rlabel metal1 25622 4182 25622 4182 0 ConfigFSM_inst._048_
rlabel metal1 26312 3910 26312 3910 0 ConfigFSM_inst._049_
rlabel metal1 24886 4114 24886 4114 0 ConfigFSM_inst._050_
rlabel metal1 24702 5542 24702 5542 0 ConfigFSM_inst._051_
rlabel metal1 24610 4046 24610 4046 0 ConfigFSM_inst._052_
rlabel metal1 24518 4114 24518 4114 0 ConfigFSM_inst._053_
rlabel metal1 25852 3978 25852 3978 0 ConfigFSM_inst._054_
rlabel metal1 28290 5270 28290 5270 0 ConfigFSM_inst._055_
rlabel metal2 25806 5270 25806 5270 0 ConfigFSM_inst._056_
rlabel metal1 28290 2414 28290 2414 0 ConfigFSM_inst._057_
rlabel metal1 28888 1530 28888 1530 0 ConfigFSM_inst._058_
rlabel metal1 29532 3094 29532 3094 0 ConfigFSM_inst._059_
rlabel metal2 27554 3604 27554 3604 0 ConfigFSM_inst._060_
rlabel metal2 19274 3910 19274 3910 0 ConfigFSM_inst._061_
rlabel metal2 2438 2652 2438 2652 0 ConfigFSM_inst._062_
rlabel metal1 26358 3162 26358 3162 0 ConfigFSM_inst._063_
rlabel metal1 26956 4114 26956 4114 0 ConfigFSM_inst._064_
rlabel metal1 26542 4080 26542 4080 0 ConfigFSM_inst._065_
rlabel metal1 26128 1802 26128 1802 0 ConfigFSM_inst._066_
rlabel metal1 29256 1190 29256 1190 0 ConfigFSM_inst._067_
rlabel metal2 29946 1700 29946 1700 0 ConfigFSM_inst._068_
rlabel metal1 31878 1802 31878 1802 0 ConfigFSM_inst._069_
rlabel metal1 31970 3400 31970 3400 0 ConfigFSM_inst._070_
rlabel metal2 36110 1377 36110 1377 0 ConfigFSM_inst._071_
rlabel metal1 26496 2074 26496 2074 0 ConfigFSM_inst._072_
rlabel metal1 28566 3910 28566 3910 0 ConfigFSM_inst._073_
rlabel metal1 28934 3468 28934 3468 0 ConfigFSM_inst._074_
rlabel metal1 31556 3434 31556 3434 0 ConfigFSM_inst._075_
rlabel metal2 31234 2567 31234 2567 0 ConfigFSM_inst._076_
rlabel metal2 33350 3502 33350 3502 0 ConfigFSM_inst._077_
rlabel metal1 32108 1326 32108 1326 0 ConfigFSM_inst._078_
rlabel metal1 31326 2822 31326 2822 0 ConfigFSM_inst._079_
rlabel metal1 33534 1190 33534 1190 0 ConfigFSM_inst._080_
rlabel metal1 33166 3162 33166 3162 0 ConfigFSM_inst._081_
rlabel metal1 30590 3706 30590 3706 0 ConfigFSM_inst._082_
rlabel metal2 29762 3638 29762 3638 0 ConfigFSM_inst._083_
rlabel metal1 28566 3536 28566 3536 0 ConfigFSM_inst._084_
rlabel metal2 28842 2482 28842 2482 0 ConfigFSM_inst._085_
rlabel metal1 28888 2414 28888 2414 0 ConfigFSM_inst._086_
rlabel metal1 1150 4624 1150 4624 0 ConfigFSM_inst._087_
rlabel metal1 1932 5202 1932 5202 0 ConfigFSM_inst._088_
rlabel metal1 2208 2414 2208 2414 0 ConfigFSM_inst._089_
rlabel metal2 3450 1938 3450 1938 0 ConfigFSM_inst._090_
rlabel metal1 4416 3026 4416 3026 0 ConfigFSM_inst._091_
rlabel metal1 4646 5202 4646 5202 0 ConfigFSM_inst._092_
rlabel metal1 5934 4182 5934 4182 0 ConfigFSM_inst._093_
rlabel metal1 6670 3502 6670 3502 0 ConfigFSM_inst._094_
rlabel metal1 7820 4590 7820 4590 0 ConfigFSM_inst._095_
rlabel metal1 14168 4046 14168 4046 0 ConfigFSM_inst._096_
rlabel metal1 8832 2618 8832 2618 0 ConfigFSM_inst._097_
rlabel metal1 9614 3706 9614 3706 0 ConfigFSM_inst._098_
rlabel metal1 9936 4590 9936 4590 0 ConfigFSM_inst._099_
rlabel metal1 11270 2006 11270 2006 0 ConfigFSM_inst._100_
rlabel metal1 11454 4148 11454 4148 0 ConfigFSM_inst._101_
rlabel metal2 12282 4998 12282 4998 0 ConfigFSM_inst._102_
rlabel metal1 12650 3060 12650 3060 0 ConfigFSM_inst._103_
rlabel metal1 13662 4114 13662 4114 0 ConfigFSM_inst._104_
rlabel metal1 15042 2992 15042 2992 0 ConfigFSM_inst._105_
rlabel metal1 15870 3060 15870 3060 0 ConfigFSM_inst._106_
rlabel metal1 21896 1870 21896 1870 0 ConfigFSM_inst._107_
rlabel metal1 17986 1972 17986 1972 0 ConfigFSM_inst._108_
rlabel metal1 18584 3502 18584 3502 0 ConfigFSM_inst._109_
rlabel metal1 19688 2414 19688 2414 0 ConfigFSM_inst._110_
rlabel metal1 20654 1972 20654 1972 0 ConfigFSM_inst._111_
rlabel metal1 20792 3026 20792 3026 0 ConfigFSM_inst._112_
rlabel metal1 23230 3468 23230 3468 0 ConfigFSM_inst._113_
rlabel metal1 22770 4250 22770 4250 0 ConfigFSM_inst._114_
rlabel metal2 23828 1870 23828 1870 0 ConfigFSM_inst._115_
rlabel metal1 23230 4794 23230 4794 0 ConfigFSM_inst._116_
rlabel metal1 23276 3026 23276 3026 0 ConfigFSM_inst._117_
rlabel metal1 24978 3502 24978 3502 0 ConfigFSM_inst._118_
rlabel metal1 26542 3060 26542 3060 0 ConfigFSM_inst._119_
rlabel metal1 25806 1530 25806 1530 0 ConfigFSM_inst.oldFrameStrobe
rlabel metal1 27140 5882 27140 5882 0 ConfigFSM_inst.old_reset
rlabel metal1 28037 5270 28037 5270 0 ConfigFSM_inst.state\[0\]
rlabel metal1 30268 2414 30268 2414 0 ConfigFSM_inst.state\[1\]
rlabel metal1 27784 4658 27784 4658 0 ConfigFSM_inst.state\[2\]
rlabel metal1 1012 22746 1012 22746 0 ConfigWriteData[0]
rlabel metal1 10212 22746 10212 22746 0 ConfigWriteData[10]
rlabel metal2 10994 23300 10994 23300 0 ConfigWriteData[11]
rlabel metal1 12052 22746 12052 22746 0 ConfigWriteData[12]
rlabel metal1 12972 22746 12972 22746 0 ConfigWriteData[13]
rlabel metal2 13754 23249 13754 23249 0 ConfigWriteData[14]
rlabel metal1 14812 22746 14812 22746 0 ConfigWriteData[15]
rlabel metal1 15916 22746 15916 22746 0 ConfigWriteData[16]
rlabel metal2 16514 23300 16514 23300 0 ConfigWriteData[17]
rlabel metal1 17572 22746 17572 22746 0 ConfigWriteData[18]
rlabel metal1 18584 22746 18584 22746 0 ConfigWriteData[19]
rlabel metal1 1932 22746 1932 22746 0 ConfigWriteData[1]
rlabel metal2 19274 23300 19274 23300 0 ConfigWriteData[20]
rlabel metal1 20332 22746 20332 22746 0 ConfigWriteData[21]
rlabel metal1 21206 22746 21206 22746 0 ConfigWriteData[22]
rlabel metal2 22034 23300 22034 23300 0 ConfigWriteData[23]
rlabel metal1 23092 22746 23092 22746 0 ConfigWriteData[24]
rlabel metal1 24012 22746 24012 22746 0 ConfigWriteData[25]
rlabel metal2 24794 23300 24794 23300 0 ConfigWriteData[26]
rlabel metal1 25852 22746 25852 22746 0 ConfigWriteData[27]
rlabel metal1 26772 22746 26772 22746 0 ConfigWriteData[28]
rlabel metal2 27554 23521 27554 23521 0 ConfigWriteData[29]
rlabel metal2 2714 23300 2714 23300 0 ConfigWriteData[2]
rlabel metal2 28474 23521 28474 23521 0 ConfigWriteData[30]
rlabel metal2 29394 23793 29394 23793 0 ConfigWriteData[31]
rlabel metal1 3772 22746 3772 22746 0 ConfigWriteData[3]
rlabel metal1 4692 22746 4692 22746 0 ConfigWriteData[4]
rlabel metal2 5474 23300 5474 23300 0 ConfigWriteData[5]
rlabel metal1 6578 22746 6578 22746 0 ConfigWriteData[6]
rlabel metal1 7452 22746 7452 22746 0 ConfigWriteData[7]
rlabel metal2 8234 23300 8234 23300 0 ConfigWriteData[8]
rlabel metal1 9292 22746 9292 22746 0 ConfigWriteData[9]
rlabel metal2 30314 23164 30314 23164 0 ConfigWriteStrobe
rlabel metal2 1203 68 1203 68 0 FrameAddressRegister[0]
rlabel metal2 9483 68 9483 68 0 FrameAddressRegister[10]
rlabel metal2 10311 68 10311 68 0 FrameAddressRegister[11]
rlabel metal2 10994 806 10994 806 0 FrameAddressRegister[12]
rlabel metal2 11967 68 11967 68 0 FrameAddressRegister[13]
rlabel metal2 12795 68 12795 68 0 FrameAddressRegister[14]
rlabel metal2 13623 68 13623 68 0 FrameAddressRegister[15]
rlabel metal2 14306 636 14306 636 0 FrameAddressRegister[16]
rlabel metal2 15134 755 15134 755 0 FrameAddressRegister[17]
rlabel metal2 15962 636 15962 636 0 FrameAddressRegister[18]
rlabel metal2 16935 68 16935 68 0 FrameAddressRegister[19]
rlabel metal2 1886 636 1886 636 0 FrameAddressRegister[1]
rlabel metal2 17618 908 17618 908 0 FrameAddressRegister[20]
rlabel metal2 18446 636 18446 636 0 FrameAddressRegister[21]
rlabel metal2 19274 755 19274 755 0 FrameAddressRegister[22]
rlabel metal2 20247 68 20247 68 0 FrameAddressRegister[23]
rlabel metal2 20983 68 20983 68 0 FrameAddressRegister[24]
rlabel metal2 21758 636 21758 636 0 FrameAddressRegister[25]
rlabel metal2 22586 636 22586 636 0 FrameAddressRegister[26]
rlabel metal2 23361 68 23361 68 0 FrameAddressRegister[27]
rlabel metal2 24242 483 24242 483 0 FrameAddressRegister[28]
rlabel metal2 25261 68 25261 68 0 FrameAddressRegister[29]
rlabel metal2 2714 806 2714 806 0 FrameAddressRegister[2]
rlabel metal2 25898 636 25898 636 0 FrameAddressRegister[30]
rlabel metal2 26917 68 26917 68 0 FrameAddressRegister[31]
rlabel metal2 3542 636 3542 636 0 FrameAddressRegister[3]
rlabel metal2 4515 68 4515 68 0 FrameAddressRegister[4]
rlabel metal2 5343 68 5343 68 0 FrameAddressRegister[5]
rlabel metal2 6026 636 6026 636 0 FrameAddressRegister[6]
rlabel metal2 6854 806 6854 806 0 FrameAddressRegister[7]
rlabel metal2 7827 68 7827 68 0 FrameAddressRegister[8]
rlabel metal2 8655 68 8655 68 0 FrameAddressRegister[9]
rlabel metal1 31418 11526 31418 11526 0 INST_config_UART.ByteWriteStrobe
rlabel metal1 19642 17612 19642 17612 0 INST_config_UART.CRCReg\[0\]
rlabel metal2 16606 20332 16606 20332 0 INST_config_UART.CRCReg\[10\]
rlabel metal1 16859 19686 16859 19686 0 INST_config_UART.CRCReg\[11\]
rlabel metal1 14743 19142 14743 19142 0 INST_config_UART.CRCReg\[12\]
rlabel metal1 14421 18598 14421 18598 0 INST_config_UART.CRCReg\[13\]
rlabel metal1 15801 17782 15801 17782 0 INST_config_UART.CRCReg\[14\]
rlabel metal1 16215 18054 16215 18054 0 INST_config_UART.CRCReg\[15\]
rlabel metal1 17848 15470 17848 15470 0 INST_config_UART.CRCReg\[16\]
rlabel metal1 17296 15878 17296 15878 0 INST_config_UART.CRCReg\[17\]
rlabel metal1 17342 16116 17342 16116 0 INST_config_UART.CRCReg\[18\]
rlabel metal1 15824 17102 15824 17102 0 INST_config_UART.CRCReg\[19\]
rlabel metal1 20010 16762 20010 16762 0 INST_config_UART.CRCReg\[1\]
rlabel metal2 21436 18258 21436 18258 0 INST_config_UART.CRCReg\[2\]
rlabel metal2 21206 19057 21206 19057 0 INST_config_UART.CRCReg\[3\]
rlabel metal1 21252 21862 21252 21862 0 INST_config_UART.CRCReg\[4\]
rlabel metal1 21620 20774 21620 20774 0 INST_config_UART.CRCReg\[5\]
rlabel metal1 19182 21930 19182 21930 0 INST_config_UART.CRCReg\[6\]
rlabel metal1 18676 20774 18676 20774 0 INST_config_UART.CRCReg\[7\]
rlabel metal1 16008 21998 16008 21998 0 INST_config_UART.CRCReg\[8\]
rlabel metal1 15640 21488 15640 21488 0 INST_config_UART.CRCReg\[9\]
rlabel metal2 20470 5474 20470 5474 0 INST_config_UART.ComCount\[0\]
rlabel metal1 17250 7514 17250 7514 0 INST_config_UART.ComCount\[10\]
rlabel metal1 18078 7344 18078 7344 0 INST_config_UART.ComCount\[11\]
rlabel metal2 20930 4794 20930 4794 0 INST_config_UART.ComCount\[1\]
rlabel metal1 20746 6154 20746 6154 0 INST_config_UART.ComCount\[2\]
rlabel metal1 18400 5338 18400 5338 0 INST_config_UART.ComCount\[3\]
rlabel metal2 17710 4964 17710 4964 0 INST_config_UART.ComCount\[4\]
rlabel metal1 17894 5678 17894 5678 0 INST_config_UART.ComCount\[5\]
rlabel metal2 15870 5202 15870 5202 0 INST_config_UART.ComCount\[6\]
rlabel metal2 16146 6137 16146 6137 0 INST_config_UART.ComCount\[7\]
rlabel metal2 16238 6154 16238 6154 0 INST_config_UART.ComCount\[8\]
rlabel metal1 15686 7480 15686 7480 0 INST_config_UART.ComCount\[9\]
rlabel metal1 23782 9588 23782 9588 0 INST_config_UART.ComState\[0\]
rlabel via1 23414 7174 23414 7174 0 INST_config_UART.ComState\[10\]
rlabel metal1 22356 8466 22356 8466 0 INST_config_UART.ComState\[1\]
rlabel metal1 20792 8534 20792 8534 0 INST_config_UART.ComState\[2\]
rlabel metal1 21758 10098 21758 10098 0 INST_config_UART.ComState\[3\]
rlabel metal1 20608 13702 20608 13702 0 INST_config_UART.ComState\[4\]
rlabel metal1 23690 8466 23690 8466 0 INST_config_UART.ComState\[5\]
rlabel metal1 19504 9622 19504 9622 0 INST_config_UART.ComState\[6\]
rlabel metal1 19320 9894 19320 9894 0 INST_config_UART.ComState\[7\]
rlabel metal1 22494 8024 22494 8024 0 INST_config_UART.ComState\[8\]
rlabel metal1 20102 8398 20102 8398 0 INST_config_UART.ComState\[9\]
rlabel metal1 22287 9622 22287 9622 0 INST_config_UART.ComTick
rlabel via1 33074 12614 33074 12614 0 INST_config_UART.Command\[0\]
rlabel metal2 32614 13702 32614 13702 0 INST_config_UART.Command\[1\]
rlabel metal1 34822 10778 34822 10778 0 INST_config_UART.Command\[2\]
rlabel metal1 35098 10234 35098 10234 0 INST_config_UART.Command\[3\]
rlabel metal1 34684 12206 34684 12206 0 INST_config_UART.Command\[4\]
rlabel metal1 35466 13158 35466 13158 0 INST_config_UART.Command\[5\]
rlabel metal1 35052 12954 35052 12954 0 INST_config_UART.Command\[6\]
rlabel metal2 24334 19346 24334 19346 0 INST_config_UART.Command\[7\]
rlabel metal1 28423 12886 28423 12886 0 INST_config_UART.Data_Reg\[0\]
rlabel metal1 27416 14382 27416 14382 0 INST_config_UART.Data_Reg\[1\]
rlabel metal1 28106 16218 28106 16218 0 INST_config_UART.Data_Reg\[2\]
rlabel metal1 28980 14790 28980 14790 0 INST_config_UART.Data_Reg\[3\]
rlabel metal1 29348 16558 29348 16558 0 INST_config_UART.Data_Reg\[4\]
rlabel metal1 27922 17850 27922 17850 0 INST_config_UART.Data_Reg\[5\]
rlabel metal1 28060 18258 28060 18258 0 INST_config_UART.Data_Reg\[6\]
rlabel metal1 29670 14246 29670 14246 0 INST_config_UART.Data_Reg\[7\]
rlabel via1 33994 6970 33994 6970 0 INST_config_UART.GetWordState\[0\]
rlabel metal1 33074 16966 33074 16966 0 INST_config_UART.GetWordState\[1\]
rlabel metal1 30314 10472 30314 10472 0 INST_config_UART.GetWordState\[2\]
rlabel metal1 29854 11730 29854 11730 0 INST_config_UART.GetWordState\[3\]
rlabel metal1 26450 12954 26450 12954 0 INST_config_UART.HexData\[0\]
rlabel metal2 26634 13872 26634 13872 0 INST_config_UART.HexData\[1\]
rlabel metal1 25990 15912 25990 15912 0 INST_config_UART.HexData\[2\]
rlabel metal1 26956 15334 26956 15334 0 INST_config_UART.HexData\[3\]
rlabel metal1 26818 17544 26818 17544 0 INST_config_UART.HexData\[4\]
rlabel metal1 28014 18938 28014 18938 0 INST_config_UART.HexData\[5\]
rlabel metal1 25438 19346 25438 19346 0 INST_config_UART.HexData\[6\]
rlabel metal1 27094 14246 27094 14246 0 INST_config_UART.HexData\[7\]
rlabel metal2 28106 11968 28106 11968 0 INST_config_UART.HexWriteStrobe
rlabel metal1 24288 17578 24288 17578 0 INST_config_UART.HighReg\[0\]
rlabel metal1 23966 19482 23966 19482 0 INST_config_UART.HighReg\[1\]
rlabel metal2 25162 18734 25162 18734 0 INST_config_UART.HighReg\[2\]
rlabel metal1 23782 16490 23782 16490 0 INST_config_UART.HighReg\[3\]
rlabel metal1 38180 16014 38180 16014 0 INST_config_UART.ID_Reg\[0\]
rlabel metal2 39238 13192 39238 13192 0 INST_config_UART.ID_Reg\[10\]
rlabel metal2 39790 13566 39790 13566 0 INST_config_UART.ID_Reg\[11\]
rlabel metal1 42182 13872 42182 13872 0 INST_config_UART.ID_Reg\[12\]
rlabel metal2 39698 13940 39698 13940 0 INST_config_UART.ID_Reg\[13\]
rlabel metal1 36662 13974 36662 13974 0 INST_config_UART.ID_Reg\[14\]
rlabel metal1 36662 13906 36662 13906 0 INST_config_UART.ID_Reg\[15\]
rlabel metal1 38180 12206 38180 12206 0 INST_config_UART.ID_Reg\[16\]
rlabel metal1 37858 12954 37858 12954 0 INST_config_UART.ID_Reg\[17\]
rlabel metal1 39606 11526 39606 11526 0 INST_config_UART.ID_Reg\[18\]
rlabel metal1 40503 12138 40503 12138 0 INST_config_UART.ID_Reg\[19\]
rlabel metal2 37674 15232 37674 15232 0 INST_config_UART.ID_Reg\[1\]
rlabel metal1 39698 10778 39698 10778 0 INST_config_UART.ID_Reg\[20\]
rlabel metal1 40664 10982 40664 10982 0 INST_config_UART.ID_Reg\[21\]
rlabel metal2 36110 10557 36110 10557 0 INST_config_UART.ID_Reg\[22\]
rlabel metal2 36294 10336 36294 10336 0 INST_config_UART.ID_Reg\[23\]
rlabel metal1 39330 16966 39330 16966 0 INST_config_UART.ID_Reg\[2\]
rlabel metal1 39238 15878 39238 15878 0 INST_config_UART.ID_Reg\[3\]
rlabel metal1 40434 16218 40434 16218 0 INST_config_UART.ID_Reg\[4\]
rlabel metal1 40526 17238 40526 17238 0 INST_config_UART.ID_Reg\[5\]
rlabel metal1 36110 16422 36110 16422 0 INST_config_UART.ID_Reg\[6\]
rlabel metal2 35742 15266 35742 15266 0 INST_config_UART.ID_Reg\[7\]
rlabel metal1 34914 15130 34914 15130 0 INST_config_UART.ID_Reg\[8\]
rlabel metal1 35696 15130 35696 15130 0 INST_config_UART.ID_Reg\[9\]
rlabel metal2 27922 11730 27922 11730 0 INST_config_UART.LocalWriteStrobe
rlabel metal1 17411 12954 17411 12954 0 INST_config_UART.PresentState\[0\]
rlabel metal1 20056 14042 20056 14042 0 INST_config_UART.PresentState\[1\]
rlabel metal1 19918 12716 19918 12716 0 INST_config_UART.PresentState\[2\]
rlabel metal1 19366 11662 19366 11662 0 INST_config_UART.PresentState\[4\]
rlabel via2 21942 13379 21942 13379 0 INST_config_UART.PresentState\[5\]
rlabel metal1 19688 14382 19688 14382 0 INST_config_UART.PresentState\[6\]
rlabel metal1 16744 9350 16744 9350 0 INST_config_UART.ReceiveLED
rlabel metal1 21574 15028 21574 15028 0 INST_config_UART.ReceiveState
rlabel metal2 24426 11662 24426 11662 0 INST_config_UART.ReceivedWord\[0\]
rlabel metal1 21666 14382 21666 14382 0 INST_config_UART.ReceivedWord\[1\]
rlabel metal1 22908 11118 22908 11118 0 INST_config_UART.ReceivedWord\[2\]
rlabel metal2 24150 13192 24150 13192 0 INST_config_UART.ReceivedWord\[3\]
rlabel metal2 42274 14824 42274 14824 0 INST_config_UART.ReceivedWord\[4\]
rlabel metal1 44114 14586 44114 14586 0 INST_config_UART.ReceivedWord\[5\]
rlabel metal1 44390 16626 44390 16626 0 INST_config_UART.ReceivedWord\[6\]
rlabel metal2 24426 9792 24426 9792 0 INST_config_UART.ReceivedWord\[7\]
rlabel metal1 16560 12410 16560 12410 0 INST_config_UART.RxLocal
rlabel metal1 17120 12342 17120 12342 0 INST_config_UART.TimeToSend
rlabel metal1 8878 9894 8878 9894 0 INST_config_UART.TimeToSendCounter\[0\]
rlabel metal2 14950 8160 14950 8160 0 INST_config_UART.TimeToSendCounter\[10\]
rlabel metal1 14674 8296 14674 8296 0 INST_config_UART.TimeToSendCounter\[11\]
rlabel metal2 14030 9146 14030 9146 0 INST_config_UART.TimeToSendCounter\[12\]
rlabel metal1 14122 11084 14122 11084 0 INST_config_UART.TimeToSendCounter\[13\]
rlabel metal1 13846 11118 13846 11118 0 INST_config_UART.TimeToSendCounter\[14\]
rlabel metal1 9108 11050 9108 11050 0 INST_config_UART.TimeToSendCounter\[1\]
rlabel metal1 9890 10234 9890 10234 0 INST_config_UART.TimeToSendCounter\[2\]
rlabel metal2 10442 9996 10442 9996 0 INST_config_UART.TimeToSendCounter\[3\]
rlabel metal1 10718 7310 10718 7310 0 INST_config_UART.TimeToSendCounter\[4\]
rlabel metal1 10672 7514 10672 7514 0 INST_config_UART.TimeToSendCounter\[5\]
rlabel metal2 11822 7548 11822 7548 0 INST_config_UART.TimeToSendCounter\[6\]
rlabel metal1 10718 10574 10718 10574 0 INST_config_UART.TimeToSendCounter\[7\]
rlabel metal1 11868 9894 11868 9894 0 INST_config_UART.TimeToSendCounter\[8\]
rlabel metal1 12466 9588 12466 9588 0 INST_config_UART.TimeToSendCounter\[9\]
rlabel metal1 27784 20026 27784 20026 0 INST_config_UART.WriteData\[0\]
rlabel metal1 33534 19482 33534 19482 0 INST_config_UART.WriteData\[10\]
rlabel metal1 32108 18938 32108 18938 0 INST_config_UART.WriteData\[11\]
rlabel metal1 33350 17850 33350 17850 0 INST_config_UART.WriteData\[12\]
rlabel metal1 32108 17102 32108 17102 0 INST_config_UART.WriteData\[13\]
rlabel metal1 33120 15878 33120 15878 0 INST_config_UART.WriteData\[14\]
rlabel metal1 32660 15334 32660 15334 0 INST_config_UART.WriteData\[15\]
rlabel metal1 32798 10098 32798 10098 0 INST_config_UART.WriteData\[16\]
rlabel metal1 33028 10506 33028 10506 0 INST_config_UART.WriteData\[17\]
rlabel metal1 30820 8806 30820 8806 0 INST_config_UART.WriteData\[18\]
rlabel metal2 28934 6800 28934 6800 0 INST_config_UART.WriteData\[19\]
rlabel metal2 28106 20502 28106 20502 0 INST_config_UART.WriteData\[1\]
rlabel metal1 28474 6698 28474 6698 0 INST_config_UART.WriteData\[20\]
rlabel metal2 30406 5576 30406 5576 0 INST_config_UART.WriteData\[21\]
rlabel metal1 31096 6426 31096 6426 0 INST_config_UART.WriteData\[22\]
rlabel via1 31786 5882 31786 5882 0 INST_config_UART.WriteData\[23\]
rlabel metal1 33074 4998 33074 4998 0 INST_config_UART.WriteData\[24\]
rlabel metal1 34086 5338 34086 5338 0 INST_config_UART.WriteData\[25\]
rlabel metal2 33442 5100 33442 5100 0 INST_config_UART.WriteData\[26\]
rlabel metal1 28520 7514 28520 7514 0 INST_config_UART.WriteData\[27\]
rlabel metal1 32660 7514 32660 7514 0 INST_config_UART.WriteData\[28\]
rlabel metal1 27830 8058 27830 8058 0 INST_config_UART.WriteData\[29\]
rlabel metal1 29302 21522 29302 21522 0 INST_config_UART.WriteData\[2\]
rlabel metal1 33396 8058 33396 8058 0 INST_config_UART.WriteData\[30\]
rlabel metal1 33672 8602 33672 8602 0 INST_config_UART.WriteData\[31\]
rlabel metal1 30636 21046 30636 21046 0 INST_config_UART.WriteData\[3\]
rlabel metal2 30682 20740 30682 20740 0 INST_config_UART.WriteData\[4\]
rlabel metal1 30314 17850 30314 17850 0 INST_config_UART.WriteData\[5\]
rlabel metal1 30912 18190 30912 18190 0 INST_config_UART.WriteData\[6\]
rlabel metal1 30682 16218 30682 16218 0 INST_config_UART.WriteData\[7\]
rlabel metal1 30866 14484 30866 14484 0 INST_config_UART.WriteData\[8\]
rlabel metal1 33028 18802 33028 18802 0 INST_config_UART.WriteData\[9\]
rlabel metal1 27370 8942 27370 8942 0 INST_config_UART.WriteStrobe
rlabel metal1 28244 11322 28244 11322 0 INST_config_UART._0000_
rlabel metal1 20010 5746 20010 5746 0 INST_config_UART._0001_
rlabel via1 15873 7718 15873 7718 0 INST_config_UART._0002_
rlabel metal1 16606 7922 16606 7922 0 INST_config_UART._0003_
rlabel metal1 18998 5814 18998 5814 0 INST_config_UART._0004_
rlabel metal2 18998 5950 18998 5950 0 INST_config_UART._0005_
rlabel metal1 17756 4794 17756 4794 0 INST_config_UART._0006_
rlabel metal2 16698 4522 16698 4522 0 INST_config_UART._0007_
rlabel metal1 16836 4522 16836 4522 0 INST_config_UART._0008_
rlabel metal1 14720 4250 14720 4250 0 INST_config_UART._0009_
rlabel metal1 14628 5882 14628 5882 0 INST_config_UART._0010_
rlabel metal1 14904 6222 14904 6222 0 INST_config_UART._0011_
rlabel via1 15127 6970 15127 6970 0 INST_config_UART._0012_
rlabel metal1 18676 7514 18676 7514 0 INST_config_UART._0013_
rlabel metal1 26266 12750 26266 12750 0 INST_config_UART._0014_
rlabel metal1 26726 11186 26726 11186 0 INST_config_UART._0015_
rlabel metal1 20240 14382 20240 14382 0 INST_config_UART._0016_
rlabel metal1 27370 19380 27370 19380 0 INST_config_UART._0017_
rlabel metal1 20884 12954 20884 12954 0 INST_config_UART._0018_
rlabel metal2 19550 10914 19550 10914 0 INST_config_UART._0019_
rlabel metal1 17848 8534 17848 8534 0 INST_config_UART._0020_
rlabel metal2 28014 9724 28014 9724 0 INST_config_UART._0021_
rlabel metal1 30268 12614 30268 12614 0 INST_config_UART._0022_
rlabel metal1 29026 10166 29026 10166 0 INST_config_UART._0023_
rlabel metal1 30958 11594 30958 11594 0 INST_config_UART._0024_
rlabel metal1 18538 12342 18538 12342 0 INST_config_UART._0025_
rlabel metal1 18676 13974 18676 13974 0 INST_config_UART._0026_
rlabel metal1 19136 13430 19136 13430 0 INST_config_UART._0027_
rlabel metal1 24472 11798 24472 11798 0 INST_config_UART._0028_
rlabel metal1 17802 11832 17802 11832 0 INST_config_UART._0029_
rlabel metal2 18262 13294 18262 13294 0 INST_config_UART._0030_
rlabel metal1 3404 10234 3404 10234 0 INST_config_UART._0031_
rlabel metal1 5244 16218 5244 16218 0 INST_config_UART._0032_
rlabel metal2 4094 17221 4094 17221 0 INST_config_UART._0033_
rlabel metal1 4094 18360 4094 18360 0 INST_config_UART._0034_
rlabel metal1 5198 17714 5198 17714 0 INST_config_UART._0035_
rlabel metal1 6854 17306 6854 17306 0 INST_config_UART._0036_
rlabel metal1 7038 18360 7038 18360 0 INST_config_UART._0037_
rlabel metal1 8602 18326 8602 18326 0 INST_config_UART._0038_
rlabel metal1 8408 18938 8408 18938 0 INST_config_UART._0039_
rlabel metal1 9062 19414 9062 19414 0 INST_config_UART._0040_
rlabel metal1 10350 18938 10350 18938 0 INST_config_UART._0041_
rlabel metal1 4278 9622 4278 9622 0 INST_config_UART._0042_
rlabel metal1 11401 19142 11401 19142 0 INST_config_UART._0043_
rlabel metal2 11638 18530 11638 18530 0 INST_config_UART._0044_
rlabel metal1 13018 17272 13018 17272 0 INST_config_UART._0045_
rlabel metal1 4416 8874 4416 8874 0 INST_config_UART._0046_
rlabel metal1 5336 10098 5336 10098 0 INST_config_UART._0047_
rlabel metal1 5888 11798 5888 11798 0 INST_config_UART._0048_
rlabel metal1 5566 12104 5566 12104 0 INST_config_UART._0049_
rlabel metal1 5428 12886 5428 12886 0 INST_config_UART._0050_
rlabel metal1 5290 14280 5290 14280 0 INST_config_UART._0051_
rlabel metal1 6026 15096 6026 15096 0 INST_config_UART._0052_
rlabel metal1 5198 15402 5198 15402 0 INST_config_UART._0053_
rlabel metal1 26082 10098 26082 10098 0 INST_config_UART._0054_
rlabel metal1 21344 11866 21344 11866 0 INST_config_UART._0055_
rlabel metal1 27232 19482 27232 19482 0 INST_config_UART._0056_
rlabel metal1 28152 19958 28152 19958 0 INST_config_UART._0057_
rlabel metal1 28612 20502 28612 20502 0 INST_config_UART._0058_
rlabel metal2 32062 20519 32062 20519 0 INST_config_UART._0059_
rlabel metal1 31326 19992 31326 19992 0 INST_config_UART._0060_
rlabel metal1 29900 17714 29900 17714 0 INST_config_UART._0061_
rlabel metal1 29532 18326 29532 18326 0 INST_config_UART._0062_
rlabel metal1 29992 15674 29992 15674 0 INST_config_UART._0063_
rlabel metal1 30866 10098 30866 10098 0 INST_config_UART._0064_
rlabel metal1 31786 10744 31786 10744 0 INST_config_UART._0065_
rlabel metal1 30038 8602 30038 8602 0 INST_config_UART._0066_
rlabel metal1 28750 7480 28750 7480 0 INST_config_UART._0067_
rlabel metal1 28704 6834 28704 6834 0 INST_config_UART._0068_
rlabel metal1 29992 4998 29992 4998 0 INST_config_UART._0069_
rlabel metal1 29854 6392 29854 6392 0 INST_config_UART._0070_
rlabel metal1 30958 5746 30958 5746 0 INST_config_UART._0071_
rlabel metal1 30215 13702 30215 13702 0 INST_config_UART._0072_
rlabel metal1 32614 18360 32614 18360 0 INST_config_UART._0073_
rlabel metal1 32936 19278 32936 19278 0 INST_config_UART._0074_
rlabel metal1 31142 18394 31142 18394 0 INST_config_UART._0075_
rlabel metal2 32246 18564 32246 18564 0 INST_config_UART._0076_
rlabel metal1 31326 16626 31326 16626 0 INST_config_UART._0077_
rlabel metal2 32706 15572 32706 15572 0 INST_config_UART._0078_
rlabel metal1 32016 15538 32016 15538 0 INST_config_UART._0079_
rlabel metal1 24472 7922 24472 7922 0 INST_config_UART._0080_
rlabel metal1 20700 11866 20700 11866 0 INST_config_UART._0081_
rlabel metal1 36846 11662 36846 11662 0 INST_config_UART._0082_
rlabel metal1 36570 11526 36570 11526 0 INST_config_UART._0083_
rlabel metal1 37582 11322 37582 11322 0 INST_config_UART._0084_
rlabel metal1 39422 10234 39422 10234 0 INST_config_UART._0085_
rlabel metal1 38134 10744 38134 10744 0 INST_config_UART._0086_
rlabel metal1 38824 10166 38824 10166 0 INST_config_UART._0087_
rlabel metal1 36662 10744 36662 10744 0 INST_config_UART._0088_
rlabel metal1 34960 9622 34960 9622 0 INST_config_UART._0089_
rlabel metal1 23138 10234 23138 10234 0 INST_config_UART._0090_
rlabel metal2 24426 7956 24426 7956 0 INST_config_UART._0091_
rlabel metal2 22034 11492 22034 11492 0 INST_config_UART._0092_
rlabel metal1 33580 15674 33580 15674 0 INST_config_UART._0093_
rlabel metal1 33902 15402 33902 15402 0 INST_config_UART._0094_
rlabel metal1 37812 13974 37812 13974 0 INST_config_UART._0095_
rlabel metal1 39790 12954 39790 12954 0 INST_config_UART._0096_
rlabel metal1 40342 14042 40342 14042 0 INST_config_UART._0097_
rlabel metal1 38870 12716 38870 12716 0 INST_config_UART._0098_
rlabel metal1 36294 14246 36294 14246 0 INST_config_UART._0099_
rlabel metal1 35558 12954 35558 12954 0 INST_config_UART._0100_
rlabel metal1 22862 17272 22862 17272 0 INST_config_UART._0101_
rlabel metal1 22770 18122 22770 18122 0 INST_config_UART._0102_
rlabel metal1 22862 18326 22862 18326 0 INST_config_UART._0103_
rlabel metal1 24196 15130 24196 15130 0 INST_config_UART._0104_
rlabel metal1 15676 12206 15676 12206 0 INST_config_UART._0105_
rlabel metal1 25714 12274 25714 12274 0 INST_config_UART._0106_
rlabel metal1 25806 13362 25806 13362 0 INST_config_UART._0107_
rlabel metal1 24656 16150 24656 16150 0 INST_config_UART._0108_
rlabel metal2 26634 15334 26634 15334 0 INST_config_UART._0109_
rlabel metal1 25070 17578 25070 17578 0 INST_config_UART._0110_
rlabel metal1 26496 18802 26496 18802 0 INST_config_UART._0111_
rlabel metal1 25208 18394 25208 18394 0 INST_config_UART._0112_
rlabel metal1 25622 14450 25622 14450 0 INST_config_UART._0113_
rlabel metal1 7774 9078 7774 9078 0 INST_config_UART._0114_
rlabel metal1 8234 9622 8234 9622 0 INST_config_UART._0115_
rlabel metal1 8556 9962 8556 9962 0 INST_config_UART._0116_
rlabel metal1 9614 10574 9614 10574 0 INST_config_UART._0117_
rlabel metal1 9108 8534 9108 8534 0 INST_config_UART._0118_
rlabel metal2 9982 8194 9982 8194 0 INST_config_UART._0119_
rlabel metal1 10626 7922 10626 7922 0 INST_config_UART._0120_
rlabel metal1 11316 10710 11316 10710 0 INST_config_UART._0121_
rlabel metal1 11224 10098 11224 10098 0 INST_config_UART._0122_
rlabel metal1 11868 8330 11868 8330 0 INST_config_UART._0123_
rlabel metal1 13754 7752 13754 7752 0 INST_config_UART._0124_
rlabel metal1 13478 9078 13478 9078 0 INST_config_UART._0125_
rlabel metal1 13064 10166 13064 10166 0 INST_config_UART._0126_
rlabel metal1 13340 10574 13340 10574 0 INST_config_UART._0127_
rlabel metal1 13018 11322 13018 11322 0 INST_config_UART._0128_
rlabel metal1 16647 9622 16647 9622 0 INST_config_UART._0129_
rlabel metal1 31786 5304 31786 5304 0 INST_config_UART._0130_
rlabel metal1 33212 4658 33212 4658 0 INST_config_UART._0131_
rlabel metal2 33258 6052 33258 6052 0 INST_config_UART._0132_
rlabel metal1 27554 7310 27554 7310 0 INST_config_UART._0133_
rlabel metal1 31809 7446 31809 7446 0 INST_config_UART._0134_
rlabel metal1 27324 7922 27324 7922 0 INST_config_UART._0135_
rlabel metal1 32338 7922 32338 7922 0 INST_config_UART._0136_
rlabel metal1 32798 8568 32798 8568 0 INST_config_UART._0137_
rlabel metal2 18446 16592 18446 16592 0 INST_config_UART._0138_
rlabel metal1 19228 16626 19228 16626 0 INST_config_UART._0139_
rlabel metal1 19412 18190 19412 18190 0 INST_config_UART._0140_
rlabel metal1 20788 18666 20788 18666 0 INST_config_UART._0141_
rlabel metal1 19780 21658 19780 21658 0 INST_config_UART._0142_
rlabel metal1 20746 20808 20746 20808 0 INST_config_UART._0143_
rlabel metal1 18722 21862 18722 21862 0 INST_config_UART._0144_
rlabel metal1 18630 21012 18630 21012 0 INST_config_UART._0145_
rlabel metal1 15410 21658 15410 21658 0 INST_config_UART._0146_
rlabel metal1 14674 20298 14674 20298 0 INST_config_UART._0147_
rlabel metal1 17020 20570 17020 20570 0 INST_config_UART._0148_
rlabel metal1 15778 19890 15778 19890 0 INST_config_UART._0149_
rlabel metal1 15732 18938 15732 18938 0 INST_config_UART._0150_
rlabel metal1 14122 18802 14122 18802 0 INST_config_UART._0151_
rlabel metal1 14490 17714 14490 17714 0 INST_config_UART._0152_
rlabel metal1 14076 18258 14076 18258 0 INST_config_UART._0153_
rlabel metal1 17250 15402 17250 15402 0 INST_config_UART._0154_
rlabel metal2 15410 14892 15410 14892 0 INST_config_UART._0155_
rlabel metal1 17158 16626 17158 16626 0 INST_config_UART._0156_
rlabel metal2 15318 16422 15318 16422 0 INST_config_UART._0157_
rlabel metal1 23818 10234 23818 10234 0 INST_config_UART._0158_
rlabel metal1 36800 16150 36800 16150 0 INST_config_UART._0159_
rlabel metal1 36386 15130 36386 15130 0 INST_config_UART._0160_
rlabel metal1 37996 16762 37996 16762 0 INST_config_UART._0161_
rlabel metal1 38686 16014 38686 16014 0 INST_config_UART._0162_
rlabel metal1 40020 15538 40020 15538 0 INST_config_UART._0163_
rlabel metal1 39330 16626 39330 16626 0 INST_config_UART._0164_
rlabel metal1 34730 17272 34730 17272 0 INST_config_UART._0165_
rlabel metal1 36110 16218 36110 16218 0 INST_config_UART._0166_
rlabel metal1 31786 12920 31786 12920 0 INST_config_UART._0167_
rlabel metal1 30820 13226 30820 13226 0 INST_config_UART._0168_
rlabel metal1 33764 10710 33764 10710 0 INST_config_UART._0169_
rlabel metal1 34076 10098 34076 10098 0 INST_config_UART._0170_
rlabel metal1 33166 14008 33166 14008 0 INST_config_UART._0171_
rlabel metal2 34362 13872 34362 13872 0 INST_config_UART._0172_
rlabel metal1 33580 12886 33580 12886 0 INST_config_UART._0173_
rlabel metal1 22816 15130 22816 15130 0 INST_config_UART._0174_
rlabel metal1 27871 13294 27871 13294 0 INST_config_UART._0175_
rlabel metal1 26767 13974 26767 13974 0 INST_config_UART._0176_
rlabel metal1 27170 16150 27170 16150 0 INST_config_UART._0177_
rlabel metal2 29670 14246 29670 14246 0 INST_config_UART._0178_
rlabel metal1 28428 16762 28428 16762 0 INST_config_UART._0179_
rlabel via1 27176 17646 27176 17646 0 INST_config_UART._0180_
rlabel metal1 26618 17238 26618 17238 0 INST_config_UART._0181_
rlabel metal1 29108 14382 29108 14382 0 INST_config_UART._0182_
rlabel metal1 22724 6358 22724 6358 0 INST_config_UART._0183_
rlabel metal2 18262 8534 18262 8534 0 INST_config_UART._0184_
rlabel metal2 20654 7446 20654 7446 0 INST_config_UART._0185_
rlabel metal1 21206 9010 21206 9010 0 INST_config_UART._0186_
rlabel metal1 22724 7446 22724 7446 0 INST_config_UART._0187_
rlabel metal1 17618 10234 17618 10234 0 INST_config_UART._0188_
rlabel metal1 17756 9622 17756 9622 0 INST_config_UART._0189_
rlabel metal1 19366 7480 19366 7480 0 INST_config_UART._0190_
rlabel metal2 21574 6562 21574 6562 0 INST_config_UART._0191_
rlabel metal1 20332 12614 20332 12614 0 INST_config_UART._0192_
rlabel metal1 26696 12886 26696 12886 0 INST_config_UART._0193_
rlabel metal1 18262 12172 18262 12172 0 INST_config_UART._0194_
rlabel metal1 20240 11594 20240 11594 0 INST_config_UART._0195_
rlabel metal1 18814 14416 18814 14416 0 INST_config_UART._0196_
rlabel metal1 18998 10166 18998 10166 0 INST_config_UART._0197_
rlabel metal1 18998 11118 18998 11118 0 INST_config_UART._0198_
rlabel metal1 18952 11322 18952 11322 0 INST_config_UART._0199_
rlabel metal1 33718 12172 33718 12172 0 INST_config_UART._0200_
rlabel metal2 36478 11424 36478 11424 0 INST_config_UART._0201_
rlabel metal1 35006 12070 35006 12070 0 INST_config_UART._0202_
rlabel metal1 36524 14518 36524 14518 0 INST_config_UART._0203_
rlabel metal1 39928 12886 39928 12886 0 INST_config_UART._0204_
rlabel metal1 38932 15402 38932 15402 0 INST_config_UART._0205_
rlabel metal1 37720 14314 37720 14314 0 INST_config_UART._0206_
rlabel metal1 39882 13362 39882 13362 0 INST_config_UART._0207_
rlabel metal1 37674 13294 37674 13294 0 INST_config_UART._0208_
rlabel metal1 37582 13498 37582 13498 0 INST_config_UART._0209_
rlabel metal2 37536 14246 37536 14246 0 INST_config_UART._0210_
rlabel metal2 33534 11917 33534 11917 0 INST_config_UART._0211_
rlabel metal1 19964 12954 19964 12954 0 INST_config_UART._0212_
rlabel metal1 18170 14246 18170 14246 0 INST_config_UART._0213_
rlabel metal1 31234 9690 31234 9690 0 INST_config_UART._0214_
rlabel metal1 32522 18870 32522 18870 0 INST_config_UART._0215_
rlabel metal3 33534 9452 33534 9452 0 INST_config_UART._0216_
rlabel metal1 31786 11696 31786 11696 0 INST_config_UART._0217_
rlabel metal1 44206 15470 44206 15470 0 INST_config_UART._0218_
rlabel metal1 21896 14314 21896 14314 0 INST_config_UART._0219_
rlabel metal1 21528 13906 21528 13906 0 INST_config_UART._0220_
rlabel metal1 43516 17578 43516 17578 0 INST_config_UART._0221_
rlabel metal1 27738 14280 27738 14280 0 INST_config_UART._0222_
rlabel metal1 28336 12954 28336 12954 0 INST_config_UART._0223_
rlabel metal1 22402 13362 22402 13362 0 INST_config_UART._0224_
rlabel metal1 24104 12750 24104 12750 0 INST_config_UART._0225_
rlabel metal1 23092 14790 23092 14790 0 INST_config_UART._0226_
rlabel metal1 23414 13872 23414 13872 0 INST_config_UART._0227_
rlabel metal1 23322 13158 23322 13158 0 INST_config_UART._0228_
rlabel metal1 24610 13906 24610 13906 0 INST_config_UART._0229_
rlabel metal1 24012 12342 24012 12342 0 INST_config_UART._0230_
rlabel metal1 24242 13940 24242 13940 0 INST_config_UART._0231_
rlabel metal1 22678 15470 22678 15470 0 INST_config_UART._0232_
rlabel metal2 22218 14110 22218 14110 0 INST_config_UART._0233_
rlabel metal1 28290 7820 28290 7820 0 INST_config_UART._0234_
rlabel metal1 29486 9146 29486 9146 0 INST_config_UART._0235_
rlabel metal1 30958 10540 30958 10540 0 INST_config_UART._0236_
rlabel metal1 30912 11866 30912 11866 0 INST_config_UART._0237_
rlabel metal1 28520 10234 28520 10234 0 INST_config_UART._0238_
rlabel metal1 29808 10778 29808 10778 0 INST_config_UART._0239_
rlabel metal1 28244 10778 28244 10778 0 INST_config_UART._0240_
rlabel metal1 30130 17204 30130 17204 0 INST_config_UART._0241_
rlabel metal1 26634 8534 26634 8534 0 INST_config_UART._0242_
rlabel metal2 26542 8687 26542 8687 0 INST_config_UART._0243_
rlabel metal1 20424 12886 20424 12886 0 INST_config_UART._0244_
rlabel metal1 20424 10438 20424 10438 0 INST_config_UART._0245_
rlabel metal2 24426 16898 24426 16898 0 INST_config_UART._0246_
rlabel metal1 29946 16626 29946 16626 0 INST_config_UART._0247_
rlabel metal1 27922 11118 27922 11118 0 INST_config_UART._0248_
rlabel metal1 26956 12206 26956 12206 0 INST_config_UART._0249_
rlabel metal1 20976 9894 20976 9894 0 INST_config_UART._0250_
rlabel metal1 21206 6426 21206 6426 0 INST_config_UART._0251_
rlabel metal2 19826 5066 19826 5066 0 INST_config_UART._0252_
rlabel metal1 18768 4590 18768 4590 0 INST_config_UART._0253_
rlabel viali 16882 5678 16882 5678 0 INST_config_UART._0254_
rlabel metal1 16514 5882 16514 5882 0 INST_config_UART._0255_
rlabel metal1 15502 7310 15502 7310 0 INST_config_UART._0256_
rlabel metal2 15870 6902 15870 6902 0 INST_config_UART._0257_
rlabel metal1 16928 6698 16928 6698 0 INST_config_UART._0258_
rlabel metal1 18906 5542 18906 5542 0 INST_config_UART._0259_
rlabel metal1 19826 6732 19826 6732 0 INST_config_UART._0260_
rlabel metal1 18906 5644 18906 5644 0 INST_config_UART._0261_
rlabel metal2 18446 6426 18446 6426 0 INST_config_UART._0262_
rlabel metal1 19642 4556 19642 4556 0 INST_config_UART._0263_
rlabel metal1 19504 5678 19504 5678 0 INST_config_UART._0264_
rlabel metal1 18124 4590 18124 4590 0 INST_config_UART._0265_
rlabel metal1 16514 5134 16514 5134 0 INST_config_UART._0266_
rlabel metal1 16330 5270 16330 5270 0 INST_config_UART._0267_
rlabel metal2 16698 5882 16698 5882 0 INST_config_UART._0268_
rlabel metal1 17434 5712 17434 5712 0 INST_config_UART._0269_
rlabel metal1 14996 4114 14996 4114 0 INST_config_UART._0270_
rlabel metal1 15318 5542 15318 5542 0 INST_config_UART._0271_
rlabel viali 15134 5684 15134 5684 0 INST_config_UART._0272_
rlabel metal2 16790 6358 16790 6358 0 INST_config_UART._0273_
rlabel metal1 15410 7344 15410 7344 0 INST_config_UART._0274_
rlabel metal2 16054 8058 16054 8058 0 INST_config_UART._0275_
rlabel metal2 17250 7548 17250 7548 0 INST_config_UART._0276_
rlabel metal1 19596 13498 19596 13498 0 INST_config_UART._0277_
rlabel metal1 19964 14586 19964 14586 0 INST_config_UART._0278_
rlabel metal1 20884 12818 20884 12818 0 INST_config_UART._0279_
rlabel metal1 5106 10506 5106 10506 0 INST_config_UART._0280_
rlabel metal1 3634 10098 3634 10098 0 INST_config_UART._0281_
rlabel metal1 5431 11730 5431 11730 0 INST_config_UART._0282_
rlabel metal1 5750 10676 5750 10676 0 INST_config_UART._0283_
rlabel metal2 5290 13090 5290 13090 0 INST_config_UART._0284_
rlabel metal1 5106 11696 5106 11696 0 INST_config_UART._0285_
rlabel metal1 4922 12784 4922 12784 0 INST_config_UART._0286_
rlabel metal1 4738 12886 4738 12886 0 INST_config_UART._0287_
rlabel metal1 5704 16082 5704 16082 0 INST_config_UART._0288_
rlabel metal1 4462 14926 4462 14926 0 INST_config_UART._0289_
rlabel metal2 5474 16150 5474 16150 0 INST_config_UART._0290_
rlabel metal1 5290 16116 5290 16116 0 INST_config_UART._0291_
rlabel metal2 4462 18326 4462 18326 0 INST_config_UART._0292_
rlabel metal1 3542 17748 3542 17748 0 INST_config_UART._0293_
rlabel metal1 6394 17306 6394 17306 0 INST_config_UART._0294_
rlabel metal1 5888 18394 5888 18394 0 INST_config_UART._0295_
rlabel metal1 7130 17136 7130 17136 0 INST_config_UART._0296_
rlabel metal2 6946 17884 6946 17884 0 INST_config_UART._0297_
rlabel metal1 7682 18836 7682 18836 0 INST_config_UART._0298_
rlabel metal1 7636 17306 7636 17306 0 INST_config_UART._0299_
rlabel metal1 10442 19312 10442 19312 0 INST_config_UART._0300_
rlabel metal2 9338 18836 9338 18836 0 INST_config_UART._0301_
rlabel metal1 11224 18938 11224 18938 0 INST_config_UART._0302_
rlabel metal1 10396 18734 10396 18734 0 INST_config_UART._0303_
rlabel metal2 12558 17986 12558 17986 0 INST_config_UART._0304_
rlabel metal1 12374 18292 12374 18292 0 INST_config_UART._0305_
rlabel metal1 21528 8874 21528 8874 0 INST_config_UART._0306_
rlabel metal1 24610 9452 24610 9452 0 INST_config_UART._0307_
rlabel metal1 24380 9350 24380 9350 0 INST_config_UART._0308_
rlabel metal1 19780 8534 19780 8534 0 INST_config_UART._0309_
rlabel metal2 20378 10370 20378 10370 0 INST_config_UART._0310_
rlabel metal1 21298 11322 21298 11322 0 INST_config_UART._0311_
rlabel metal1 21850 16490 21850 16490 0 INST_config_UART._0312_
rlabel metal1 29210 12954 29210 12954 0 INST_config_UART._0313_
rlabel via1 34002 9622 34002 9622 0 INST_config_UART._0314_
rlabel metal1 27508 12818 27508 12818 0 INST_config_UART._0315_
rlabel metal3 29394 19380 29394 19380 0 INST_config_UART._0316_
rlabel metal1 28842 16116 28842 16116 0 INST_config_UART._0317_
rlabel via2 34270 18309 34270 18309 0 INST_config_UART._0318_
rlabel metal1 28106 15028 28106 15028 0 INST_config_UART._0319_
rlabel metal2 33534 10047 33534 10047 0 INST_config_UART._0320_
rlabel metal1 30406 16762 30406 16762 0 INST_config_UART._0321_
rlabel metal2 34684 7310 34684 7310 0 INST_config_UART._0322_
rlabel metal1 28336 16558 28336 16558 0 INST_config_UART._0323_
rlabel metal1 30920 8534 30920 8534 0 INST_config_UART._0324_
rlabel viali 29948 17170 29948 17170 0 INST_config_UART._0325_
rlabel via1 36854 9622 36854 9622 0 INST_config_UART._0326_
rlabel metal2 30682 15334 30682 15334 0 INST_config_UART._0327_
rlabel metal1 36494 8874 36494 8874 0 INST_config_UART._0328_
rlabel metal1 33626 9690 33626 9690 0 INST_config_UART._0329_
rlabel metal2 31786 10710 31786 10710 0 INST_config_UART._0330_
rlabel metal1 30636 8466 30636 8466 0 INST_config_UART._0331_
rlabel metal1 29854 7922 29854 7922 0 INST_config_UART._0332_
rlabel metal1 28658 6732 28658 6732 0 INST_config_UART._0333_
rlabel metal1 31234 5236 31234 5236 0 INST_config_UART._0334_
rlabel metal1 35788 8874 35788 8874 0 INST_config_UART._0335_
rlabel metal1 32154 6902 32154 6902 0 INST_config_UART._0336_
rlabel via1 31786 7973 31786 7973 0 INST_config_UART._0337_
rlabel metal1 31326 14450 31326 14450 0 INST_config_UART._0338_
rlabel metal1 33534 9146 33534 9146 0 INST_config_UART._0339_
rlabel metal2 31234 18003 31234 18003 0 INST_config_UART._0340_
rlabel metal2 34546 18836 34546 18836 0 INST_config_UART._0341_
rlabel metal1 31970 18156 31970 18156 0 INST_config_UART._0342_
rlabel metal1 32936 17034 32936 17034 0 INST_config_UART._0343_
rlabel metal1 31556 17306 31556 17306 0 INST_config_UART._0344_
rlabel metal2 33166 15334 33166 15334 0 INST_config_UART._0345_
rlabel metal2 32798 15062 32798 15062 0 INST_config_UART._0346_
rlabel metal1 22586 7718 22586 7718 0 INST_config_UART._0347_
rlabel metal1 23782 7922 23782 7922 0 INST_config_UART._0348_
rlabel metal1 24380 8058 24380 8058 0 INST_config_UART._0349_
rlabel metal1 19274 8976 19274 8976 0 INST_config_UART._0350_
rlabel metal2 25254 8772 25254 8772 0 INST_config_UART._0351_
rlabel metal1 20608 10166 20608 10166 0 INST_config_UART._0352_
rlabel metal1 20976 11322 20976 11322 0 INST_config_UART._0353_
rlabel metal1 20516 10234 20516 10234 0 INST_config_UART._0354_
rlabel via2 20010 11611 20010 11611 0 INST_config_UART._0355_
rlabel metal2 38870 11254 38870 11254 0 INST_config_UART._0356_
rlabel metal1 36110 11798 36110 11798 0 INST_config_UART._0357_
rlabel metal1 36386 11764 36386 11764 0 INST_config_UART._0358_
rlabel metal1 37858 11118 37858 11118 0 INST_config_UART._0359_
rlabel metal1 39100 10030 39100 10030 0 INST_config_UART._0360_
rlabel metal1 37628 10642 37628 10642 0 INST_config_UART._0361_
rlabel metal1 38778 10064 38778 10064 0 INST_config_UART._0362_
rlabel metal1 36846 10574 36846 10574 0 INST_config_UART._0363_
rlabel metal2 35926 10982 35926 10982 0 INST_config_UART._0364_
rlabel metal1 23322 9690 23322 9690 0 INST_config_UART._0365_
rlabel metal1 23690 10098 23690 10098 0 INST_config_UART._0366_
rlabel metal2 23322 9369 23322 9369 0 INST_config_UART._0367_
rlabel metal1 23874 8398 23874 8398 0 INST_config_UART._0368_
rlabel metal1 24472 7174 24472 7174 0 INST_config_UART._0369_
rlabel metal1 24610 7446 24610 7446 0 INST_config_UART._0370_
rlabel metal2 22494 10438 22494 10438 0 INST_config_UART._0371_
rlabel metal1 22540 10778 22540 10778 0 INST_config_UART._0372_
rlabel metal2 22218 10948 22218 10948 0 INST_config_UART._0373_
rlabel metal1 28474 12240 28474 12240 0 INST_config_UART._0374_
rlabel metal1 42366 13770 42366 13770 0 INST_config_UART._0375_
rlabel metal1 34132 15130 34132 15130 0 INST_config_UART._0376_
rlabel metal1 35282 15130 35282 15130 0 INST_config_UART._0377_
rlabel metal1 38088 13498 38088 13498 0 INST_config_UART._0378_
rlabel metal1 40204 12818 40204 12818 0 INST_config_UART._0379_
rlabel metal1 41814 13974 41814 13974 0 INST_config_UART._0380_
rlabel metal1 39008 12818 39008 12818 0 INST_config_UART._0381_
rlabel metal1 35880 14042 35880 14042 0 INST_config_UART._0382_
rlabel metal1 35512 12818 35512 12818 0 INST_config_UART._0383_
rlabel metal1 24060 12818 24060 12818 0 INST_config_UART._0384_
rlabel metal1 23598 12852 23598 12852 0 INST_config_UART._0385_
rlabel metal1 23828 12954 23828 12954 0 INST_config_UART._0386_
rlabel via1 23782 12835 23782 12835 0 INST_config_UART._0387_
rlabel metal1 22586 15096 22586 15096 0 INST_config_UART._0388_
rlabel metal2 23414 15334 23414 15334 0 INST_config_UART._0389_
rlabel metal1 22770 17714 22770 17714 0 INST_config_UART._0390_
rlabel metal1 21068 14858 21068 14858 0 INST_config_UART._0391_
rlabel metal1 22816 14382 22816 14382 0 INST_config_UART._0392_
rlabel metal1 21574 16592 21574 16592 0 INST_config_UART._0393_
rlabel metal1 22816 17850 22816 17850 0 INST_config_UART._0394_
rlabel metal1 25116 16626 25116 16626 0 INST_config_UART._0395_
rlabel metal1 23736 18394 23736 18394 0 INST_config_UART._0396_
rlabel metal1 24518 15028 24518 15028 0 INST_config_UART._0397_
rlabel metal1 17618 11322 17618 11322 0 INST_config_UART._0398_
rlabel metal1 15502 10710 15502 10710 0 INST_config_UART._0399_
rlabel metal2 10166 9860 10166 9860 0 INST_config_UART._0400_
rlabel metal1 11178 8602 11178 8602 0 INST_config_UART._0401_
rlabel metal2 12374 10676 12374 10676 0 INST_config_UART._0402_
rlabel metal1 13156 7922 13156 7922 0 INST_config_UART._0403_
rlabel metal1 14490 8874 14490 8874 0 INST_config_UART._0404_
rlabel metal1 14306 9962 14306 9962 0 INST_config_UART._0405_
rlabel metal1 14352 10982 14352 10982 0 INST_config_UART._0406_
rlabel metal1 15502 10642 15502 10642 0 INST_config_UART._0407_
rlabel metal1 16928 11798 16928 11798 0 INST_config_UART._0408_
rlabel metal1 15916 11866 15916 11866 0 INST_config_UART._0409_
rlabel metal1 25576 12614 25576 12614 0 INST_config_UART._0410_
rlabel via2 24610 14603 24610 14603 0 INST_config_UART._0411_
rlabel metal1 24794 16762 24794 16762 0 INST_config_UART._0412_
rlabel metal1 26772 14994 26772 14994 0 INST_config_UART._0413_
rlabel metal1 25024 17306 25024 17306 0 INST_config_UART._0414_
rlabel metal1 25806 19380 25806 19380 0 INST_config_UART._0415_
rlabel metal1 25714 18292 25714 18292 0 INST_config_UART._0416_
rlabel metal1 25070 15028 25070 15028 0 INST_config_UART._0417_
rlabel metal1 14398 10234 14398 10234 0 INST_config_UART._0418_
rlabel metal1 8740 10438 8740 10438 0 INST_config_UART._0419_
rlabel metal2 9338 9928 9338 9928 0 INST_config_UART._0420_
rlabel metal1 8602 10608 8602 10608 0 INST_config_UART._0421_
rlabel metal2 10534 9350 10534 9350 0 INST_config_UART._0422_
rlabel metal1 9338 8942 9338 8942 0 INST_config_UART._0423_
rlabel metal1 10396 10234 10396 10234 0 INST_config_UART._0424_
rlabel metal1 10672 9622 10672 9622 0 INST_config_UART._0425_
rlabel metal1 9246 7718 9246 7718 0 INST_config_UART._0426_
rlabel metal1 9062 7888 9062 7888 0 INST_config_UART._0427_
rlabel metal2 10166 8432 10166 8432 0 INST_config_UART._0428_
rlabel metal1 10304 6630 10304 6630 0 INST_config_UART._0429_
rlabel metal1 11178 8500 11178 8500 0 INST_config_UART._0430_
rlabel metal1 11086 10778 11086 10778 0 INST_config_UART._0431_
rlabel metal1 11592 11254 11592 11254 0 INST_config_UART._0432_
rlabel metal1 12236 11186 12236 11186 0 INST_config_UART._0433_
rlabel metal1 11730 9622 11730 9622 0 INST_config_UART._0434_
rlabel metal1 12282 8500 12282 8500 0 INST_config_UART._0435_
rlabel metal1 12880 8466 12880 8466 0 INST_config_UART._0436_
rlabel metal1 12880 8058 12880 8058 0 INST_config_UART._0437_
rlabel metal1 13294 8058 13294 8058 0 INST_config_UART._0438_
rlabel metal1 13156 9690 13156 9690 0 INST_config_UART._0439_
rlabel metal1 14214 9894 14214 9894 0 INST_config_UART._0440_
rlabel metal1 13754 10064 13754 10064 0 INST_config_UART._0441_
rlabel metal1 15364 18734 15364 18734 0 INST_config_UART._0442_
rlabel metal1 17618 18122 17618 18122 0 INST_config_UART._0443_
rlabel metal1 21252 19482 21252 19482 0 INST_config_UART._0444_
rlabel metal1 17618 17612 17618 17612 0 INST_config_UART._0445_
rlabel metal1 18262 17782 18262 17782 0 INST_config_UART._0446_
rlabel metal1 17250 19822 17250 19822 0 INST_config_UART._0447_
rlabel metal1 16974 16218 16974 16218 0 INST_config_UART._0448_
rlabel metal1 17066 13906 17066 13906 0 INST_config_UART._0449_
rlabel metal1 16790 13498 16790 13498 0 INST_config_UART._0450_
rlabel metal2 16606 13129 16606 13129 0 INST_config_UART._0451_
rlabel metal1 32890 5746 32890 5746 0 INST_config_UART._0452_
rlabel metal2 34546 6579 34546 6579 0 INST_config_UART._0453_
rlabel metal1 33856 5678 33856 5678 0 INST_config_UART._0454_
rlabel metal2 31786 9180 31786 9180 0 INST_config_UART._0455_
rlabel metal2 34454 7344 34454 7344 0 INST_config_UART._0456_
rlabel metal1 28520 7922 28520 7922 0 INST_config_UART._0457_
rlabel metal3 32614 10268 32614 10268 0 INST_config_UART._0458_
rlabel metal1 32982 9044 32982 9044 0 INST_config_UART._0459_
rlabel metal1 19458 15368 19458 15368 0 INST_config_UART._0460_
rlabel metal1 19642 15674 19642 15674 0 INST_config_UART._0461_
rlabel metal1 19090 17272 19090 17272 0 INST_config_UART._0462_
rlabel metal1 20838 15504 20838 15504 0 INST_config_UART._0463_
rlabel metal1 20010 15912 20010 15912 0 INST_config_UART._0464_
rlabel metal1 16652 17306 16652 17306 0 INST_config_UART._0465_
rlabel metal1 18676 21930 18676 21930 0 INST_config_UART._0466_
rlabel metal1 17388 15062 17388 15062 0 INST_config_UART._0467_
rlabel via1 15597 17170 15597 17170 0 INST_config_UART._0468_
rlabel metal1 16514 17272 16514 17272 0 INST_config_UART._0469_
rlabel metal1 21574 15674 21574 15674 0 INST_config_UART._0470_
rlabel metal1 21114 17510 21114 17510 0 INST_config_UART._0471_
rlabel metal1 20654 15674 20654 15674 0 INST_config_UART._0472_
rlabel metal1 20332 16490 20332 16490 0 INST_config_UART._0473_
rlabel metal2 20654 17442 20654 17442 0 INST_config_UART._0474_
rlabel metal1 20194 16218 20194 16218 0 INST_config_UART._0475_
rlabel metal2 21206 17986 21206 17986 0 INST_config_UART._0476_
rlabel metal1 20286 17782 20286 17782 0 INST_config_UART._0477_
rlabel metal2 20516 18258 20516 18258 0 INST_config_UART._0478_
rlabel metal1 20240 17850 20240 17850 0 INST_config_UART._0479_
rlabel metal1 21482 18224 21482 18224 0 INST_config_UART._0480_
rlabel metal2 20654 18768 20654 18768 0 INST_config_UART._0481_
rlabel viali 20389 19346 20389 19346 0 INST_config_UART._0482_
rlabel metal1 19550 18836 19550 18836 0 INST_config_UART._0483_
rlabel metal1 19274 18700 19274 18700 0 INST_config_UART._0484_
rlabel metal1 19320 18802 19320 18802 0 INST_config_UART._0485_
rlabel metal1 19964 18734 19964 18734 0 INST_config_UART._0486_
rlabel metal1 20884 20434 20884 20434 0 INST_config_UART._0487_
rlabel metal1 23644 18938 23644 18938 0 INST_config_UART._0488_
rlabel metal1 22954 20570 22954 20570 0 INST_config_UART._0489_
rlabel metal2 20838 21012 20838 21012 0 INST_config_UART._0490_
rlabel metal1 21206 20536 21206 20536 0 INST_config_UART._0491_
rlabel metal1 20102 20570 20102 20570 0 INST_config_UART._0492_
rlabel metal1 21482 21556 21482 21556 0 INST_config_UART._0493_
rlabel metal1 21850 19890 21850 19890 0 INST_config_UART._0494_
rlabel metal1 21252 21522 21252 21522 0 INST_config_UART._0495_
rlabel metal2 20562 21726 20562 21726 0 INST_config_UART._0496_
rlabel metal1 19826 20910 19826 20910 0 INST_config_UART._0497_
rlabel metal1 20562 20570 20562 20570 0 INST_config_UART._0498_
rlabel metal1 19596 19754 19596 19754 0 INST_config_UART._0499_
rlabel metal1 19412 19346 19412 19346 0 INST_config_UART._0500_
rlabel metal1 18831 20434 18831 20434 0 INST_config_UART._0501_
rlabel metal1 19182 20366 19182 20366 0 INST_config_UART._0502_
rlabel metal1 21620 19822 21620 19822 0 INST_config_UART._0503_
rlabel metal1 19274 19142 19274 19142 0 INST_config_UART._0504_
rlabel metal2 20286 20298 20286 20298 0 INST_config_UART._0505_
rlabel metal2 18170 20502 18170 20502 0 INST_config_UART._0506_
rlabel metal1 19320 20366 19320 20366 0 INST_config_UART._0507_
rlabel metal1 18630 22032 18630 22032 0 INST_config_UART._0508_
rlabel metal1 18262 20570 18262 20570 0 INST_config_UART._0509_
rlabel metal1 18630 18768 18630 18768 0 INST_config_UART._0510_
rlabel metal1 18584 20026 18584 20026 0 INST_config_UART._0511_
rlabel metal1 18630 19856 18630 19856 0 INST_config_UART._0512_
rlabel metal1 18630 19380 18630 19380 0 INST_config_UART._0513_
rlabel metal1 17572 20298 17572 20298 0 INST_config_UART._0514_
rlabel metal1 18906 20944 18906 20944 0 INST_config_UART._0515_
rlabel metal2 19964 20230 19964 20230 0 INST_config_UART._0516_
rlabel metal1 18308 19346 18308 19346 0 INST_config_UART._0517_
rlabel metal1 18630 19482 18630 19482 0 INST_config_UART._0518_
rlabel metal1 17986 19380 17986 19380 0 INST_config_UART._0519_
rlabel metal2 17986 20264 17986 20264 0 INST_config_UART._0520_
rlabel metal1 16100 21590 16100 21590 0 INST_config_UART._0521_
rlabel metal1 16238 21454 16238 21454 0 INST_config_UART._0522_
rlabel metal2 15226 20689 15226 20689 0 INST_config_UART._0523_
rlabel metal1 15134 20502 15134 20502 0 INST_config_UART._0524_
rlabel metal1 16813 20298 16813 20298 0 INST_config_UART._0525_
rlabel metal1 15962 20230 15962 20230 0 INST_config_UART._0526_
rlabel metal1 17250 20468 17250 20468 0 INST_config_UART._0527_
rlabel metal2 16974 19074 16974 19074 0 INST_config_UART._0528_
rlabel metal1 15410 19142 15410 19142 0 INST_config_UART._0529_
rlabel metal1 17940 17850 17940 17850 0 INST_config_UART._0530_
rlabel metal2 16514 19584 16514 19584 0 INST_config_UART._0531_
rlabel metal1 15456 19210 15456 19210 0 INST_config_UART._0532_
rlabel metal1 13892 18938 13892 18938 0 INST_config_UART._0533_
rlabel metal2 14858 19652 14858 19652 0 INST_config_UART._0534_
rlabel metal1 16422 18224 16422 18224 0 INST_config_UART._0535_
rlabel metal1 16100 18326 16100 18326 0 INST_config_UART._0536_
rlabel metal1 16237 17578 16237 17578 0 INST_config_UART._0537_
rlabel metal1 14398 17850 14398 17850 0 INST_config_UART._0538_
rlabel metal2 16422 17697 16422 17697 0 INST_config_UART._0539_
rlabel metal1 17388 14858 17388 14858 0 INST_config_UART._0540_
rlabel metal1 17572 15470 17572 15470 0 INST_config_UART._0541_
rlabel metal1 16422 15130 16422 15130 0 INST_config_UART._0542_
rlabel metal1 14996 15130 14996 15130 0 INST_config_UART._0543_
rlabel metal2 16790 17442 16790 17442 0 INST_config_UART._0544_
rlabel metal1 16560 17510 16560 17510 0 INST_config_UART._0545_
rlabel metal1 17066 16150 17066 16150 0 INST_config_UART._0546_
rlabel metal2 15502 16524 15502 16524 0 INST_config_UART._0547_
rlabel metal1 15870 16082 15870 16082 0 INST_config_UART._0548_
rlabel metal1 23322 8942 23322 8942 0 INST_config_UART._0549_
rlabel metal1 23598 9146 23598 9146 0 INST_config_UART._0550_
rlabel metal1 24334 8840 24334 8840 0 INST_config_UART._0551_
rlabel metal2 21574 13889 21574 13889 0 INST_config_UART._0552_
rlabel metal1 35696 16014 35696 16014 0 INST_config_UART._0553_
rlabel metal1 36800 16762 36800 16762 0 INST_config_UART._0554_
rlabel metal1 36570 14994 36570 14994 0 INST_config_UART._0555_
rlabel metal1 37950 16524 37950 16524 0 INST_config_UART._0556_
rlabel metal2 38318 16116 38318 16116 0 INST_config_UART._0557_
rlabel metal1 41354 16014 41354 16014 0 INST_config_UART._0558_
rlabel metal1 39054 17646 39054 17646 0 INST_config_UART._0559_
rlabel metal2 35926 17170 35926 17170 0 INST_config_UART._0560_
rlabel metal1 36386 16014 36386 16014 0 INST_config_UART._0561_
rlabel metal1 21390 14008 21390 14008 0 INST_config_UART._0562_
rlabel metal1 32154 13804 32154 13804 0 INST_config_UART._0563_
rlabel metal1 32430 13192 32430 13192 0 INST_config_UART._0564_
rlabel metal1 30682 13294 30682 13294 0 INST_config_UART._0565_
rlabel metal1 34178 11118 34178 11118 0 INST_config_UART._0566_
rlabel metal1 33212 11254 33212 11254 0 INST_config_UART._0567_
rlabel metal2 33902 14484 33902 14484 0 INST_config_UART._0568_
rlabel metal1 34270 14042 34270 14042 0 INST_config_UART._0569_
rlabel metal1 33856 13294 33856 13294 0 INST_config_UART._0570_
rlabel metal1 23138 15028 23138 15028 0 INST_config_UART._0571_
rlabel metal2 27094 13702 27094 13702 0 INST_config_UART._0572_
rlabel metal1 27830 14484 27830 14484 0 INST_config_UART._0573_
rlabel metal1 27738 12954 27738 12954 0 INST_config_UART._0574_
rlabel metal1 27186 14586 27186 14586 0 INST_config_UART._0575_
rlabel metal1 27462 15674 27462 15674 0 INST_config_UART._0576_
rlabel metal1 29808 13294 29808 13294 0 INST_config_UART._0577_
rlabel metal1 28750 16626 28750 16626 0 INST_config_UART._0578_
rlabel metal1 26956 18258 26956 18258 0 INST_config_UART._0579_
rlabel metal1 26634 18292 26634 18292 0 INST_config_UART._0580_
rlabel metal1 28566 14042 28566 14042 0 INST_config_UART._0581_
rlabel metal1 22126 7514 22126 7514 0 INST_config_UART._0582_
rlabel metal2 18446 8330 18446 8330 0 INST_config_UART._0583_
rlabel metal1 20838 6800 20838 6800 0 INST_config_UART._0584_
rlabel metal2 22862 7412 22862 7412 0 INST_config_UART._0585_
rlabel metal1 17894 9996 17894 9996 0 INST_config_UART._0586_
rlabel metal2 19366 10302 19366 10302 0 INST_config_UART._0587_
rlabel metal1 21758 6358 21758 6358 0 INST_config_UART._0588_
rlabel metal2 5198 10217 5198 10217 0 INST_config_UART.blink\[0\]
rlabel metal2 6578 16218 6578 16218 0 INST_config_UART.blink\[10\]
rlabel metal1 5612 17306 5612 17306 0 INST_config_UART.blink\[11\]
rlabel metal1 5520 18394 5520 18394 0 INST_config_UART.blink\[12\]
rlabel metal1 6072 17510 6072 17510 0 INST_config_UART.blink\[13\]
rlabel metal1 8142 17680 8142 17680 0 INST_config_UART.blink\[14\]
rlabel metal1 8188 18394 8188 18394 0 INST_config_UART.blink\[15\]
rlabel metal1 8694 17714 8694 17714 0 INST_config_UART.blink\[16\]
rlabel metal2 9154 18224 9154 18224 0 INST_config_UART.blink\[17\]
rlabel metal2 9614 18666 9614 18666 0 INST_config_UART.blink\[18\]
rlabel metal1 10764 19346 10764 19346 0 INST_config_UART.blink\[19\]
rlabel metal1 5658 9350 5658 9350 0 INST_config_UART.blink\[1\]
rlabel metal1 11960 19822 11960 19822 0 INST_config_UART.blink\[20\]
rlabel metal2 12098 18326 12098 18326 0 INST_config_UART.blink\[21\]
rlabel metal1 14720 17306 14720 17306 0 INST_config_UART.blink\[22\]
rlabel metal1 6026 9486 6026 9486 0 INST_config_UART.blink\[2\]
rlabel metal1 6026 9894 6026 9894 0 INST_config_UART.blink\[3\]
rlabel metal2 5566 11814 5566 11814 0 INST_config_UART.blink\[4\]
rlabel metal2 5658 13396 5658 13396 0 INST_config_UART.blink\[5\]
rlabel metal1 7222 12954 7222 12954 0 INST_config_UART.blink\[6\]
rlabel viali 5290 14996 5290 14996 0 INST_config_UART.blink\[7\]
rlabel metal1 5290 14824 5290 14824 0 INST_config_UART.blink\[8\]
rlabel metal2 5842 15844 5842 15844 0 INST_config_UART.blink\[9\]
rlabel metal1 14398 11832 14398 11832 0 Inst_bitbang._000_
rlabel metal1 16008 10098 16008 10098 0 Inst_bitbang._001_
rlabel metal2 14214 15844 14214 15844 0 Inst_bitbang._002_
rlabel metal1 23460 21862 23460 21862 0 Inst_bitbang._003_
rlabel metal1 26496 22406 26496 22406 0 Inst_bitbang._004_
rlabel metal2 33166 22304 33166 22304 0 Inst_bitbang._005_
rlabel metal2 32890 21250 32890 21250 0 Inst_bitbang._006_
rlabel metal1 33718 21896 33718 21896 0 Inst_bitbang._007_
rlabel metal1 35052 17850 35052 17850 0 Inst_bitbang._008_
rlabel metal1 36478 21590 36478 21590 0 Inst_bitbang._009_
rlabel metal2 36110 20978 36110 20978 0 Inst_bitbang._010_
rlabel metal1 37858 20536 37858 20536 0 Inst_bitbang._011_
rlabel metal1 37582 19448 37582 19448 0 Inst_bitbang._012_
rlabel metal1 39192 20842 39192 20842 0 Inst_bitbang._013_
rlabel metal1 40112 22066 40112 22066 0 Inst_bitbang._014_
rlabel metal1 42596 19890 42596 19890 0 Inst_bitbang._015_
rlabel metal1 42090 18360 42090 18360 0 Inst_bitbang._016_
rlabel metal1 41768 16150 41768 16150 0 Inst_bitbang._017_
rlabel metal1 42090 15096 42090 15096 0 Inst_bitbang._018_
rlabel metal1 37352 9622 37352 9622 0 Inst_bitbang._019_
rlabel metal2 37030 9452 37030 9452 0 Inst_bitbang._020_
rlabel metal2 34914 8585 34914 8585 0 Inst_bitbang._021_
rlabel metal1 34776 5882 34776 5882 0 Inst_bitbang._022_
rlabel metal1 35834 5134 35834 5134 0 Inst_bitbang._023_
rlabel metal1 34592 3706 34592 3706 0 Inst_bitbang._024_
rlabel metal2 34132 2006 34132 2006 0 Inst_bitbang._025_
rlabel metal1 39514 1530 39514 1530 0 Inst_bitbang._026_
rlabel metal1 39652 1462 39652 1462 0 Inst_bitbang._027_
rlabel metal1 40066 1870 40066 1870 0 Inst_bitbang._028_
rlabel metal1 39514 3400 39514 3400 0 Inst_bitbang._029_
rlabel metal1 39192 4794 39192 4794 0 Inst_bitbang._030_
rlabel metal1 37352 6358 37352 6358 0 Inst_bitbang._031_
rlabel via1 41347 6970 41347 6970 0 Inst_bitbang._032_
rlabel metal1 41170 5746 41170 5746 0 Inst_bitbang._033_
rlabel metal1 42090 8568 42090 8568 0 Inst_bitbang._034_
rlabel metal2 22034 21284 22034 21284 0 Inst_bitbang._035_
rlabel via1 23867 21318 23867 21318 0 Inst_bitbang._036_
rlabel metal2 25622 21250 25622 21250 0 Inst_bitbang._037_
rlabel metal1 32430 21114 32430 21114 0 Inst_bitbang._038_
rlabel metal2 33442 20706 33442 20706 0 Inst_bitbang._039_
rlabel metal2 34730 19244 34730 19244 0 Inst_bitbang._040_
rlabel metal1 36386 18802 36386 18802 0 Inst_bitbang._041_
rlabel metal1 36386 21658 36386 21658 0 Inst_bitbang._042_
rlabel metal1 38088 21658 38088 21658 0 Inst_bitbang._043_
rlabel metal1 37168 18326 37168 18326 0 Inst_bitbang._044_
rlabel metal1 38962 17850 38962 17850 0 Inst_bitbang._045_
rlabel metal1 40296 19278 40296 19278 0 Inst_bitbang._046_
rlabel metal1 41124 19482 41124 19482 0 Inst_bitbang._047_
rlabel metal1 40802 17578 40802 17578 0 Inst_bitbang._048_
rlabel metal1 40986 16626 40986 16626 0 Inst_bitbang._049_
rlabel metal1 40158 15096 40158 15096 0 Inst_bitbang._050_
rlabel metal1 41814 10166 41814 10166 0 Inst_bitbang._051_
rlabel metal1 38817 8262 38817 8262 0 Inst_bitbang._052_
rlabel metal1 37023 8262 37023 8262 0 Inst_bitbang._053_
rlabel metal1 36110 7922 36110 7922 0 Inst_bitbang._054_
rlabel metal1 35880 5746 35880 5746 0 Inst_bitbang._055_
rlabel metal1 34408 4658 34408 4658 0 Inst_bitbang._056_
rlabel metal2 34362 2621 34362 2621 0 Inst_bitbang._057_
rlabel metal1 36018 2482 36018 2482 0 Inst_bitbang._058_
rlabel metal1 36846 2958 36846 2958 0 Inst_bitbang._059_
rlabel metal1 38916 2618 38916 2618 0 Inst_bitbang._060_
rlabel metal1 38456 3706 38456 3706 0 Inst_bitbang._061_
rlabel metal1 38134 4794 38134 4794 0 Inst_bitbang._062_
rlabel metal1 38410 6120 38410 6120 0 Inst_bitbang._063_
rlabel metal1 39691 6970 39691 6970 0 Inst_bitbang._064_
rlabel metal1 39974 7752 39974 7752 0 Inst_bitbang._065_
rlabel metal1 40158 8840 40158 8840 0 Inst_bitbang._066_
rlabel metal1 10534 17238 10534 17238 0 Inst_bitbang._067_
rlabel metal1 10856 15402 10856 15402 0 Inst_bitbang._068_
rlabel metal1 10764 15334 10764 15334 0 Inst_bitbang._069_
rlabel metal1 10028 16626 10028 16626 0 Inst_bitbang._070_
rlabel metal1 8418 16150 8418 16150 0 Inst_bitbang._071_
rlabel metal1 8188 15062 8188 15062 0 Inst_bitbang._072_
rlabel metal1 7866 15402 7866 15402 0 Inst_bitbang._073_
rlabel metal1 8142 14314 8142 14314 0 Inst_bitbang._074_
rlabel metal1 8464 13974 8464 13974 0 Inst_bitbang._075_
rlabel metal1 8786 12886 8786 12886 0 Inst_bitbang._076_
rlabel metal2 9982 12308 9982 12308 0 Inst_bitbang._077_
rlabel metal1 10212 13362 10212 13362 0 Inst_bitbang._078_
rlabel metal1 11684 12410 11684 12410 0 Inst_bitbang._079_
rlabel metal2 12466 13056 12466 13056 0 Inst_bitbang._080_
rlabel metal1 13616 13362 13616 13362 0 Inst_bitbang._081_
rlabel metal1 13701 13702 13701 13702 0 Inst_bitbang._082_
rlabel metal1 14030 14994 14030 14994 0 Inst_bitbang._083_
rlabel metal2 13202 13940 13202 13940 0 Inst_bitbang._084_
rlabel metal2 13110 15164 13110 15164 0 Inst_bitbang._085_
rlabel metal1 12190 14994 12190 14994 0 Inst_bitbang._086_
rlabel metal1 38042 7344 38042 7344 0 Inst_bitbang._087_
rlabel metal1 43746 20842 43746 20842 0 Inst_bitbang._088_
rlabel metal1 16790 10608 16790 10608 0 Inst_bitbang._089_
rlabel viali 13201 15538 13201 15538 0 Inst_bitbang._090_
rlabel metal1 12880 15538 12880 15538 0 Inst_bitbang._091_
rlabel metal1 14122 15402 14122 15402 0 Inst_bitbang._092_
rlabel metal1 24518 21658 24518 21658 0 Inst_bitbang._093_
rlabel metal2 26542 21862 26542 21862 0 Inst_bitbang._094_
rlabel metal1 33350 22678 33350 22678 0 Inst_bitbang._095_
rlabel metal1 33120 20910 33120 20910 0 Inst_bitbang._096_
rlabel metal1 34546 21658 34546 21658 0 Inst_bitbang._097_
rlabel metal1 35328 17646 35328 17646 0 Inst_bitbang._098_
rlabel metal1 35834 20570 35834 20570 0 Inst_bitbang._099_
rlabel metal1 37536 21114 37536 21114 0 Inst_bitbang._100_
rlabel metal2 41630 19958 41630 19958 0 Inst_bitbang._101_
rlabel metal2 38134 21495 38134 21495 0 Inst_bitbang._102_
rlabel metal1 38318 18938 38318 18938 0 Inst_bitbang._103_
rlabel metal1 39054 20944 39054 20944 0 Inst_bitbang._104_
rlabel metal1 41768 20230 41768 20230 0 Inst_bitbang._105_
rlabel metal2 41814 19924 41814 19924 0 Inst_bitbang._106_
rlabel metal1 42412 18734 42412 18734 0 Inst_bitbang._107_
rlabel metal2 41814 16763 41814 16763 0 Inst_bitbang._108_
rlabel metal1 42274 14586 42274 14586 0 Inst_bitbang._109_
rlabel metal1 38824 9690 38824 9690 0 Inst_bitbang._110_
rlabel metal1 37214 10064 37214 10064 0 Inst_bitbang._111_
rlabel metal1 39790 4692 39790 4692 0 Inst_bitbang._112_
rlabel metal1 35052 7514 35052 7514 0 Inst_bitbang._113_
rlabel metal1 35098 5780 35098 5780 0 Inst_bitbang._114_
rlabel metal1 36984 5202 36984 5202 0 Inst_bitbang._115_
rlabel metal1 35006 3502 35006 3502 0 Inst_bitbang._116_
rlabel metal1 34776 1190 34776 1190 0 Inst_bitbang._117_
rlabel metal1 37858 1224 37858 1224 0 Inst_bitbang._118_
rlabel metal1 40434 1326 40434 1326 0 Inst_bitbang._119_
rlabel metal1 39836 1190 39836 1190 0 Inst_bitbang._120_
rlabel metal1 39054 3536 39054 3536 0 Inst_bitbang._121_
rlabel metal1 39146 4590 39146 4590 0 Inst_bitbang._122_
rlabel metal1 37812 6766 37812 6766 0 Inst_bitbang._123_
rlabel metal1 41676 6426 41676 6426 0 Inst_bitbang._124_
rlabel metal1 41354 7378 41354 7378 0 Inst_bitbang._125_
rlabel metal1 41492 8058 41492 8058 0 Inst_bitbang._126_
rlabel metal2 44942 20672 44942 20672 0 Inst_bitbang._127_
rlabel metal1 26542 20978 26542 20978 0 Inst_bitbang._128_
rlabel metal1 23460 20570 23460 20570 0 Inst_bitbang._129_
rlabel metal1 24104 21862 24104 21862 0 Inst_bitbang._130_
rlabel metal1 25760 20434 25760 20434 0 Inst_bitbang._131_
rlabel metal1 32292 20910 32292 20910 0 Inst_bitbang._132_
rlabel metal1 33672 20434 33672 20434 0 Inst_bitbang._133_
rlabel metal1 34730 19482 34730 19482 0 Inst_bitbang._134_
rlabel metal1 35880 17850 35880 17850 0 Inst_bitbang._135_
rlabel metal1 36570 20570 36570 20570 0 Inst_bitbang._136_
rlabel metal1 37168 20026 37168 20026 0 Inst_bitbang._137_
rlabel metal1 37214 19426 37214 19426 0 Inst_bitbang._138_
rlabel metal1 41446 18258 41446 18258 0 Inst_bitbang._139_
rlabel metal1 38594 17680 38594 17680 0 Inst_bitbang._140_
rlabel metal1 41032 19346 41032 19346 0 Inst_bitbang._141_
rlabel metal2 41538 19142 41538 19142 0 Inst_bitbang._142_
rlabel metal1 40848 18258 40848 18258 0 Inst_bitbang._143_
rlabel metal1 40848 17170 40848 17170 0 Inst_bitbang._144_
rlabel metal1 41308 15470 41308 15470 0 Inst_bitbang._145_
rlabel metal2 41998 10948 41998 10948 0 Inst_bitbang._146_
rlabel metal1 39054 8976 39054 8976 0 Inst_bitbang._147_
rlabel metal1 37582 7514 37582 7514 0 Inst_bitbang._148_
rlabel metal1 36984 8058 36984 8058 0 Inst_bitbang._149_
rlabel metal1 35190 2958 35190 2958 0 Inst_bitbang._150_
rlabel metal1 36432 6290 36432 6290 0 Inst_bitbang._151_
rlabel metal1 35650 4794 35650 4794 0 Inst_bitbang._152_
rlabel metal1 34822 3162 34822 3162 0 Inst_bitbang._153_
rlabel metal1 36018 2958 36018 2958 0 Inst_bitbang._154_
rlabel metal1 36478 3060 36478 3060 0 Inst_bitbang._155_
rlabel metal1 39146 2414 39146 2414 0 Inst_bitbang._156_
rlabel metal1 38824 3502 38824 3502 0 Inst_bitbang._157_
rlabel metal1 38410 4624 38410 4624 0 Inst_bitbang._158_
rlabel via2 40802 6171 40802 6171 0 Inst_bitbang._159_
rlabel metal1 39882 7378 39882 7378 0 Inst_bitbang._160_
rlabel metal1 39882 7514 39882 7514 0 Inst_bitbang._161_
rlabel metal1 40112 8330 40112 8330 0 Inst_bitbang._162_
rlabel metal1 15088 13838 15088 13838 0 Inst_bitbang._163_
rlabel metal2 8050 14688 8050 14688 0 Inst_bitbang._164_
rlabel metal1 10074 17136 10074 17136 0 Inst_bitbang._165_
rlabel metal1 11546 16762 11546 16762 0 Inst_bitbang._166_
rlabel metal1 10534 15572 10534 15572 0 Inst_bitbang._167_
rlabel metal1 10166 16218 10166 16218 0 Inst_bitbang._168_
rlabel metal1 8832 16558 8832 16558 0 Inst_bitbang._169_
rlabel metal2 8510 16762 8510 16762 0 Inst_bitbang._170_
rlabel metal1 7360 15470 7360 15470 0 Inst_bitbang._171_
rlabel metal1 7866 14416 7866 14416 0 Inst_bitbang._172_
rlabel metal1 7774 14042 7774 14042 0 Inst_bitbang._173_
rlabel metal1 9108 13294 9108 13294 0 Inst_bitbang._174_
rlabel metal1 9522 13498 9522 13498 0 Inst_bitbang._175_
rlabel metal1 10718 13974 10718 13974 0 Inst_bitbang._176_
rlabel metal2 11822 12410 11822 12410 0 Inst_bitbang._177_
rlabel metal2 12558 13333 12558 13333 0 Inst_bitbang._178_
rlabel metal1 14766 13872 14766 13872 0 Inst_bitbang._179_
rlabel metal1 14720 14382 14720 14382 0 Inst_bitbang._180_
rlabel metal1 44942 17102 44942 17102 0 Inst_bitbang.active
rlabel metal1 26956 22542 26956 22542 0 Inst_bitbang.data\[0\]
rlabel metal1 41469 20978 41469 20978 0 Inst_bitbang.data\[10\]
rlabel metal1 42320 20570 42320 20570 0 Inst_bitbang.data\[11\]
rlabel metal1 43562 19482 43562 19482 0 Inst_bitbang.data\[12\]
rlabel metal1 43286 18394 43286 18394 0 Inst_bitbang.data\[13\]
rlabel metal1 42826 17170 42826 17170 0 Inst_bitbang.data\[14\]
rlabel metal2 42642 14858 42642 14858 0 Inst_bitbang.data\[15\]
rlabel metal1 38042 9486 38042 9486 0 Inst_bitbang.data\[16\]
rlabel metal1 37674 9146 37674 9146 0 Inst_bitbang.data\[17\]
rlabel metal1 36110 8602 36110 8602 0 Inst_bitbang.data\[18\]
rlabel metal1 35696 6426 35696 6426 0 Inst_bitbang.data\[19\]
rlabel metal1 27554 21318 27554 21318 0 Inst_bitbang.data\[1\]
rlabel metal1 36662 5338 36662 5338 0 Inst_bitbang.data\[20\]
rlabel metal1 35558 3604 35558 3604 0 Inst_bitbang.data\[21\]
rlabel metal1 35926 1870 35926 1870 0 Inst_bitbang.data\[22\]
rlabel metal1 38180 2482 38180 2482 0 Inst_bitbang.data\[23\]
rlabel metal1 40342 2346 40342 2346 0 Inst_bitbang.data\[24\]
rlabel metal1 40572 2074 40572 2074 0 Inst_bitbang.data\[25\]
rlabel metal1 40894 4250 40894 4250 0 Inst_bitbang.data\[26\]
rlabel metal2 40894 4828 40894 4828 0 Inst_bitbang.data\[27\]
rlabel metal2 38870 6528 38870 6528 0 Inst_bitbang.data\[28\]
rlabel metal1 43102 6834 43102 6834 0 Inst_bitbang.data\[29\]
rlabel metal1 32292 22134 32292 22134 0 Inst_bitbang.data\[2\]
rlabel metal2 43102 6902 43102 6902 0 Inst_bitbang.data\[30\]
rlabel metal2 42826 8092 42826 8092 0 Inst_bitbang.data\[31\]
rlabel metal1 34270 21318 34270 21318 0 Inst_bitbang.data\[3\]
rlabel metal1 35328 21454 35328 21454 0 Inst_bitbang.data\[4\]
rlabel metal2 35834 18836 35834 18836 0 Inst_bitbang.data\[5\]
rlabel metal1 36570 20434 36570 20434 0 Inst_bitbang.data\[6\]
rlabel metal1 38226 21012 38226 21012 0 Inst_bitbang.data\[7\]
rlabel metal1 39514 20570 39514 20570 0 Inst_bitbang.data\[8\]
rlabel metal1 38824 18734 38824 18734 0 Inst_bitbang.data\[9\]
rlabel metal1 15548 11050 15548 11050 0 Inst_bitbang.local_strobe
rlabel metal1 16468 10710 16468 10710 0 Inst_bitbang.old_local_strobe
rlabel metal1 4094 14008 4094 14008 0 Inst_bitbang.s_clk_sample\[0\]
rlabel metal1 6072 13226 6072 13226 0 Inst_bitbang.s_clk_sample\[1\]
rlabel metal1 8050 13192 8050 13192 0 Inst_bitbang.s_clk_sample\[2\]
rlabel metal1 15548 12614 15548 12614 0 Inst_bitbang.s_clk_sample\[3\]
rlabel metal1 3864 20502 3864 20502 0 Inst_bitbang.s_data_sample\[0\]
rlabel metal1 6118 20570 6118 20570 0 Inst_bitbang.s_data_sample\[1\]
rlabel metal1 8694 20978 8694 20978 0 Inst_bitbang.s_data_sample\[2\]
rlabel metal1 17250 19992 17250 19992 0 Inst_bitbang.s_data_sample\[3\]
rlabel metal1 12604 16422 12604 16422 0 Inst_bitbang.serial_control\[0\]
rlabel metal1 10994 12852 10994 12852 0 Inst_bitbang.serial_control\[10\]
rlabel metal1 11408 13498 11408 13498 0 Inst_bitbang.serial_control\[11\]
rlabel metal1 13064 13498 13064 13498 0 Inst_bitbang.serial_control\[12\]
rlabel metal1 13202 14042 13202 14042 0 Inst_bitbang.serial_control\[13\]
rlabel metal1 13892 12886 13892 12886 0 Inst_bitbang.serial_control\[14\]
rlabel metal2 13938 13600 13938 13600 0 Inst_bitbang.serial_control\[15\]
rlabel metal1 12098 15334 12098 15334 0 Inst_bitbang.serial_control\[1\]
rlabel metal2 12650 15776 12650 15776 0 Inst_bitbang.serial_control\[2\]
rlabel metal2 13294 15266 13294 15266 0 Inst_bitbang.serial_control\[3\]
rlabel metal2 9706 15232 9706 15232 0 Inst_bitbang.serial_control\[4\]
rlabel metal1 9522 14960 9522 14960 0 Inst_bitbang.serial_control\[5\]
rlabel metal1 8970 15334 8970 15334 0 Inst_bitbang.serial_control\[6\]
rlabel metal2 10074 14144 10074 14144 0 Inst_bitbang.serial_control\[7\]
rlabel metal1 9062 13838 9062 13838 0 Inst_bitbang.serial_control\[8\]
rlabel metal1 9844 12750 9844 12750 0 Inst_bitbang.serial_control\[9\]
rlabel metal1 24978 21930 24978 21930 0 Inst_bitbang.serial_data\[0\]
rlabel metal2 40986 19856 40986 19856 0 Inst_bitbang.serial_data\[10\]
rlabel metal2 41446 19584 41446 19584 0 Inst_bitbang.serial_data\[11\]
rlabel metal2 42182 19584 42182 19584 0 Inst_bitbang.serial_data\[12\]
rlabel metal1 42366 17850 42366 17850 0 Inst_bitbang.serial_data\[13\]
rlabel metal2 41584 16252 41584 16252 0 Inst_bitbang.serial_data\[14\]
rlabel metal1 41814 14246 41814 14246 0 Inst_bitbang.serial_data\[15\]
rlabel metal1 39744 9622 39744 9622 0 Inst_bitbang.serial_data\[16\]
rlabel metal1 40204 9486 40204 9486 0 Inst_bitbang.serial_data\[17\]
rlabel metal1 37904 7854 37904 7854 0 Inst_bitbang.serial_data\[18\]
rlabel metal1 37214 7718 37214 7718 0 Inst_bitbang.serial_data\[19\]
rlabel metal1 25346 21522 25346 21522 0 Inst_bitbang.serial_data\[1\]
rlabel metal1 36938 5882 36938 5882 0 Inst_bitbang.serial_data\[20\]
rlabel metal1 36524 4454 36524 4454 0 Inst_bitbang.serial_data\[21\]
rlabel metal1 35006 3094 35006 3094 0 Inst_bitbang.serial_data\[22\]
rlabel metal1 37490 2618 37490 2618 0 Inst_bitbang.serial_data\[23\]
rlabel metal1 39514 2414 39514 2414 0 Inst_bitbang.serial_data\[24\]
rlabel metal1 39698 2516 39698 2516 0 Inst_bitbang.serial_data\[25\]
rlabel metal1 39928 4250 39928 4250 0 Inst_bitbang.serial_data\[26\]
rlabel metal1 40342 5338 40342 5338 0 Inst_bitbang.serial_data\[27\]
rlabel metal1 39284 7378 39284 7378 0 Inst_bitbang.serial_data\[28\]
rlabel metal1 40020 7446 40020 7446 0 Inst_bitbang.serial_data\[29\]
rlabel metal1 32016 20842 32016 20842 0 Inst_bitbang.serial_data\[2\]
rlabel metal1 41354 7922 41354 7922 0 Inst_bitbang.serial_data\[30\]
rlabel metal1 41768 8806 41768 8806 0 Inst_bitbang.serial_data\[31\]
rlabel metal1 33810 20774 33810 20774 0 Inst_bitbang.serial_data\[3\]
rlabel metal1 35696 21114 35696 21114 0 Inst_bitbang.serial_data\[4\]
rlabel metal1 35374 19346 35374 19346 0 Inst_bitbang.serial_data\[5\]
rlabel metal1 36938 20502 36938 20502 0 Inst_bitbang.serial_data\[6\]
rlabel metal1 37950 20774 37950 20774 0 Inst_bitbang.serial_data\[7\]
rlabel metal1 39376 21318 39376 21318 0 Inst_bitbang.serial_data\[8\]
rlabel metal1 38226 18734 38226 18734 0 Inst_bitbang.serial_data\[9\]
rlabel metal1 16606 8874 16606 8874 0 Inst_bitbang.strobe
rlabel metal2 27554 823 27554 823 0 LongFrameStrobe
rlabel metal3 544 8772 544 8772 0 ReceiveLED
rlabel metal2 28619 68 28619 68 0 RowSelect[0]
rlabel metal2 29210 1180 29210 1180 0 RowSelect[1]
rlabel metal2 30038 806 30038 806 0 RowSelect[2]
rlabel metal2 30866 908 30866 908 0 RowSelect[3]
rlabel metal1 32154 1496 32154 1496 0 RowSelect[4]
rlabel metal3 45548 14756 45548 14756 0 Rx
rlabel metal2 31234 23589 31234 23589 0 SelfWriteData[0]
rlabel metal2 40434 23232 40434 23232 0 SelfWriteData[10]
rlabel metal2 41446 23800 41446 23800 0 SelfWriteData[11]
rlabel metal2 42274 23232 42274 23232 0 SelfWriteData[12]
rlabel metal2 43194 23232 43194 23232 0 SelfWriteData[13]
rlabel metal2 44114 23232 44114 23232 0 SelfWriteData[14]
rlabel metal2 45034 23232 45034 23232 0 SelfWriteData[15]
rlabel metal2 32522 415 32522 415 0 SelfWriteData[16]
rlabel metal2 33350 347 33350 347 0 SelfWriteData[17]
rlabel metal2 34178 143 34178 143 0 SelfWriteData[18]
rlabel metal2 35006 806 35006 806 0 SelfWriteData[19]
rlabel metal2 32154 23793 32154 23793 0 SelfWriteData[1]
rlabel metal1 38594 2414 38594 2414 0 SelfWriteData[20]
rlabel metal1 40756 1938 40756 1938 0 SelfWriteData[21]
rlabel metal2 37681 68 37681 68 0 SelfWriteData[22]
rlabel metal2 38318 534 38318 534 0 SelfWriteData[23]
rlabel metal2 39146 143 39146 143 0 SelfWriteData[24]
rlabel metal1 41630 1292 41630 1292 0 SelfWriteData[25]
rlabel metal2 41998 986 41998 986 0 SelfWriteData[26]
rlabel metal2 41630 670 41630 670 0 SelfWriteData[27]
rlabel metal2 42603 68 42603 68 0 SelfWriteData[28]
rlabel metal2 43431 68 43431 68 0 SelfWriteData[29]
rlabel metal1 33350 21998 33350 21998 0 SelfWriteData[2]
rlabel metal2 44351 68 44351 68 0 SelfWriteData[30]
rlabel metal2 45087 68 45087 68 0 SelfWriteData[31]
rlabel metal2 33994 23538 33994 23538 0 SelfWriteData[3]
rlabel metal2 34914 23266 34914 23266 0 SelfWriteData[4]
rlabel metal2 35834 23232 35834 23232 0 SelfWriteData[5]
rlabel metal2 36754 23538 36754 23538 0 SelfWriteData[6]
rlabel metal2 37674 23793 37674 23793 0 SelfWriteData[7]
rlabel metal2 38594 23538 38594 23538 0 SelfWriteData[8]
rlabel metal2 39514 23232 39514 23232 0 SelfWriteData[9]
rlabel metal3 452 2788 452 2788 0 SelfWriteStrobe
rlabel metal1 37950 17850 37950 17850 0 _000_
rlabel metal1 28336 19142 28336 19142 0 _001_
rlabel metal1 28336 18870 28336 18870 0 _002_
rlabel metal2 27554 22202 27554 22202 0 _003_
rlabel metal1 27186 21896 27186 21896 0 _004_
rlabel metal2 28014 21386 28014 21386 0 _005_
rlabel metal1 25162 20400 25162 20400 0 _006_
rlabel metal2 32614 21760 32614 21760 0 _007_
rlabel metal1 28474 21522 28474 21522 0 _008_
rlabel metal1 29946 21998 29946 21998 0 _009_
rlabel metal2 29394 22372 29394 22372 0 _010_
rlabel metal1 34638 20298 34638 20298 0 _011_
rlabel metal1 29256 21658 29256 21658 0 _012_
rlabel metal2 35190 19261 35190 19261 0 _013_
rlabel metal1 29210 18938 29210 18938 0 _014_
rlabel metal2 36662 21981 36662 21981 0 _015_
rlabel metal1 30222 22610 30222 22610 0 _016_
rlabel metal2 37858 21641 37858 21641 0 _017_
rlabel metal2 30774 21250 30774 21250 0 _018_
rlabel metal2 38824 20842 38824 20842 0 _019_
rlabel metal2 30958 22345 30958 22345 0 _020_
rlabel metal1 42458 20910 42458 20910 0 _021_
rlabel metal1 36570 18224 36570 18224 0 _022_
rlabel metal1 32614 14926 32614 14926 0 _023_
rlabel metal1 33856 18734 33856 18734 0 _024_
rlabel metal1 40342 21420 40342 21420 0 _025_
rlabel metal1 32384 20434 32384 20434 0 _026_
rlabel metal2 41906 20825 41906 20825 0 _027_
rlabel metal1 31464 19346 31464 19346 0 _028_
rlabel metal1 42642 19312 42642 19312 0 _029_
rlabel metal1 32522 19822 32522 19822 0 _030_
rlabel metal1 32430 17238 32430 17238 0 _031_
rlabel metal1 31740 17238 31740 17238 0 _032_
rlabel metal2 42918 16320 42918 16320 0 _033_
rlabel metal1 33120 16558 33120 16558 0 _034_
rlabel metal1 41630 14994 41630 14994 0 _035_
rlabel metal1 31809 15130 31809 15130 0 _036_
rlabel metal2 32982 9792 32982 9792 0 _037_
rlabel metal1 32430 8942 32430 8942 0 _038_
rlabel metal1 33856 8806 33856 8806 0 _039_
rlabel metal1 31648 8534 31648 8534 0 _040_
rlabel metal1 31924 8942 31924 8942 0 _041_
rlabel metal1 30912 7786 30912 7786 0 _042_
rlabel metal1 36478 1870 36478 1870 0 _043_
rlabel metal2 34730 6528 34730 6528 0 _044_
rlabel metal1 33534 6834 33534 6834 0 _045_
rlabel metal1 28566 6392 28566 6392 0 _046_
rlabel metal1 35650 4726 35650 4726 0 _047_
rlabel metal2 29118 5474 29118 5474 0 _048_
rlabel metal1 35558 3366 35558 3366 0 _049_
rlabel metal1 29394 5270 29394 5270 0 _050_
rlabel metal1 35650 2074 35650 2074 0 _051_
rlabel metal1 29992 4522 29992 4522 0 _052_
rlabel metal2 37674 3145 37674 3145 0 _053_
rlabel metal1 30774 4216 30774 4216 0 _054_
rlabel metal2 40894 2329 40894 2329 0 _055_
rlabel metal2 32430 3944 32430 3944 0 _056_
rlabel metal1 40250 2890 40250 2890 0 _057_
rlabel metal1 33810 4216 33810 4216 0 _058_
rlabel metal1 40710 3978 40710 3978 0 _059_
rlabel metal1 31970 4012 31970 4012 0 _060_
rlabel metal1 37214 6188 37214 6188 0 _061_
rlabel metal1 26864 6426 26864 6426 0 _062_
rlabel metal2 38134 6103 38134 6103 0 _063_
rlabel metal1 31832 6834 31832 6834 0 _064_
rlabel metal2 30498 8177 30498 8177 0 _065_
rlabel metal1 26358 7412 26358 7412 0 _066_
rlabel metal1 41262 6256 41262 6256 0 _067_
rlabel metal1 33166 7208 33166 7208 0 _068_
rlabel metal1 34454 7378 34454 7378 0 _069_
rlabel metal1 33902 7514 33902 7514 0 _070_
rlabel metal2 15870 8857 15870 8857 0 _071_
rlabel metal1 26450 9146 26450 9146 0 _072_
rlabel metal1 2622 3604 2622 3604 0 net1
rlabel metal1 36202 1394 36202 1394 0 net10
rlabel metal1 6164 1326 6164 1326 0 net100
rlabel metal1 6946 1326 6946 1326 0 net101
rlabel metal2 7774 1530 7774 1530 0 net102
rlabel metal1 8786 1326 8786 1326 0 net103
rlabel metal1 27922 1326 27922 1326 0 net104
rlabel metal1 13110 9044 13110 9044 0 net105
rlabel metal1 30774 1292 30774 1292 0 net106
rlabel metal1 30544 2414 30544 2414 0 net107
rlabel metal2 34362 1054 34362 1054 0 net108
rlabel metal1 31694 1938 31694 1938 0 net109
rlabel metal1 36340 1190 36340 1190 0 net11
rlabel via1 32881 1258 32881 1258 0 net110
rlabel metal1 13570 19686 13570 19686 0 net111
rlabel metal1 2622 4073 2622 4073 0 net112
rlabel metal1 17848 1870 17848 1870 0 net113
rlabel metal1 36938 1224 36938 1224 0 net12
rlabel metal1 38502 1836 38502 1836 0 net13
rlabel metal2 33488 22406 33488 22406 0 net14
rlabel metal1 38134 2550 38134 2550 0 net15
rlabel metal3 38732 3060 38732 3060 0 net16
rlabel metal1 40434 1530 40434 1530 0 net17
rlabel metal1 40802 1190 40802 1190 0 net18
rlabel metal1 41078 1530 41078 1530 0 net19
rlabel metal1 44896 11730 44896 11730 0 net2
rlabel metal1 41078 3026 41078 3026 0 net20
rlabel metal1 41492 4182 41492 4182 0 net21
rlabel metal1 41446 5202 41446 5202 0 net22
rlabel metal2 42550 1020 42550 1020 0 net23
rlabel metal1 43332 1190 43332 1190 0 net24
rlabel metal1 33442 21896 33442 21896 0 net25
rlabel metal1 44390 1258 44390 1258 0 net26
rlabel metal1 45034 1258 45034 1258 0 net27
rlabel metal1 34684 22610 34684 22610 0 net28
rlabel metal1 35052 20570 35052 20570 0 net29
rlabel metal2 27922 22882 27922 22882 0 net3
rlabel metal1 35696 19822 35696 19822 0 net30
rlabel metal1 37398 22746 37398 22746 0 net31
rlabel metal1 38594 21998 38594 21998 0 net32
rlabel metal1 39422 21998 39422 21998 0 net33
rlabel metal1 39238 18326 39238 18326 0 net34
rlabel metal1 1150 3162 1150 3162 0 net35
rlabel metal2 2254 2312 2254 2312 0 net36
rlabel metal1 1978 13838 1978 13838 0 net37
rlabel metal1 1472 20502 1472 20502 0 net38
rlabel metal1 44390 20026 44390 20026 0 net39
rlabel metal1 40618 21658 40618 21658 0 net4
rlabel metal1 1196 22202 1196 22202 0 net40
rlabel metal2 10166 22406 10166 22406 0 net41
rlabel metal1 11040 22202 11040 22202 0 net42
rlabel metal1 11914 22202 11914 22202 0 net43
rlabel metal1 12880 22202 12880 22202 0 net44
rlabel metal1 13524 22202 13524 22202 0 net45
rlabel metal1 14444 22202 14444 22202 0 net46
rlabel metal1 16054 22644 16054 22644 0 net47
rlabel metal2 16790 22406 16790 22406 0 net48
rlabel metal1 17388 22202 17388 22202 0 net49
rlabel metal1 41860 20910 41860 20910 0 net5
rlabel metal2 18262 22406 18262 22406 0 net50
rlabel metal1 1978 22202 1978 22202 0 net51
rlabel metal2 19734 22406 19734 22406 0 net52
rlabel metal1 20148 22202 20148 22202 0 net53
rlabel metal1 21390 22610 21390 22610 0 net54
rlabel metal1 22172 22202 22172 22202 0 net55
rlabel metal1 22908 22202 22908 22202 0 net56
rlabel metal2 23138 22406 23138 22406 0 net57
rlabel metal1 24886 22202 24886 22202 0 net58
rlabel metal1 25806 22644 25806 22644 0 net59
rlabel metal1 42872 19414 42872 19414 0 net6
rlabel metal1 26910 22610 26910 22610 0 net60
rlabel metal2 29026 21488 29026 21488 0 net61
rlabel metal1 3036 22202 3036 22202 0 net62
rlabel metal1 29578 22576 29578 22576 0 net63
rlabel metal1 30268 20298 30268 20298 0 net64
rlabel metal1 3956 22202 3956 22202 0 net65
rlabel metal2 4646 22406 4646 22406 0 net66
rlabel metal1 5658 22202 5658 22202 0 net67
rlabel metal2 6486 22406 6486 22406 0 net68
rlabel metal1 7360 22202 7360 22202 0 net69
rlabel metal1 43102 17646 43102 17646 0 net7
rlabel metal1 8372 22202 8372 22202 0 net70
rlabel metal1 9338 22202 9338 22202 0 net71
rlabel metal2 42826 22848 42826 22848 0 net72
rlabel metal1 1242 1326 1242 1326 0 net73
rlabel metal1 9568 1326 9568 1326 0 net74
rlabel metal1 10304 1326 10304 1326 0 net75
rlabel metal1 11086 1326 11086 1326 0 net76
rlabel metal1 11960 1326 11960 1326 0 net77
rlabel metal2 12282 1530 12282 1530 0 net78
rlabel metal1 13524 1326 13524 1326 0 net79
rlabel metal1 43838 16558 43838 16558 0 net8
rlabel metal2 14398 1530 14398 1530 0 net80
rlabel metal1 15272 1326 15272 1326 0 net81
rlabel metal1 16146 1326 16146 1326 0 net82
rlabel metal1 17618 1326 17618 1326 0 net83
rlabel metal1 2070 1326 2070 1326 0 net84
rlabel metal1 18538 1326 18538 1326 0 net85
rlabel metal1 19504 1326 19504 1326 0 net86
rlabel metal2 20194 1530 20194 1530 0 net87
rlabel metal1 21022 1326 21022 1326 0 net88
rlabel metal1 21850 1292 21850 1292 0 net89
rlabel metal1 43792 15402 43792 15402 0 net9
rlabel metal1 22678 1360 22678 1360 0 net90
rlabel metal1 23506 1258 23506 1258 0 net91
rlabel metal1 22402 1224 22402 1224 0 net92
rlabel metal1 26358 1326 26358 1326 0 net93
rlabel metal1 3128 1326 3128 1326 0 net94
rlabel metal1 27094 1326 27094 1326 0 net95
rlabel metal1 28198 1292 28198 1292 0 net96
rlabel metal1 3864 1326 3864 1326 0 net97
rlabel metal1 4508 1326 4508 1326 0 net98
rlabel metal1 5244 1326 5244 1326 0 net99
rlabel metal3 45272 8772 45272 8772 0 resetn
rlabel metal3 544 14756 544 14756 0 s_clk
rlabel metal3 544 20740 544 20740 0 s_data
<< properties >>
string FIXED_BBOX 0 0 46000 24000
<< end >>
