magic
tech sky130A
magscale 1 2
timestamp 1733618896
<< viali >>
rect 4997 7497 5031 7531
rect 5549 7497 5583 7531
rect 6377 7497 6411 7531
rect 7021 7497 7055 7531
rect 7573 7497 7607 7531
rect 8125 7497 8159 7531
rect 8677 7497 8711 7531
rect 10057 7497 10091 7531
rect 10609 7497 10643 7531
rect 12081 7497 12115 7531
rect 12633 7497 12667 7531
rect 13277 7497 13311 7531
rect 13829 7497 13863 7531
rect 14749 7497 14783 7531
rect 15301 7497 15335 7531
rect 15853 7497 15887 7531
rect 16681 7497 16715 7531
rect 17141 7497 17175 7531
rect 17693 7497 17727 7531
rect 18245 7497 18279 7531
rect 18797 7497 18831 7531
rect 19441 7497 19475 7531
rect 19993 7497 20027 7531
rect 21465 7497 21499 7531
rect 22017 7497 22051 7531
rect 23029 7497 23063 7531
rect 23949 7497 23983 7531
rect 25697 7497 25731 7531
rect 26065 7497 26099 7531
rect 31401 7497 31435 7531
rect 33701 7497 33735 7531
rect 34069 7497 34103 7531
rect 34897 7497 34931 7531
rect 35449 7497 35483 7531
rect 36553 7497 36587 7531
rect 36921 7497 36955 7531
rect 40601 7497 40635 7531
rect 5273 7429 5307 7463
rect 10701 7429 10735 7463
rect 13001 7429 13035 7463
rect 13553 7429 13587 7463
rect 16129 7429 16163 7463
rect 38301 7429 38335 7463
rect 38485 7429 38519 7463
rect 40325 7429 40359 7463
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 7297 7361 7331 7395
rect 7849 7361 7883 7395
rect 8401 7361 8435 7395
rect 9137 7361 9171 7395
rect 9689 7361 9723 7395
rect 11253 7361 11287 7395
rect 11713 7361 11747 7395
rect 12173 7361 12207 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 15025 7361 15059 7395
rect 15577 7361 15611 7395
rect 16497 7361 16531 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 17601 7361 17635 7395
rect 18153 7361 18187 7395
rect 18705 7361 18739 7395
rect 19349 7361 19383 7395
rect 19901 7361 19935 7395
rect 20361 7361 20395 7395
rect 20637 7361 20671 7395
rect 21097 7361 21131 7395
rect 21189 7361 21223 7395
rect 21649 7361 21683 7395
rect 22201 7361 22235 7395
rect 22477 7361 22511 7395
rect 22753 7361 22787 7395
rect 22845 7361 22879 7395
rect 23305 7361 23339 7395
rect 23581 7361 23615 7395
rect 23857 7361 23891 7395
rect 24133 7361 24167 7395
rect 24593 7361 24627 7395
rect 24869 7361 24903 7395
rect 24961 7361 24995 7395
rect 25421 7361 25455 7395
rect 25513 7361 25547 7395
rect 25973 7361 26007 7395
rect 26249 7361 26283 7395
rect 26525 7361 26559 7395
rect 26801 7361 26835 7395
rect 27169 7361 27203 7395
rect 27445 7361 27479 7395
rect 27721 7361 27755 7395
rect 27997 7361 28031 7395
rect 28273 7361 28307 7395
rect 28549 7361 28583 7395
rect 28825 7361 28859 7395
rect 29101 7361 29135 7395
rect 29377 7361 29411 7395
rect 29745 7361 29779 7395
rect 30021 7361 30055 7395
rect 30113 7361 30147 7395
rect 30389 7361 30423 7395
rect 30665 7361 30699 7395
rect 30941 7361 30975 7395
rect 31217 7361 31251 7395
rect 31493 7361 31527 7395
rect 31769 7361 31803 7395
rect 32137 7361 32171 7395
rect 32413 7361 32447 7395
rect 32689 7361 32723 7395
rect 32965 7361 32999 7395
rect 33241 7361 33275 7395
rect 33517 7361 33551 7395
rect 33977 7361 34011 7395
rect 34805 7361 34839 7395
rect 35357 7361 35391 7395
rect 35909 7361 35943 7395
rect 36461 7361 36495 7395
rect 37105 7361 37139 7395
rect 37381 7361 37415 7395
rect 37933 7361 37967 7395
rect 39037 7361 39071 7395
rect 39957 7361 39991 7395
rect 40509 7361 40543 7395
rect 6101 7293 6135 7327
rect 10977 7293 11011 7327
rect 8953 7225 8987 7259
rect 14105 7225 14139 7259
rect 22293 7225 22327 7259
rect 22569 7225 22603 7259
rect 25789 7225 25823 7259
rect 26985 7225 27019 7259
rect 31677 7225 31711 7259
rect 32597 7225 32631 7259
rect 33149 7225 33183 7259
rect 38669 7225 38703 7259
rect 4353 7157 4387 7191
rect 11529 7157 11563 7191
rect 20545 7157 20579 7191
rect 20821 7157 20855 7191
rect 20913 7157 20947 7191
rect 21373 7157 21407 7191
rect 23121 7157 23155 7191
rect 23397 7157 23431 7191
rect 23673 7157 23707 7191
rect 24409 7157 24443 7191
rect 24685 7157 24719 7191
rect 25145 7157 25179 7191
rect 25237 7157 25271 7191
rect 26341 7157 26375 7191
rect 26617 7157 26651 7191
rect 27261 7157 27295 7191
rect 27537 7157 27571 7191
rect 27813 7157 27847 7191
rect 28089 7157 28123 7191
rect 28365 7157 28399 7191
rect 28641 7157 28675 7191
rect 28917 7157 28951 7191
rect 29193 7157 29227 7191
rect 29561 7157 29595 7191
rect 29837 7157 29871 7191
rect 30297 7157 30331 7191
rect 30573 7157 30607 7191
rect 30849 7157 30883 7191
rect 31125 7157 31159 7191
rect 31953 7157 31987 7191
rect 32321 7157 32355 7191
rect 32873 7157 32907 7191
rect 33425 7157 33459 7191
rect 36001 7157 36035 7191
rect 37473 7157 37507 7191
rect 39129 7157 39163 7191
rect 5181 6953 5215 6987
rect 5733 6953 5767 6987
rect 10885 6953 10919 6987
rect 11437 6953 11471 6987
rect 11989 6953 12023 6987
rect 18889 6953 18923 6987
rect 19441 6885 19475 6919
rect 22017 6885 22051 6919
rect 6469 6817 6503 6851
rect 7021 6817 7055 6851
rect 7573 6817 7607 6851
rect 8125 6817 8159 6851
rect 8677 6817 8711 6851
rect 9597 6817 9631 6851
rect 10149 6817 10183 6851
rect 13277 6817 13311 6851
rect 13829 6817 13863 6851
rect 14657 6817 14691 6851
rect 15209 6817 15243 6851
rect 15761 6817 15795 6851
rect 16313 6817 16347 6851
rect 16865 6817 16899 6851
rect 17417 6817 17451 6851
rect 17969 6817 18003 6851
rect 18521 6817 18555 6851
rect 34345 6817 34379 6851
rect 35633 6817 35667 6851
rect 36185 6817 36219 6851
rect 37841 6817 37875 6851
rect 40785 6817 40819 6851
rect 5089 6749 5123 6783
rect 6745 6749 6779 6783
rect 7297 6749 7331 6783
rect 11345 6749 11379 6783
rect 14381 6749 14415 6783
rect 14933 6749 14967 6783
rect 19073 6749 19107 6783
rect 19257 6749 19291 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 20085 6749 20119 6783
rect 20361 6749 20395 6783
rect 20637 6749 20671 6783
rect 20913 6749 20947 6783
rect 21189 6749 21223 6783
rect 21465 6749 21499 6783
rect 22201 6749 22235 6783
rect 22293 6749 22327 6783
rect 22661 6749 22695 6783
rect 22937 6749 22971 6783
rect 25053 6749 25087 6783
rect 25329 6749 25363 6783
rect 25789 6749 25823 6783
rect 26157 6749 26191 6783
rect 26525 6749 26559 6783
rect 26893 6749 26927 6783
rect 27261 6749 27295 6783
rect 27537 6749 27571 6783
rect 27813 6749 27847 6783
rect 28365 6749 28399 6783
rect 28825 6749 28859 6783
rect 28917 6749 28951 6783
rect 29561 6749 29595 6783
rect 29837 6749 29871 6783
rect 30113 6749 30147 6783
rect 33057 6749 33091 6783
rect 33333 6749 33367 6783
rect 33609 6749 33643 6783
rect 36461 6749 36495 6783
rect 38669 6749 38703 6783
rect 5641 6681 5675 6715
rect 6193 6681 6227 6715
rect 7849 6681 7883 6715
rect 8401 6681 8435 6715
rect 9321 6681 9355 6715
rect 9873 6681 9907 6715
rect 10793 6681 10827 6715
rect 11897 6681 11931 6715
rect 12449 6681 12483 6715
rect 12817 6681 12851 6715
rect 13001 6681 13035 6715
rect 13553 6681 13587 6715
rect 15485 6681 15519 6715
rect 16037 6681 16071 6715
rect 16589 6681 16623 6715
rect 17141 6681 17175 6715
rect 17693 6681 17727 6715
rect 18245 6681 18279 6715
rect 35357 6681 35391 6715
rect 35909 6681 35943 6715
rect 37013 6681 37047 6715
rect 37565 6681 37599 6715
rect 38117 6681 38151 6715
rect 39221 6681 39255 6715
rect 39957 6681 39991 6715
rect 40509 6681 40543 6715
rect 19717 6613 19751 6647
rect 19993 6613 20027 6647
rect 20269 6613 20303 6647
rect 20545 6613 20579 6647
rect 20821 6613 20855 6647
rect 21097 6613 21131 6647
rect 21373 6613 21407 6647
rect 21649 6613 21683 6647
rect 22477 6613 22511 6647
rect 22845 6613 22879 6647
rect 23121 6613 23155 6647
rect 25237 6613 25271 6647
rect 25513 6613 25547 6647
rect 25973 6613 26007 6647
rect 26341 6613 26375 6647
rect 26709 6613 26743 6647
rect 27077 6613 27111 6647
rect 27445 6613 27479 6647
rect 27721 6613 27755 6647
rect 27997 6613 28031 6647
rect 28549 6613 28583 6647
rect 28641 6613 28675 6647
rect 29101 6613 29135 6647
rect 29745 6613 29779 6647
rect 30021 6613 30055 6647
rect 30297 6613 30331 6647
rect 33241 6613 33275 6647
rect 33517 6613 33551 6647
rect 33793 6613 33827 6647
rect 36553 6613 36587 6647
rect 37105 6613 37139 6647
rect 38209 6613 38243 6647
rect 38761 6613 38795 6647
rect 39313 6613 39347 6647
rect 40049 6613 40083 6647
rect 6377 6409 6411 6443
rect 7021 6409 7055 6443
rect 9229 6409 9263 6443
rect 9781 6409 9815 6443
rect 10333 6409 10367 6443
rect 10701 6409 10735 6443
rect 12541 6409 12575 6443
rect 12909 6409 12943 6443
rect 14197 6409 14231 6443
rect 14749 6409 14783 6443
rect 15485 6409 15519 6443
rect 15945 6409 15979 6443
rect 16313 6409 16347 6443
rect 16865 6409 16899 6443
rect 17601 6409 17635 6443
rect 18061 6409 18095 6443
rect 18429 6409 18463 6443
rect 18797 6409 18831 6443
rect 19533 6409 19567 6443
rect 9137 6341 9171 6375
rect 5917 6273 5951 6307
rect 6561 6273 6595 6307
rect 6929 6273 6963 6307
rect 9689 6273 9723 6307
rect 10241 6273 10275 6307
rect 10885 6273 10919 6307
rect 12449 6273 12483 6307
rect 13093 6273 13127 6307
rect 14105 6273 14139 6307
rect 14933 6273 14967 6307
rect 15209 6273 15243 6307
rect 15669 6273 15703 6307
rect 16129 6273 16163 6307
rect 16497 6273 16531 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 17785 6273 17819 6307
rect 18245 6273 18279 6307
rect 18613 6273 18647 6307
rect 18981 6273 19015 6307
rect 19349 6273 19383 6307
rect 19717 6273 19751 6307
rect 23213 6273 23247 6307
rect 23857 6273 23891 6307
rect 24225 6273 24259 6307
rect 5733 6137 5767 6171
rect 15025 6137 15059 6171
rect 17141 6137 17175 6171
rect 24041 6137 24075 6171
rect 24409 6137 24443 6171
rect 19165 6069 19199 6103
rect 23397 6069 23431 6103
rect 9781 5865 9815 5899
rect 9689 5661 9723 5695
rect 33977 3689 34011 3723
rect 34161 3485 34195 3519
rect 16865 3145 16899 3179
rect 33333 3145 33367 3179
rect 37841 3145 37875 3179
rect 16681 3009 16715 3043
rect 18613 3009 18647 3043
rect 20729 3009 20763 3043
rect 22661 3009 22695 3043
rect 24961 3009 24995 3043
rect 33517 3009 33551 3043
rect 38025 3009 38059 3043
rect 22845 2873 22879 2907
rect 25145 2873 25179 2907
rect 18797 2805 18831 2839
rect 20913 2805 20947 2839
rect 5641 2601 5675 2635
rect 16037 2601 16071 2635
rect 18153 2601 18187 2635
rect 20269 2601 20303 2635
rect 22385 2601 22419 2635
rect 24501 2601 24535 2635
rect 33425 2601 33459 2635
rect 33793 2601 33827 2635
rect 34713 2601 34747 2635
rect 37289 2601 37323 2635
rect 37841 2601 37875 2635
rect 39037 2601 39071 2635
rect 40141 2601 40175 2635
rect 42441 2601 42475 2635
rect 14749 2533 14783 2567
rect 33149 2533 33183 2567
rect 34253 2533 34287 2567
rect 37565 2533 37599 2567
rect 42993 2533 43027 2567
rect 12449 2465 12483 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 5457 2397 5491 2431
rect 7573 2397 7607 2431
rect 9689 2397 9723 2431
rect 11989 2397 12023 2431
rect 14289 2397 14323 2431
rect 16221 2397 16255 2431
rect 18337 2397 18371 2431
rect 20453 2397 20487 2431
rect 22569 2397 22603 2431
rect 24685 2397 24719 2431
rect 26617 2397 26651 2431
rect 28733 2397 28767 2431
rect 31033 2397 31067 2431
rect 33333 2397 33367 2431
rect 33609 2397 33643 2431
rect 33977 2397 34011 2431
rect 34437 2397 34471 2431
rect 34897 2397 34931 2431
rect 35265 2397 35299 2431
rect 35725 2397 35759 2431
rect 37473 2397 37507 2431
rect 37749 2397 37783 2431
rect 38025 2397 38059 2431
rect 39221 2397 39255 2431
rect 39497 2397 39531 2431
rect 40325 2397 40359 2431
rect 41613 2397 41647 2431
rect 42625 2397 42659 2431
rect 43177 2397 43211 2431
rect 12265 2329 12299 2363
rect 14565 2329 14599 2363
rect 7757 2261 7791 2295
rect 9873 2261 9907 2295
rect 11805 2261 11839 2295
rect 14105 2261 14139 2295
rect 26801 2261 26835 2295
rect 28917 2261 28951 2295
rect 30849 2261 30883 2295
rect 35081 2261 35115 2295
rect 35541 2261 35575 2295
rect 39313 2261 39347 2295
rect 41429 2261 41463 2295
<< metal1 >>
rect 16206 8508 16212 8560
rect 16264 8548 16270 8560
rect 33318 8548 33324 8560
rect 16264 8520 33324 8548
rect 16264 8508 16270 8520
rect 33318 8508 33324 8520
rect 33376 8508 33382 8560
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 33594 8480 33600 8492
rect 15804 8452 33600 8480
rect 15804 8440 15810 8452
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 15654 8372 15660 8424
rect 15712 8412 15718 8424
rect 33686 8412 33692 8424
rect 15712 8384 33692 8412
rect 15712 8372 15718 8384
rect 33686 8372 33692 8384
rect 33744 8372 33750 8424
rect 10502 8304 10508 8356
rect 10560 8344 10566 8356
rect 29270 8344 29276 8356
rect 10560 8316 29276 8344
rect 10560 8304 10566 8316
rect 29270 8304 29276 8316
rect 29328 8304 29334 8356
rect 24946 8236 24952 8288
rect 25004 8276 25010 8288
rect 25958 8276 25964 8288
rect 25004 8248 25964 8276
rect 25004 8236 25010 8248
rect 25958 8236 25964 8248
rect 26016 8236 26022 8288
rect 30190 8236 30196 8288
rect 30248 8276 30254 8288
rect 30650 8276 30656 8288
rect 30248 8248 30656 8276
rect 30248 8236 30254 8248
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 7190 8168 7196 8220
rect 7248 8208 7254 8220
rect 22830 8208 22836 8220
rect 7248 8180 22836 8208
rect 7248 8168 7254 8180
rect 22830 8168 22836 8180
rect 22888 8168 22894 8220
rect 25222 8168 25228 8220
rect 25280 8208 25286 8220
rect 26050 8208 26056 8220
rect 25280 8180 26056 8208
rect 25280 8168 25286 8180
rect 26050 8168 26056 8180
rect 26108 8168 26114 8220
rect 26160 8180 31432 8208
rect 15194 8140 15200 8152
rect 12544 8112 15200 8140
rect 11330 7964 11336 8016
rect 11388 8004 11394 8016
rect 12544 8004 12572 8112
rect 15194 8100 15200 8112
rect 15252 8100 15258 8152
rect 24486 8100 24492 8152
rect 24544 8140 24550 8152
rect 26160 8140 26188 8180
rect 24544 8112 26188 8140
rect 24544 8100 24550 8112
rect 27614 8100 27620 8152
rect 27672 8140 27678 8152
rect 28534 8140 28540 8152
rect 27672 8112 28540 8140
rect 27672 8100 27678 8112
rect 28534 8100 28540 8112
rect 28592 8100 28598 8152
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 20714 8072 20720 8084
rect 12676 8044 20720 8072
rect 12676 8032 12682 8044
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 24578 8032 24584 8084
rect 24636 8072 24642 8084
rect 24636 8044 30604 8072
rect 24636 8032 24642 8044
rect 30576 8016 30604 8044
rect 11388 7976 12572 8004
rect 11388 7964 11394 7976
rect 14366 7964 14372 8016
rect 14424 8004 14430 8016
rect 25682 8004 25688 8016
rect 14424 7976 25688 8004
rect 14424 7964 14430 7976
rect 25682 7964 25688 7976
rect 25740 7964 25746 8016
rect 27706 7964 27712 8016
rect 27764 8004 27770 8016
rect 28626 8004 28632 8016
rect 27764 7976 28632 8004
rect 27764 7964 27770 7976
rect 28626 7964 28632 7976
rect 28684 7964 28690 8016
rect 30558 7964 30564 8016
rect 30616 7964 30622 8016
rect 15102 7936 15108 7948
rect 7760 7908 15108 7936
rect 7760 7744 7788 7908
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 22002 7896 22008 7948
rect 22060 7936 22066 7948
rect 22060 7908 31156 7936
rect 22060 7896 22066 7908
rect 31128 7880 31156 7908
rect 31404 7880 31432 8180
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 20990 7868 20996 7880
rect 14056 7840 20996 7868
rect 14056 7828 14062 7840
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 30098 7868 30104 7880
rect 23808 7840 30104 7868
rect 23808 7828 23814 7840
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 31110 7828 31116 7880
rect 31168 7828 31174 7880
rect 31386 7828 31392 7880
rect 31444 7828 31450 7880
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 21266 7800 21272 7812
rect 12952 7772 21272 7800
rect 12952 7760 12958 7772
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 32398 7800 32404 7812
rect 22066 7772 32404 7800
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 16298 7732 16304 7744
rect 8352 7704 16304 7732
rect 8352 7692 8358 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 22066 7732 22094 7772
rect 32398 7760 32404 7772
rect 32456 7760 32462 7812
rect 16908 7704 22094 7732
rect 16908 7692 16914 7704
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 30834 7732 30840 7744
rect 22980 7704 30840 7732
rect 22980 7692 22986 7704
rect 30834 7692 30840 7704
rect 30892 7692 30898 7744
rect 1104 7642 43675 7664
rect 1104 7590 11552 7642
rect 11604 7590 11616 7642
rect 11668 7590 11680 7642
rect 11732 7590 11744 7642
rect 11796 7590 11808 7642
rect 11860 7590 22155 7642
rect 22207 7590 22219 7642
rect 22271 7590 22283 7642
rect 22335 7590 22347 7642
rect 22399 7590 22411 7642
rect 22463 7590 32758 7642
rect 32810 7590 32822 7642
rect 32874 7590 32886 7642
rect 32938 7590 32950 7642
rect 33002 7590 33014 7642
rect 33066 7590 43361 7642
rect 43413 7590 43425 7642
rect 43477 7590 43489 7642
rect 43541 7590 43553 7642
rect 43605 7590 43617 7642
rect 43669 7590 43675 7642
rect 1104 7568 43675 7590
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5350 7528 5356 7540
rect 5031 7500 5356 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5537 7531 5595 7537
rect 5537 7497 5549 7531
rect 5583 7528 5595 7531
rect 5902 7528 5908 7540
rect 5583 7500 5908 7528
rect 5583 7497 5595 7500
rect 5537 7491 5595 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7282 7528 7288 7540
rect 7055 7500 7288 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 6380 7460 6408 7491
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 7834 7528 7840 7540
rect 7607 7500 7840 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8386 7528 8392 7540
rect 8159 7500 8392 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7528 8723 7531
rect 8938 7528 8944 7540
rect 8711 7500 8944 7528
rect 8711 7497 8723 7500
rect 8665 7491 8723 7497
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10502 7528 10508 7540
rect 10091 7500 10508 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 10597 7531 10655 7537
rect 10597 7497 10609 7531
rect 10643 7528 10655 7531
rect 11146 7528 11152 7540
rect 10643 7500 11152 7528
rect 10643 7497 10655 7500
rect 10597 7491 10655 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 12526 7528 12532 7540
rect 12115 7500 12532 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13630 7528 13636 7540
rect 13311 7500 13636 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7528 13875 7531
rect 14182 7528 14188 7540
rect 13863 7500 14188 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15010 7528 15016 7540
rect 14783 7500 15016 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15562 7528 15568 7540
rect 15335 7500 15568 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 16022 7528 16028 7540
rect 15887 7500 16028 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 10520 7460 10548 7488
rect 10689 7463 10747 7469
rect 10689 7460 10701 7463
rect 5307 7432 6408 7460
rect 8404 7432 10456 7460
rect 10520 7432 10701 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 5534 7392 5540 7404
rect 4755 7364 5540 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6822 7392 6828 7404
rect 6779 7364 6828 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7324 6147 7327
rect 6454 7324 6460 7336
rect 6135 7296 6460 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 4338 7148 4344 7200
rect 4396 7148 4402 7200
rect 6564 7188 6592 7355
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7742 7392 7748 7404
rect 7331 7364 7748 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8294 7392 8300 7404
rect 7883 7364 8300 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8404 7401 8432 7432
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 10428 7392 10456 7432
rect 10689 7429 10701 7432
rect 10735 7429 10747 7463
rect 12894 7460 12900 7472
rect 10689 7423 10747 7429
rect 10796 7432 12900 7460
rect 10796 7392 10824 7432
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7429 13047 7463
rect 12989 7423 13047 7429
rect 13541 7463 13599 7469
rect 13541 7429 13553 7463
rect 13587 7460 13599 7463
rect 15930 7460 15936 7472
rect 13587 7432 15936 7460
rect 13587 7429 13599 7432
rect 13541 7423 13599 7429
rect 11241 7395 11299 7401
rect 11241 7392 11253 7395
rect 10428 7364 10824 7392
rect 10888 7364 11253 7392
rect 9677 7355 9735 7361
rect 9692 7324 9720 7355
rect 10888 7324 10916 7364
rect 11241 7361 11253 7364
rect 11287 7392 11299 7395
rect 11330 7392 11336 7404
rect 11287 7364 11336 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12066 7392 12072 7404
rect 11747 7364 12072 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12618 7392 12624 7404
rect 12207 7364 12624 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 9692 7296 10916 7324
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11882 7324 11888 7336
rect 11011 7296 11888 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12894 7324 12900 7336
rect 12406 7296 12900 7324
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 9858 7256 9864 7268
rect 8987 7228 9864 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 12406 7256 12434 7296
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 10980 7228 12434 7256
rect 10980 7188 11008 7228
rect 6564 7160 11008 7188
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11112 7160 11529 7188
rect 11112 7148 11118 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 13004 7188 13032 7423
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16684 7460 16712 7491
rect 17126 7488 17132 7540
rect 17184 7488 17190 7540
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 18230 7488 18236 7540
rect 18288 7488 18294 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 19208 7500 19441 7528
rect 19208 7488 19214 7500
rect 19429 7497 19441 7500
rect 19475 7497 19487 7531
rect 19429 7491 19487 7497
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7497 20039 7531
rect 19981 7491 20039 7497
rect 16163 7432 16712 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 18874 7420 18880 7472
rect 18932 7460 18938 7472
rect 19996 7460 20024 7491
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20588 7500 21465 7528
rect 20588 7488 20594 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 22005 7531 22063 7537
rect 22005 7497 22017 7531
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22020 7460 22048 7491
rect 22830 7488 22836 7540
rect 22888 7528 22894 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22888 7500 23029 7528
rect 22888 7488 22894 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 23937 7531 23995 7537
rect 23937 7497 23949 7531
rect 23983 7497 23995 7531
rect 24486 7528 24492 7540
rect 23937 7491 23995 7497
rect 24044 7500 24492 7528
rect 22554 7460 22560 7472
rect 18932 7432 20024 7460
rect 20364 7432 22048 7460
rect 22388 7432 22560 7460
rect 18932 7420 18938 7432
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14568 7364 15025 7392
rect 14093 7259 14151 7265
rect 14093 7225 14105 7259
rect 14139 7256 14151 7259
rect 14568 7256 14596 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16666 7392 16672 7404
rect 16531 7364 16672 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16850 7352 16856 7404
rect 16908 7352 16914 7404
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17218 7392 17224 7404
rect 17083 7364 17224 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17862 7392 17868 7404
rect 17635 7364 17868 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18506 7392 18512 7404
rect 18187 7364 18512 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18690 7352 18696 7404
rect 18748 7352 18754 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 20364 7401 20392 7432
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 20640 7324 20668 7355
rect 21082 7352 21088 7404
rect 21140 7352 21146 7404
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 21192 7324 21220 7355
rect 21634 7352 21640 7404
rect 21692 7352 21698 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22388 7392 22416 7432
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 23952 7460 23980 7491
rect 22848 7432 23980 7460
rect 22235 7364 22416 7392
rect 22465 7395 22523 7401
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22465 7361 22477 7395
rect 22511 7392 22523 7395
rect 22646 7392 22652 7404
rect 22511 7364 22652 7392
rect 22511 7361 22523 7364
rect 22465 7355 22523 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 22848 7401 22876 7432
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 23014 7352 23020 7404
rect 23072 7392 23078 7404
rect 23293 7395 23351 7401
rect 23293 7392 23305 7395
rect 23072 7364 23305 7392
rect 23072 7352 23078 7364
rect 23293 7361 23305 7364
rect 23339 7361 23351 7395
rect 23293 7355 23351 7361
rect 23566 7352 23572 7404
rect 23624 7352 23630 7404
rect 23658 7352 23664 7404
rect 23716 7392 23722 7404
rect 23845 7395 23903 7401
rect 23845 7392 23857 7395
rect 23716 7364 23857 7392
rect 23716 7352 23722 7364
rect 23845 7361 23857 7364
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 24044 7324 24072 7500
rect 24486 7488 24492 7500
rect 24544 7488 24550 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 24728 7500 25452 7528
rect 24728 7488 24734 7500
rect 24394 7420 24400 7472
rect 24452 7460 24458 7472
rect 24452 7432 24900 7460
rect 24452 7420 24458 7432
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24302 7352 24308 7404
rect 24360 7392 24366 7404
rect 24872 7401 24900 7432
rect 25424 7401 25452 7500
rect 25682 7488 25688 7540
rect 25740 7488 25746 7540
rect 26053 7531 26111 7537
rect 26053 7497 26065 7531
rect 26099 7497 26111 7531
rect 26053 7491 26111 7497
rect 26068 7460 26096 7491
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 26292 7500 27200 7528
rect 26292 7488 26298 7500
rect 25516 7432 26096 7460
rect 25516 7401 25544 7432
rect 26142 7420 26148 7472
rect 26200 7460 26206 7472
rect 26200 7432 26832 7460
rect 26200 7420 26206 7432
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24360 7364 24593 7392
rect 24360 7352 24366 7364
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24857 7395 24915 7401
rect 24857 7361 24869 7395
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 20640 7296 21128 7324
rect 21192 7296 22600 7324
rect 14139 7228 14596 7256
rect 14139 7225 14151 7228
rect 14093 7219 14151 7225
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 21100 7256 21128 7296
rect 22572 7265 22600 7296
rect 22756 7296 24072 7324
rect 24964 7324 24992 7355
rect 25590 7352 25596 7404
rect 25648 7392 25654 7404
rect 25648 7364 25912 7392
rect 25648 7352 25654 7364
rect 25884 7324 25912 7364
rect 25958 7352 25964 7404
rect 26016 7352 26022 7404
rect 26050 7352 26056 7404
rect 26108 7392 26114 7404
rect 26804 7401 26832 7432
rect 27172 7401 27200 7500
rect 27430 7488 27436 7540
rect 27488 7528 27494 7540
rect 27488 7500 27844 7528
rect 27488 7488 27494 7500
rect 27246 7420 27252 7472
rect 27304 7460 27310 7472
rect 27304 7432 27752 7460
rect 27304 7420 27310 7432
rect 27724 7401 27752 7432
rect 26237 7395 26295 7401
rect 26237 7392 26249 7395
rect 26108 7364 26249 7392
rect 26108 7352 26114 7364
rect 26237 7361 26249 7364
rect 26283 7361 26295 7395
rect 26237 7355 26295 7361
rect 26513 7395 26571 7401
rect 26513 7361 26525 7395
rect 26559 7361 26571 7395
rect 26513 7355 26571 7361
rect 26789 7395 26847 7401
rect 26789 7361 26801 7395
rect 26835 7361 26847 7395
rect 26789 7355 26847 7361
rect 27157 7395 27215 7401
rect 27157 7361 27169 7395
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27816 7392 27844 7500
rect 28718 7488 28724 7540
rect 28776 7528 28782 7540
rect 28776 7500 29408 7528
rect 28776 7488 28782 7500
rect 28350 7420 28356 7472
rect 28408 7460 28414 7472
rect 28408 7432 29132 7460
rect 28408 7420 28414 7432
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 27816 7364 27997 7392
rect 27709 7355 27767 7361
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28261 7395 28319 7401
rect 28261 7361 28273 7395
rect 28307 7361 28319 7395
rect 28261 7355 28319 7361
rect 26528 7324 26556 7355
rect 24964 7296 25820 7324
rect 25884 7296 26556 7324
rect 22756 7268 22784 7296
rect 22281 7259 22339 7265
rect 22281 7256 22293 7259
rect 16356 7228 20668 7256
rect 21100 7228 22293 7256
rect 16356 7216 16362 7228
rect 16482 7188 16488 7200
rect 13004 7160 16488 7188
rect 11517 7151 11575 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 16632 7160 20545 7188
rect 16632 7148 16638 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 20640 7188 20668 7228
rect 22281 7225 22293 7228
rect 22327 7225 22339 7259
rect 22281 7219 22339 7225
rect 22557 7259 22615 7265
rect 22557 7225 22569 7259
rect 22603 7225 22615 7259
rect 22557 7219 22615 7225
rect 22738 7216 22744 7268
rect 22796 7216 22802 7268
rect 23290 7216 23296 7268
rect 23348 7256 23354 7268
rect 25792 7265 25820 7296
rect 26694 7284 26700 7336
rect 26752 7324 26758 7336
rect 27448 7324 27476 7355
rect 26752 7296 27476 7324
rect 26752 7284 26758 7296
rect 25777 7259 25835 7265
rect 23348 7228 25176 7256
rect 23348 7216 23354 7228
rect 20809 7191 20867 7197
rect 20809 7188 20821 7191
rect 20640 7160 20821 7188
rect 20533 7151 20591 7157
rect 20809 7157 20821 7160
rect 20855 7157 20867 7191
rect 20809 7151 20867 7157
rect 20901 7191 20959 7197
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 20990 7188 20996 7200
rect 20947 7160 20996 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21232 7160 21373 7188
rect 21232 7148 21238 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 23106 7148 23112 7200
rect 23164 7148 23170 7200
rect 23382 7148 23388 7200
rect 23440 7148 23446 7200
rect 23658 7148 23664 7200
rect 23716 7148 23722 7200
rect 23842 7148 23848 7200
rect 23900 7188 23906 7200
rect 24397 7191 24455 7197
rect 24397 7188 24409 7191
rect 23900 7160 24409 7188
rect 23900 7148 23906 7160
rect 24397 7157 24409 7160
rect 24443 7157 24455 7191
rect 24397 7151 24455 7157
rect 24670 7148 24676 7200
rect 24728 7148 24734 7200
rect 25148 7197 25176 7228
rect 25777 7225 25789 7259
rect 25823 7225 25835 7259
rect 25777 7219 25835 7225
rect 26418 7216 26424 7268
rect 26476 7256 26482 7268
rect 26973 7259 27031 7265
rect 26973 7256 26985 7259
rect 26476 7228 26985 7256
rect 26476 7216 26482 7228
rect 26973 7225 26985 7228
rect 27019 7225 27031 7259
rect 26973 7219 27031 7225
rect 27430 7216 27436 7268
rect 27488 7256 27494 7268
rect 28276 7256 28304 7355
rect 28534 7352 28540 7404
rect 28592 7352 28598 7404
rect 28626 7352 28632 7404
rect 28684 7392 28690 7404
rect 29104 7401 29132 7432
rect 29380 7401 29408 7500
rect 30466 7488 30472 7540
rect 30524 7528 30530 7540
rect 30524 7500 31248 7528
rect 30524 7488 30530 7500
rect 29454 7420 29460 7472
rect 29512 7460 29518 7472
rect 29512 7432 30144 7460
rect 29512 7420 29518 7432
rect 30116 7401 30144 7432
rect 30282 7420 30288 7472
rect 30340 7460 30346 7472
rect 30340 7432 30972 7460
rect 30340 7420 30346 7432
rect 28813 7395 28871 7401
rect 28813 7392 28825 7395
rect 28684 7364 28825 7392
rect 28684 7352 28690 7364
rect 28813 7361 28825 7364
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 29365 7395 29423 7401
rect 29365 7361 29377 7395
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 29733 7395 29791 7401
rect 29733 7361 29745 7395
rect 29779 7361 29791 7395
rect 29733 7355 29791 7361
rect 30009 7395 30067 7401
rect 30009 7361 30021 7395
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 30101 7395 30159 7401
rect 30101 7361 30113 7395
rect 30147 7361 30159 7395
rect 30101 7355 30159 7361
rect 28994 7284 29000 7336
rect 29052 7324 29058 7336
rect 29748 7324 29776 7355
rect 29052 7296 29776 7324
rect 29052 7284 29058 7296
rect 27488 7228 28304 7256
rect 27488 7216 27494 7228
rect 29086 7216 29092 7268
rect 29144 7256 29150 7268
rect 30024 7256 30052 7355
rect 30190 7352 30196 7404
rect 30248 7392 30254 7404
rect 30377 7395 30435 7401
rect 30377 7392 30389 7395
rect 30248 7364 30389 7392
rect 30248 7352 30254 7364
rect 30377 7361 30389 7364
rect 30423 7361 30435 7395
rect 30377 7355 30435 7361
rect 30650 7352 30656 7404
rect 30708 7352 30714 7404
rect 30944 7401 30972 7432
rect 31220 7401 31248 7500
rect 31386 7488 31392 7540
rect 31444 7488 31450 7540
rect 31662 7488 31668 7540
rect 31720 7528 31726 7540
rect 31720 7500 32444 7528
rect 31720 7488 31726 7500
rect 31294 7420 31300 7472
rect 31352 7460 31358 7472
rect 31352 7432 31800 7460
rect 31352 7420 31358 7432
rect 31772 7401 31800 7432
rect 30929 7395 30987 7401
rect 30929 7361 30941 7395
rect 30975 7361 30987 7395
rect 30929 7355 30987 7361
rect 31205 7395 31263 7401
rect 31205 7361 31217 7395
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7361 31539 7395
rect 31481 7355 31539 7361
rect 31757 7395 31815 7401
rect 31757 7361 31769 7395
rect 31803 7361 31815 7395
rect 31757 7355 31815 7361
rect 30742 7284 30748 7336
rect 30800 7324 30806 7336
rect 31496 7324 31524 7355
rect 31846 7352 31852 7404
rect 31904 7392 31910 7404
rect 32416 7401 32444 7500
rect 32766 7488 32772 7540
rect 32824 7528 32830 7540
rect 32824 7500 33548 7528
rect 32824 7488 32830 7500
rect 32490 7420 32496 7472
rect 32548 7460 32554 7472
rect 32548 7432 32996 7460
rect 32548 7420 32554 7432
rect 32968 7401 32996 7432
rect 33520 7401 33548 7500
rect 33686 7488 33692 7540
rect 33744 7488 33750 7540
rect 33778 7488 33784 7540
rect 33836 7528 33842 7540
rect 34057 7531 34115 7537
rect 34057 7528 34069 7531
rect 33836 7500 34069 7528
rect 33836 7488 33842 7500
rect 34057 7497 34069 7500
rect 34103 7497 34115 7531
rect 34057 7491 34115 7497
rect 34330 7488 34336 7540
rect 34388 7528 34394 7540
rect 34885 7531 34943 7537
rect 34885 7528 34897 7531
rect 34388 7500 34897 7528
rect 34388 7488 34394 7500
rect 34885 7497 34897 7500
rect 34931 7497 34943 7531
rect 34885 7491 34943 7497
rect 35437 7531 35495 7537
rect 35437 7497 35449 7531
rect 35483 7497 35495 7531
rect 35437 7491 35495 7497
rect 34606 7420 34612 7472
rect 34664 7460 34670 7472
rect 35452 7460 35480 7491
rect 35618 7488 35624 7540
rect 35676 7528 35682 7540
rect 36541 7531 36599 7537
rect 36541 7528 36553 7531
rect 35676 7500 36553 7528
rect 35676 7488 35682 7500
rect 36541 7497 36553 7500
rect 36587 7497 36599 7531
rect 36541 7491 36599 7497
rect 36909 7531 36967 7537
rect 36909 7497 36921 7531
rect 36955 7528 36967 7531
rect 36955 7500 38516 7528
rect 36955 7497 36967 7500
rect 36909 7491 36967 7497
rect 34664 7432 35480 7460
rect 34664 7420 34670 7432
rect 36998 7420 37004 7472
rect 37056 7460 37062 7472
rect 38488 7469 38516 7500
rect 39482 7488 39488 7540
rect 39540 7528 39546 7540
rect 40589 7531 40647 7537
rect 40589 7528 40601 7531
rect 39540 7500 40601 7528
rect 39540 7488 39546 7500
rect 40589 7497 40601 7500
rect 40635 7497 40647 7531
rect 40589 7491 40647 7497
rect 38289 7463 38347 7469
rect 38289 7460 38301 7463
rect 37056 7432 38301 7460
rect 37056 7420 37062 7432
rect 38289 7429 38301 7432
rect 38335 7429 38347 7463
rect 38289 7423 38347 7429
rect 38473 7463 38531 7469
rect 38473 7429 38485 7463
rect 38519 7429 38531 7463
rect 38473 7423 38531 7429
rect 38930 7420 38936 7472
rect 38988 7460 38994 7472
rect 40313 7463 40371 7469
rect 40313 7460 40325 7463
rect 38988 7432 40325 7460
rect 38988 7420 38994 7432
rect 40313 7429 40325 7432
rect 40359 7429 40371 7463
rect 40313 7423 40371 7429
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31904 7364 32137 7392
rect 31904 7352 31910 7364
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 32401 7395 32459 7401
rect 32401 7361 32413 7395
rect 32447 7361 32459 7395
rect 32401 7355 32459 7361
rect 32677 7395 32735 7401
rect 32677 7361 32689 7395
rect 32723 7361 32735 7395
rect 32677 7355 32735 7361
rect 32953 7395 33011 7401
rect 32953 7361 32965 7395
rect 32999 7361 33011 7395
rect 32953 7355 33011 7361
rect 33229 7395 33287 7401
rect 33229 7361 33241 7395
rect 33275 7361 33287 7395
rect 33229 7355 33287 7361
rect 33505 7395 33563 7401
rect 33505 7361 33517 7395
rect 33551 7361 33563 7395
rect 33505 7355 33563 7361
rect 33965 7395 34023 7401
rect 33965 7361 33977 7395
rect 34011 7361 34023 7395
rect 33965 7355 34023 7361
rect 30800 7296 31524 7324
rect 30800 7284 30806 7296
rect 31938 7284 31944 7336
rect 31996 7324 32002 7336
rect 32692 7324 32720 7355
rect 31996 7296 32720 7324
rect 31996 7284 32002 7296
rect 32858 7284 32864 7336
rect 32916 7324 32922 7336
rect 33244 7324 33272 7355
rect 32916 7296 33272 7324
rect 32916 7284 32922 7296
rect 33318 7284 33324 7336
rect 33376 7284 33382 7336
rect 33410 7284 33416 7336
rect 33468 7324 33474 7336
rect 33980 7324 34008 7355
rect 34146 7352 34152 7404
rect 34204 7392 34210 7404
rect 34793 7395 34851 7401
rect 34793 7392 34805 7395
rect 34204 7364 34805 7392
rect 34204 7352 34210 7364
rect 34793 7361 34805 7364
rect 34839 7361 34851 7395
rect 34793 7355 34851 7361
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 35897 7395 35955 7401
rect 35897 7361 35909 7395
rect 35943 7361 35955 7395
rect 35897 7355 35955 7361
rect 33468 7296 34008 7324
rect 33468 7284 33474 7296
rect 34422 7284 34428 7336
rect 34480 7324 34486 7336
rect 35360 7324 35388 7355
rect 34480 7296 35388 7324
rect 34480 7284 34486 7296
rect 29144 7228 30052 7256
rect 29144 7216 29150 7228
rect 30098 7216 30104 7268
rect 30156 7256 30162 7268
rect 30156 7228 30328 7256
rect 30156 7216 30162 7228
rect 25133 7191 25191 7197
rect 25133 7157 25145 7191
rect 25179 7157 25191 7191
rect 25133 7151 25191 7157
rect 25222 7148 25228 7200
rect 25280 7148 25286 7200
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 25924 7160 26341 7188
rect 25924 7148 25930 7160
rect 26329 7157 26341 7160
rect 26375 7157 26387 7191
rect 26329 7151 26387 7157
rect 26602 7148 26608 7200
rect 26660 7148 26666 7200
rect 27062 7148 27068 7200
rect 27120 7188 27126 7200
rect 27249 7191 27307 7197
rect 27249 7188 27261 7191
rect 27120 7160 27261 7188
rect 27120 7148 27126 7160
rect 27249 7157 27261 7160
rect 27295 7157 27307 7191
rect 27249 7151 27307 7157
rect 27338 7148 27344 7200
rect 27396 7188 27402 7200
rect 27525 7191 27583 7197
rect 27525 7188 27537 7191
rect 27396 7160 27537 7188
rect 27396 7148 27402 7160
rect 27525 7157 27537 7160
rect 27571 7157 27583 7191
rect 27525 7151 27583 7157
rect 27798 7148 27804 7200
rect 27856 7148 27862 7200
rect 28074 7148 28080 7200
rect 28132 7148 28138 7200
rect 28166 7148 28172 7200
rect 28224 7188 28230 7200
rect 28353 7191 28411 7197
rect 28353 7188 28365 7191
rect 28224 7160 28365 7188
rect 28224 7148 28230 7160
rect 28353 7157 28365 7160
rect 28399 7157 28411 7191
rect 28353 7151 28411 7157
rect 28626 7148 28632 7200
rect 28684 7148 28690 7200
rect 28718 7148 28724 7200
rect 28776 7188 28782 7200
rect 28905 7191 28963 7197
rect 28905 7188 28917 7191
rect 28776 7160 28917 7188
rect 28776 7148 28782 7160
rect 28905 7157 28917 7160
rect 28951 7157 28963 7191
rect 28905 7151 28963 7157
rect 29178 7148 29184 7200
rect 29236 7148 29242 7200
rect 29549 7191 29607 7197
rect 29549 7157 29561 7191
rect 29595 7188 29607 7191
rect 29730 7188 29736 7200
rect 29595 7160 29736 7188
rect 29595 7157 29607 7160
rect 29549 7151 29607 7157
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 29825 7191 29883 7197
rect 29825 7157 29837 7191
rect 29871 7188 29883 7191
rect 30006 7188 30012 7200
rect 29871 7160 30012 7188
rect 29871 7157 29883 7160
rect 29825 7151 29883 7157
rect 30006 7148 30012 7160
rect 30064 7148 30070 7200
rect 30300 7197 30328 7228
rect 30374 7216 30380 7268
rect 30432 7256 30438 7268
rect 31665 7259 31723 7265
rect 31665 7256 31677 7259
rect 30432 7228 31677 7256
rect 30432 7216 30438 7228
rect 31665 7225 31677 7228
rect 31711 7225 31723 7259
rect 31665 7219 31723 7225
rect 31754 7216 31760 7268
rect 31812 7256 31818 7268
rect 32585 7259 32643 7265
rect 32585 7256 32597 7259
rect 31812 7228 32597 7256
rect 31812 7216 31818 7228
rect 32585 7225 32597 7228
rect 32631 7225 32643 7259
rect 32585 7219 32643 7225
rect 33137 7259 33195 7265
rect 33137 7225 33149 7259
rect 33183 7256 33195 7259
rect 33336 7256 33364 7284
rect 33183 7228 33364 7256
rect 33183 7225 33195 7228
rect 33137 7219 33195 7225
rect 33594 7216 33600 7268
rect 33652 7216 33658 7268
rect 34790 7216 34796 7268
rect 34848 7256 34854 7268
rect 35912 7256 35940 7355
rect 36078 7352 36084 7404
rect 36136 7392 36142 7404
rect 36449 7395 36507 7401
rect 36449 7392 36461 7395
rect 36136 7364 36461 7392
rect 36136 7352 36142 7364
rect 36449 7361 36461 7364
rect 36495 7361 36507 7395
rect 36449 7355 36507 7361
rect 36906 7352 36912 7404
rect 36964 7392 36970 7404
rect 37093 7395 37151 7401
rect 37093 7392 37105 7395
rect 36964 7364 37105 7392
rect 36964 7352 36970 7364
rect 37093 7361 37105 7364
rect 37139 7361 37151 7395
rect 37093 7355 37151 7361
rect 37366 7352 37372 7404
rect 37424 7352 37430 7404
rect 37826 7352 37832 7404
rect 37884 7392 37890 7404
rect 37921 7395 37979 7401
rect 37921 7392 37933 7395
rect 37884 7364 37933 7392
rect 37884 7352 37890 7364
rect 37921 7361 37933 7364
rect 37967 7361 37979 7395
rect 37921 7355 37979 7361
rect 38746 7352 38752 7404
rect 38804 7392 38810 7404
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 38804 7364 39037 7392
rect 38804 7352 38810 7364
rect 39025 7361 39037 7364
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 39945 7395 40003 7401
rect 39945 7361 39957 7395
rect 39991 7361 40003 7395
rect 39945 7355 40003 7361
rect 38562 7284 38568 7336
rect 38620 7324 38626 7336
rect 39960 7324 39988 7355
rect 40494 7352 40500 7404
rect 40552 7352 40558 7404
rect 38620 7296 39988 7324
rect 38620 7284 38626 7296
rect 34848 7228 35940 7256
rect 34848 7216 34854 7228
rect 38654 7216 38660 7268
rect 38712 7216 38718 7268
rect 30285 7191 30343 7197
rect 30285 7157 30297 7191
rect 30331 7157 30343 7191
rect 30285 7151 30343 7157
rect 30558 7148 30564 7200
rect 30616 7148 30622 7200
rect 30834 7148 30840 7200
rect 30892 7148 30898 7200
rect 31110 7148 31116 7200
rect 31168 7148 31174 7200
rect 31941 7191 31999 7197
rect 31941 7157 31953 7191
rect 31987 7188 31999 7191
rect 32122 7188 32128 7200
rect 31987 7160 32128 7188
rect 31987 7157 31999 7160
rect 31941 7151 31999 7157
rect 32122 7148 32128 7160
rect 32180 7148 32186 7200
rect 32306 7148 32312 7200
rect 32364 7148 32370 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32456 7160 32873 7188
rect 32456 7148 32462 7160
rect 32861 7157 32873 7160
rect 32907 7157 32919 7191
rect 32861 7151 32919 7157
rect 33413 7191 33471 7197
rect 33413 7157 33425 7191
rect 33459 7188 33471 7191
rect 33612 7188 33640 7216
rect 33459 7160 33640 7188
rect 33459 7157 33471 7160
rect 33413 7151 33471 7157
rect 35066 7148 35072 7200
rect 35124 7188 35130 7200
rect 35989 7191 36047 7197
rect 35989 7188 36001 7191
rect 35124 7160 36001 7188
rect 35124 7148 35130 7160
rect 35989 7157 36001 7160
rect 36035 7157 36047 7191
rect 35989 7151 36047 7157
rect 36446 7148 36452 7200
rect 36504 7188 36510 7200
rect 37461 7191 37519 7197
rect 37461 7188 37473 7191
rect 36504 7160 37473 7188
rect 36504 7148 36510 7160
rect 37461 7157 37473 7160
rect 37507 7157 37519 7191
rect 37461 7151 37519 7157
rect 39114 7148 39120 7200
rect 39172 7148 39178 7200
rect 1104 7098 43516 7120
rect 1104 7046 6251 7098
rect 6303 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 16854 7098
rect 16906 7046 16918 7098
rect 16970 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 27457 7098
rect 27509 7046 27521 7098
rect 27573 7046 27585 7098
rect 27637 7046 27649 7098
rect 27701 7046 27713 7098
rect 27765 7046 38060 7098
rect 38112 7046 38124 7098
rect 38176 7046 38188 7098
rect 38240 7046 38252 7098
rect 38304 7046 38316 7098
rect 38368 7046 43516 7098
rect 1104 7024 43516 7046
rect 5166 6944 5172 6996
rect 5224 6944 5230 6996
rect 5718 6944 5724 6996
rect 5776 6944 5782 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9180 6956 10824 6984
rect 9180 6944 9186 6956
rect 10796 6916 10824 6956
rect 10870 6944 10876 6996
rect 10928 6944 10934 6996
rect 11422 6944 11428 6996
rect 11480 6944 11486 6996
rect 11974 6944 11980 6996
rect 12032 6944 12038 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 18598 6984 18604 6996
rect 12124 6956 18604 6984
rect 12124 6944 12130 6956
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18748 6956 18889 6984
rect 18748 6944 18754 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 18966 6944 18972 6996
rect 19024 6984 19030 6996
rect 20806 6984 20812 6996
rect 19024 6956 20812 6984
rect 19024 6944 19030 6956
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 22922 6984 22928 6996
rect 21008 6956 22928 6984
rect 12342 6916 12348 6928
rect 8588 6888 8800 6916
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6236 6820 6469 6848
rect 6236 6808 6242 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 7006 6808 7012 6860
rect 7064 6808 7070 6860
rect 7558 6808 7564 6860
rect 7616 6808 7622 6860
rect 8110 6808 8116 6860
rect 8168 6808 8174 6860
rect 8588 6848 8616 6888
rect 8312 6820 8616 6848
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4396 6752 5089 6780
rect 4396 6740 4402 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7190 6780 7196 6792
rect 6779 6752 7196 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 8312 6780 8340 6820
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8772 6848 8800 6888
rect 9508 6888 10732 6916
rect 10796 6888 12348 6916
rect 9508 6848 9536 6888
rect 8772 6820 9536 6848
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 10042 6848 10048 6860
rect 9631 6820 10048 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10594 6848 10600 6860
rect 10183 6820 10600 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10704 6848 10732 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 19429 6919 19487 6925
rect 19429 6916 19441 6919
rect 12952 6888 19441 6916
rect 12952 6876 12958 6888
rect 19429 6885 19441 6888
rect 19475 6885 19487 6919
rect 19429 6879 19487 6885
rect 12158 6848 12164 6860
rect 10704 6820 12164 6848
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12860 6820 13277 6848
rect 12860 6808 12866 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13412 6820 13829 6848
rect 13412 6808 13418 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 14642 6808 14648 6860
rect 14700 6808 14706 6860
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15197 6851 15255 6857
rect 15197 6848 15209 6851
rect 14792 6820 15209 6848
rect 14792 6808 14798 6820
rect 15197 6817 15209 6820
rect 15243 6817 15255 6851
rect 15197 6811 15255 6817
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15344 6820 15761 6848
rect 15344 6808 15350 6820
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 15749 6811 15807 6817
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15896 6820 16313 6848
rect 15896 6808 15902 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16853 6851 16911 6857
rect 16853 6848 16865 6851
rect 16448 6820 16865 6848
rect 16448 6808 16454 6820
rect 16853 6817 16865 6820
rect 16899 6817 16911 6851
rect 16853 6811 16911 6817
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17000 6820 17417 6848
rect 17000 6808 17006 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17552 6820 17969 6848
rect 17552 6808 17558 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 18104 6820 18521 6848
rect 18104 6808 18110 6820
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 21008 6848 21036 6956
rect 22922 6944 22928 6956
rect 22980 6944 22986 6996
rect 23106 6944 23112 6996
rect 23164 6944 23170 6996
rect 23658 6944 23664 6996
rect 23716 6944 23722 6996
rect 25866 6944 25872 6996
rect 25924 6944 25930 6996
rect 26602 6944 26608 6996
rect 26660 6944 26666 6996
rect 27062 6944 27068 6996
rect 27120 6944 27126 6996
rect 27798 6984 27804 6996
rect 27172 6956 27804 6984
rect 22005 6919 22063 6925
rect 22005 6885 22017 6919
rect 22051 6885 22063 6919
rect 23124 6916 23152 6944
rect 22005 6879 22063 6885
rect 22296 6888 23152 6916
rect 22020 6848 22048 6879
rect 18509 6811 18567 6817
rect 19076 6820 21036 6848
rect 21192 6820 22048 6848
rect 11333 6783 11391 6789
rect 7331 6752 8340 6780
rect 8404 6752 11284 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 5626 6672 5632 6724
rect 5684 6672 5690 6724
rect 6178 6672 6184 6724
rect 6236 6672 6242 6724
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 8404 6721 8432 6752
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6681 8447 6715
rect 8389 6675 8447 6681
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6681 9367 6715
rect 9309 6675 9367 6681
rect 9861 6715 9919 6721
rect 9861 6681 9873 6715
rect 9907 6712 9919 6715
rect 10594 6712 10600 6724
rect 9907 6684 10600 6712
rect 9907 6681 9919 6684
rect 9861 6675 9919 6681
rect 9324 6644 9352 6675
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 11256 6712 11284 6752
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 12618 6780 12624 6792
rect 11379 6752 12624 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13078 6780 13084 6792
rect 12820 6752 13084 6780
rect 11606 6712 11612 6724
rect 11256 6684 11612 6712
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 11882 6672 11888 6724
rect 11940 6672 11946 6724
rect 12437 6715 12495 6721
rect 12437 6681 12449 6715
rect 12483 6712 12495 6715
rect 12710 6712 12716 6724
rect 12483 6684 12716 6712
rect 12483 6681 12495 6684
rect 12437 6675 12495 6681
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 12820 6721 12848 6752
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 14182 6780 14188 6792
rect 13464 6752 14188 6780
rect 12805 6715 12863 6721
rect 12805 6681 12817 6715
rect 12851 6681 12863 6715
rect 12805 6675 12863 6681
rect 12989 6715 13047 6721
rect 12989 6681 13001 6715
rect 13035 6712 13047 6715
rect 13464 6712 13492 6752
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6780 14979 6783
rect 18414 6780 18420 6792
rect 14967 6752 18420 6780
rect 14967 6749 14979 6752
rect 14921 6743 14979 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 19076 6789 19104 6820
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6749 19119 6783
rect 19061 6743 19119 6749
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6780 19303 6783
rect 19426 6780 19432 6792
rect 19291 6752 19432 6780
rect 19291 6749 19303 6752
rect 19245 6743 19303 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 13035 6684 13492 6712
rect 13541 6715 13599 6721
rect 13035 6681 13047 6684
rect 12989 6675 13047 6681
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 15010 6712 15016 6724
rect 13587 6684 15016 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15473 6715 15531 6721
rect 15473 6712 15485 6715
rect 15160 6684 15485 6712
rect 15160 6672 15166 6684
rect 15473 6681 15485 6684
rect 15519 6681 15531 6715
rect 15473 6675 15531 6681
rect 16022 6672 16028 6724
rect 16080 6672 16086 6724
rect 16574 6672 16580 6724
rect 16632 6672 16638 6724
rect 17126 6672 17132 6724
rect 17184 6672 17190 6724
rect 17678 6672 17684 6724
rect 17736 6672 17742 6724
rect 18230 6672 18236 6724
rect 18288 6672 18294 6724
rect 19610 6712 19616 6724
rect 18340 6684 19616 6712
rect 10686 6644 10692 6656
rect 9324 6616 10692 6644
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 18340 6644 18368 6684
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 19812 6712 19840 6743
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 20346 6740 20352 6792
rect 20404 6740 20410 6792
rect 20530 6740 20536 6792
rect 20588 6740 20594 6792
rect 20622 6740 20628 6792
rect 20680 6740 20686 6792
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 21192 6789 21220 6820
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22296 6789 22324 6888
rect 23676 6848 23704 6944
rect 25884 6916 25912 6944
rect 26620 6916 26648 6944
rect 22940 6820 23704 6848
rect 25056 6888 25912 6916
rect 26068 6888 26648 6916
rect 22940 6789 22968 6820
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21968 6752 22201 6780
rect 21968 6740 21974 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6749 22339 6783
rect 22281 6743 22339 6749
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 22925 6783 22983 6789
rect 22925 6749 22937 6783
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 20548 6712 20576 6740
rect 19812 6684 20576 6712
rect 20824 6712 20852 6740
rect 22664 6712 22692 6743
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 25056 6789 25084 6888
rect 26068 6848 26096 6888
rect 27080 6848 27108 6944
rect 25332 6820 26096 6848
rect 26160 6820 27108 6848
rect 25332 6789 25360 6820
rect 26160 6789 26188 6820
rect 25041 6783 25099 6789
rect 23256 6752 23612 6780
rect 23256 6740 23262 6752
rect 23382 6712 23388 6724
rect 20824 6684 21680 6712
rect 22664 6684 23388 6712
rect 10928 6616 18368 6644
rect 10928 6604 10934 6616
rect 18414 6604 18420 6656
rect 18472 6644 18478 6656
rect 19705 6647 19763 6653
rect 19705 6644 19717 6647
rect 18472 6616 19717 6644
rect 18472 6604 18478 6616
rect 19705 6613 19717 6616
rect 19751 6613 19763 6647
rect 19705 6607 19763 6613
rect 19978 6604 19984 6656
rect 20036 6604 20042 6656
rect 20254 6604 20260 6656
rect 20312 6604 20318 6656
rect 20530 6604 20536 6656
rect 20588 6604 20594 6656
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 20680 6616 20821 6644
rect 20680 6604 20686 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 21082 6604 21088 6656
rect 21140 6604 21146 6656
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21652 6653 21680 6684
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 21361 6647 21419 6653
rect 21361 6644 21373 6647
rect 21324 6616 21373 6644
rect 21324 6604 21330 6616
rect 21361 6613 21373 6616
rect 21407 6613 21419 6647
rect 21361 6607 21419 6613
rect 21637 6647 21695 6653
rect 21637 6613 21649 6647
rect 21683 6613 21695 6647
rect 21637 6607 21695 6613
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 22465 6647 22523 6653
rect 22465 6644 22477 6647
rect 21784 6616 22477 6644
rect 21784 6604 21790 6616
rect 22465 6613 22477 6616
rect 22511 6613 22523 6647
rect 22465 6607 22523 6613
rect 22830 6604 22836 6656
rect 22888 6604 22894 6656
rect 23106 6604 23112 6656
rect 23164 6604 23170 6656
rect 23584 6644 23612 6752
rect 25041 6749 25053 6783
rect 25087 6749 25099 6783
rect 25041 6743 25099 6749
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 25777 6783 25835 6789
rect 25777 6749 25789 6783
rect 25823 6749 25835 6783
rect 25777 6743 25835 6749
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 25792 6712 25820 6743
rect 26418 6740 26424 6792
rect 26476 6740 26482 6792
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6749 26571 6783
rect 26513 6743 26571 6749
rect 26881 6783 26939 6789
rect 26881 6749 26893 6783
rect 26927 6780 26939 6783
rect 27172 6780 27200 6956
rect 27798 6944 27804 6956
rect 27856 6944 27862 6996
rect 28074 6944 28080 6996
rect 28132 6944 28138 6996
rect 28626 6944 28632 6996
rect 28684 6944 28690 6996
rect 28092 6916 28120 6944
rect 27632 6888 28120 6916
rect 27632 6848 27660 6888
rect 28644 6848 28672 6944
rect 37550 6876 37556 6928
rect 37608 6916 37614 6928
rect 37608 6888 37964 6916
rect 37608 6876 37614 6888
rect 27264 6820 27660 6848
rect 27816 6820 28672 6848
rect 27264 6789 27292 6820
rect 26927 6752 27200 6780
rect 27249 6783 27307 6789
rect 26927 6749 26939 6752
rect 26881 6743 26939 6749
rect 27249 6749 27261 6783
rect 27295 6749 27307 6783
rect 27249 6743 27307 6749
rect 26436 6712 26464 6740
rect 25792 6684 26464 6712
rect 26528 6712 26556 6743
rect 27338 6740 27344 6792
rect 27396 6740 27402 6792
rect 27816 6789 27844 6820
rect 34054 6808 34060 6860
rect 34112 6848 34118 6860
rect 34333 6851 34391 6857
rect 34333 6848 34345 6851
rect 34112 6820 34345 6848
rect 34112 6808 34118 6820
rect 34333 6817 34345 6820
rect 34379 6817 34391 6851
rect 34333 6811 34391 6817
rect 35158 6808 35164 6860
rect 35216 6848 35222 6860
rect 35621 6851 35679 6857
rect 35621 6848 35633 6851
rect 35216 6820 35633 6848
rect 35216 6808 35222 6820
rect 35621 6817 35633 6820
rect 35667 6817 35679 6851
rect 35621 6811 35679 6817
rect 35710 6808 35716 6860
rect 35768 6848 35774 6860
rect 36173 6851 36231 6857
rect 36173 6848 36185 6851
rect 35768 6820 36185 6848
rect 35768 6808 35774 6820
rect 36173 6817 36185 6820
rect 36219 6817 36231 6851
rect 36173 6811 36231 6817
rect 37090 6808 37096 6860
rect 37148 6848 37154 6860
rect 37829 6851 37887 6857
rect 37829 6848 37841 6851
rect 37148 6820 37841 6848
rect 37148 6808 37154 6820
rect 37829 6817 37841 6820
rect 37875 6817 37887 6851
rect 37936 6848 37964 6888
rect 38286 6848 38292 6860
rect 37936 6820 38292 6848
rect 37829 6811 37887 6817
rect 38286 6808 38292 6820
rect 38344 6808 38350 6860
rect 39574 6808 39580 6860
rect 39632 6848 39638 6860
rect 40773 6851 40831 6857
rect 40773 6848 40785 6851
rect 39632 6820 40785 6848
rect 39632 6808 39638 6820
rect 40773 6817 40785 6820
rect 40819 6817 40831 6851
rect 40773 6811 40831 6817
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6749 27859 6783
rect 27801 6743 27859 6749
rect 27356 6712 27384 6740
rect 26528 6684 27384 6712
rect 27540 6712 27568 6743
rect 28166 6740 28172 6792
rect 28224 6740 28230 6792
rect 28353 6783 28411 6789
rect 28353 6749 28365 6783
rect 28399 6780 28411 6783
rect 28718 6780 28724 6792
rect 28399 6752 28724 6780
rect 28399 6749 28411 6752
rect 28353 6743 28411 6749
rect 28718 6740 28724 6752
rect 28776 6740 28782 6792
rect 28810 6740 28816 6792
rect 28868 6740 28874 6792
rect 28905 6783 28963 6789
rect 28905 6749 28917 6783
rect 28951 6780 28963 6783
rect 29178 6780 29184 6792
rect 28951 6752 29184 6780
rect 28951 6749 28963 6752
rect 28905 6743 28963 6749
rect 29178 6740 29184 6752
rect 29236 6740 29242 6792
rect 29549 6783 29607 6789
rect 29549 6749 29561 6783
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 28184 6712 28212 6740
rect 29564 6712 29592 6743
rect 29730 6740 29736 6792
rect 29788 6780 29794 6792
rect 29825 6783 29883 6789
rect 29825 6780 29837 6783
rect 29788 6752 29837 6780
rect 29788 6740 29794 6752
rect 29825 6749 29837 6752
rect 29871 6749 29883 6783
rect 29825 6743 29883 6749
rect 30006 6740 30012 6792
rect 30064 6780 30070 6792
rect 30101 6783 30159 6789
rect 30101 6780 30113 6783
rect 30064 6752 30113 6780
rect 30064 6740 30070 6752
rect 30101 6749 30113 6752
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 33042 6740 33048 6792
rect 33100 6740 33106 6792
rect 33318 6740 33324 6792
rect 33376 6740 33382 6792
rect 33594 6740 33600 6792
rect 33652 6740 33658 6792
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 36449 6783 36507 6789
rect 36449 6780 36461 6783
rect 33744 6752 36461 6780
rect 33744 6740 33750 6752
rect 36449 6749 36461 6752
rect 36495 6749 36507 6783
rect 36449 6743 36507 6749
rect 36722 6740 36728 6792
rect 36780 6780 36786 6792
rect 38657 6783 38715 6789
rect 36780 6752 37596 6780
rect 36780 6740 36786 6752
rect 27540 6684 28212 6712
rect 28644 6684 29592 6712
rect 25225 6647 25283 6653
rect 25225 6644 25237 6647
rect 23584 6616 25237 6644
rect 25225 6613 25237 6616
rect 25271 6613 25283 6647
rect 25225 6607 25283 6613
rect 25498 6604 25504 6656
rect 25556 6604 25562 6656
rect 25958 6604 25964 6656
rect 26016 6604 26022 6656
rect 26326 6604 26332 6656
rect 26384 6604 26390 6656
rect 26694 6604 26700 6656
rect 26752 6604 26758 6656
rect 27062 6604 27068 6656
rect 27120 6604 27126 6656
rect 27154 6604 27160 6656
rect 27212 6644 27218 6656
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 27212 6616 27445 6644
rect 27212 6604 27218 6616
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 27433 6607 27491 6613
rect 27522 6604 27528 6656
rect 27580 6644 27586 6656
rect 27709 6647 27767 6653
rect 27709 6644 27721 6647
rect 27580 6616 27721 6644
rect 27580 6604 27586 6616
rect 27709 6613 27721 6616
rect 27755 6613 27767 6647
rect 27709 6607 27767 6613
rect 27982 6604 27988 6656
rect 28040 6604 28046 6656
rect 28534 6604 28540 6656
rect 28592 6604 28598 6656
rect 28644 6653 28672 6684
rect 35342 6672 35348 6724
rect 35400 6672 35406 6724
rect 35894 6672 35900 6724
rect 35952 6672 35958 6724
rect 36998 6672 37004 6724
rect 37056 6672 37062 6724
rect 37568 6721 37596 6752
rect 38657 6749 38669 6783
rect 38703 6780 38715 6783
rect 38838 6780 38844 6792
rect 38703 6752 38844 6780
rect 38703 6749 38715 6752
rect 38657 6743 38715 6749
rect 38838 6740 38844 6752
rect 38896 6740 38902 6792
rect 39022 6740 39028 6792
rect 39080 6780 39086 6792
rect 39080 6752 40080 6780
rect 39080 6740 39086 6752
rect 37553 6715 37611 6721
rect 37553 6681 37565 6715
rect 37599 6681 37611 6715
rect 37553 6675 37611 6681
rect 37734 6672 37740 6724
rect 37792 6712 37798 6724
rect 38105 6715 38163 6721
rect 38105 6712 38117 6715
rect 37792 6684 38117 6712
rect 37792 6672 37798 6684
rect 38105 6681 38117 6684
rect 38151 6681 38163 6715
rect 38105 6675 38163 6681
rect 38470 6672 38476 6724
rect 38528 6712 38534 6724
rect 38528 6684 38884 6712
rect 38528 6672 38534 6684
rect 28629 6647 28687 6653
rect 28629 6613 28641 6647
rect 28675 6613 28687 6647
rect 28629 6607 28687 6613
rect 29086 6604 29092 6656
rect 29144 6604 29150 6656
rect 29270 6604 29276 6656
rect 29328 6644 29334 6656
rect 29733 6647 29791 6653
rect 29733 6644 29745 6647
rect 29328 6616 29745 6644
rect 29328 6604 29334 6616
rect 29733 6613 29745 6616
rect 29779 6613 29791 6647
rect 29733 6607 29791 6613
rect 30006 6604 30012 6656
rect 30064 6604 30070 6656
rect 30282 6604 30288 6656
rect 30340 6604 30346 6656
rect 33226 6604 33232 6656
rect 33284 6604 33290 6656
rect 33502 6604 33508 6656
rect 33560 6604 33566 6656
rect 33778 6604 33784 6656
rect 33836 6604 33842 6656
rect 35986 6604 35992 6656
rect 36044 6644 36050 6656
rect 36541 6647 36599 6653
rect 36541 6644 36553 6647
rect 36044 6616 36553 6644
rect 36044 6604 36050 6616
rect 36541 6613 36553 6616
rect 36587 6613 36599 6647
rect 36541 6607 36599 6613
rect 36630 6604 36636 6656
rect 36688 6644 36694 6656
rect 37093 6647 37151 6653
rect 37093 6644 37105 6647
rect 36688 6616 37105 6644
rect 36688 6604 36694 6616
rect 37093 6613 37105 6616
rect 37139 6613 37151 6647
rect 37093 6607 37151 6613
rect 37642 6604 37648 6656
rect 37700 6644 37706 6656
rect 38197 6647 38255 6653
rect 38197 6644 38209 6647
rect 37700 6616 38209 6644
rect 37700 6604 37706 6616
rect 38197 6613 38209 6616
rect 38243 6613 38255 6647
rect 38197 6607 38255 6613
rect 38378 6604 38384 6656
rect 38436 6644 38442 6656
rect 38749 6647 38807 6653
rect 38749 6644 38761 6647
rect 38436 6616 38761 6644
rect 38436 6604 38442 6616
rect 38749 6613 38761 6616
rect 38795 6613 38807 6647
rect 38856 6644 38884 6684
rect 38930 6672 38936 6724
rect 38988 6712 38994 6724
rect 39209 6715 39267 6721
rect 39209 6712 39221 6715
rect 38988 6684 39221 6712
rect 38988 6672 38994 6684
rect 39209 6681 39221 6684
rect 39255 6681 39267 6715
rect 39209 6675 39267 6681
rect 39942 6672 39948 6724
rect 40000 6672 40006 6724
rect 40052 6653 40080 6752
rect 40497 6715 40555 6721
rect 40497 6681 40509 6715
rect 40543 6712 40555 6715
rect 41322 6712 41328 6724
rect 40543 6684 41328 6712
rect 40543 6681 40555 6684
rect 40497 6675 40555 6681
rect 41322 6672 41328 6684
rect 41380 6672 41386 6724
rect 39301 6647 39359 6653
rect 39301 6644 39313 6647
rect 38856 6616 39313 6644
rect 38749 6607 38807 6613
rect 39301 6613 39313 6616
rect 39347 6613 39359 6647
rect 39301 6607 39359 6613
rect 40037 6647 40095 6653
rect 40037 6613 40049 6647
rect 40083 6613 40095 6647
rect 40037 6607 40095 6613
rect 1104 6554 43675 6576
rect 1104 6502 11552 6554
rect 11604 6502 11616 6554
rect 11668 6502 11680 6554
rect 11732 6502 11744 6554
rect 11796 6502 11808 6554
rect 11860 6502 22155 6554
rect 22207 6502 22219 6554
rect 22271 6502 22283 6554
rect 22335 6502 22347 6554
rect 22399 6502 22411 6554
rect 22463 6502 32758 6554
rect 32810 6502 32822 6554
rect 32874 6502 32886 6554
rect 32938 6502 32950 6554
rect 33002 6502 33014 6554
rect 33066 6502 43361 6554
rect 43413 6502 43425 6554
rect 43477 6502 43489 6554
rect 43541 6502 43553 6554
rect 43605 6502 43617 6554
rect 43669 6502 43675 6554
rect 1104 6480 43675 6502
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5684 6412 6377 6440
rect 5684 6400 5690 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6788 6412 7021 6440
rect 6788 6400 6794 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 7009 6403 7067 6409
rect 9214 6400 9220 6452
rect 9272 6400 9278 6452
rect 9766 6400 9772 6452
rect 9824 6400 9830 6452
rect 10318 6400 10324 6452
rect 10376 6400 10382 6452
rect 10686 6400 10692 6452
rect 10744 6400 10750 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12529 6443 12587 6449
rect 12529 6440 12541 6443
rect 12308 6412 12541 6440
rect 12308 6400 12314 6412
rect 12529 6409 12541 6412
rect 12575 6409 12587 6443
rect 12529 6403 12587 6409
rect 12897 6443 12955 6449
rect 12897 6409 12909 6443
rect 12943 6409 12955 6443
rect 12897 6403 12955 6409
rect 9125 6375 9183 6381
rect 9125 6341 9137 6375
rect 9171 6372 9183 6375
rect 11974 6372 11980 6384
rect 9171 6344 11980 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 5552 6168 5580 6196
rect 5721 6171 5779 6177
rect 5721 6168 5733 6171
rect 5552 6140 5733 6168
rect 5721 6137 5733 6140
rect 5767 6137 5779 6171
rect 5721 6131 5779 6137
rect 6564 6100 6592 6267
rect 6932 6168 6960 6267
rect 9692 6236 9720 6267
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9916 6276 10241 6304
rect 9916 6264 9922 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 12912 6236 12940 6403
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13964 6412 14197 6440
rect 13964 6400 13970 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15102 6440 15108 6452
rect 14783 6412 15108 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 15473 6443 15531 6449
rect 15473 6409 15485 6443
rect 15519 6409 15531 6443
rect 15473 6403 15531 6409
rect 13998 6372 14004 6384
rect 13096 6344 14004 6372
rect 13096 6313 13124 6344
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 15378 6372 15384 6384
rect 14108 6344 15384 6372
rect 14108 6313 14136 6344
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 15488 6372 15516 6403
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15620 6412 15945 6440
rect 15620 6400 15626 6412
rect 15933 6409 15945 6412
rect 15979 6409 15991 6443
rect 15933 6403 15991 6409
rect 16022 6400 16028 6452
rect 16080 6400 16086 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 16574 6440 16580 6452
rect 16347 6412 16580 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 17126 6440 17132 6452
rect 16899 6412 17132 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17402 6440 17408 6452
rect 17236 6412 17408 6440
rect 16040 6372 16068 6400
rect 15488 6344 16068 6372
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14458 6264 14464 6316
rect 14516 6264 14522 6316
rect 14918 6264 14924 6316
rect 14976 6264 14982 6316
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 15068 6276 15148 6304
rect 15068 6264 15074 6276
rect 9692 6208 12940 6236
rect 9674 6168 9680 6180
rect 6932 6140 9680 6168
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 14476 6168 14504 6264
rect 15120 6236 15148 6276
rect 15194 6264 15200 6316
rect 15252 6264 15258 6316
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16117 6307 16175 6313
rect 16117 6304 16129 6307
rect 15804 6276 16129 6304
rect 15804 6264 15810 6276
rect 16117 6273 16129 6276
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 16264 6276 16497 6304
rect 16264 6264 16270 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17236 6304 17264 6412
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 17678 6440 17684 6452
rect 17635 6412 17684 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17920 6412 18061 6440
rect 17920 6400 17926 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 18288 6412 18429 6440
rect 18288 6400 18294 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 18506 6400 18512 6452
rect 18564 6440 18570 6452
rect 18785 6443 18843 6449
rect 18785 6440 18797 6443
rect 18564 6412 18797 6440
rect 18564 6400 18570 6412
rect 18785 6409 18797 6412
rect 18831 6409 18843 6443
rect 18785 6403 18843 6409
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19521 6443 19579 6449
rect 19521 6440 19533 6443
rect 19392 6412 19533 6440
rect 19392 6400 19398 6412
rect 19521 6409 19533 6412
rect 19567 6409 19579 6443
rect 19521 6403 19579 6409
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 21082 6440 21088 6452
rect 19668 6412 21088 6440
rect 19668 6400 19674 6412
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 23106 6440 23112 6452
rect 22066 6412 23112 6440
rect 17328 6344 19656 6372
rect 17328 6313 17356 6344
rect 17083 6276 17264 6304
rect 17313 6307 17371 6313
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17313 6273 17325 6307
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 17770 6264 17776 6316
rect 17828 6264 17834 6316
rect 18230 6264 18236 6316
rect 18288 6264 18294 6316
rect 18598 6264 18604 6316
rect 18656 6264 18662 6316
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6304 19027 6307
rect 19015 6276 19288 6304
rect 19015 6273 19027 6276
rect 18969 6267 19027 6273
rect 16758 6236 16764 6248
rect 15120 6208 16764 6236
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17218 6196 17224 6248
rect 17276 6196 17282 6248
rect 15013 6171 15071 6177
rect 15013 6168 15025 6171
rect 14476 6140 15025 6168
rect 15013 6137 15025 6140
rect 15059 6137 15071 6171
rect 15013 6131 15071 6137
rect 17129 6171 17187 6177
rect 17129 6137 17141 6171
rect 17175 6168 17187 6171
rect 17236 6168 17264 6196
rect 17175 6140 17264 6168
rect 19260 6168 19288 6276
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 19628 6236 19656 6344
rect 19794 6332 19800 6384
rect 19852 6372 19858 6384
rect 22066 6372 22094 6412
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 24670 6400 24676 6452
rect 24728 6400 24734 6452
rect 25222 6400 25228 6452
rect 25280 6400 25286 6452
rect 25590 6400 25596 6452
rect 25648 6440 25654 6452
rect 29086 6440 29092 6452
rect 25648 6412 29092 6440
rect 25648 6400 25654 6412
rect 29086 6400 29092 6412
rect 29144 6400 29150 6452
rect 31754 6400 31760 6452
rect 31812 6440 31818 6452
rect 36722 6440 36728 6452
rect 31812 6412 36728 6440
rect 31812 6400 31818 6412
rect 36722 6400 36728 6412
rect 36780 6400 36786 6452
rect 36998 6400 37004 6452
rect 37056 6400 37062 6452
rect 37918 6400 37924 6452
rect 37976 6440 37982 6452
rect 39114 6440 39120 6452
rect 37976 6412 39120 6440
rect 37976 6400 37982 6412
rect 39114 6400 39120 6412
rect 39172 6400 39178 6452
rect 24688 6372 24716 6400
rect 19852 6344 22094 6372
rect 23124 6344 23796 6372
rect 19852 6332 19858 6344
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 23124 6304 23152 6344
rect 23768 6316 23796 6344
rect 23860 6344 24716 6372
rect 19751 6276 23152 6304
rect 23201 6308 23259 6313
rect 23201 6307 23336 6308
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 23201 6273 23213 6307
rect 23247 6304 23336 6307
rect 23658 6304 23664 6316
rect 23247 6280 23664 6304
rect 23247 6273 23259 6280
rect 23308 6276 23664 6280
rect 23201 6267 23259 6273
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 23750 6264 23756 6316
rect 23808 6264 23814 6316
rect 23860 6313 23888 6344
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6273 23903 6307
rect 23845 6267 23903 6273
rect 24213 6307 24271 6313
rect 24213 6273 24225 6307
rect 24259 6304 24271 6307
rect 25240 6304 25268 6400
rect 30374 6332 30380 6384
rect 30432 6372 30438 6384
rect 37016 6372 37044 6400
rect 30432 6344 37044 6372
rect 30432 6332 30438 6344
rect 38286 6332 38292 6384
rect 38344 6372 38350 6384
rect 38654 6372 38660 6384
rect 38344 6344 38660 6372
rect 38344 6332 38350 6344
rect 38654 6332 38660 6344
rect 38712 6332 38718 6384
rect 24259 6276 25268 6304
rect 24259 6273 24271 6276
rect 24213 6267 24271 6273
rect 19628 6208 31754 6236
rect 22002 6168 22008 6180
rect 19260 6140 22008 6168
rect 17175 6137 17187 6140
rect 17129 6131 17187 6137
rect 22002 6128 22008 6140
rect 22060 6128 22066 6180
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 23072 6140 23980 6168
rect 23072 6128 23078 6140
rect 14366 6100 14372 6112
rect 6564 6072 14372 6100
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 19153 6103 19211 6109
rect 19153 6069 19165 6103
rect 19199 6100 19211 6103
rect 19886 6100 19892 6112
rect 19199 6072 19892 6100
rect 19199 6069 19211 6072
rect 19153 6063 19211 6069
rect 19886 6060 19892 6072
rect 19944 6060 19950 6112
rect 23382 6060 23388 6112
rect 23440 6060 23446 6112
rect 23952 6100 23980 6140
rect 24026 6128 24032 6180
rect 24084 6128 24090 6180
rect 24302 6128 24308 6180
rect 24360 6168 24366 6180
rect 24397 6171 24455 6177
rect 24397 6168 24409 6171
rect 24360 6140 24409 6168
rect 24360 6128 24366 6140
rect 24397 6137 24409 6140
rect 24443 6137 24455 6171
rect 24397 6131 24455 6137
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 28534 6168 28540 6180
rect 24820 6140 28540 6168
rect 24820 6128 24826 6140
rect 28534 6128 28540 6140
rect 28592 6128 28598 6180
rect 31726 6168 31754 6208
rect 32306 6168 32312 6180
rect 31726 6140 32312 6168
rect 32306 6128 32312 6140
rect 32364 6128 32370 6180
rect 25958 6100 25964 6112
rect 23952 6072 25964 6100
rect 25958 6060 25964 6072
rect 26016 6060 26022 6112
rect 1104 6010 43516 6032
rect 1104 5958 6251 6010
rect 6303 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 16854 6010
rect 16906 5958 16918 6010
rect 16970 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 27457 6010
rect 27509 5958 27521 6010
rect 27573 5958 27585 6010
rect 27637 5958 27649 6010
rect 27701 5958 27713 6010
rect 27765 5958 38060 6010
rect 38112 5958 38124 6010
rect 38176 5958 38188 6010
rect 38240 5958 38252 6010
rect 38304 5958 38316 6010
rect 38368 5958 43516 6010
rect 1104 5936 43516 5958
rect 5902 5856 5908 5908
rect 5960 5856 5966 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9769 5899 9827 5905
rect 9769 5896 9781 5899
rect 9548 5868 9781 5896
rect 9548 5856 9554 5868
rect 9769 5865 9781 5868
rect 9815 5865 9827 5899
rect 9769 5859 9827 5865
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 17218 5896 17224 5908
rect 12768 5868 17224 5896
rect 12768 5856 12774 5868
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 20254 5896 20260 5908
rect 17328 5868 20260 5896
rect 5920 5828 5948 5856
rect 17328 5828 17356 5868
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 27154 5896 27160 5908
rect 20772 5868 27160 5896
rect 20772 5856 20778 5868
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 5920 5800 17356 5828
rect 23198 5788 23204 5840
rect 23256 5828 23262 5840
rect 30282 5828 30288 5840
rect 23256 5800 30288 5828
rect 23256 5788 23262 5800
rect 30282 5788 30288 5800
rect 30340 5788 30346 5840
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4580 5732 16528 5760
rect 4580 5720 4586 5732
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 11054 5692 11060 5704
rect 9723 5664 11060 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 15102 5692 15108 5704
rect 11940 5664 15108 5692
rect 11940 5652 11946 5664
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 7852 5624 7880 5652
rect 13722 5624 13728 5636
rect 7852 5596 13728 5624
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 16500 5624 16528 5732
rect 18598 5720 18604 5772
rect 18656 5760 18662 5772
rect 22738 5760 22744 5772
rect 18656 5732 22744 5760
rect 18656 5720 18662 5732
rect 22738 5720 22744 5732
rect 22796 5720 22802 5772
rect 23290 5720 23296 5772
rect 23348 5760 23354 5772
rect 25498 5760 25504 5772
rect 23348 5732 25504 5760
rect 23348 5720 23354 5732
rect 25498 5720 25504 5732
rect 25556 5720 25562 5772
rect 20530 5624 20536 5636
rect 16500 5596 20536 5624
rect 20530 5584 20536 5596
rect 20588 5584 20594 5636
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 24578 5556 24584 5568
rect 19392 5528 24584 5556
rect 19392 5516 19398 5528
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 1104 5466 43675 5488
rect 1104 5414 11552 5466
rect 11604 5414 11616 5466
rect 11668 5414 11680 5466
rect 11732 5414 11744 5466
rect 11796 5414 11808 5466
rect 11860 5414 22155 5466
rect 22207 5414 22219 5466
rect 22271 5414 22283 5466
rect 22335 5414 22347 5466
rect 22399 5414 22411 5466
rect 22463 5414 32758 5466
rect 32810 5414 32822 5466
rect 32874 5414 32886 5466
rect 32938 5414 32950 5466
rect 33002 5414 33014 5466
rect 33066 5414 43361 5466
rect 43413 5414 43425 5466
rect 43477 5414 43489 5466
rect 43541 5414 43553 5466
rect 43605 5414 43617 5466
rect 43669 5414 43675 5466
rect 1104 5392 43675 5414
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 26326 5352 26332 5364
rect 16816 5324 26332 5352
rect 16816 5312 16822 5324
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 15378 5244 15384 5296
rect 15436 5284 15442 5296
rect 23290 5284 23296 5296
rect 15436 5256 23296 5284
rect 15436 5244 15442 5256
rect 23290 5244 23296 5256
rect 23348 5244 23354 5296
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 26694 5216 26700 5228
rect 17276 5188 26700 5216
rect 17276 5176 17282 5188
rect 26694 5176 26700 5188
rect 26752 5176 26758 5228
rect 15102 5108 15108 5160
rect 15160 5148 15166 5160
rect 27982 5148 27988 5160
rect 15160 5120 27988 5148
rect 15160 5108 15166 5120
rect 27982 5108 27988 5120
rect 28040 5108 28046 5160
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 25590 5080 25596 5092
rect 12676 5052 25596 5080
rect 12676 5040 12682 5052
rect 25590 5040 25596 5052
rect 25648 5040 25654 5092
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 30006 5012 30012 5024
rect 10836 4984 30012 5012
rect 10836 4972 10842 4984
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 1104 4922 43516 4944
rect 1104 4870 6251 4922
rect 6303 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 16854 4922
rect 16906 4870 16918 4922
rect 16970 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 27457 4922
rect 27509 4870 27521 4922
rect 27573 4870 27585 4922
rect 27637 4870 27649 4922
rect 27701 4870 27713 4922
rect 27765 4870 38060 4922
rect 38112 4870 38124 4922
rect 38176 4870 38188 4922
rect 38240 4870 38252 4922
rect 38304 4870 38316 4922
rect 38368 4870 43516 4922
rect 1104 4848 43516 4870
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 27338 4808 27344 4820
rect 12492 4780 27344 4808
rect 12492 4768 12498 4780
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 19794 4740 19800 4752
rect 6880 4712 19800 4740
rect 6880 4700 6886 4712
rect 19794 4700 19800 4712
rect 19852 4700 19858 4752
rect 1104 4378 43675 4400
rect 1104 4326 11552 4378
rect 11604 4326 11616 4378
rect 11668 4326 11680 4378
rect 11732 4326 11744 4378
rect 11796 4326 11808 4378
rect 11860 4326 22155 4378
rect 22207 4326 22219 4378
rect 22271 4326 22283 4378
rect 22335 4326 22347 4378
rect 22399 4326 22411 4378
rect 22463 4326 32758 4378
rect 32810 4326 32822 4378
rect 32874 4326 32886 4378
rect 32938 4326 32950 4378
rect 33002 4326 33014 4378
rect 33066 4326 43361 4378
rect 43413 4326 43425 4378
rect 43477 4326 43489 4378
rect 43541 4326 43553 4378
rect 43605 4326 43617 4378
rect 43669 4326 43675 4378
rect 1104 4304 43675 4326
rect 30834 3884 30840 3936
rect 30892 3924 30898 3936
rect 35894 3924 35900 3936
rect 30892 3896 35900 3924
rect 30892 3884 30898 3896
rect 35894 3884 35900 3896
rect 35952 3884 35958 3936
rect 1104 3834 43516 3856
rect 1104 3782 6251 3834
rect 6303 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 16854 3834
rect 16906 3782 16918 3834
rect 16970 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 27457 3834
rect 27509 3782 27521 3834
rect 27573 3782 27585 3834
rect 27637 3782 27649 3834
rect 27701 3782 27713 3834
rect 27765 3782 38060 3834
rect 38112 3782 38124 3834
rect 38176 3782 38188 3834
rect 38240 3782 38252 3834
rect 38304 3782 38316 3834
rect 38368 3782 43516 3834
rect 1104 3760 43516 3782
rect 33965 3723 34023 3729
rect 33965 3689 33977 3723
rect 34011 3720 34023 3723
rect 34422 3720 34428 3732
rect 34011 3692 34428 3720
rect 34011 3689 34023 3692
rect 33965 3683 34023 3689
rect 34422 3680 34428 3692
rect 34480 3680 34486 3732
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 34149 3519 34207 3525
rect 34149 3516 34161 3519
rect 5684 3488 34161 3516
rect 5684 3476 5690 3488
rect 34149 3485 34161 3488
rect 34195 3485 34207 3519
rect 34149 3479 34207 3485
rect 1104 3290 43675 3312
rect 1104 3238 11552 3290
rect 11604 3238 11616 3290
rect 11668 3238 11680 3290
rect 11732 3238 11744 3290
rect 11796 3238 11808 3290
rect 11860 3238 22155 3290
rect 22207 3238 22219 3290
rect 22271 3238 22283 3290
rect 22335 3238 22347 3290
rect 22399 3238 22411 3290
rect 22463 3238 32758 3290
rect 32810 3238 32822 3290
rect 32874 3238 32886 3290
rect 32938 3238 32950 3290
rect 33002 3238 33014 3290
rect 33066 3238 43361 3290
rect 43413 3238 43425 3290
rect 43477 3238 43489 3290
rect 43541 3238 43553 3290
rect 43605 3238 43617 3290
rect 43669 3238 43675 3290
rect 1104 3216 43675 3238
rect 16853 3179 16911 3185
rect 16853 3145 16865 3179
rect 16899 3176 16911 3179
rect 24946 3176 24952 3188
rect 16899 3148 24952 3176
rect 16899 3145 16911 3148
rect 16853 3139 16911 3145
rect 24946 3136 24952 3148
rect 25004 3136 25010 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 33321 3179 33379 3185
rect 25280 3148 31754 3176
rect 25280 3136 25286 3148
rect 31726 3108 31754 3148
rect 33321 3145 33333 3179
rect 33367 3176 33379 3179
rect 37829 3179 37887 3185
rect 33367 3148 37228 3176
rect 33367 3145 33379 3148
rect 33321 3139 33379 3145
rect 37200 3108 37228 3148
rect 37829 3145 37841 3179
rect 37875 3176 37887 3179
rect 38562 3176 38568 3188
rect 37875 3148 38568 3176
rect 37875 3145 37887 3148
rect 37829 3139 37887 3145
rect 38562 3136 38568 3148
rect 38620 3136 38626 3188
rect 38838 3136 38844 3188
rect 38896 3136 38902 3188
rect 38856 3108 38884 3136
rect 31726 3080 35894 3108
rect 37200 3080 38884 3108
rect 16666 3000 16672 3052
rect 16724 3000 16730 3052
rect 18598 3000 18604 3052
rect 18656 3000 18662 3052
rect 20714 3000 20720 3052
rect 20772 3000 20778 3052
rect 22646 3000 22652 3052
rect 22704 3000 22710 3052
rect 24854 3040 24860 3052
rect 22756 3012 24860 3040
rect 22756 2972 22784 3012
rect 24854 3000 24860 3012
rect 24912 3000 24918 3052
rect 24946 3000 24952 3052
rect 25004 3000 25010 3052
rect 31754 3040 31760 3052
rect 25148 3012 31760 3040
rect 19306 2944 22784 2972
rect 18785 2839 18843 2845
rect 18785 2805 18797 2839
rect 18831 2836 18843 2839
rect 19306 2836 19334 2944
rect 22833 2907 22891 2913
rect 22833 2873 22845 2907
rect 22879 2904 22891 2907
rect 25038 2904 25044 2916
rect 22879 2876 25044 2904
rect 22879 2873 22891 2876
rect 22833 2867 22891 2873
rect 25038 2864 25044 2876
rect 25096 2864 25102 2916
rect 25148 2913 25176 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 33502 3000 33508 3052
rect 33560 3000 33566 3052
rect 35866 3040 35894 3080
rect 37274 3040 37280 3052
rect 35866 3012 37280 3040
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 37826 3000 37832 3052
rect 37884 3040 37890 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37884 3012 38025 3040
rect 37884 3000 37890 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 25314 2932 25320 2984
rect 25372 2972 25378 2984
rect 37918 2972 37924 2984
rect 25372 2944 37924 2972
rect 25372 2932 25378 2944
rect 37918 2932 37924 2944
rect 37976 2932 37982 2984
rect 25133 2907 25191 2913
rect 25133 2873 25145 2907
rect 25179 2873 25191 2907
rect 25133 2867 25191 2873
rect 25222 2864 25228 2916
rect 25280 2904 25286 2916
rect 33686 2904 33692 2916
rect 25280 2876 33692 2904
rect 25280 2864 25286 2876
rect 33686 2864 33692 2876
rect 33744 2864 33750 2916
rect 18831 2808 19334 2836
rect 20901 2839 20959 2845
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 20901 2805 20913 2839
rect 20947 2836 20959 2839
rect 30374 2836 30380 2848
rect 20947 2808 30380 2836
rect 20947 2805 20959 2808
rect 20901 2799 20959 2805
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 1104 2746 43516 2768
rect 1104 2694 6251 2746
rect 6303 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 16854 2746
rect 16906 2694 16918 2746
rect 16970 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 27457 2746
rect 27509 2694 27521 2746
rect 27573 2694 27585 2746
rect 27637 2694 27649 2746
rect 27701 2694 27713 2746
rect 27765 2694 38060 2746
rect 38112 2694 38124 2746
rect 38176 2694 38188 2746
rect 38240 2694 38252 2746
rect 38304 2694 38316 2746
rect 38368 2694 43516 2746
rect 1104 2672 43516 2694
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 16025 2635 16083 2641
rect 16025 2601 16037 2635
rect 16071 2632 16083 2635
rect 16666 2632 16672 2644
rect 16071 2604 16672 2632
rect 16071 2601 16083 2604
rect 16025 2595 16083 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 18598 2632 18604 2644
rect 18187 2604 18604 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 20257 2635 20315 2641
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20714 2632 20720 2644
rect 20303 2604 20720 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22373 2635 22431 2641
rect 22373 2601 22385 2635
rect 22419 2632 22431 2635
rect 22646 2632 22652 2644
rect 22419 2604 22652 2632
rect 22419 2601 22431 2604
rect 22373 2595 22431 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 24489 2635 24547 2641
rect 24489 2601 24501 2635
rect 24535 2632 24547 2635
rect 24946 2632 24952 2644
rect 24535 2604 24952 2632
rect 24535 2601 24547 2604
rect 24489 2595 24547 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 33226 2632 33232 2644
rect 33152 2604 33232 2632
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 30834 2564 30840 2576
rect 14783 2536 30840 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 30834 2524 30840 2536
rect 30892 2524 30898 2576
rect 33152 2573 33180 2604
rect 33226 2592 33232 2604
rect 33284 2592 33290 2644
rect 33413 2635 33471 2641
rect 33413 2601 33425 2635
rect 33459 2632 33471 2635
rect 33502 2632 33508 2644
rect 33459 2604 33508 2632
rect 33459 2601 33471 2604
rect 33413 2595 33471 2601
rect 33502 2592 33508 2604
rect 33560 2592 33566 2644
rect 33781 2635 33839 2641
rect 33781 2601 33793 2635
rect 33827 2632 33839 2635
rect 34146 2632 34152 2644
rect 33827 2604 34152 2632
rect 33827 2601 33839 2604
rect 33781 2595 33839 2601
rect 34146 2592 34152 2604
rect 34204 2592 34210 2644
rect 34701 2635 34759 2641
rect 34701 2601 34713 2635
rect 34747 2632 34759 2635
rect 35342 2632 35348 2644
rect 34747 2604 35348 2632
rect 34747 2601 34759 2604
rect 34701 2595 34759 2601
rect 35342 2592 35348 2604
rect 35400 2592 35406 2644
rect 37277 2635 37335 2641
rect 37277 2601 37289 2635
rect 37323 2632 37335 2635
rect 37734 2632 37740 2644
rect 37323 2604 37740 2632
rect 37323 2601 37335 2604
rect 37277 2595 37335 2601
rect 37734 2592 37740 2604
rect 37792 2592 37798 2644
rect 37826 2592 37832 2644
rect 37884 2592 37890 2644
rect 38746 2592 38752 2644
rect 38804 2592 38810 2644
rect 39025 2635 39083 2641
rect 39025 2601 39037 2635
rect 39071 2632 39083 2635
rect 39942 2632 39948 2644
rect 39071 2604 39948 2632
rect 39071 2601 39083 2604
rect 39025 2595 39083 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 40129 2635 40187 2641
rect 40129 2601 40141 2635
rect 40175 2632 40187 2635
rect 40494 2632 40500 2644
rect 40175 2604 40500 2632
rect 40175 2601 40187 2604
rect 40129 2595 40187 2601
rect 40494 2592 40500 2604
rect 40552 2592 40558 2644
rect 41322 2592 41328 2644
rect 41380 2632 41386 2644
rect 42429 2635 42487 2641
rect 42429 2632 42441 2635
rect 41380 2604 42441 2632
rect 41380 2592 41386 2604
rect 42429 2601 42441 2604
rect 42475 2601 42487 2635
rect 42429 2595 42487 2601
rect 33137 2567 33195 2573
rect 30944 2536 31156 2564
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 12483 2468 28856 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 1118 2388 1124 2440
rect 1176 2428 1182 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1176 2400 1409 2428
rect 1176 2388 1182 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 9674 2388 9680 2440
rect 9732 2388 9738 2440
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13872 2400 14289 2428
rect 13872 2388 13878 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 18322 2388 18328 2440
rect 18380 2388 18386 2440
rect 20438 2388 20444 2440
rect 20496 2388 20502 2440
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 26602 2388 26608 2440
rect 26660 2388 26666 2440
rect 28718 2388 28724 2440
rect 28776 2388 28782 2440
rect 12253 2363 12311 2369
rect 12253 2329 12265 2363
rect 12299 2329 12311 2363
rect 12253 2323 12311 2329
rect 14553 2363 14611 2369
rect 14553 2329 14565 2363
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 9858 2252 9864 2304
rect 9916 2252 9922 2304
rect 11793 2295 11851 2301
rect 11793 2261 11805 2295
rect 11839 2292 11851 2295
rect 12268 2292 12296 2323
rect 11839 2264 12296 2292
rect 14093 2295 14151 2301
rect 11839 2261 11851 2264
rect 11793 2255 11851 2261
rect 14093 2261 14105 2295
rect 14139 2292 14151 2295
rect 14568 2292 14596 2323
rect 28828 2304 28856 2468
rect 29822 2456 29828 2508
rect 29880 2496 29886 2508
rect 30944 2496 30972 2536
rect 29880 2468 30972 2496
rect 31128 2496 31156 2536
rect 33137 2533 33149 2567
rect 33183 2533 33195 2567
rect 34241 2567 34299 2573
rect 33137 2527 33195 2533
rect 33244 2536 33456 2564
rect 33244 2496 33272 2536
rect 31128 2468 33272 2496
rect 33428 2496 33456 2536
rect 34241 2533 34253 2567
rect 34287 2564 34299 2567
rect 34790 2564 34796 2576
rect 34287 2536 34796 2564
rect 34287 2533 34299 2536
rect 34241 2527 34299 2533
rect 34790 2524 34796 2536
rect 34848 2524 34854 2576
rect 37553 2567 37611 2573
rect 37553 2533 37565 2567
rect 37599 2564 37611 2567
rect 38764 2564 38792 2592
rect 37599 2536 38792 2564
rect 42981 2567 43039 2573
rect 37599 2533 37611 2536
rect 37553 2527 37611 2533
rect 42981 2533 42993 2567
rect 43027 2533 43039 2567
rect 42981 2527 43039 2533
rect 33428 2468 34928 2496
rect 29880 2456 29886 2468
rect 31018 2388 31024 2440
rect 31076 2388 31082 2440
rect 33318 2388 33324 2440
rect 33376 2388 33382 2440
rect 33594 2388 33600 2440
rect 33652 2388 33658 2440
rect 33962 2388 33968 2440
rect 34020 2388 34026 2440
rect 34422 2388 34428 2440
rect 34480 2388 34486 2440
rect 34900 2437 34928 2468
rect 37182 2456 37188 2508
rect 37240 2496 37246 2508
rect 37240 2468 38056 2496
rect 37240 2456 37246 2468
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35250 2388 35256 2440
rect 35308 2388 35314 2440
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 35728 2360 35756 2391
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 38028 2437 38056 2468
rect 37737 2431 37795 2437
rect 37737 2397 37749 2431
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38013 2431 38071 2437
rect 38013 2397 38025 2431
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2428 39267 2431
rect 39255 2400 39344 2428
rect 39255 2397 39267 2400
rect 39209 2391 39267 2397
rect 28920 2332 33180 2360
rect 14139 2264 14596 2292
rect 14139 2261 14151 2264
rect 14093 2255 14151 2261
rect 26786 2252 26792 2304
rect 26844 2252 26850 2304
rect 28810 2252 28816 2304
rect 28868 2252 28874 2304
rect 28920 2301 28948 2332
rect 28905 2295 28963 2301
rect 28905 2261 28917 2295
rect 28951 2261 28963 2295
rect 28905 2255 28963 2261
rect 30837 2295 30895 2301
rect 30837 2261 30849 2295
rect 30883 2292 30895 2295
rect 32674 2292 32680 2304
rect 30883 2264 32680 2292
rect 30883 2261 30895 2264
rect 30837 2255 30895 2261
rect 32674 2252 32680 2264
rect 32732 2252 32738 2304
rect 33152 2292 33180 2332
rect 35084 2332 35756 2360
rect 33410 2292 33416 2304
rect 33152 2264 33416 2292
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 35084 2301 35112 2332
rect 36814 2320 36820 2372
rect 36872 2360 36878 2372
rect 37752 2360 37780 2391
rect 36872 2332 37780 2360
rect 36872 2320 36878 2332
rect 38930 2320 38936 2372
rect 38988 2320 38994 2372
rect 35069 2295 35127 2301
rect 35069 2261 35081 2295
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 35529 2295 35587 2301
rect 35529 2261 35541 2295
rect 35575 2292 35587 2295
rect 38948 2292 38976 2320
rect 39316 2301 39344 2400
rect 39482 2388 39488 2440
rect 39540 2388 39546 2440
rect 40313 2431 40371 2437
rect 40313 2397 40325 2431
rect 40359 2428 40371 2431
rect 40359 2400 41460 2428
rect 40359 2397 40371 2400
rect 40313 2391 40371 2397
rect 41432 2301 41460 2400
rect 41598 2388 41604 2440
rect 41656 2388 41662 2440
rect 42613 2431 42671 2437
rect 42613 2397 42625 2431
rect 42659 2428 42671 2431
rect 42996 2428 43024 2527
rect 42659 2400 43024 2428
rect 42659 2397 42671 2400
rect 42613 2391 42671 2397
rect 43162 2388 43168 2440
rect 43220 2388 43226 2440
rect 35575 2264 38976 2292
rect 39301 2295 39359 2301
rect 35575 2261 35587 2264
rect 35529 2255 35587 2261
rect 39301 2261 39313 2295
rect 39347 2261 39359 2295
rect 39301 2255 39359 2261
rect 41417 2295 41475 2301
rect 41417 2261 41429 2295
rect 41463 2261 41475 2295
rect 41417 2255 41475 2261
rect 1104 2202 43675 2224
rect 1104 2150 11552 2202
rect 11604 2150 11616 2202
rect 11668 2150 11680 2202
rect 11732 2150 11744 2202
rect 11796 2150 11808 2202
rect 11860 2150 22155 2202
rect 22207 2150 22219 2202
rect 22271 2150 22283 2202
rect 22335 2150 22347 2202
rect 22399 2150 22411 2202
rect 22463 2150 32758 2202
rect 32810 2150 32822 2202
rect 32874 2150 32886 2202
rect 32938 2150 32950 2202
rect 33002 2150 33014 2202
rect 33066 2150 43361 2202
rect 43413 2150 43425 2202
rect 43477 2150 43489 2202
rect 43541 2150 43553 2202
rect 43605 2150 43617 2202
rect 43669 2150 43675 2202
rect 1104 2128 43675 2150
rect 1670 2048 1676 2100
rect 1728 2048 1734 2100
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 4120 2060 6914 2088
rect 4120 2048 4126 2060
rect 1688 1748 1716 2048
rect 6886 1816 6914 2060
rect 7742 2048 7748 2100
rect 7800 2048 7806 2100
rect 9858 2048 9864 2100
rect 9916 2088 9922 2100
rect 29822 2088 29828 2100
rect 9916 2060 29828 2088
rect 9916 2048 9922 2060
rect 29822 2048 29828 2060
rect 29880 2048 29886 2100
rect 34422 2088 34428 2100
rect 30116 2060 34428 2088
rect 7760 1884 7788 2048
rect 30116 1952 30144 2060
rect 34422 2048 34428 2060
rect 34480 2048 34486 2100
rect 34514 2048 34520 2100
rect 34572 2088 34578 2100
rect 36078 2088 36084 2100
rect 34572 2060 36084 2088
rect 34572 2048 34578 2060
rect 36078 2048 36084 2060
rect 36136 2048 36142 2100
rect 36814 2048 36820 2100
rect 36872 2048 36878 2100
rect 37458 2048 37464 2100
rect 37516 2048 37522 2100
rect 32674 1980 32680 2032
rect 32732 2020 32738 2032
rect 36832 2020 36860 2048
rect 32732 1992 36860 2020
rect 32732 1980 32738 1992
rect 26206 1924 30144 1952
rect 26206 1884 26234 1924
rect 33410 1912 33416 1964
rect 33468 1952 33474 1964
rect 37476 1952 37504 2048
rect 33468 1924 37504 1952
rect 33468 1912 33474 1924
rect 33962 1884 33968 1896
rect 7760 1856 26234 1884
rect 30116 1856 33968 1884
rect 30116 1816 30144 1856
rect 33962 1844 33968 1856
rect 34020 1844 34026 1896
rect 6886 1788 30144 1816
rect 33318 1776 33324 1828
rect 33376 1776 33382 1828
rect 33336 1748 33364 1776
rect 1688 1720 33364 1748
rect 26786 1640 26792 1692
rect 26844 1680 26850 1692
rect 36906 1680 36912 1692
rect 26844 1652 36912 1680
rect 26844 1640 26850 1652
rect 36906 1640 36912 1652
rect 36964 1640 36970 1692
rect 28810 1572 28816 1624
rect 28868 1612 28874 1624
rect 34514 1612 34520 1624
rect 28868 1584 34520 1612
rect 28868 1572 28874 1584
rect 34514 1572 34520 1584
rect 34572 1572 34578 1624
rect 32858 1368 32864 1420
rect 32916 1408 32922 1420
rect 33594 1408 33600 1420
rect 32916 1380 33600 1408
rect 32916 1368 32922 1380
rect 33594 1368 33600 1380
rect 33652 1368 33658 1420
<< via1 >>
rect 16212 8508 16264 8560
rect 33324 8508 33376 8560
rect 15752 8440 15804 8492
rect 33600 8440 33652 8492
rect 15660 8372 15712 8424
rect 33692 8372 33744 8424
rect 10508 8304 10560 8356
rect 29276 8304 29328 8356
rect 24952 8236 25004 8288
rect 25964 8236 26016 8288
rect 30196 8236 30248 8288
rect 30656 8236 30708 8288
rect 7196 8168 7248 8220
rect 22836 8168 22888 8220
rect 25228 8168 25280 8220
rect 26056 8168 26108 8220
rect 11336 7964 11388 8016
rect 15200 8100 15252 8152
rect 24492 8100 24544 8152
rect 27620 8100 27672 8152
rect 28540 8100 28592 8152
rect 12624 8032 12676 8084
rect 20720 8032 20772 8084
rect 24584 8032 24636 8084
rect 14372 7964 14424 8016
rect 25688 7964 25740 8016
rect 27712 7964 27764 8016
rect 28632 7964 28684 8016
rect 30564 7964 30616 8016
rect 15108 7896 15160 7948
rect 22008 7896 22060 7948
rect 14004 7828 14056 7880
rect 20996 7828 21048 7880
rect 23756 7828 23808 7880
rect 30104 7828 30156 7880
rect 31116 7828 31168 7880
rect 31392 7828 31444 7880
rect 12900 7760 12952 7812
rect 21272 7760 21324 7812
rect 7748 7692 7800 7744
rect 8300 7692 8352 7744
rect 16304 7692 16356 7744
rect 16856 7692 16908 7744
rect 32404 7760 32456 7812
rect 22928 7692 22980 7744
rect 30840 7692 30892 7744
rect 11552 7590 11604 7642
rect 11616 7590 11668 7642
rect 11680 7590 11732 7642
rect 11744 7590 11796 7642
rect 11808 7590 11860 7642
rect 22155 7590 22207 7642
rect 22219 7590 22271 7642
rect 22283 7590 22335 7642
rect 22347 7590 22399 7642
rect 22411 7590 22463 7642
rect 32758 7590 32810 7642
rect 32822 7590 32874 7642
rect 32886 7590 32938 7642
rect 32950 7590 33002 7642
rect 33014 7590 33066 7642
rect 43361 7590 43413 7642
rect 43425 7590 43477 7642
rect 43489 7590 43541 7642
rect 43553 7590 43605 7642
rect 43617 7590 43669 7642
rect 5356 7488 5408 7540
rect 5908 7488 5960 7540
rect 7288 7488 7340 7540
rect 7840 7488 7892 7540
rect 8392 7488 8444 7540
rect 8944 7488 8996 7540
rect 10508 7488 10560 7540
rect 11152 7488 11204 7540
rect 12532 7488 12584 7540
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13636 7488 13688 7540
rect 14188 7488 14240 7540
rect 15016 7488 15068 7540
rect 15568 7488 15620 7540
rect 16028 7488 16080 7540
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5540 7352 5592 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6460 7284 6512 7336
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 6828 7352 6880 7404
rect 7748 7352 7800 7404
rect 8300 7352 8352 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 12900 7420 12952 7472
rect 11336 7352 11388 7404
rect 12072 7352 12124 7404
rect 12624 7352 12676 7404
rect 11888 7284 11940 7336
rect 9864 7216 9916 7268
rect 12900 7284 12952 7336
rect 11060 7148 11112 7200
rect 15936 7420 15988 7472
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 19156 7488 19208 7540
rect 18880 7420 18932 7472
rect 20536 7488 20588 7540
rect 22836 7488 22888 7540
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16672 7352 16724 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17224 7352 17276 7404
rect 17868 7352 17920 7404
rect 18512 7352 18564 7404
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22560 7420 22612 7472
rect 22652 7352 22704 7404
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 23020 7352 23072 7404
rect 23572 7395 23624 7404
rect 23572 7361 23581 7395
rect 23581 7361 23615 7395
rect 23615 7361 23624 7395
rect 23572 7352 23624 7361
rect 23664 7352 23716 7404
rect 24492 7488 24544 7540
rect 24676 7488 24728 7540
rect 24400 7420 24452 7472
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24308 7352 24360 7404
rect 25688 7531 25740 7540
rect 25688 7497 25697 7531
rect 25697 7497 25731 7531
rect 25731 7497 25740 7531
rect 25688 7488 25740 7497
rect 26240 7488 26292 7540
rect 26148 7420 26200 7472
rect 16304 7216 16356 7268
rect 25596 7352 25648 7404
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 26056 7352 26108 7404
rect 27436 7488 27488 7540
rect 27252 7420 27304 7472
rect 28724 7488 28776 7540
rect 28356 7420 28408 7472
rect 16488 7148 16540 7200
rect 16580 7148 16632 7200
rect 22744 7216 22796 7268
rect 23296 7216 23348 7268
rect 26700 7284 26752 7336
rect 20996 7148 21048 7200
rect 21180 7148 21232 7200
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 23848 7148 23900 7200
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 26424 7216 26476 7268
rect 27436 7216 27488 7268
rect 28540 7395 28592 7404
rect 28540 7361 28549 7395
rect 28549 7361 28583 7395
rect 28583 7361 28592 7395
rect 28540 7352 28592 7361
rect 28632 7352 28684 7404
rect 30472 7488 30524 7540
rect 29460 7420 29512 7472
rect 30288 7420 30340 7472
rect 29000 7284 29052 7336
rect 29092 7216 29144 7268
rect 30196 7352 30248 7404
rect 30656 7395 30708 7404
rect 30656 7361 30665 7395
rect 30665 7361 30699 7395
rect 30699 7361 30708 7395
rect 30656 7352 30708 7361
rect 31392 7531 31444 7540
rect 31392 7497 31401 7531
rect 31401 7497 31435 7531
rect 31435 7497 31444 7531
rect 31392 7488 31444 7497
rect 31668 7488 31720 7540
rect 31300 7420 31352 7472
rect 30748 7284 30800 7336
rect 31852 7352 31904 7404
rect 32772 7488 32824 7540
rect 32496 7420 32548 7472
rect 33692 7531 33744 7540
rect 33692 7497 33701 7531
rect 33701 7497 33735 7531
rect 33735 7497 33744 7531
rect 33692 7488 33744 7497
rect 33784 7488 33836 7540
rect 34336 7488 34388 7540
rect 34612 7420 34664 7472
rect 35624 7488 35676 7540
rect 37004 7420 37056 7472
rect 39488 7488 39540 7540
rect 38936 7420 38988 7472
rect 31944 7284 31996 7336
rect 32864 7284 32916 7336
rect 33324 7284 33376 7336
rect 33416 7284 33468 7336
rect 34152 7352 34204 7404
rect 34428 7284 34480 7336
rect 30104 7216 30156 7268
rect 25228 7191 25280 7200
rect 25228 7157 25237 7191
rect 25237 7157 25271 7191
rect 25271 7157 25280 7191
rect 25228 7148 25280 7157
rect 25872 7148 25924 7200
rect 26608 7191 26660 7200
rect 26608 7157 26617 7191
rect 26617 7157 26651 7191
rect 26651 7157 26660 7191
rect 26608 7148 26660 7157
rect 27068 7148 27120 7200
rect 27344 7148 27396 7200
rect 27804 7191 27856 7200
rect 27804 7157 27813 7191
rect 27813 7157 27847 7191
rect 27847 7157 27856 7191
rect 27804 7148 27856 7157
rect 28080 7191 28132 7200
rect 28080 7157 28089 7191
rect 28089 7157 28123 7191
rect 28123 7157 28132 7191
rect 28080 7148 28132 7157
rect 28172 7148 28224 7200
rect 28632 7191 28684 7200
rect 28632 7157 28641 7191
rect 28641 7157 28675 7191
rect 28675 7157 28684 7191
rect 28632 7148 28684 7157
rect 28724 7148 28776 7200
rect 29184 7191 29236 7200
rect 29184 7157 29193 7191
rect 29193 7157 29227 7191
rect 29227 7157 29236 7191
rect 29184 7148 29236 7157
rect 29736 7148 29788 7200
rect 30012 7148 30064 7200
rect 30380 7216 30432 7268
rect 31760 7216 31812 7268
rect 33600 7216 33652 7268
rect 34796 7216 34848 7268
rect 36084 7352 36136 7404
rect 36912 7352 36964 7404
rect 37372 7395 37424 7404
rect 37372 7361 37381 7395
rect 37381 7361 37415 7395
rect 37415 7361 37424 7395
rect 37372 7352 37424 7361
rect 37832 7352 37884 7404
rect 38752 7352 38804 7404
rect 38568 7284 38620 7336
rect 40500 7395 40552 7404
rect 40500 7361 40509 7395
rect 40509 7361 40543 7395
rect 40543 7361 40552 7395
rect 40500 7352 40552 7361
rect 38660 7259 38712 7268
rect 38660 7225 38669 7259
rect 38669 7225 38703 7259
rect 38703 7225 38712 7259
rect 38660 7216 38712 7225
rect 30564 7191 30616 7200
rect 30564 7157 30573 7191
rect 30573 7157 30607 7191
rect 30607 7157 30616 7191
rect 30564 7148 30616 7157
rect 30840 7191 30892 7200
rect 30840 7157 30849 7191
rect 30849 7157 30883 7191
rect 30883 7157 30892 7191
rect 30840 7148 30892 7157
rect 31116 7191 31168 7200
rect 31116 7157 31125 7191
rect 31125 7157 31159 7191
rect 31159 7157 31168 7191
rect 31116 7148 31168 7157
rect 32128 7148 32180 7200
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 32404 7148 32456 7200
rect 35072 7148 35124 7200
rect 36452 7148 36504 7200
rect 39120 7191 39172 7200
rect 39120 7157 39129 7191
rect 39129 7157 39163 7191
rect 39163 7157 39172 7191
rect 39120 7148 39172 7157
rect 6251 7046 6303 7098
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 16854 7046 16906 7098
rect 16918 7046 16970 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 27457 7046 27509 7098
rect 27521 7046 27573 7098
rect 27585 7046 27637 7098
rect 27649 7046 27701 7098
rect 27713 7046 27765 7098
rect 38060 7046 38112 7098
rect 38124 7046 38176 7098
rect 38188 7046 38240 7098
rect 38252 7046 38304 7098
rect 38316 7046 38368 7098
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 5724 6987 5776 6996
rect 5724 6953 5733 6987
rect 5733 6953 5767 6987
rect 5767 6953 5776 6987
rect 5724 6944 5776 6953
rect 9128 6944 9180 6996
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 12072 6944 12124 6996
rect 18604 6944 18656 6996
rect 18696 6944 18748 6996
rect 18972 6944 19024 6996
rect 20812 6944 20864 6996
rect 6184 6808 6236 6860
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 4344 6740 4396 6792
rect 7196 6740 7248 6792
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 10048 6808 10100 6860
rect 10600 6808 10652 6860
rect 12348 6876 12400 6928
rect 12900 6876 12952 6928
rect 12164 6808 12216 6860
rect 12808 6808 12860 6860
rect 13360 6808 13412 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 14740 6808 14792 6860
rect 15292 6808 15344 6860
rect 15844 6808 15896 6860
rect 16396 6808 16448 6860
rect 16948 6808 17000 6860
rect 17500 6808 17552 6860
rect 18052 6808 18104 6860
rect 22928 6944 22980 6996
rect 23112 6944 23164 6996
rect 23664 6944 23716 6996
rect 25872 6944 25924 6996
rect 26608 6944 26660 6996
rect 27068 6944 27120 6996
rect 5632 6715 5684 6724
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 7840 6715 7892 6724
rect 7840 6681 7849 6715
rect 7849 6681 7883 6715
rect 7883 6681 7892 6715
rect 7840 6672 7892 6681
rect 10600 6672 10652 6724
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 12624 6740 12676 6792
rect 11612 6672 11664 6724
rect 11888 6715 11940 6724
rect 11888 6681 11897 6715
rect 11897 6681 11931 6715
rect 11931 6681 11940 6715
rect 11888 6672 11940 6681
rect 12716 6672 12768 6724
rect 13084 6740 13136 6792
rect 14188 6740 14240 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 18420 6740 18472 6792
rect 19432 6740 19484 6792
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 15016 6672 15068 6724
rect 15108 6672 15160 6724
rect 16028 6715 16080 6724
rect 16028 6681 16037 6715
rect 16037 6681 16071 6715
rect 16071 6681 16080 6715
rect 16028 6672 16080 6681
rect 16580 6715 16632 6724
rect 16580 6681 16589 6715
rect 16589 6681 16623 6715
rect 16623 6681 16632 6715
rect 16580 6672 16632 6681
rect 17132 6715 17184 6724
rect 17132 6681 17141 6715
rect 17141 6681 17175 6715
rect 17175 6681 17184 6715
rect 17132 6672 17184 6681
rect 17684 6715 17736 6724
rect 17684 6681 17693 6715
rect 17693 6681 17727 6715
rect 17727 6681 17736 6715
rect 17684 6672 17736 6681
rect 18236 6715 18288 6724
rect 18236 6681 18245 6715
rect 18245 6681 18279 6715
rect 18279 6681 18288 6715
rect 18236 6672 18288 6681
rect 10692 6604 10744 6656
rect 10876 6604 10928 6656
rect 19616 6672 19668 6724
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 20536 6740 20588 6792
rect 20628 6783 20680 6792
rect 20628 6749 20637 6783
rect 20637 6749 20671 6783
rect 20671 6749 20680 6783
rect 20628 6740 20680 6749
rect 20812 6740 20864 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21916 6740 21968 6792
rect 23204 6740 23256 6792
rect 18420 6604 18472 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 20628 6604 20680 6656
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 21272 6604 21324 6656
rect 23388 6672 23440 6724
rect 21732 6604 21784 6656
rect 22836 6647 22888 6656
rect 22836 6613 22845 6647
rect 22845 6613 22879 6647
rect 22879 6613 22888 6647
rect 22836 6604 22888 6613
rect 23112 6647 23164 6656
rect 23112 6613 23121 6647
rect 23121 6613 23155 6647
rect 23155 6613 23164 6647
rect 23112 6604 23164 6613
rect 26424 6740 26476 6792
rect 27804 6944 27856 6996
rect 28080 6944 28132 6996
rect 28632 6944 28684 6996
rect 37556 6876 37608 6928
rect 27344 6740 27396 6792
rect 34060 6808 34112 6860
rect 35164 6808 35216 6860
rect 35716 6808 35768 6860
rect 37096 6808 37148 6860
rect 38292 6808 38344 6860
rect 39580 6808 39632 6860
rect 28172 6740 28224 6792
rect 28724 6740 28776 6792
rect 28816 6783 28868 6792
rect 28816 6749 28825 6783
rect 28825 6749 28859 6783
rect 28859 6749 28868 6783
rect 28816 6740 28868 6749
rect 29184 6740 29236 6792
rect 29736 6740 29788 6792
rect 30012 6740 30064 6792
rect 33048 6783 33100 6792
rect 33048 6749 33057 6783
rect 33057 6749 33091 6783
rect 33091 6749 33100 6783
rect 33048 6740 33100 6749
rect 33324 6783 33376 6792
rect 33324 6749 33333 6783
rect 33333 6749 33367 6783
rect 33367 6749 33376 6783
rect 33324 6740 33376 6749
rect 33600 6783 33652 6792
rect 33600 6749 33609 6783
rect 33609 6749 33643 6783
rect 33643 6749 33652 6783
rect 33600 6740 33652 6749
rect 33692 6740 33744 6792
rect 36728 6740 36780 6792
rect 25504 6647 25556 6656
rect 25504 6613 25513 6647
rect 25513 6613 25547 6647
rect 25547 6613 25556 6647
rect 25504 6604 25556 6613
rect 25964 6647 26016 6656
rect 25964 6613 25973 6647
rect 25973 6613 26007 6647
rect 26007 6613 26016 6647
rect 25964 6604 26016 6613
rect 26332 6647 26384 6656
rect 26332 6613 26341 6647
rect 26341 6613 26375 6647
rect 26375 6613 26384 6647
rect 26332 6604 26384 6613
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 27068 6647 27120 6656
rect 27068 6613 27077 6647
rect 27077 6613 27111 6647
rect 27111 6613 27120 6647
rect 27068 6604 27120 6613
rect 27160 6604 27212 6656
rect 27528 6604 27580 6656
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 28540 6647 28592 6656
rect 28540 6613 28549 6647
rect 28549 6613 28583 6647
rect 28583 6613 28592 6647
rect 28540 6604 28592 6613
rect 35348 6715 35400 6724
rect 35348 6681 35357 6715
rect 35357 6681 35391 6715
rect 35391 6681 35400 6715
rect 35348 6672 35400 6681
rect 35900 6715 35952 6724
rect 35900 6681 35909 6715
rect 35909 6681 35943 6715
rect 35943 6681 35952 6715
rect 35900 6672 35952 6681
rect 37004 6715 37056 6724
rect 37004 6681 37013 6715
rect 37013 6681 37047 6715
rect 37047 6681 37056 6715
rect 37004 6672 37056 6681
rect 38844 6740 38896 6792
rect 39028 6740 39080 6792
rect 37740 6672 37792 6724
rect 38476 6672 38528 6724
rect 29092 6647 29144 6656
rect 29092 6613 29101 6647
rect 29101 6613 29135 6647
rect 29135 6613 29144 6647
rect 29092 6604 29144 6613
rect 29276 6604 29328 6656
rect 30012 6647 30064 6656
rect 30012 6613 30021 6647
rect 30021 6613 30055 6647
rect 30055 6613 30064 6647
rect 30012 6604 30064 6613
rect 30288 6647 30340 6656
rect 30288 6613 30297 6647
rect 30297 6613 30331 6647
rect 30331 6613 30340 6647
rect 30288 6604 30340 6613
rect 33232 6647 33284 6656
rect 33232 6613 33241 6647
rect 33241 6613 33275 6647
rect 33275 6613 33284 6647
rect 33232 6604 33284 6613
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 33784 6647 33836 6656
rect 33784 6613 33793 6647
rect 33793 6613 33827 6647
rect 33827 6613 33836 6647
rect 33784 6604 33836 6613
rect 35992 6604 36044 6656
rect 36636 6604 36688 6656
rect 37648 6604 37700 6656
rect 38384 6604 38436 6656
rect 38936 6672 38988 6724
rect 39948 6715 40000 6724
rect 39948 6681 39957 6715
rect 39957 6681 39991 6715
rect 39991 6681 40000 6715
rect 39948 6672 40000 6681
rect 41328 6672 41380 6724
rect 11552 6502 11604 6554
rect 11616 6502 11668 6554
rect 11680 6502 11732 6554
rect 11744 6502 11796 6554
rect 11808 6502 11860 6554
rect 22155 6502 22207 6554
rect 22219 6502 22271 6554
rect 22283 6502 22335 6554
rect 22347 6502 22399 6554
rect 22411 6502 22463 6554
rect 32758 6502 32810 6554
rect 32822 6502 32874 6554
rect 32886 6502 32938 6554
rect 32950 6502 33002 6554
rect 33014 6502 33066 6554
rect 43361 6502 43413 6554
rect 43425 6502 43477 6554
rect 43489 6502 43541 6554
rect 43553 6502 43605 6554
rect 43617 6502 43669 6554
rect 5632 6400 5684 6452
rect 6736 6400 6788 6452
rect 9220 6443 9272 6452
rect 9220 6409 9229 6443
rect 9229 6409 9263 6443
rect 9263 6409 9272 6443
rect 9220 6400 9272 6409
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 12256 6400 12308 6452
rect 11980 6332 12032 6384
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 5540 6196 5592 6248
rect 9864 6264 9916 6316
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 13912 6400 13964 6452
rect 15108 6400 15160 6452
rect 14004 6332 14056 6384
rect 15384 6332 15436 6384
rect 15568 6400 15620 6452
rect 16028 6400 16080 6452
rect 16580 6400 16632 6452
rect 17132 6400 17184 6452
rect 14464 6264 14516 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15016 6264 15068 6316
rect 9680 6128 9732 6180
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 15752 6264 15804 6316
rect 16212 6264 16264 6316
rect 17408 6400 17460 6452
rect 17684 6400 17736 6452
rect 17868 6400 17920 6452
rect 18236 6400 18288 6452
rect 18512 6400 18564 6452
rect 19340 6400 19392 6452
rect 19616 6400 19668 6452
rect 21088 6400 21140 6452
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 16764 6196 16816 6248
rect 17224 6196 17276 6248
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 19800 6332 19852 6384
rect 23112 6400 23164 6452
rect 24676 6400 24728 6452
rect 25228 6400 25280 6452
rect 25596 6400 25648 6452
rect 29092 6400 29144 6452
rect 31760 6400 31812 6452
rect 36728 6400 36780 6452
rect 37004 6400 37056 6452
rect 37924 6400 37976 6452
rect 39120 6400 39172 6452
rect 23664 6264 23716 6316
rect 23756 6264 23808 6316
rect 30380 6332 30432 6384
rect 38292 6332 38344 6384
rect 38660 6332 38712 6384
rect 22008 6128 22060 6180
rect 23020 6128 23072 6180
rect 14372 6060 14424 6112
rect 19892 6060 19944 6112
rect 23388 6103 23440 6112
rect 23388 6069 23397 6103
rect 23397 6069 23431 6103
rect 23431 6069 23440 6103
rect 23388 6060 23440 6069
rect 24032 6171 24084 6180
rect 24032 6137 24041 6171
rect 24041 6137 24075 6171
rect 24075 6137 24084 6171
rect 24032 6128 24084 6137
rect 24308 6128 24360 6180
rect 24768 6128 24820 6180
rect 28540 6128 28592 6180
rect 32312 6128 32364 6180
rect 25964 6060 26016 6112
rect 6251 5958 6303 6010
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 16854 5958 16906 6010
rect 16918 5958 16970 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 27457 5958 27509 6010
rect 27521 5958 27573 6010
rect 27585 5958 27637 6010
rect 27649 5958 27701 6010
rect 27713 5958 27765 6010
rect 38060 5958 38112 6010
rect 38124 5958 38176 6010
rect 38188 5958 38240 6010
rect 38252 5958 38304 6010
rect 38316 5958 38368 6010
rect 5908 5856 5960 5908
rect 9496 5856 9548 5908
rect 12716 5856 12768 5908
rect 17224 5856 17276 5908
rect 20260 5856 20312 5908
rect 20720 5856 20772 5908
rect 27160 5856 27212 5908
rect 23204 5788 23256 5840
rect 30288 5788 30340 5840
rect 4528 5720 4580 5772
rect 7840 5652 7892 5704
rect 11060 5652 11112 5704
rect 11888 5652 11940 5704
rect 15108 5652 15160 5704
rect 13728 5584 13780 5636
rect 18604 5720 18656 5772
rect 22744 5720 22796 5772
rect 23296 5720 23348 5772
rect 25504 5720 25556 5772
rect 20536 5584 20588 5636
rect 19340 5516 19392 5568
rect 24584 5516 24636 5568
rect 11552 5414 11604 5466
rect 11616 5414 11668 5466
rect 11680 5414 11732 5466
rect 11744 5414 11796 5466
rect 11808 5414 11860 5466
rect 22155 5414 22207 5466
rect 22219 5414 22271 5466
rect 22283 5414 22335 5466
rect 22347 5414 22399 5466
rect 22411 5414 22463 5466
rect 32758 5414 32810 5466
rect 32822 5414 32874 5466
rect 32886 5414 32938 5466
rect 32950 5414 33002 5466
rect 33014 5414 33066 5466
rect 43361 5414 43413 5466
rect 43425 5414 43477 5466
rect 43489 5414 43541 5466
rect 43553 5414 43605 5466
rect 43617 5414 43669 5466
rect 16764 5312 16816 5364
rect 26332 5312 26384 5364
rect 15384 5244 15436 5296
rect 23296 5244 23348 5296
rect 17224 5176 17276 5228
rect 26700 5176 26752 5228
rect 15108 5108 15160 5160
rect 27988 5108 28040 5160
rect 12624 5040 12676 5092
rect 25596 5040 25648 5092
rect 10784 4972 10836 5024
rect 30012 4972 30064 5024
rect 6251 4870 6303 4922
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 16854 4870 16906 4922
rect 16918 4870 16970 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 27457 4870 27509 4922
rect 27521 4870 27573 4922
rect 27585 4870 27637 4922
rect 27649 4870 27701 4922
rect 27713 4870 27765 4922
rect 38060 4870 38112 4922
rect 38124 4870 38176 4922
rect 38188 4870 38240 4922
rect 38252 4870 38304 4922
rect 38316 4870 38368 4922
rect 12440 4768 12492 4820
rect 27344 4768 27396 4820
rect 6828 4700 6880 4752
rect 19800 4700 19852 4752
rect 11552 4326 11604 4378
rect 11616 4326 11668 4378
rect 11680 4326 11732 4378
rect 11744 4326 11796 4378
rect 11808 4326 11860 4378
rect 22155 4326 22207 4378
rect 22219 4326 22271 4378
rect 22283 4326 22335 4378
rect 22347 4326 22399 4378
rect 22411 4326 22463 4378
rect 32758 4326 32810 4378
rect 32822 4326 32874 4378
rect 32886 4326 32938 4378
rect 32950 4326 33002 4378
rect 33014 4326 33066 4378
rect 43361 4326 43413 4378
rect 43425 4326 43477 4378
rect 43489 4326 43541 4378
rect 43553 4326 43605 4378
rect 43617 4326 43669 4378
rect 30840 3884 30892 3936
rect 35900 3884 35952 3936
rect 6251 3782 6303 3834
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 16854 3782 16906 3834
rect 16918 3782 16970 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 27457 3782 27509 3834
rect 27521 3782 27573 3834
rect 27585 3782 27637 3834
rect 27649 3782 27701 3834
rect 27713 3782 27765 3834
rect 38060 3782 38112 3834
rect 38124 3782 38176 3834
rect 38188 3782 38240 3834
rect 38252 3782 38304 3834
rect 38316 3782 38368 3834
rect 34428 3680 34480 3732
rect 5632 3476 5684 3528
rect 11552 3238 11604 3290
rect 11616 3238 11668 3290
rect 11680 3238 11732 3290
rect 11744 3238 11796 3290
rect 11808 3238 11860 3290
rect 22155 3238 22207 3290
rect 22219 3238 22271 3290
rect 22283 3238 22335 3290
rect 22347 3238 22399 3290
rect 22411 3238 22463 3290
rect 32758 3238 32810 3290
rect 32822 3238 32874 3290
rect 32886 3238 32938 3290
rect 32950 3238 33002 3290
rect 33014 3238 33066 3290
rect 43361 3238 43413 3290
rect 43425 3238 43477 3290
rect 43489 3238 43541 3290
rect 43553 3238 43605 3290
rect 43617 3238 43669 3290
rect 24952 3136 25004 3188
rect 25228 3136 25280 3188
rect 38568 3136 38620 3188
rect 38844 3136 38896 3188
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 22652 3043 22704 3052
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 24860 3000 24912 3052
rect 24952 3043 25004 3052
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 25044 2864 25096 2916
rect 31760 3000 31812 3052
rect 33508 3043 33560 3052
rect 33508 3009 33517 3043
rect 33517 3009 33551 3043
rect 33551 3009 33560 3043
rect 33508 3000 33560 3009
rect 37280 3000 37332 3052
rect 37832 3000 37884 3052
rect 25320 2932 25372 2984
rect 37924 2932 37976 2984
rect 25228 2864 25280 2916
rect 33692 2864 33744 2916
rect 30380 2796 30432 2848
rect 6251 2694 6303 2746
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 16854 2694 16906 2746
rect 16918 2694 16970 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 27457 2694 27509 2746
rect 27521 2694 27573 2746
rect 27585 2694 27637 2746
rect 27649 2694 27701 2746
rect 27713 2694 27765 2746
rect 38060 2694 38112 2746
rect 38124 2694 38176 2746
rect 38188 2694 38240 2746
rect 38252 2694 38304 2746
rect 38316 2694 38368 2746
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 16672 2592 16724 2644
rect 18604 2592 18656 2644
rect 20720 2592 20772 2644
rect 22652 2592 22704 2644
rect 24952 2592 25004 2644
rect 30840 2524 30892 2576
rect 33232 2592 33284 2644
rect 33508 2592 33560 2644
rect 34152 2592 34204 2644
rect 35348 2592 35400 2644
rect 37740 2592 37792 2644
rect 37832 2635 37884 2644
rect 37832 2601 37841 2635
rect 37841 2601 37875 2635
rect 37875 2601 37884 2635
rect 37832 2592 37884 2601
rect 38752 2592 38804 2644
rect 39948 2592 40000 2644
rect 40500 2592 40552 2644
rect 41328 2592 41380 2644
rect 1124 2388 1176 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3240 2388 3292 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 13820 2388 13872 2440
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 20444 2431 20496 2440
rect 20444 2397 20453 2431
rect 20453 2397 20487 2431
rect 20487 2397 20496 2431
rect 20444 2388 20496 2397
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 26608 2431 26660 2440
rect 26608 2397 26617 2431
rect 26617 2397 26651 2431
rect 26651 2397 26660 2431
rect 26608 2388 26660 2397
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 29828 2456 29880 2508
rect 34796 2524 34848 2576
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 33600 2431 33652 2440
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 33968 2431 34020 2440
rect 33968 2397 33977 2431
rect 33977 2397 34011 2431
rect 34011 2397 34020 2431
rect 33968 2388 34020 2397
rect 34428 2431 34480 2440
rect 34428 2397 34437 2431
rect 34437 2397 34471 2431
rect 34471 2397 34480 2431
rect 34428 2388 34480 2397
rect 37188 2456 37240 2508
rect 35256 2431 35308 2440
rect 35256 2397 35265 2431
rect 35265 2397 35299 2431
rect 35299 2397 35308 2431
rect 35256 2388 35308 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 26792 2295 26844 2304
rect 26792 2261 26801 2295
rect 26801 2261 26835 2295
rect 26835 2261 26844 2295
rect 26792 2252 26844 2261
rect 28816 2252 28868 2304
rect 32680 2252 32732 2304
rect 33416 2252 33468 2304
rect 36820 2320 36872 2372
rect 38936 2320 38988 2372
rect 39488 2431 39540 2440
rect 39488 2397 39497 2431
rect 39497 2397 39531 2431
rect 39531 2397 39540 2431
rect 39488 2388 39540 2397
rect 41604 2431 41656 2440
rect 41604 2397 41613 2431
rect 41613 2397 41647 2431
rect 41647 2397 41656 2431
rect 41604 2388 41656 2397
rect 43168 2431 43220 2440
rect 43168 2397 43177 2431
rect 43177 2397 43211 2431
rect 43211 2397 43220 2431
rect 43168 2388 43220 2397
rect 11552 2150 11604 2202
rect 11616 2150 11668 2202
rect 11680 2150 11732 2202
rect 11744 2150 11796 2202
rect 11808 2150 11860 2202
rect 22155 2150 22207 2202
rect 22219 2150 22271 2202
rect 22283 2150 22335 2202
rect 22347 2150 22399 2202
rect 22411 2150 22463 2202
rect 32758 2150 32810 2202
rect 32822 2150 32874 2202
rect 32886 2150 32938 2202
rect 32950 2150 33002 2202
rect 33014 2150 33066 2202
rect 43361 2150 43413 2202
rect 43425 2150 43477 2202
rect 43489 2150 43541 2202
rect 43553 2150 43605 2202
rect 43617 2150 43669 2202
rect 1676 2048 1728 2100
rect 4068 2048 4120 2100
rect 7748 2048 7800 2100
rect 9864 2048 9916 2100
rect 29828 2048 29880 2100
rect 34428 2048 34480 2100
rect 34520 2048 34572 2100
rect 36084 2048 36136 2100
rect 36820 2048 36872 2100
rect 37464 2048 37516 2100
rect 32680 1980 32732 2032
rect 33416 1912 33468 1964
rect 33968 1844 34020 1896
rect 33324 1776 33376 1828
rect 26792 1640 26844 1692
rect 36912 1640 36964 1692
rect 28816 1572 28868 1624
rect 34520 1572 34572 1624
rect 32864 1368 32916 1420
rect 33600 1368 33652 1420
<< metal2 >>
rect 5078 9840 5134 10300
rect 5354 9840 5410 10300
rect 5630 9840 5686 10300
rect 5906 9840 5962 10300
rect 6182 9840 6238 10300
rect 6458 9840 6514 10300
rect 6734 9840 6790 10300
rect 7010 9840 7066 10300
rect 7286 9840 7342 10300
rect 7562 9840 7618 10300
rect 7838 9840 7894 10300
rect 8114 9840 8170 10300
rect 8390 9840 8446 10300
rect 8666 9840 8722 10300
rect 8942 9840 8998 10300
rect 9218 9840 9274 10300
rect 9494 9840 9550 10300
rect 9770 9840 9826 10300
rect 10046 9840 10102 10300
rect 10322 9840 10378 10300
rect 10598 9840 10654 10300
rect 10874 9840 10930 10300
rect 11150 9840 11206 10300
rect 11426 9840 11482 10300
rect 11702 9840 11758 10300
rect 11978 9840 12034 10300
rect 12254 9840 12310 10300
rect 12530 9840 12586 10300
rect 12806 9840 12862 10300
rect 13082 9840 13138 10300
rect 13358 9840 13414 10300
rect 13634 9840 13690 10300
rect 13910 9840 13966 10300
rect 14186 9840 14242 10300
rect 14462 9840 14518 10300
rect 14738 9840 14794 10300
rect 15014 9840 15070 10300
rect 15290 9840 15346 10300
rect 15566 9840 15622 10300
rect 15842 9840 15898 10300
rect 16118 9840 16174 10300
rect 16394 9840 16450 10300
rect 16670 9840 16726 10300
rect 16946 9840 17002 10300
rect 17222 9840 17278 10300
rect 17498 9840 17554 10300
rect 17774 9840 17830 10300
rect 18050 9840 18106 10300
rect 18326 9840 18382 10300
rect 18602 9840 18658 10300
rect 18878 9840 18934 10300
rect 19154 9840 19210 10300
rect 19430 9840 19486 10300
rect 19706 9840 19762 10300
rect 19982 9840 20038 10300
rect 20258 9840 20314 10300
rect 20534 9840 20590 10300
rect 20810 9840 20866 10300
rect 21086 9840 21142 10300
rect 21362 9840 21418 10300
rect 21638 9840 21694 10300
rect 21914 9840 21970 10300
rect 22190 9840 22246 10300
rect 22466 9840 22522 10300
rect 22742 9840 22798 10300
rect 23018 9840 23074 10300
rect 23294 9840 23350 10300
rect 23570 9840 23626 10300
rect 23846 9840 23902 10300
rect 24122 9840 24178 10300
rect 24398 9840 24454 10300
rect 24674 9840 24730 10300
rect 24950 9840 25006 10300
rect 25226 9840 25282 10300
rect 25502 9840 25558 10300
rect 25778 9840 25834 10300
rect 26054 9840 26110 10300
rect 26330 9840 26386 10300
rect 26606 9840 26662 10300
rect 26882 9840 26938 10300
rect 27158 9840 27214 10300
rect 27434 9840 27490 10300
rect 27710 9840 27766 10300
rect 27986 9840 28042 10300
rect 28262 9840 28318 10300
rect 28538 9840 28594 10300
rect 28814 9840 28870 10300
rect 29090 9840 29146 10300
rect 29366 9840 29422 10300
rect 29642 9840 29698 10300
rect 29918 9840 29974 10300
rect 30194 9840 30250 10300
rect 30470 9840 30526 10300
rect 30746 9840 30802 10300
rect 31022 9840 31078 10300
rect 31298 9840 31354 10300
rect 31574 9840 31630 10300
rect 31850 9840 31906 10300
rect 32126 9840 32182 10300
rect 32402 9840 32458 10300
rect 32678 9840 32734 10300
rect 32954 9840 33010 10300
rect 33230 9840 33286 10300
rect 33506 9840 33562 10300
rect 33782 9840 33838 10300
rect 34058 9840 34114 10300
rect 34334 9840 34390 10300
rect 34610 9840 34666 10300
rect 34886 9840 34942 10300
rect 35162 9840 35218 10300
rect 35438 9840 35494 10300
rect 35714 9840 35770 10300
rect 35990 9840 36046 10300
rect 36266 9840 36322 10300
rect 36542 9840 36598 10300
rect 36818 9840 36874 10300
rect 37094 9840 37150 10300
rect 37370 9840 37426 10300
rect 37646 9840 37702 10300
rect 37922 9840 37978 10300
rect 38198 9840 38254 10300
rect 38474 9840 38530 10300
rect 38750 9840 38806 10300
rect 39026 9840 39082 10300
rect 39302 9840 39358 10300
rect 39578 9840 39634 10300
rect 5092 8242 5120 9840
rect 5092 8214 5212 8242
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4356 6798 4384 7142
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4540 5778 4568 7346
rect 5184 7002 5212 8214
rect 5368 7546 5396 9840
rect 5644 8242 5672 9840
rect 5644 8214 5764 8242
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5552 6254 5580 7346
rect 5736 7002 5764 8214
rect 5920 7546 5948 9840
rect 6196 8242 6224 9840
rect 6104 8214 6224 8242
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5644 6458 5672 6666
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 6248 5592 6254
rect 5828 6225 5856 7346
rect 6104 6848 6132 8214
rect 6472 7342 6500 9840
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6251 7100 6559 7109
rect 6251 7098 6257 7100
rect 6313 7098 6337 7100
rect 6393 7098 6417 7100
rect 6473 7098 6497 7100
rect 6553 7098 6559 7100
rect 6313 7046 6315 7098
rect 6495 7046 6497 7098
rect 6251 7044 6257 7046
rect 6313 7044 6337 7046
rect 6393 7044 6417 7046
rect 6473 7044 6497 7046
rect 6553 7044 6559 7046
rect 6251 7035 6559 7044
rect 6184 6860 6236 6866
rect 6104 6820 6184 6848
rect 6184 6802 6236 6808
rect 6182 6760 6238 6769
rect 6182 6695 6184 6704
rect 6236 6695 6238 6704
rect 6184 6666 6236 6672
rect 6748 6458 6776 9840
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5540 6190 5592 6196
rect 5814 6216 5870 6225
rect 5814 6151 5870 6160
rect 5920 5914 5948 6258
rect 6251 6012 6559 6021
rect 6251 6010 6257 6012
rect 6313 6010 6337 6012
rect 6393 6010 6417 6012
rect 6473 6010 6497 6012
rect 6553 6010 6559 6012
rect 6313 5958 6315 6010
rect 6495 5958 6497 6010
rect 6251 5956 6257 5958
rect 6313 5956 6337 5958
rect 6393 5956 6417 5958
rect 6473 5956 6497 5958
rect 6553 5956 6559 5958
rect 6251 5947 6559 5956
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 6251 4924 6559 4933
rect 6251 4922 6257 4924
rect 6313 4922 6337 4924
rect 6393 4922 6417 4924
rect 6473 4922 6497 4924
rect 6553 4922 6559 4924
rect 6313 4870 6315 4922
rect 6495 4870 6497 4922
rect 6251 4868 6257 4870
rect 6313 4868 6337 4870
rect 6393 4868 6417 4870
rect 6473 4868 6497 4870
rect 6553 4868 6559 4870
rect 6251 4859 6559 4868
rect 6840 4758 6868 7346
rect 7024 6866 7052 9840
rect 7196 8220 7248 8226
rect 7196 8162 7248 8168
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7208 6798 7236 8162
rect 7300 7546 7328 9840
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7576 6866 7604 9840
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 7410 7788 7686
rect 7852 7546 7880 9840
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8128 6866 8156 9840
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7410 8340 7686
rect 8404 7546 8432 9840
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8680 6866 8708 9840
rect 8956 7546 8984 9840
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9140 7002 9168 7346
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 5710 7880 6666
rect 9232 6458 9260 9840
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9508 5914 9536 9840
rect 9784 6458 9812 9840
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 6322 9904 7210
rect 10060 6866 10088 9840
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10336 6458 10364 9840
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10520 7546 10548 8298
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 6866 10640 9840
rect 10888 7002 10916 9840
rect 11164 7546 11192 9840
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11348 7410 11376 7958
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 7840 5704 7892 5710
rect 9692 5681 9720 6122
rect 7840 5646 7892 5652
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 10612 5273 10640 6666
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6458 10732 6598
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10598 5264 10654 5273
rect 10598 5199 10654 5208
rect 10796 5030 10824 6666
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6322 10916 6598
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11072 5710 11100 7142
rect 11440 7002 11468 9840
rect 11716 7834 11744 9840
rect 11716 7806 11928 7834
rect 11552 7644 11860 7653
rect 11552 7642 11558 7644
rect 11614 7642 11638 7644
rect 11694 7642 11718 7644
rect 11774 7642 11798 7644
rect 11854 7642 11860 7644
rect 11614 7590 11616 7642
rect 11796 7590 11798 7642
rect 11552 7588 11558 7590
rect 11614 7588 11638 7590
rect 11694 7588 11718 7590
rect 11774 7588 11798 7590
rect 11854 7588 11860 7590
rect 11552 7579 11860 7588
rect 11900 7342 11928 7806
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11610 7032 11666 7041
rect 11428 6996 11480 7002
rect 11992 7002 12020 9840
rect 12162 8256 12218 8265
rect 12162 8191 12218 8200
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7002 12112 7346
rect 11610 6967 11666 6976
rect 11980 6996 12032 7002
rect 11428 6938 11480 6944
rect 11624 6730 11652 6967
rect 11980 6938 12032 6944
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12176 6866 12204 8191
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11552 6556 11860 6565
rect 11552 6554 11558 6556
rect 11614 6554 11638 6556
rect 11694 6554 11718 6556
rect 11774 6554 11798 6556
rect 11854 6554 11860 6556
rect 11614 6502 11616 6554
rect 11796 6502 11798 6554
rect 11552 6500 11558 6502
rect 11614 6500 11638 6502
rect 11694 6500 11718 6502
rect 11774 6500 11798 6502
rect 11854 6500 11860 6502
rect 11552 6491 11860 6500
rect 11900 5710 11928 6666
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11992 6390 12020 6559
rect 12268 6458 12296 9840
rect 12544 7546 12572 9840
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12636 7546 12664 8026
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12636 7410 12664 7482
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 12360 5545 12388 6870
rect 12820 6866 12848 9840
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12912 7478 12940 7754
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12912 6934 12940 7278
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 13096 6798 13124 9840
rect 13372 6866 13400 9840
rect 13648 7546 13676 9840
rect 13726 8392 13782 8401
rect 13726 8327 13782 8336
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12346 5536 12402 5545
rect 11552 5468 11860 5477
rect 12346 5471 12402 5480
rect 11552 5466 11558 5468
rect 11614 5466 11638 5468
rect 11694 5466 11718 5468
rect 11774 5466 11798 5468
rect 11854 5466 11860 5468
rect 11614 5414 11616 5466
rect 11796 5414 11798 5466
rect 11552 5412 11558 5414
rect 11614 5412 11638 5414
rect 11694 5412 11718 5414
rect 11774 5412 11798 5414
rect 11854 5412 11860 5414
rect 11552 5403 11860 5412
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 12452 4826 12480 6258
rect 12636 5098 12664 6734
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 5914 12756 6666
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 13740 5642 13768 8327
rect 13924 6458 13952 9840
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14016 6390 14044 7822
rect 14200 7546 14228 9840
rect 14476 8242 14504 9840
rect 14476 8214 14688 8242
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14188 6792 14240 6798
rect 14292 6769 14320 7346
rect 14384 6798 14412 7958
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 6792 14424 6798
rect 14188 6734 14240 6740
rect 14278 6760 14334 6769
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 6828 4752 6880 4758
rect 14200 4729 14228 6734
rect 14372 6734 14424 6740
rect 14278 6695 14334 6704
rect 14370 6488 14426 6497
rect 14370 6423 14426 6432
rect 14384 6118 14412 6423
rect 14476 6322 14504 7346
rect 14660 6866 14688 8214
rect 14752 6866 14780 9840
rect 15028 7546 15056 9840
rect 15106 8528 15162 8537
rect 15106 8463 15162 8472
rect 15120 7954 15148 8463
rect 15200 8152 15252 8158
rect 15200 8094 15252 8100
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 15212 6746 15240 8094
rect 15304 6866 15332 9840
rect 15580 7546 15608 9840
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 15108 6724 15160 6730
rect 15212 6718 15332 6746
rect 15108 6666 15160 6672
rect 15028 6322 15056 6666
rect 15120 6458 15148 6666
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15198 6352 15254 6361
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15016 6316 15068 6322
rect 15198 6287 15200 6296
rect 15016 6258 15068 6264
rect 15252 6287 15254 6296
rect 15200 6258 15252 6264
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14936 5137 14964 6258
rect 15304 5817 15332 6718
rect 15580 6458 15608 7346
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15290 5808 15346 5817
rect 15290 5743 15346 5752
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 5166 15148 5646
rect 15396 5302 15424 6326
rect 15672 6322 15700 8366
rect 15764 6322 15792 8434
rect 15856 6866 15884 9840
rect 15934 7848 15990 7857
rect 15934 7783 15990 7792
rect 15948 7478 15976 7783
rect 16132 7562 16160 9840
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16040 7546 16160 7562
rect 16028 7540 16160 7546
rect 16080 7534 16160 7540
rect 16028 7482 16080 7488
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16040 6458 16068 6666
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16224 6322 16252 8502
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7274 16344 7686
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16408 6866 16436 9840
rect 16486 8120 16542 8129
rect 16486 8055 16542 8064
rect 16500 7206 16528 8055
rect 16684 7410 16712 9840
rect 16960 8242 16988 9840
rect 17236 8514 17264 9840
rect 16776 8214 16988 8242
rect 17144 8486 17264 8514
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16592 7041 16620 7142
rect 16578 7032 16634 7041
rect 16578 6967 16634 6976
rect 16776 6984 16804 8214
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7410 16896 7686
rect 17144 7546 17172 8486
rect 17314 7984 17370 7993
rect 17314 7919 17370 7928
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 16854 7100 17162 7109
rect 16854 7098 16860 7100
rect 16916 7098 16940 7100
rect 16996 7098 17020 7100
rect 17076 7098 17100 7100
rect 17156 7098 17162 7100
rect 16916 7046 16918 7098
rect 17098 7046 17100 7098
rect 16854 7044 16860 7046
rect 16916 7044 16940 7046
rect 16996 7044 17020 7046
rect 17076 7044 17100 7046
rect 17156 7044 17162 7046
rect 16854 7035 17162 7044
rect 16776 6956 16988 6984
rect 16960 6866 16988 6956
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16592 6458 16620 6666
rect 17144 6458 17172 6666
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 17236 6254 17264 7346
rect 17328 7177 17356 7919
rect 17406 7304 17462 7313
rect 17406 7239 17462 7248
rect 17314 7168 17370 7177
rect 17314 7103 17370 7112
rect 17420 6458 17448 7239
rect 17512 6866 17540 9840
rect 17788 8514 17816 9840
rect 17696 8486 17816 8514
rect 17696 7546 17724 8486
rect 17774 7984 17830 7993
rect 17774 7919 17830 7928
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17696 6458 17724 6666
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17788 6322 17816 7919
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 6458 17908 7346
rect 18064 6866 18092 9840
rect 18340 8514 18368 9840
rect 18248 8486 18368 8514
rect 18616 8514 18644 9840
rect 18616 8486 18828 8514
rect 18248 7546 18276 8486
rect 18800 7546 18828 8486
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18892 7478 18920 9840
rect 19168 7546 19196 9840
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 18880 7472 18932 7478
rect 18326 7440 18382 7449
rect 18880 7414 18932 7420
rect 18326 7375 18382 7384
rect 18512 7404 18564 7410
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18248 6458 18276 6666
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18340 6338 18368 7375
rect 18512 7346 18564 7352
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 18418 7032 18474 7041
rect 18418 6967 18474 6976
rect 18432 6798 18460 6967
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6497 18460 6598
rect 18418 6488 18474 6497
rect 18524 6458 18552 7346
rect 18708 7002 18736 7346
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18696 6996 18748 7002
rect 18972 6996 19024 7002
rect 18696 6938 18748 6944
rect 18892 6956 18972 6984
rect 18616 6882 18644 6938
rect 18892 6882 18920 6956
rect 18972 6938 19024 6944
rect 18616 6854 18920 6882
rect 19352 6458 19380 7346
rect 19444 6798 19472 9840
rect 19720 8378 19748 9840
rect 19536 8350 19748 8378
rect 19996 8378 20024 9840
rect 20272 9738 20300 9840
rect 20272 9710 20392 9738
rect 19996 8350 20116 8378
rect 19536 6798 19564 8350
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19628 6458 19656 6666
rect 18418 6423 18474 6432
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 18248 6322 18368 6338
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 18236 6316 18368 6322
rect 18288 6310 18368 6316
rect 18604 6316 18656 6322
rect 18236 6258 18288 6264
rect 18604 6258 18656 6264
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16776 5370 16804 6190
rect 16854 6012 17162 6021
rect 16854 6010 16860 6012
rect 16916 6010 16940 6012
rect 16996 6010 17020 6012
rect 17076 6010 17100 6012
rect 17156 6010 17162 6012
rect 16916 5958 16918 6010
rect 17098 5958 17100 6010
rect 16854 5956 16860 5958
rect 16916 5956 16940 5958
rect 16996 5956 17020 5958
rect 17076 5956 17100 5958
rect 17156 5956 17162 5958
rect 16854 5947 17162 5956
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 17236 5234 17264 5850
rect 18616 5778 18644 6258
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 19352 5574 19380 6258
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 15108 5160 15160 5166
rect 14922 5128 14978 5137
rect 15108 5102 15160 5108
rect 14922 5063 14978 5072
rect 16854 4924 17162 4933
rect 16854 4922 16860 4924
rect 16916 4922 16940 4924
rect 16996 4922 17020 4924
rect 17076 4922 17100 4924
rect 17156 4922 17162 4924
rect 16916 4870 16918 4922
rect 17098 4870 17100 4922
rect 16854 4868 16860 4870
rect 16916 4868 16940 4870
rect 16996 4868 17020 4870
rect 17076 4868 17100 4870
rect 17156 4868 17162 4870
rect 16854 4859 17162 4868
rect 19812 4758 19840 6326
rect 19904 6118 19932 7346
rect 20088 6798 20116 8350
rect 20364 6798 20392 9710
rect 20548 8378 20576 9840
rect 20824 8378 20852 9840
rect 20548 8350 20668 8378
rect 20824 8350 20944 8378
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20548 6798 20576 7482
rect 20640 6798 20668 8350
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 19984 6656 20036 6662
rect 19982 6624 19984 6633
rect 20260 6656 20312 6662
rect 20036 6624 20038 6633
rect 20260 6598 20312 6604
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 19982 6559 20038 6568
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 20272 5914 20300 6598
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20548 5642 20576 6598
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 20640 5545 20668 6598
rect 20732 5914 20760 8026
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20824 6798 20852 6938
rect 20916 6798 20944 8350
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21008 7206 21036 7822
rect 21100 7410 21128 9840
rect 21178 8392 21234 8401
rect 21376 8378 21404 9840
rect 21376 8350 21496 8378
rect 21178 8327 21234 8336
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21192 7206 21220 8327
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21284 6662 21312 7754
rect 21468 6798 21496 8350
rect 21652 7410 21680 9840
rect 21730 8528 21786 8537
rect 21730 8463 21786 8472
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21744 6662 21772 8463
rect 21928 6798 21956 9840
rect 22204 8650 22232 9840
rect 22480 8786 22508 9840
rect 22480 8758 22692 8786
rect 22204 8622 22600 8650
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21100 6458 21128 6598
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 22020 6186 22048 7890
rect 22155 7644 22463 7653
rect 22155 7642 22161 7644
rect 22217 7642 22241 7644
rect 22297 7642 22321 7644
rect 22377 7642 22401 7644
rect 22457 7642 22463 7644
rect 22217 7590 22219 7642
rect 22399 7590 22401 7642
rect 22155 7588 22161 7590
rect 22217 7588 22241 7590
rect 22297 7588 22321 7590
rect 22377 7588 22401 7590
rect 22457 7588 22463 7590
rect 22155 7579 22463 7588
rect 22572 7478 22600 8622
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22664 7410 22692 8758
rect 22756 7410 22784 9840
rect 22836 8220 22888 8226
rect 22836 8162 22888 8168
rect 22848 7546 22876 8162
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22155 6556 22463 6565
rect 22155 6554 22161 6556
rect 22217 6554 22241 6556
rect 22297 6554 22321 6556
rect 22377 6554 22401 6556
rect 22457 6554 22463 6556
rect 22217 6502 22219 6554
rect 22399 6502 22401 6554
rect 22155 6500 22161 6502
rect 22217 6500 22241 6502
rect 22297 6500 22321 6502
rect 22377 6500 22401 6502
rect 22457 6500 22463 6502
rect 22155 6491 22463 6500
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 22756 5778 22784 7210
rect 22834 7168 22890 7177
rect 22834 7103 22890 7112
rect 22848 6662 22876 7103
rect 22940 7002 22968 7686
rect 23032 7410 23060 9840
rect 23202 8120 23258 8129
rect 23124 8078 23202 8106
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23124 7290 23152 8078
rect 23202 8055 23258 8064
rect 23202 7848 23258 7857
rect 23202 7783 23258 7792
rect 23032 7262 23152 7290
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 23032 6186 23060 7262
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23124 7002 23152 7142
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23216 6798 23244 7783
rect 23308 7392 23336 9840
rect 23584 7834 23612 9840
rect 23860 8650 23888 9840
rect 24136 8650 24164 9840
rect 23860 8622 23980 8650
rect 24136 8622 24256 8650
rect 23756 7880 23808 7886
rect 23584 7806 23704 7834
rect 23756 7822 23808 7828
rect 23676 7410 23704 7806
rect 23572 7404 23624 7410
rect 23308 7364 23572 7392
rect 23572 7346 23624 7352
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 23308 7041 23336 7210
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23294 7032 23350 7041
rect 23294 6967 23350 6976
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23400 6730 23428 7142
rect 23676 7002 23704 7142
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23124 6458 23152 6598
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23768 6322 23796 7822
rect 23952 7392 23980 8622
rect 24124 7404 24176 7410
rect 23952 7364 24124 7392
rect 24228 7392 24256 8622
rect 24412 7478 24440 9840
rect 24492 8152 24544 8158
rect 24492 8094 24544 8100
rect 24504 7546 24532 8094
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24308 7404 24360 7410
rect 24228 7364 24308 7392
rect 24124 7346 24176 7352
rect 24308 7346 24360 7352
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23676 6202 23704 6258
rect 23860 6202 23888 7142
rect 24306 6896 24362 6905
rect 24306 6831 24362 6840
rect 23020 6180 23072 6186
rect 23676 6174 23888 6202
rect 24030 6216 24086 6225
rect 24320 6186 24348 6831
rect 24030 6151 24032 6160
rect 23020 6122 23072 6128
rect 24084 6151 24086 6160
rect 24308 6180 24360 6186
rect 24032 6122 24084 6128
rect 24308 6122 24360 6128
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 20626 5536 20682 5545
rect 20626 5471 20682 5480
rect 22155 5468 22463 5477
rect 22155 5466 22161 5468
rect 22217 5466 22241 5468
rect 22297 5466 22321 5468
rect 22377 5466 22401 5468
rect 22457 5466 22463 5468
rect 22217 5414 22219 5466
rect 22399 5414 22401 5466
rect 22155 5412 22161 5414
rect 22217 5412 22241 5414
rect 22297 5412 22321 5414
rect 22377 5412 22401 5414
rect 22457 5412 22463 5414
rect 22155 5403 22463 5412
rect 23216 5273 23244 5782
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23308 5302 23336 5714
rect 23400 5681 23428 6054
rect 23386 5672 23442 5681
rect 23386 5607 23442 5616
rect 24596 5574 24624 8026
rect 24688 7546 24716 9840
rect 24964 8294 24992 9840
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 25240 8226 25268 9840
rect 25228 8220 25280 8226
rect 25228 8162 25280 8168
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 25516 7392 25544 9840
rect 25792 8650 25820 9840
rect 26068 8786 26096 9840
rect 26068 8758 26280 8786
rect 25792 8622 26188 8650
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25688 8016 25740 8022
rect 25688 7958 25740 7964
rect 25700 7546 25728 7958
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25976 7410 26004 8230
rect 26056 8220 26108 8226
rect 26056 8162 26108 8168
rect 26068 7410 26096 8162
rect 26160 7478 26188 8622
rect 26252 7546 26280 8758
rect 26344 8650 26372 9840
rect 26620 8650 26648 9840
rect 26896 8786 26924 9840
rect 27172 8922 27200 9840
rect 27448 9058 27476 9840
rect 27448 9030 27660 9058
rect 27172 8894 27568 8922
rect 26896 8758 27476 8786
rect 26344 8622 26556 8650
rect 26620 8622 27292 8650
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26148 7472 26200 7478
rect 26148 7414 26200 7420
rect 25596 7404 25648 7410
rect 25516 7364 25596 7392
rect 25596 7346 25648 7352
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26528 7324 26556 8622
rect 27264 7478 27292 8622
rect 27448 7546 27476 8758
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 26700 7336 26752 7342
rect 26528 7296 26700 7324
rect 26700 7278 26752 7284
rect 26424 7268 26476 7274
rect 26424 7210 26476 7216
rect 27436 7268 27488 7274
rect 27540 7256 27568 8894
rect 27632 8158 27660 9030
rect 27620 8152 27672 8158
rect 27620 8094 27672 8100
rect 27724 8022 27752 9840
rect 28000 8650 28028 9840
rect 28276 8786 28304 9840
rect 28276 8758 28488 8786
rect 28000 8622 28396 8650
rect 27712 8016 27764 8022
rect 27712 7958 27764 7964
rect 28368 7478 28396 8622
rect 28460 8242 28488 8758
rect 28552 8378 28580 9840
rect 28828 8650 28856 9840
rect 28828 8622 28948 8650
rect 28552 8350 28856 8378
rect 28460 8214 28764 8242
rect 28540 8152 28592 8158
rect 28540 8094 28592 8100
rect 28356 7472 28408 7478
rect 28356 7414 28408 7420
rect 28552 7410 28580 8094
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28644 7410 28672 7958
rect 28736 7546 28764 8214
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28632 7404 28684 7410
rect 28632 7346 28684 7352
rect 27488 7228 27568 7256
rect 27436 7210 27488 7216
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 24688 6458 24716 7142
rect 25240 6458 25268 7142
rect 25884 7002 25912 7142
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 26436 6798 26464 7210
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 27068 7200 27120 7206
rect 27068 7142 27120 7148
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 28080 7200 28132 7206
rect 28080 7142 28132 7148
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28724 7200 28776 7206
rect 28724 7142 28776 7148
rect 26620 7002 26648 7142
rect 27080 7002 27108 7142
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 27068 6996 27120 7002
rect 27068 6938 27120 6944
rect 27356 6798 27384 7142
rect 27457 7100 27765 7109
rect 27457 7098 27463 7100
rect 27519 7098 27543 7100
rect 27599 7098 27623 7100
rect 27679 7098 27703 7100
rect 27759 7098 27765 7100
rect 27519 7046 27521 7098
rect 27701 7046 27703 7098
rect 27457 7044 27463 7046
rect 27519 7044 27543 7046
rect 27599 7044 27623 7046
rect 27679 7044 27703 7046
rect 27759 7044 27765 7046
rect 27457 7035 27765 7044
rect 27816 7002 27844 7142
rect 28092 7002 28120 7142
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 28080 6996 28132 7002
rect 28080 6938 28132 6944
rect 28184 6798 28212 7142
rect 28644 7002 28672 7142
rect 28632 6996 28684 7002
rect 28632 6938 28684 6944
rect 28736 6798 28764 7142
rect 28828 6798 28856 8350
rect 28920 7324 28948 8622
rect 29000 7336 29052 7342
rect 28920 7296 29000 7324
rect 29000 7278 29052 7284
rect 29104 7274 29132 9840
rect 29380 8650 29408 9840
rect 29380 8622 29500 8650
rect 29276 8356 29328 8362
rect 29276 8298 29328 8304
rect 29092 7268 29144 7274
rect 29092 7210 29144 7216
rect 29184 7200 29236 7206
rect 29184 7142 29236 7148
rect 29196 6798 29224 7142
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29288 6662 29316 8298
rect 29472 7478 29500 8622
rect 29656 8106 29684 9840
rect 29932 8514 29960 9840
rect 30208 8650 30236 9840
rect 30208 8622 30328 8650
rect 29932 8486 30236 8514
rect 30208 8294 30236 8486
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 29656 8078 30236 8106
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 29460 7472 29512 7478
rect 29460 7414 29512 7420
rect 30116 7274 30144 7822
rect 30208 7410 30236 8078
rect 30300 7478 30328 8622
rect 30484 7546 30512 9840
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30288 7472 30340 7478
rect 30288 7414 30340 7420
rect 30378 7440 30434 7449
rect 30196 7404 30248 7410
rect 30378 7375 30434 7384
rect 30196 7346 30248 7352
rect 30392 7274 30420 7375
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 30576 7206 30604 7958
rect 30668 7410 30696 8230
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30760 7342 30788 9840
rect 31036 8378 31064 9840
rect 31312 8650 31340 9840
rect 31588 8650 31616 9840
rect 31864 8650 31892 9840
rect 31312 8622 31432 8650
rect 31588 8622 31708 8650
rect 31864 8622 31984 8650
rect 31404 8378 31432 8622
rect 31036 8350 31340 8378
rect 31404 8350 31524 8378
rect 31116 7880 31168 7886
rect 31116 7822 31168 7828
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30852 7206 30880 7686
rect 31128 7206 31156 7822
rect 31312 7478 31340 8350
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31404 7546 31432 7822
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31300 7472 31352 7478
rect 31300 7414 31352 7420
rect 31496 7392 31524 8350
rect 31680 7546 31708 8622
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31852 7404 31904 7410
rect 31496 7364 31852 7392
rect 31852 7346 31904 7352
rect 31956 7342 31984 8622
rect 32140 8514 32168 9840
rect 32416 8650 32444 9840
rect 32416 8622 32628 8650
rect 32140 8486 32536 8514
rect 32034 7984 32090 7993
rect 32034 7919 32090 7928
rect 32048 7392 32076 7919
rect 32404 7812 32456 7818
rect 32404 7754 32456 7760
rect 32048 7364 32168 7392
rect 31944 7336 31996 7342
rect 31758 7304 31814 7313
rect 31944 7278 31996 7284
rect 31758 7239 31760 7248
rect 31812 7239 31814 7248
rect 31760 7210 31812 7216
rect 32140 7206 32168 7364
rect 32416 7206 32444 7754
rect 32508 7478 32536 8486
rect 32496 7472 32548 7478
rect 32496 7414 32548 7420
rect 32600 7324 32628 8622
rect 32692 7426 32720 9840
rect 32968 7732 32996 9840
rect 32968 7704 33180 7732
rect 32758 7644 33066 7653
rect 32758 7642 32764 7644
rect 32820 7642 32844 7644
rect 32900 7642 32924 7644
rect 32980 7642 33004 7644
rect 33060 7642 33066 7644
rect 32820 7590 32822 7642
rect 33002 7590 33004 7642
rect 32758 7588 32764 7590
rect 32820 7588 32844 7590
rect 32900 7588 32924 7590
rect 32980 7588 33004 7590
rect 33060 7588 33066 7590
rect 32758 7579 33066 7588
rect 32772 7540 32824 7546
rect 32772 7482 32824 7488
rect 32784 7426 32812 7482
rect 33152 7460 33180 7704
rect 32692 7398 32812 7426
rect 33060 7432 33180 7460
rect 32864 7336 32916 7342
rect 32600 7296 32864 7324
rect 32864 7278 32916 7284
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 30012 7200 30064 7206
rect 30012 7142 30064 7148
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 31116 7200 31168 7206
rect 31116 7142 31168 7148
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 29748 6798 29776 7142
rect 30024 6798 30052 7142
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 27160 6656 27212 6662
rect 27528 6656 27580 6662
rect 27160 6598 27212 6604
rect 27356 6616 27528 6644
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24780 5817 24808 6122
rect 24766 5808 24822 5817
rect 25516 5778 25544 6598
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 24766 5743 24822 5752
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 23296 5296 23348 5302
rect 23202 5264 23258 5273
rect 23296 5238 23348 5244
rect 23202 5199 23258 5208
rect 25608 5098 25636 6394
rect 25976 6118 26004 6598
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 26344 5370 26372 6598
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26712 5234 26740 6598
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 25596 5092 25648 5098
rect 25596 5034 25648 5040
rect 19800 4752 19852 4758
rect 6828 4694 6880 4700
rect 14186 4720 14242 4729
rect 27080 4729 27108 6598
rect 27172 5914 27200 6598
rect 27160 5908 27212 5914
rect 27160 5850 27212 5856
rect 27356 4826 27384 6616
rect 27528 6598 27580 6604
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28540 6656 28592 6662
rect 28540 6598 28592 6604
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 27457 6012 27765 6021
rect 27457 6010 27463 6012
rect 27519 6010 27543 6012
rect 27599 6010 27623 6012
rect 27679 6010 27703 6012
rect 27759 6010 27765 6012
rect 27519 5958 27521 6010
rect 27701 5958 27703 6010
rect 27457 5956 27463 5958
rect 27519 5956 27543 5958
rect 27599 5956 27623 5958
rect 27679 5956 27703 5958
rect 27759 5956 27765 5958
rect 27457 5947 27765 5956
rect 28000 5166 28028 6598
rect 28552 6186 28580 6598
rect 29104 6458 29132 6598
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 28540 6180 28592 6186
rect 28540 6122 28592 6128
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 30024 5030 30052 6598
rect 30300 5846 30328 6598
rect 31760 6452 31812 6458
rect 31760 6394 31812 6400
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 30288 5840 30340 5846
rect 30288 5782 30340 5788
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 27457 4924 27765 4933
rect 27457 4922 27463 4924
rect 27519 4922 27543 4924
rect 27599 4922 27623 4924
rect 27679 4922 27703 4924
rect 27759 4922 27765 4924
rect 27519 4870 27521 4922
rect 27701 4870 27703 4922
rect 27457 4868 27463 4870
rect 27519 4868 27543 4870
rect 27599 4868 27623 4870
rect 27679 4868 27703 4870
rect 27759 4868 27765 4870
rect 27457 4859 27765 4868
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 19800 4694 19852 4700
rect 27066 4720 27122 4729
rect 14186 4655 14242 4664
rect 27066 4655 27122 4664
rect 11552 4380 11860 4389
rect 11552 4378 11558 4380
rect 11614 4378 11638 4380
rect 11694 4378 11718 4380
rect 11774 4378 11798 4380
rect 11854 4378 11860 4380
rect 11614 4326 11616 4378
rect 11796 4326 11798 4378
rect 11552 4324 11558 4326
rect 11614 4324 11638 4326
rect 11694 4324 11718 4326
rect 11774 4324 11798 4326
rect 11854 4324 11860 4326
rect 11552 4315 11860 4324
rect 22155 4380 22463 4389
rect 22155 4378 22161 4380
rect 22217 4378 22241 4380
rect 22297 4378 22321 4380
rect 22377 4378 22401 4380
rect 22457 4378 22463 4380
rect 22217 4326 22219 4378
rect 22399 4326 22401 4378
rect 22155 4324 22161 4326
rect 22217 4324 22241 4326
rect 22297 4324 22321 4326
rect 22377 4324 22401 4326
rect 22457 4324 22463 4326
rect 22155 4315 22463 4324
rect 6251 3836 6559 3845
rect 6251 3834 6257 3836
rect 6313 3834 6337 3836
rect 6393 3834 6417 3836
rect 6473 3834 6497 3836
rect 6553 3834 6559 3836
rect 6313 3782 6315 3834
rect 6495 3782 6497 3834
rect 6251 3780 6257 3782
rect 6313 3780 6337 3782
rect 6393 3780 6417 3782
rect 6473 3780 6497 3782
rect 6553 3780 6559 3782
rect 6251 3771 6559 3780
rect 16854 3836 17162 3845
rect 16854 3834 16860 3836
rect 16916 3834 16940 3836
rect 16996 3834 17020 3836
rect 17076 3834 17100 3836
rect 17156 3834 17162 3836
rect 16916 3782 16918 3834
rect 17098 3782 17100 3834
rect 16854 3780 16860 3782
rect 16916 3780 16940 3782
rect 16996 3780 17020 3782
rect 17076 3780 17100 3782
rect 17156 3780 17162 3782
rect 16854 3771 17162 3780
rect 27457 3836 27765 3845
rect 27457 3834 27463 3836
rect 27519 3834 27543 3836
rect 27599 3834 27623 3836
rect 27679 3834 27703 3836
rect 27759 3834 27765 3836
rect 27519 3782 27521 3834
rect 27701 3782 27703 3834
rect 27457 3780 27463 3782
rect 27519 3780 27543 3782
rect 27599 3780 27623 3782
rect 27679 3780 27703 3782
rect 27759 3780 27765 3782
rect 27457 3771 27765 3780
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 2650 5672 3470
rect 24872 3318 25268 3346
rect 11552 3292 11860 3301
rect 11552 3290 11558 3292
rect 11614 3290 11638 3292
rect 11694 3290 11718 3292
rect 11774 3290 11798 3292
rect 11854 3290 11860 3292
rect 11614 3238 11616 3290
rect 11796 3238 11798 3290
rect 11552 3236 11558 3238
rect 11614 3236 11638 3238
rect 11694 3236 11718 3238
rect 11774 3236 11798 3238
rect 11854 3236 11860 3238
rect 11552 3227 11860 3236
rect 22155 3292 22463 3301
rect 22155 3290 22161 3292
rect 22217 3290 22241 3292
rect 22297 3290 22321 3292
rect 22377 3290 22401 3292
rect 22457 3290 22463 3292
rect 22217 3238 22219 3290
rect 22399 3238 22401 3290
rect 22155 3236 22161 3238
rect 22217 3236 22241 3238
rect 22297 3236 22321 3238
rect 22377 3236 22401 3238
rect 22457 3236 22463 3238
rect 22155 3227 22463 3236
rect 24872 3058 24900 3318
rect 25240 3194 25268 3318
rect 24952 3188 25004 3194
rect 25228 3188 25280 3194
rect 25004 3148 25176 3176
rect 24952 3130 25004 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 6251 2748 6559 2757
rect 6251 2746 6257 2748
rect 6313 2746 6337 2748
rect 6393 2746 6417 2748
rect 6473 2746 6497 2748
rect 6553 2746 6559 2748
rect 6313 2694 6315 2746
rect 6495 2694 6497 2746
rect 6251 2692 6257 2694
rect 6313 2692 6337 2694
rect 6393 2692 6417 2694
rect 6473 2692 6497 2694
rect 6553 2692 6559 2694
rect 6251 2683 6559 2692
rect 16684 2650 16712 2994
rect 16854 2748 17162 2757
rect 16854 2746 16860 2748
rect 16916 2746 16940 2748
rect 16996 2746 17020 2748
rect 17076 2746 17100 2748
rect 17156 2746 17162 2748
rect 16916 2694 16918 2746
rect 17098 2694 17100 2746
rect 16854 2692 16860 2694
rect 16916 2692 16940 2694
rect 16996 2692 17020 2694
rect 17076 2692 17100 2694
rect 17156 2692 17162 2694
rect 16854 2683 17162 2692
rect 18616 2650 18644 2994
rect 20732 2650 20760 2994
rect 22664 2650 22692 2994
rect 24964 2650 24992 2994
rect 25044 2916 25096 2922
rect 25148 2904 25176 3148
rect 25228 3130 25280 3136
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25228 2916 25280 2922
rect 25148 2876 25228 2904
rect 25044 2858 25096 2864
rect 25228 2858 25280 2864
rect 25056 2802 25084 2858
rect 25332 2802 25360 2926
rect 30392 2854 30420 6326
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 25056 2774 25360 2802
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 27457 2748 27765 2757
rect 27457 2746 27463 2748
rect 27519 2746 27543 2748
rect 27599 2746 27623 2748
rect 27679 2746 27703 2748
rect 27759 2746 27765 2748
rect 27519 2694 27521 2746
rect 27701 2694 27703 2746
rect 27457 2692 27463 2694
rect 27519 2692 27543 2694
rect 27599 2692 27623 2694
rect 27679 2692 27703 2694
rect 27759 2692 27765 2694
rect 27457 2683 27765 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 30852 2582 30880 3878
rect 31772 3058 31800 6394
rect 32324 6186 32352 7142
rect 33060 6798 33088 7432
rect 33244 6914 33272 9840
rect 33324 8560 33376 8566
rect 33324 8502 33376 8508
rect 33336 7342 33364 8502
rect 33324 7336 33376 7342
rect 33324 7278 33376 7284
rect 33416 7336 33468 7342
rect 33416 7278 33468 7284
rect 33244 6886 33364 6914
rect 33336 6798 33364 6886
rect 33048 6792 33100 6798
rect 33324 6792 33376 6798
rect 33048 6734 33100 6740
rect 33230 6760 33286 6769
rect 33324 6734 33376 6740
rect 33230 6695 33286 6704
rect 33244 6662 33272 6695
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 32758 6556 33066 6565
rect 32758 6554 32764 6556
rect 32820 6554 32844 6556
rect 32900 6554 32924 6556
rect 32980 6554 33004 6556
rect 33060 6554 33066 6556
rect 32820 6502 32822 6554
rect 33002 6502 33004 6554
rect 32758 6500 32764 6502
rect 32820 6500 32844 6502
rect 32900 6500 32924 6502
rect 32980 6500 33004 6502
rect 33060 6500 33066 6502
rect 32758 6491 33066 6500
rect 32312 6180 32364 6186
rect 32312 6122 32364 6128
rect 32758 5468 33066 5477
rect 32758 5466 32764 5468
rect 32820 5466 32844 5468
rect 32900 5466 32924 5468
rect 32980 5466 33004 5468
rect 33060 5466 33066 5468
rect 32820 5414 32822 5466
rect 33002 5414 33004 5466
rect 32758 5412 32764 5414
rect 32820 5412 32844 5414
rect 32900 5412 32924 5414
rect 32980 5412 33004 5414
rect 33060 5412 33066 5414
rect 32758 5403 33066 5412
rect 32758 4380 33066 4389
rect 32758 4378 32764 4380
rect 32820 4378 32844 4380
rect 32900 4378 32924 4380
rect 32980 4378 33004 4380
rect 33060 4378 33066 4380
rect 32820 4326 32822 4378
rect 33002 4326 33004 4378
rect 32758 4324 32764 4326
rect 32820 4324 32844 4326
rect 32900 4324 32924 4326
rect 32980 4324 33004 4326
rect 33060 4324 33066 4326
rect 32758 4315 33066 4324
rect 32758 3292 33066 3301
rect 32758 3290 32764 3292
rect 32820 3290 32844 3292
rect 32900 3290 32924 3292
rect 32980 3290 33004 3292
rect 33060 3290 33066 3292
rect 32820 3238 32822 3290
rect 33002 3238 33004 3290
rect 32758 3236 32764 3238
rect 32820 3236 32844 3238
rect 32900 3236 32924 3238
rect 32980 3236 33004 3238
rect 33060 3236 33066 3238
rect 32758 3227 33066 3236
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 33428 2802 33456 7278
rect 33520 6914 33548 9840
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33612 7274 33640 8434
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33704 7546 33732 8366
rect 33796 7546 33824 9840
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33520 6886 33640 6914
rect 33612 6798 33640 6886
rect 34072 6866 34100 9840
rect 34348 7546 34376 9840
rect 34336 7540 34388 7546
rect 34336 7482 34388 7488
rect 34624 7478 34652 9840
rect 34900 8514 34928 9840
rect 34900 8486 35112 8514
rect 34612 7472 34664 7478
rect 34612 7414 34664 7420
rect 34152 7404 34204 7410
rect 34152 7346 34204 7352
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33520 5137 33548 6598
rect 33506 5128 33562 5137
rect 33506 5063 33562 5072
rect 33508 3052 33560 3058
rect 33508 2994 33560 3000
rect 33244 2774 33456 2802
rect 33244 2650 33272 2774
rect 33520 2650 33548 2994
rect 33704 2922 33732 6734
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33796 6361 33824 6598
rect 33782 6352 33838 6361
rect 33782 6287 33838 6296
rect 33692 2916 33744 2922
rect 33692 2858 33744 2864
rect 34164 2650 34192 7346
rect 34428 7336 34480 7342
rect 34428 7278 34480 7284
rect 34440 3738 34468 7278
rect 34796 7268 34848 7274
rect 34796 7210 34848 7216
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 33232 2644 33284 2650
rect 33232 2586 33284 2592
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 34808 2582 34836 7210
rect 35084 7206 35112 8486
rect 35072 7200 35124 7206
rect 35072 7142 35124 7148
rect 35176 6866 35204 9840
rect 35452 8650 35480 9840
rect 35452 8622 35664 8650
rect 35636 7546 35664 8622
rect 35624 7540 35676 7546
rect 35624 7482 35676 7488
rect 35728 6866 35756 9840
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 35716 6860 35768 6866
rect 35716 6802 35768 6808
rect 35348 6724 35400 6730
rect 35348 6666 35400 6672
rect 35900 6724 35952 6730
rect 35900 6666 35952 6672
rect 35360 2650 35388 6666
rect 35912 3942 35940 6666
rect 36004 6662 36032 9840
rect 36280 8514 36308 9840
rect 36280 8486 36492 8514
rect 36084 7404 36136 7410
rect 36084 7346 36136 7352
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 30840 2576 30892 2582
rect 30840 2518 30892 2524
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 29828 2508 29880 2514
rect 29828 2450 29880 2456
rect 1124 2440 1176 2446
rect 1124 2382 1176 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 1136 160 1164 2382
rect 1688 2106 1716 2382
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 3252 160 3280 2382
rect 4080 2106 4108 2382
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 1122 -300 1178 160
rect 3238 -300 3294 160
rect 5354 82 5410 160
rect 5460 82 5488 2382
rect 5354 54 5488 82
rect 7470 82 7526 160
rect 7576 82 7604 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 2106 7788 2246
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 9692 1442 9720 2382
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9876 2106 9904 2246
rect 11552 2204 11860 2213
rect 11552 2202 11558 2204
rect 11614 2202 11638 2204
rect 11694 2202 11718 2204
rect 11774 2202 11798 2204
rect 11854 2202 11860 2204
rect 11614 2150 11616 2202
rect 11796 2150 11798 2202
rect 11552 2148 11558 2150
rect 11614 2148 11638 2150
rect 11694 2148 11718 2150
rect 11774 2148 11798 2150
rect 11854 2148 11860 2150
rect 11552 2139 11860 2148
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9600 1414 9720 1442
rect 9600 160 9628 1414
rect 7470 54 7604 82
rect 5354 -300 5410 54
rect 7470 -300 7526 54
rect 9586 -300 9642 160
rect 11702 82 11758 160
rect 11992 82 12020 2382
rect 13832 160 13860 2382
rect 11702 54 12020 82
rect 11702 -300 11758 54
rect 13818 -300 13874 160
rect 15934 82 15990 160
rect 16224 82 16252 2382
rect 15934 54 16252 82
rect 18050 82 18106 160
rect 18340 82 18368 2382
rect 18050 54 18368 82
rect 20166 82 20222 160
rect 20456 82 20484 2382
rect 22155 2204 22463 2213
rect 22155 2202 22161 2204
rect 22217 2202 22241 2204
rect 22297 2202 22321 2204
rect 22377 2202 22401 2204
rect 22457 2202 22463 2204
rect 22217 2150 22219 2202
rect 22399 2150 22401 2202
rect 22155 2148 22161 2150
rect 22217 2148 22241 2150
rect 22297 2148 22321 2150
rect 22377 2148 22401 2150
rect 22457 2148 22463 2150
rect 22155 2139 22463 2148
rect 22296 190 22416 218
rect 22296 160 22324 190
rect 20166 54 20484 82
rect 15934 -300 15990 54
rect 18050 -300 18106 54
rect 20166 -300 20222 54
rect 22282 -300 22338 160
rect 22388 82 22416 190
rect 22572 82 22600 2382
rect 22388 54 22600 82
rect 24398 82 24454 160
rect 24688 82 24716 2382
rect 26620 1306 26648 2382
rect 26792 2304 26844 2310
rect 26792 2246 26844 2252
rect 26804 1698 26832 2246
rect 26792 1692 26844 1698
rect 26792 1634 26844 1640
rect 26528 1278 26648 1306
rect 26528 160 26556 1278
rect 24398 54 24716 82
rect 24398 -300 24454 54
rect 26514 -300 26570 160
rect 28630 82 28686 160
rect 28736 82 28764 2382
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 28828 1630 28856 2246
rect 29840 2106 29868 2450
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 29828 2100 29880 2106
rect 29828 2042 29880 2048
rect 28816 1624 28868 1630
rect 28816 1566 28868 1572
rect 28630 54 28764 82
rect 30746 82 30802 160
rect 31036 82 31064 2382
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 32692 2038 32720 2246
rect 32758 2204 33066 2213
rect 32758 2202 32764 2204
rect 32820 2202 32844 2204
rect 32900 2202 32924 2204
rect 32980 2202 33004 2204
rect 33060 2202 33066 2204
rect 32820 2150 32822 2202
rect 33002 2150 33004 2202
rect 32758 2148 32764 2150
rect 32820 2148 32844 2150
rect 32900 2148 32924 2150
rect 32980 2148 33004 2150
rect 33060 2148 33066 2150
rect 32758 2139 33066 2148
rect 32680 2032 32732 2038
rect 32680 1974 32732 1980
rect 33336 1834 33364 2382
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 33428 1970 33456 2246
rect 33416 1964 33468 1970
rect 33416 1906 33468 1912
rect 33324 1828 33376 1834
rect 33324 1770 33376 1776
rect 33612 1426 33640 2382
rect 33980 1902 34008 2382
rect 34440 2106 34468 2382
rect 34428 2100 34480 2106
rect 34428 2042 34480 2048
rect 34520 2100 34572 2106
rect 34520 2042 34572 2048
rect 33968 1896 34020 1902
rect 33968 1838 34020 1844
rect 34532 1630 34560 2042
rect 34520 1624 34572 1630
rect 34520 1566 34572 1572
rect 32864 1420 32916 1426
rect 32864 1362 32916 1368
rect 33600 1420 33652 1426
rect 33600 1362 33652 1368
rect 32876 160 32904 1362
rect 30746 54 31064 82
rect 28630 -300 28686 54
rect 30746 -300 30802 54
rect 32862 -300 32918 160
rect 34978 82 35034 160
rect 35268 82 35296 2382
rect 36096 2106 36124 7346
rect 36464 7206 36492 8486
rect 36452 7200 36504 7206
rect 36452 7142 36504 7148
rect 36556 6914 36584 9840
rect 36832 8514 36860 9840
rect 36832 8486 37044 8514
rect 37016 7478 37044 8486
rect 37004 7472 37056 7478
rect 37004 7414 37056 7420
rect 36912 7404 36964 7410
rect 36912 7346 36964 7352
rect 36556 6886 36676 6914
rect 36648 6662 36676 6886
rect 36728 6792 36780 6798
rect 36728 6734 36780 6740
rect 36636 6656 36688 6662
rect 36636 6598 36688 6604
rect 36740 6458 36768 6734
rect 36728 6452 36780 6458
rect 36728 6394 36780 6400
rect 36820 2372 36872 2378
rect 36820 2314 36872 2320
rect 36832 2106 36860 2314
rect 36084 2100 36136 2106
rect 36084 2042 36136 2048
rect 36820 2100 36872 2106
rect 36820 2042 36872 2048
rect 36924 1698 36952 7346
rect 37108 6866 37136 9840
rect 37384 8378 37412 9840
rect 37384 8350 37596 8378
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37384 6914 37412 7346
rect 37568 6934 37596 8350
rect 37292 6886 37412 6914
rect 37556 6928 37608 6934
rect 37096 6860 37148 6866
rect 37096 6802 37148 6808
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 37016 6458 37044 6666
rect 37004 6452 37056 6458
rect 37004 6394 37056 6400
rect 37292 3058 37320 6886
rect 37556 6870 37608 6876
rect 37660 6662 37688 9840
rect 37832 7404 37884 7410
rect 37832 7346 37884 7352
rect 37740 6724 37792 6730
rect 37740 6666 37792 6672
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37752 2650 37780 6666
rect 37844 3210 37872 7346
rect 37936 6458 37964 9840
rect 38212 8378 38240 9840
rect 38212 8350 38424 8378
rect 38060 7100 38368 7109
rect 38060 7098 38066 7100
rect 38122 7098 38146 7100
rect 38202 7098 38226 7100
rect 38282 7098 38306 7100
rect 38362 7098 38368 7100
rect 38122 7046 38124 7098
rect 38304 7046 38306 7098
rect 38060 7044 38066 7046
rect 38122 7044 38146 7046
rect 38202 7044 38226 7046
rect 38282 7044 38306 7046
rect 38362 7044 38368 7046
rect 38060 7035 38368 7044
rect 38292 6860 38344 6866
rect 38292 6802 38344 6808
rect 37924 6452 37976 6458
rect 37924 6394 37976 6400
rect 38304 6390 38332 6802
rect 38396 6662 38424 8350
rect 38488 6730 38516 9840
rect 38764 8514 38792 9840
rect 38764 8486 38976 8514
rect 38948 7478 38976 8486
rect 38936 7472 38988 7478
rect 38936 7414 38988 7420
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 38568 7336 38620 7342
rect 38568 7278 38620 7284
rect 38476 6724 38528 6730
rect 38476 6666 38528 6672
rect 38384 6656 38436 6662
rect 38384 6598 38436 6604
rect 38292 6384 38344 6390
rect 38292 6326 38344 6332
rect 38060 6012 38368 6021
rect 38060 6010 38066 6012
rect 38122 6010 38146 6012
rect 38202 6010 38226 6012
rect 38282 6010 38306 6012
rect 38362 6010 38368 6012
rect 38122 5958 38124 6010
rect 38304 5958 38306 6010
rect 38060 5956 38066 5958
rect 38122 5956 38146 5958
rect 38202 5956 38226 5958
rect 38282 5956 38306 5958
rect 38362 5956 38368 5958
rect 38060 5947 38368 5956
rect 38060 4924 38368 4933
rect 38060 4922 38066 4924
rect 38122 4922 38146 4924
rect 38202 4922 38226 4924
rect 38282 4922 38306 4924
rect 38362 4922 38368 4924
rect 38122 4870 38124 4922
rect 38304 4870 38306 4922
rect 38060 4868 38066 4870
rect 38122 4868 38146 4870
rect 38202 4868 38226 4870
rect 38282 4868 38306 4870
rect 38362 4868 38368 4870
rect 38060 4859 38368 4868
rect 38060 3836 38368 3845
rect 38060 3834 38066 3836
rect 38122 3834 38146 3836
rect 38202 3834 38226 3836
rect 38282 3834 38306 3836
rect 38362 3834 38368 3836
rect 38122 3782 38124 3834
rect 38304 3782 38306 3834
rect 38060 3780 38066 3782
rect 38122 3780 38146 3782
rect 38202 3780 38226 3782
rect 38282 3780 38306 3782
rect 38362 3780 38368 3782
rect 38060 3771 38368 3780
rect 37844 3182 37964 3210
rect 38580 3194 38608 7278
rect 38660 7268 38712 7274
rect 38660 7210 38712 7216
rect 38672 6390 38700 7210
rect 38660 6384 38712 6390
rect 38660 6326 38712 6332
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 37844 2650 37872 2994
rect 37936 2990 37964 3182
rect 38568 3188 38620 3194
rect 38568 3130 38620 3136
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 38060 2748 38368 2757
rect 38060 2746 38066 2748
rect 38122 2746 38146 2748
rect 38202 2746 38226 2748
rect 38282 2746 38306 2748
rect 38362 2746 38368 2748
rect 38122 2694 38124 2746
rect 38304 2694 38306 2746
rect 38060 2692 38066 2694
rect 38122 2692 38146 2694
rect 38202 2692 38226 2694
rect 38282 2692 38306 2694
rect 38362 2692 38368 2694
rect 38060 2683 38368 2692
rect 38764 2650 38792 7346
rect 39040 6798 39068 9840
rect 39316 7528 39344 9840
rect 39488 7540 39540 7546
rect 39316 7500 39488 7528
rect 39488 7482 39540 7488
rect 39120 7200 39172 7206
rect 39120 7142 39172 7148
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 39028 6792 39080 6798
rect 39028 6734 39080 6740
rect 38856 3194 38884 6734
rect 38936 6724 38988 6730
rect 38936 6666 38988 6672
rect 38844 3188 38896 3194
rect 38844 3130 38896 3136
rect 37740 2644 37792 2650
rect 37740 2586 37792 2592
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 37108 2514 37228 2530
rect 37108 2508 37240 2514
rect 37108 2502 37188 2508
rect 36912 1692 36964 1698
rect 36912 1634 36964 1640
rect 37108 160 37136 2502
rect 37188 2450 37240 2456
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37476 2106 37504 2382
rect 38948 2378 38976 6666
rect 39132 6458 39160 7142
rect 39592 6866 39620 9840
rect 43361 7644 43669 7653
rect 43361 7642 43367 7644
rect 43423 7642 43447 7644
rect 43503 7642 43527 7644
rect 43583 7642 43607 7644
rect 43663 7642 43669 7644
rect 43423 7590 43425 7642
rect 43605 7590 43607 7642
rect 43361 7588 43367 7590
rect 43423 7588 43447 7590
rect 43503 7588 43527 7590
rect 43583 7588 43607 7590
rect 43663 7588 43669 7590
rect 43361 7579 43669 7588
rect 40500 7404 40552 7410
rect 40500 7346 40552 7352
rect 39580 6860 39632 6866
rect 39580 6802 39632 6808
rect 39948 6724 40000 6730
rect 39948 6666 40000 6672
rect 39120 6452 39172 6458
rect 39120 6394 39172 6400
rect 39960 2650 39988 6666
rect 40512 2650 40540 7346
rect 41328 6724 41380 6730
rect 41328 6666 41380 6672
rect 41340 2650 41368 6666
rect 43361 6556 43669 6565
rect 43361 6554 43367 6556
rect 43423 6554 43447 6556
rect 43503 6554 43527 6556
rect 43583 6554 43607 6556
rect 43663 6554 43669 6556
rect 43423 6502 43425 6554
rect 43605 6502 43607 6554
rect 43361 6500 43367 6502
rect 43423 6500 43447 6502
rect 43503 6500 43527 6502
rect 43583 6500 43607 6502
rect 43663 6500 43669 6502
rect 43361 6491 43669 6500
rect 43361 5468 43669 5477
rect 43361 5466 43367 5468
rect 43423 5466 43447 5468
rect 43503 5466 43527 5468
rect 43583 5466 43607 5468
rect 43663 5466 43669 5468
rect 43423 5414 43425 5466
rect 43605 5414 43607 5466
rect 43361 5412 43367 5414
rect 43423 5412 43447 5414
rect 43503 5412 43527 5414
rect 43583 5412 43607 5414
rect 43663 5412 43669 5414
rect 43361 5403 43669 5412
rect 43361 4380 43669 4389
rect 43361 4378 43367 4380
rect 43423 4378 43447 4380
rect 43503 4378 43527 4380
rect 43583 4378 43607 4380
rect 43663 4378 43669 4380
rect 43423 4326 43425 4378
rect 43605 4326 43607 4378
rect 43361 4324 43367 4326
rect 43423 4324 43447 4326
rect 43503 4324 43527 4326
rect 43583 4324 43607 4326
rect 43663 4324 43669 4326
rect 43361 4315 43669 4324
rect 43361 3292 43669 3301
rect 43361 3290 43367 3292
rect 43423 3290 43447 3292
rect 43503 3290 43527 3292
rect 43583 3290 43607 3292
rect 43663 3290 43669 3292
rect 43423 3238 43425 3290
rect 43605 3238 43607 3290
rect 43361 3236 43367 3238
rect 43423 3236 43447 3238
rect 43503 3236 43527 3238
rect 43583 3236 43607 3238
rect 43663 3236 43669 3238
rect 43361 3227 43669 3236
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 40500 2644 40552 2650
rect 40500 2586 40552 2592
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 39488 2440 39540 2446
rect 39488 2382 39540 2388
rect 41604 2440 41656 2446
rect 41604 2382 41656 2388
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 38936 2372 38988 2378
rect 38936 2314 38988 2320
rect 37464 2100 37516 2106
rect 37464 2042 37516 2048
rect 39224 190 39344 218
rect 39224 160 39252 190
rect 34978 54 35296 82
rect 34978 -300 35034 54
rect 37094 -300 37150 160
rect 39210 -300 39266 160
rect 39316 82 39344 190
rect 39500 82 39528 2382
rect 41616 1442 41644 2382
rect 41340 1414 41644 1442
rect 41340 160 41368 1414
rect 39316 54 39528 82
rect 41326 -300 41382 160
rect 43180 82 43208 2382
rect 43361 2204 43669 2213
rect 43361 2202 43367 2204
rect 43423 2202 43447 2204
rect 43503 2202 43527 2204
rect 43583 2202 43607 2204
rect 43663 2202 43669 2204
rect 43423 2150 43425 2202
rect 43605 2150 43607 2202
rect 43361 2148 43367 2150
rect 43423 2148 43447 2150
rect 43503 2148 43527 2150
rect 43583 2148 43607 2150
rect 43663 2148 43669 2150
rect 43361 2139 43669 2148
rect 43442 82 43498 160
rect 43180 54 43498 82
rect 43442 -300 43498 54
<< via2 >>
rect 6257 7098 6313 7100
rect 6337 7098 6393 7100
rect 6417 7098 6473 7100
rect 6497 7098 6553 7100
rect 6257 7046 6303 7098
rect 6303 7046 6313 7098
rect 6337 7046 6367 7098
rect 6367 7046 6379 7098
rect 6379 7046 6393 7098
rect 6417 7046 6431 7098
rect 6431 7046 6443 7098
rect 6443 7046 6473 7098
rect 6497 7046 6507 7098
rect 6507 7046 6553 7098
rect 6257 7044 6313 7046
rect 6337 7044 6393 7046
rect 6417 7044 6473 7046
rect 6497 7044 6553 7046
rect 6182 6724 6238 6760
rect 6182 6704 6184 6724
rect 6184 6704 6236 6724
rect 6236 6704 6238 6724
rect 5814 6160 5870 6216
rect 6257 6010 6313 6012
rect 6337 6010 6393 6012
rect 6417 6010 6473 6012
rect 6497 6010 6553 6012
rect 6257 5958 6303 6010
rect 6303 5958 6313 6010
rect 6337 5958 6367 6010
rect 6367 5958 6379 6010
rect 6379 5958 6393 6010
rect 6417 5958 6431 6010
rect 6431 5958 6443 6010
rect 6443 5958 6473 6010
rect 6497 5958 6507 6010
rect 6507 5958 6553 6010
rect 6257 5956 6313 5958
rect 6337 5956 6393 5958
rect 6417 5956 6473 5958
rect 6497 5956 6553 5958
rect 6257 4922 6313 4924
rect 6337 4922 6393 4924
rect 6417 4922 6473 4924
rect 6497 4922 6553 4924
rect 6257 4870 6303 4922
rect 6303 4870 6313 4922
rect 6337 4870 6367 4922
rect 6367 4870 6379 4922
rect 6379 4870 6393 4922
rect 6417 4870 6431 4922
rect 6431 4870 6443 4922
rect 6443 4870 6473 4922
rect 6497 4870 6507 4922
rect 6507 4870 6553 4922
rect 6257 4868 6313 4870
rect 6337 4868 6393 4870
rect 6417 4868 6473 4870
rect 6497 4868 6553 4870
rect 9678 5616 9734 5672
rect 10598 5208 10654 5264
rect 11558 7642 11614 7644
rect 11638 7642 11694 7644
rect 11718 7642 11774 7644
rect 11798 7642 11854 7644
rect 11558 7590 11604 7642
rect 11604 7590 11614 7642
rect 11638 7590 11668 7642
rect 11668 7590 11680 7642
rect 11680 7590 11694 7642
rect 11718 7590 11732 7642
rect 11732 7590 11744 7642
rect 11744 7590 11774 7642
rect 11798 7590 11808 7642
rect 11808 7590 11854 7642
rect 11558 7588 11614 7590
rect 11638 7588 11694 7590
rect 11718 7588 11774 7590
rect 11798 7588 11854 7590
rect 11610 6976 11666 7032
rect 12162 8200 12218 8256
rect 11558 6554 11614 6556
rect 11638 6554 11694 6556
rect 11718 6554 11774 6556
rect 11798 6554 11854 6556
rect 11558 6502 11604 6554
rect 11604 6502 11614 6554
rect 11638 6502 11668 6554
rect 11668 6502 11680 6554
rect 11680 6502 11694 6554
rect 11718 6502 11732 6554
rect 11732 6502 11744 6554
rect 11744 6502 11774 6554
rect 11798 6502 11808 6554
rect 11808 6502 11854 6554
rect 11558 6500 11614 6502
rect 11638 6500 11694 6502
rect 11718 6500 11774 6502
rect 11798 6500 11854 6502
rect 11978 6568 12034 6624
rect 13726 8336 13782 8392
rect 12346 5480 12402 5536
rect 11558 5466 11614 5468
rect 11638 5466 11694 5468
rect 11718 5466 11774 5468
rect 11798 5466 11854 5468
rect 11558 5414 11604 5466
rect 11604 5414 11614 5466
rect 11638 5414 11668 5466
rect 11668 5414 11680 5466
rect 11680 5414 11694 5466
rect 11718 5414 11732 5466
rect 11732 5414 11744 5466
rect 11744 5414 11774 5466
rect 11798 5414 11808 5466
rect 11808 5414 11854 5466
rect 11558 5412 11614 5414
rect 11638 5412 11694 5414
rect 11718 5412 11774 5414
rect 11798 5412 11854 5414
rect 14278 6704 14334 6760
rect 14370 6432 14426 6488
rect 15106 8472 15162 8528
rect 15198 6316 15254 6352
rect 15198 6296 15200 6316
rect 15200 6296 15252 6316
rect 15252 6296 15254 6316
rect 15290 5752 15346 5808
rect 15934 7792 15990 7848
rect 16486 8064 16542 8120
rect 16578 6976 16634 7032
rect 17314 7928 17370 7984
rect 16860 7098 16916 7100
rect 16940 7098 16996 7100
rect 17020 7098 17076 7100
rect 17100 7098 17156 7100
rect 16860 7046 16906 7098
rect 16906 7046 16916 7098
rect 16940 7046 16970 7098
rect 16970 7046 16982 7098
rect 16982 7046 16996 7098
rect 17020 7046 17034 7098
rect 17034 7046 17046 7098
rect 17046 7046 17076 7098
rect 17100 7046 17110 7098
rect 17110 7046 17156 7098
rect 16860 7044 16916 7046
rect 16940 7044 16996 7046
rect 17020 7044 17076 7046
rect 17100 7044 17156 7046
rect 17406 7248 17462 7304
rect 17314 7112 17370 7168
rect 17774 7928 17830 7984
rect 18326 7384 18382 7440
rect 18418 6976 18474 7032
rect 18418 6432 18474 6488
rect 16860 6010 16916 6012
rect 16940 6010 16996 6012
rect 17020 6010 17076 6012
rect 17100 6010 17156 6012
rect 16860 5958 16906 6010
rect 16906 5958 16916 6010
rect 16940 5958 16970 6010
rect 16970 5958 16982 6010
rect 16982 5958 16996 6010
rect 17020 5958 17034 6010
rect 17034 5958 17046 6010
rect 17046 5958 17076 6010
rect 17100 5958 17110 6010
rect 17110 5958 17156 6010
rect 16860 5956 16916 5958
rect 16940 5956 16996 5958
rect 17020 5956 17076 5958
rect 17100 5956 17156 5958
rect 14922 5072 14978 5128
rect 16860 4922 16916 4924
rect 16940 4922 16996 4924
rect 17020 4922 17076 4924
rect 17100 4922 17156 4924
rect 16860 4870 16906 4922
rect 16906 4870 16916 4922
rect 16940 4870 16970 4922
rect 16970 4870 16982 4922
rect 16982 4870 16996 4922
rect 17020 4870 17034 4922
rect 17034 4870 17046 4922
rect 17046 4870 17076 4922
rect 17100 4870 17110 4922
rect 17110 4870 17156 4922
rect 16860 4868 16916 4870
rect 16940 4868 16996 4870
rect 17020 4868 17076 4870
rect 17100 4868 17156 4870
rect 19982 6604 19984 6624
rect 19984 6604 20036 6624
rect 20036 6604 20038 6624
rect 19982 6568 20038 6604
rect 21178 8336 21234 8392
rect 21730 8472 21786 8528
rect 22161 7642 22217 7644
rect 22241 7642 22297 7644
rect 22321 7642 22377 7644
rect 22401 7642 22457 7644
rect 22161 7590 22207 7642
rect 22207 7590 22217 7642
rect 22241 7590 22271 7642
rect 22271 7590 22283 7642
rect 22283 7590 22297 7642
rect 22321 7590 22335 7642
rect 22335 7590 22347 7642
rect 22347 7590 22377 7642
rect 22401 7590 22411 7642
rect 22411 7590 22457 7642
rect 22161 7588 22217 7590
rect 22241 7588 22297 7590
rect 22321 7588 22377 7590
rect 22401 7588 22457 7590
rect 22161 6554 22217 6556
rect 22241 6554 22297 6556
rect 22321 6554 22377 6556
rect 22401 6554 22457 6556
rect 22161 6502 22207 6554
rect 22207 6502 22217 6554
rect 22241 6502 22271 6554
rect 22271 6502 22283 6554
rect 22283 6502 22297 6554
rect 22321 6502 22335 6554
rect 22335 6502 22347 6554
rect 22347 6502 22377 6554
rect 22401 6502 22411 6554
rect 22411 6502 22457 6554
rect 22161 6500 22217 6502
rect 22241 6500 22297 6502
rect 22321 6500 22377 6502
rect 22401 6500 22457 6502
rect 22834 7112 22890 7168
rect 23202 8064 23258 8120
rect 23202 7792 23258 7848
rect 23294 6976 23350 7032
rect 24306 6840 24362 6896
rect 24030 6180 24086 6216
rect 24030 6160 24032 6180
rect 24032 6160 24084 6180
rect 24084 6160 24086 6180
rect 20626 5480 20682 5536
rect 22161 5466 22217 5468
rect 22241 5466 22297 5468
rect 22321 5466 22377 5468
rect 22401 5466 22457 5468
rect 22161 5414 22207 5466
rect 22207 5414 22217 5466
rect 22241 5414 22271 5466
rect 22271 5414 22283 5466
rect 22283 5414 22297 5466
rect 22321 5414 22335 5466
rect 22335 5414 22347 5466
rect 22347 5414 22377 5466
rect 22401 5414 22411 5466
rect 22411 5414 22457 5466
rect 22161 5412 22217 5414
rect 22241 5412 22297 5414
rect 22321 5412 22377 5414
rect 22401 5412 22457 5414
rect 23386 5616 23442 5672
rect 27463 7098 27519 7100
rect 27543 7098 27599 7100
rect 27623 7098 27679 7100
rect 27703 7098 27759 7100
rect 27463 7046 27509 7098
rect 27509 7046 27519 7098
rect 27543 7046 27573 7098
rect 27573 7046 27585 7098
rect 27585 7046 27599 7098
rect 27623 7046 27637 7098
rect 27637 7046 27649 7098
rect 27649 7046 27679 7098
rect 27703 7046 27713 7098
rect 27713 7046 27759 7098
rect 27463 7044 27519 7046
rect 27543 7044 27599 7046
rect 27623 7044 27679 7046
rect 27703 7044 27759 7046
rect 30378 7384 30434 7440
rect 32034 7928 32090 7984
rect 31758 7268 31814 7304
rect 31758 7248 31760 7268
rect 31760 7248 31812 7268
rect 31812 7248 31814 7268
rect 32764 7642 32820 7644
rect 32844 7642 32900 7644
rect 32924 7642 32980 7644
rect 33004 7642 33060 7644
rect 32764 7590 32810 7642
rect 32810 7590 32820 7642
rect 32844 7590 32874 7642
rect 32874 7590 32886 7642
rect 32886 7590 32900 7642
rect 32924 7590 32938 7642
rect 32938 7590 32950 7642
rect 32950 7590 32980 7642
rect 33004 7590 33014 7642
rect 33014 7590 33060 7642
rect 32764 7588 32820 7590
rect 32844 7588 32900 7590
rect 32924 7588 32980 7590
rect 33004 7588 33060 7590
rect 24766 5752 24822 5808
rect 23202 5208 23258 5264
rect 14186 4664 14242 4720
rect 27463 6010 27519 6012
rect 27543 6010 27599 6012
rect 27623 6010 27679 6012
rect 27703 6010 27759 6012
rect 27463 5958 27509 6010
rect 27509 5958 27519 6010
rect 27543 5958 27573 6010
rect 27573 5958 27585 6010
rect 27585 5958 27599 6010
rect 27623 5958 27637 6010
rect 27637 5958 27649 6010
rect 27649 5958 27679 6010
rect 27703 5958 27713 6010
rect 27713 5958 27759 6010
rect 27463 5956 27519 5958
rect 27543 5956 27599 5958
rect 27623 5956 27679 5958
rect 27703 5956 27759 5958
rect 27463 4922 27519 4924
rect 27543 4922 27599 4924
rect 27623 4922 27679 4924
rect 27703 4922 27759 4924
rect 27463 4870 27509 4922
rect 27509 4870 27519 4922
rect 27543 4870 27573 4922
rect 27573 4870 27585 4922
rect 27585 4870 27599 4922
rect 27623 4870 27637 4922
rect 27637 4870 27649 4922
rect 27649 4870 27679 4922
rect 27703 4870 27713 4922
rect 27713 4870 27759 4922
rect 27463 4868 27519 4870
rect 27543 4868 27599 4870
rect 27623 4868 27679 4870
rect 27703 4868 27759 4870
rect 27066 4664 27122 4720
rect 11558 4378 11614 4380
rect 11638 4378 11694 4380
rect 11718 4378 11774 4380
rect 11798 4378 11854 4380
rect 11558 4326 11604 4378
rect 11604 4326 11614 4378
rect 11638 4326 11668 4378
rect 11668 4326 11680 4378
rect 11680 4326 11694 4378
rect 11718 4326 11732 4378
rect 11732 4326 11744 4378
rect 11744 4326 11774 4378
rect 11798 4326 11808 4378
rect 11808 4326 11854 4378
rect 11558 4324 11614 4326
rect 11638 4324 11694 4326
rect 11718 4324 11774 4326
rect 11798 4324 11854 4326
rect 22161 4378 22217 4380
rect 22241 4378 22297 4380
rect 22321 4378 22377 4380
rect 22401 4378 22457 4380
rect 22161 4326 22207 4378
rect 22207 4326 22217 4378
rect 22241 4326 22271 4378
rect 22271 4326 22283 4378
rect 22283 4326 22297 4378
rect 22321 4326 22335 4378
rect 22335 4326 22347 4378
rect 22347 4326 22377 4378
rect 22401 4326 22411 4378
rect 22411 4326 22457 4378
rect 22161 4324 22217 4326
rect 22241 4324 22297 4326
rect 22321 4324 22377 4326
rect 22401 4324 22457 4326
rect 6257 3834 6313 3836
rect 6337 3834 6393 3836
rect 6417 3834 6473 3836
rect 6497 3834 6553 3836
rect 6257 3782 6303 3834
rect 6303 3782 6313 3834
rect 6337 3782 6367 3834
rect 6367 3782 6379 3834
rect 6379 3782 6393 3834
rect 6417 3782 6431 3834
rect 6431 3782 6443 3834
rect 6443 3782 6473 3834
rect 6497 3782 6507 3834
rect 6507 3782 6553 3834
rect 6257 3780 6313 3782
rect 6337 3780 6393 3782
rect 6417 3780 6473 3782
rect 6497 3780 6553 3782
rect 16860 3834 16916 3836
rect 16940 3834 16996 3836
rect 17020 3834 17076 3836
rect 17100 3834 17156 3836
rect 16860 3782 16906 3834
rect 16906 3782 16916 3834
rect 16940 3782 16970 3834
rect 16970 3782 16982 3834
rect 16982 3782 16996 3834
rect 17020 3782 17034 3834
rect 17034 3782 17046 3834
rect 17046 3782 17076 3834
rect 17100 3782 17110 3834
rect 17110 3782 17156 3834
rect 16860 3780 16916 3782
rect 16940 3780 16996 3782
rect 17020 3780 17076 3782
rect 17100 3780 17156 3782
rect 27463 3834 27519 3836
rect 27543 3834 27599 3836
rect 27623 3834 27679 3836
rect 27703 3834 27759 3836
rect 27463 3782 27509 3834
rect 27509 3782 27519 3834
rect 27543 3782 27573 3834
rect 27573 3782 27585 3834
rect 27585 3782 27599 3834
rect 27623 3782 27637 3834
rect 27637 3782 27649 3834
rect 27649 3782 27679 3834
rect 27703 3782 27713 3834
rect 27713 3782 27759 3834
rect 27463 3780 27519 3782
rect 27543 3780 27599 3782
rect 27623 3780 27679 3782
rect 27703 3780 27759 3782
rect 11558 3290 11614 3292
rect 11638 3290 11694 3292
rect 11718 3290 11774 3292
rect 11798 3290 11854 3292
rect 11558 3238 11604 3290
rect 11604 3238 11614 3290
rect 11638 3238 11668 3290
rect 11668 3238 11680 3290
rect 11680 3238 11694 3290
rect 11718 3238 11732 3290
rect 11732 3238 11744 3290
rect 11744 3238 11774 3290
rect 11798 3238 11808 3290
rect 11808 3238 11854 3290
rect 11558 3236 11614 3238
rect 11638 3236 11694 3238
rect 11718 3236 11774 3238
rect 11798 3236 11854 3238
rect 22161 3290 22217 3292
rect 22241 3290 22297 3292
rect 22321 3290 22377 3292
rect 22401 3290 22457 3292
rect 22161 3238 22207 3290
rect 22207 3238 22217 3290
rect 22241 3238 22271 3290
rect 22271 3238 22283 3290
rect 22283 3238 22297 3290
rect 22321 3238 22335 3290
rect 22335 3238 22347 3290
rect 22347 3238 22377 3290
rect 22401 3238 22411 3290
rect 22411 3238 22457 3290
rect 22161 3236 22217 3238
rect 22241 3236 22297 3238
rect 22321 3236 22377 3238
rect 22401 3236 22457 3238
rect 6257 2746 6313 2748
rect 6337 2746 6393 2748
rect 6417 2746 6473 2748
rect 6497 2746 6553 2748
rect 6257 2694 6303 2746
rect 6303 2694 6313 2746
rect 6337 2694 6367 2746
rect 6367 2694 6379 2746
rect 6379 2694 6393 2746
rect 6417 2694 6431 2746
rect 6431 2694 6443 2746
rect 6443 2694 6473 2746
rect 6497 2694 6507 2746
rect 6507 2694 6553 2746
rect 6257 2692 6313 2694
rect 6337 2692 6393 2694
rect 6417 2692 6473 2694
rect 6497 2692 6553 2694
rect 16860 2746 16916 2748
rect 16940 2746 16996 2748
rect 17020 2746 17076 2748
rect 17100 2746 17156 2748
rect 16860 2694 16906 2746
rect 16906 2694 16916 2746
rect 16940 2694 16970 2746
rect 16970 2694 16982 2746
rect 16982 2694 16996 2746
rect 17020 2694 17034 2746
rect 17034 2694 17046 2746
rect 17046 2694 17076 2746
rect 17100 2694 17110 2746
rect 17110 2694 17156 2746
rect 16860 2692 16916 2694
rect 16940 2692 16996 2694
rect 17020 2692 17076 2694
rect 17100 2692 17156 2694
rect 27463 2746 27519 2748
rect 27543 2746 27599 2748
rect 27623 2746 27679 2748
rect 27703 2746 27759 2748
rect 27463 2694 27509 2746
rect 27509 2694 27519 2746
rect 27543 2694 27573 2746
rect 27573 2694 27585 2746
rect 27585 2694 27599 2746
rect 27623 2694 27637 2746
rect 27637 2694 27649 2746
rect 27649 2694 27679 2746
rect 27703 2694 27713 2746
rect 27713 2694 27759 2746
rect 27463 2692 27519 2694
rect 27543 2692 27599 2694
rect 27623 2692 27679 2694
rect 27703 2692 27759 2694
rect 33230 6704 33286 6760
rect 32764 6554 32820 6556
rect 32844 6554 32900 6556
rect 32924 6554 32980 6556
rect 33004 6554 33060 6556
rect 32764 6502 32810 6554
rect 32810 6502 32820 6554
rect 32844 6502 32874 6554
rect 32874 6502 32886 6554
rect 32886 6502 32900 6554
rect 32924 6502 32938 6554
rect 32938 6502 32950 6554
rect 32950 6502 32980 6554
rect 33004 6502 33014 6554
rect 33014 6502 33060 6554
rect 32764 6500 32820 6502
rect 32844 6500 32900 6502
rect 32924 6500 32980 6502
rect 33004 6500 33060 6502
rect 32764 5466 32820 5468
rect 32844 5466 32900 5468
rect 32924 5466 32980 5468
rect 33004 5466 33060 5468
rect 32764 5414 32810 5466
rect 32810 5414 32820 5466
rect 32844 5414 32874 5466
rect 32874 5414 32886 5466
rect 32886 5414 32900 5466
rect 32924 5414 32938 5466
rect 32938 5414 32950 5466
rect 32950 5414 32980 5466
rect 33004 5414 33014 5466
rect 33014 5414 33060 5466
rect 32764 5412 32820 5414
rect 32844 5412 32900 5414
rect 32924 5412 32980 5414
rect 33004 5412 33060 5414
rect 32764 4378 32820 4380
rect 32844 4378 32900 4380
rect 32924 4378 32980 4380
rect 33004 4378 33060 4380
rect 32764 4326 32810 4378
rect 32810 4326 32820 4378
rect 32844 4326 32874 4378
rect 32874 4326 32886 4378
rect 32886 4326 32900 4378
rect 32924 4326 32938 4378
rect 32938 4326 32950 4378
rect 32950 4326 32980 4378
rect 33004 4326 33014 4378
rect 33014 4326 33060 4378
rect 32764 4324 32820 4326
rect 32844 4324 32900 4326
rect 32924 4324 32980 4326
rect 33004 4324 33060 4326
rect 32764 3290 32820 3292
rect 32844 3290 32900 3292
rect 32924 3290 32980 3292
rect 33004 3290 33060 3292
rect 32764 3238 32810 3290
rect 32810 3238 32820 3290
rect 32844 3238 32874 3290
rect 32874 3238 32886 3290
rect 32886 3238 32900 3290
rect 32924 3238 32938 3290
rect 32938 3238 32950 3290
rect 32950 3238 32980 3290
rect 33004 3238 33014 3290
rect 33014 3238 33060 3290
rect 32764 3236 32820 3238
rect 32844 3236 32900 3238
rect 32924 3236 32980 3238
rect 33004 3236 33060 3238
rect 33506 5072 33562 5128
rect 33782 6296 33838 6352
rect 11558 2202 11614 2204
rect 11638 2202 11694 2204
rect 11718 2202 11774 2204
rect 11798 2202 11854 2204
rect 11558 2150 11604 2202
rect 11604 2150 11614 2202
rect 11638 2150 11668 2202
rect 11668 2150 11680 2202
rect 11680 2150 11694 2202
rect 11718 2150 11732 2202
rect 11732 2150 11744 2202
rect 11744 2150 11774 2202
rect 11798 2150 11808 2202
rect 11808 2150 11854 2202
rect 11558 2148 11614 2150
rect 11638 2148 11694 2150
rect 11718 2148 11774 2150
rect 11798 2148 11854 2150
rect 22161 2202 22217 2204
rect 22241 2202 22297 2204
rect 22321 2202 22377 2204
rect 22401 2202 22457 2204
rect 22161 2150 22207 2202
rect 22207 2150 22217 2202
rect 22241 2150 22271 2202
rect 22271 2150 22283 2202
rect 22283 2150 22297 2202
rect 22321 2150 22335 2202
rect 22335 2150 22347 2202
rect 22347 2150 22377 2202
rect 22401 2150 22411 2202
rect 22411 2150 22457 2202
rect 22161 2148 22217 2150
rect 22241 2148 22297 2150
rect 22321 2148 22377 2150
rect 22401 2148 22457 2150
rect 32764 2202 32820 2204
rect 32844 2202 32900 2204
rect 32924 2202 32980 2204
rect 33004 2202 33060 2204
rect 32764 2150 32810 2202
rect 32810 2150 32820 2202
rect 32844 2150 32874 2202
rect 32874 2150 32886 2202
rect 32886 2150 32900 2202
rect 32924 2150 32938 2202
rect 32938 2150 32950 2202
rect 32950 2150 32980 2202
rect 33004 2150 33014 2202
rect 33014 2150 33060 2202
rect 32764 2148 32820 2150
rect 32844 2148 32900 2150
rect 32924 2148 32980 2150
rect 33004 2148 33060 2150
rect 38066 7098 38122 7100
rect 38146 7098 38202 7100
rect 38226 7098 38282 7100
rect 38306 7098 38362 7100
rect 38066 7046 38112 7098
rect 38112 7046 38122 7098
rect 38146 7046 38176 7098
rect 38176 7046 38188 7098
rect 38188 7046 38202 7098
rect 38226 7046 38240 7098
rect 38240 7046 38252 7098
rect 38252 7046 38282 7098
rect 38306 7046 38316 7098
rect 38316 7046 38362 7098
rect 38066 7044 38122 7046
rect 38146 7044 38202 7046
rect 38226 7044 38282 7046
rect 38306 7044 38362 7046
rect 38066 6010 38122 6012
rect 38146 6010 38202 6012
rect 38226 6010 38282 6012
rect 38306 6010 38362 6012
rect 38066 5958 38112 6010
rect 38112 5958 38122 6010
rect 38146 5958 38176 6010
rect 38176 5958 38188 6010
rect 38188 5958 38202 6010
rect 38226 5958 38240 6010
rect 38240 5958 38252 6010
rect 38252 5958 38282 6010
rect 38306 5958 38316 6010
rect 38316 5958 38362 6010
rect 38066 5956 38122 5958
rect 38146 5956 38202 5958
rect 38226 5956 38282 5958
rect 38306 5956 38362 5958
rect 38066 4922 38122 4924
rect 38146 4922 38202 4924
rect 38226 4922 38282 4924
rect 38306 4922 38362 4924
rect 38066 4870 38112 4922
rect 38112 4870 38122 4922
rect 38146 4870 38176 4922
rect 38176 4870 38188 4922
rect 38188 4870 38202 4922
rect 38226 4870 38240 4922
rect 38240 4870 38252 4922
rect 38252 4870 38282 4922
rect 38306 4870 38316 4922
rect 38316 4870 38362 4922
rect 38066 4868 38122 4870
rect 38146 4868 38202 4870
rect 38226 4868 38282 4870
rect 38306 4868 38362 4870
rect 38066 3834 38122 3836
rect 38146 3834 38202 3836
rect 38226 3834 38282 3836
rect 38306 3834 38362 3836
rect 38066 3782 38112 3834
rect 38112 3782 38122 3834
rect 38146 3782 38176 3834
rect 38176 3782 38188 3834
rect 38188 3782 38202 3834
rect 38226 3782 38240 3834
rect 38240 3782 38252 3834
rect 38252 3782 38282 3834
rect 38306 3782 38316 3834
rect 38316 3782 38362 3834
rect 38066 3780 38122 3782
rect 38146 3780 38202 3782
rect 38226 3780 38282 3782
rect 38306 3780 38362 3782
rect 38066 2746 38122 2748
rect 38146 2746 38202 2748
rect 38226 2746 38282 2748
rect 38306 2746 38362 2748
rect 38066 2694 38112 2746
rect 38112 2694 38122 2746
rect 38146 2694 38176 2746
rect 38176 2694 38188 2746
rect 38188 2694 38202 2746
rect 38226 2694 38240 2746
rect 38240 2694 38252 2746
rect 38252 2694 38282 2746
rect 38306 2694 38316 2746
rect 38316 2694 38362 2746
rect 38066 2692 38122 2694
rect 38146 2692 38202 2694
rect 38226 2692 38282 2694
rect 38306 2692 38362 2694
rect 43367 7642 43423 7644
rect 43447 7642 43503 7644
rect 43527 7642 43583 7644
rect 43607 7642 43663 7644
rect 43367 7590 43413 7642
rect 43413 7590 43423 7642
rect 43447 7590 43477 7642
rect 43477 7590 43489 7642
rect 43489 7590 43503 7642
rect 43527 7590 43541 7642
rect 43541 7590 43553 7642
rect 43553 7590 43583 7642
rect 43607 7590 43617 7642
rect 43617 7590 43663 7642
rect 43367 7588 43423 7590
rect 43447 7588 43503 7590
rect 43527 7588 43583 7590
rect 43607 7588 43663 7590
rect 43367 6554 43423 6556
rect 43447 6554 43503 6556
rect 43527 6554 43583 6556
rect 43607 6554 43663 6556
rect 43367 6502 43413 6554
rect 43413 6502 43423 6554
rect 43447 6502 43477 6554
rect 43477 6502 43489 6554
rect 43489 6502 43503 6554
rect 43527 6502 43541 6554
rect 43541 6502 43553 6554
rect 43553 6502 43583 6554
rect 43607 6502 43617 6554
rect 43617 6502 43663 6554
rect 43367 6500 43423 6502
rect 43447 6500 43503 6502
rect 43527 6500 43583 6502
rect 43607 6500 43663 6502
rect 43367 5466 43423 5468
rect 43447 5466 43503 5468
rect 43527 5466 43583 5468
rect 43607 5466 43663 5468
rect 43367 5414 43413 5466
rect 43413 5414 43423 5466
rect 43447 5414 43477 5466
rect 43477 5414 43489 5466
rect 43489 5414 43503 5466
rect 43527 5414 43541 5466
rect 43541 5414 43553 5466
rect 43553 5414 43583 5466
rect 43607 5414 43617 5466
rect 43617 5414 43663 5466
rect 43367 5412 43423 5414
rect 43447 5412 43503 5414
rect 43527 5412 43583 5414
rect 43607 5412 43663 5414
rect 43367 4378 43423 4380
rect 43447 4378 43503 4380
rect 43527 4378 43583 4380
rect 43607 4378 43663 4380
rect 43367 4326 43413 4378
rect 43413 4326 43423 4378
rect 43447 4326 43477 4378
rect 43477 4326 43489 4378
rect 43489 4326 43503 4378
rect 43527 4326 43541 4378
rect 43541 4326 43553 4378
rect 43553 4326 43583 4378
rect 43607 4326 43617 4378
rect 43617 4326 43663 4378
rect 43367 4324 43423 4326
rect 43447 4324 43503 4326
rect 43527 4324 43583 4326
rect 43607 4324 43663 4326
rect 43367 3290 43423 3292
rect 43447 3290 43503 3292
rect 43527 3290 43583 3292
rect 43607 3290 43663 3292
rect 43367 3238 43413 3290
rect 43413 3238 43423 3290
rect 43447 3238 43477 3290
rect 43477 3238 43489 3290
rect 43489 3238 43503 3290
rect 43527 3238 43541 3290
rect 43541 3238 43553 3290
rect 43553 3238 43583 3290
rect 43607 3238 43617 3290
rect 43617 3238 43663 3290
rect 43367 3236 43423 3238
rect 43447 3236 43503 3238
rect 43527 3236 43583 3238
rect 43607 3236 43663 3238
rect 43367 2202 43423 2204
rect 43447 2202 43503 2204
rect 43527 2202 43583 2204
rect 43607 2202 43663 2204
rect 43367 2150 43413 2202
rect 43413 2150 43423 2202
rect 43447 2150 43477 2202
rect 43477 2150 43489 2202
rect 43489 2150 43503 2202
rect 43527 2150 43541 2202
rect 43541 2150 43553 2202
rect 43553 2150 43583 2202
rect 43607 2150 43617 2202
rect 43617 2150 43663 2202
rect 43367 2148 43423 2150
rect 43447 2148 43503 2150
rect 43527 2148 43583 2150
rect 43607 2148 43663 2150
<< metal3 >>
rect 15101 8530 15167 8533
rect 21725 8530 21791 8533
rect 15101 8528 21791 8530
rect 15101 8472 15106 8528
rect 15162 8472 21730 8528
rect 21786 8472 21791 8528
rect 15101 8470 21791 8472
rect 15101 8467 15167 8470
rect 21725 8467 21791 8470
rect 13721 8394 13787 8397
rect 21173 8394 21239 8397
rect 13721 8392 21239 8394
rect 13721 8336 13726 8392
rect 13782 8336 21178 8392
rect 21234 8336 21239 8392
rect 13721 8334 21239 8336
rect 13721 8331 13787 8334
rect 21173 8331 21239 8334
rect 12157 8258 12223 8261
rect 12157 8256 16314 8258
rect 12157 8200 12162 8256
rect 12218 8200 16314 8256
rect 12157 8198 16314 8200
rect 12157 8195 12223 8198
rect 16254 7986 16314 8198
rect 16481 8122 16547 8125
rect 23197 8122 23263 8125
rect 16481 8120 23263 8122
rect 16481 8064 16486 8120
rect 16542 8064 23202 8120
rect 23258 8064 23263 8120
rect 16481 8062 23263 8064
rect 16481 8059 16547 8062
rect 23197 8059 23263 8062
rect 17309 7986 17375 7989
rect 16254 7984 17375 7986
rect 16254 7928 17314 7984
rect 17370 7928 17375 7984
rect 16254 7926 17375 7928
rect 17309 7923 17375 7926
rect 17769 7986 17835 7989
rect 32029 7986 32095 7989
rect 17769 7984 32095 7986
rect 17769 7928 17774 7984
rect 17830 7928 32034 7984
rect 32090 7928 32095 7984
rect 17769 7926 32095 7928
rect 17769 7923 17835 7926
rect 32029 7923 32095 7926
rect 15929 7850 15995 7853
rect 23197 7850 23263 7853
rect 15929 7848 23263 7850
rect 15929 7792 15934 7848
rect 15990 7792 23202 7848
rect 23258 7792 23263 7848
rect 15929 7790 23263 7792
rect 15929 7787 15995 7790
rect 23197 7787 23263 7790
rect 11548 7648 11864 7649
rect 11548 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11864 7648
rect 11548 7583 11864 7584
rect 22151 7648 22467 7649
rect 22151 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22467 7648
rect 22151 7583 22467 7584
rect 32754 7648 33070 7649
rect 32754 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33070 7648
rect 32754 7583 33070 7584
rect 43357 7648 43673 7649
rect 43357 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43673 7648
rect 43357 7583 43673 7584
rect 18321 7442 18387 7445
rect 30373 7442 30439 7445
rect 18321 7440 30439 7442
rect 18321 7384 18326 7440
rect 18382 7384 30378 7440
rect 30434 7384 30439 7440
rect 18321 7382 30439 7384
rect 18321 7379 18387 7382
rect 30373 7379 30439 7382
rect 17401 7306 17467 7309
rect 31753 7306 31819 7309
rect 17401 7304 31819 7306
rect 17401 7248 17406 7304
rect 17462 7248 31758 7304
rect 31814 7248 31819 7304
rect 17401 7246 31819 7248
rect 17401 7243 17467 7246
rect 31753 7243 31819 7246
rect 17309 7170 17375 7173
rect 22829 7170 22895 7173
rect 17309 7168 22895 7170
rect 17309 7112 17314 7168
rect 17370 7112 22834 7168
rect 22890 7112 22895 7168
rect 17309 7110 22895 7112
rect 17309 7107 17375 7110
rect 22829 7107 22895 7110
rect 6247 7104 6563 7105
rect 6247 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6563 7104
rect 6247 7039 6563 7040
rect 16850 7104 17166 7105
rect 16850 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17166 7104
rect 16850 7039 17166 7040
rect 27453 7104 27769 7105
rect 27453 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27769 7104
rect 27453 7039 27769 7040
rect 38056 7104 38372 7105
rect 38056 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38372 7104
rect 38056 7039 38372 7040
rect 11605 7034 11671 7037
rect 16573 7034 16639 7037
rect 11605 7032 16639 7034
rect 11605 6976 11610 7032
rect 11666 6976 16578 7032
rect 16634 6976 16639 7032
rect 11605 6974 16639 6976
rect 11605 6971 11671 6974
rect 16573 6971 16639 6974
rect 18413 7034 18479 7037
rect 23289 7034 23355 7037
rect 18413 7032 23355 7034
rect 18413 6976 18418 7032
rect 18474 6976 23294 7032
rect 23350 6976 23355 7032
rect 18413 6974 23355 6976
rect 18413 6971 18479 6974
rect 23289 6971 23355 6974
rect 24301 6898 24367 6901
rect 12390 6896 24367 6898
rect 12390 6840 24306 6896
rect 24362 6840 24367 6896
rect 12390 6838 24367 6840
rect 6177 6762 6243 6765
rect 12390 6762 12450 6838
rect 24301 6835 24367 6838
rect 6177 6760 12450 6762
rect 6177 6704 6182 6760
rect 6238 6704 12450 6760
rect 6177 6702 12450 6704
rect 14273 6762 14339 6765
rect 33225 6762 33291 6765
rect 14273 6760 33291 6762
rect 14273 6704 14278 6760
rect 14334 6704 33230 6760
rect 33286 6704 33291 6760
rect 14273 6702 33291 6704
rect 6177 6699 6243 6702
rect 14273 6699 14339 6702
rect 33225 6699 33291 6702
rect 11973 6626 12039 6629
rect 19977 6626 20043 6629
rect 11973 6624 20043 6626
rect 11973 6568 11978 6624
rect 12034 6568 19982 6624
rect 20038 6568 20043 6624
rect 11973 6566 20043 6568
rect 11973 6563 12039 6566
rect 19977 6563 20043 6566
rect 11548 6560 11864 6561
rect 11548 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11864 6560
rect 11548 6495 11864 6496
rect 22151 6560 22467 6561
rect 22151 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22467 6560
rect 22151 6495 22467 6496
rect 32754 6560 33070 6561
rect 32754 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33070 6560
rect 32754 6495 33070 6496
rect 43357 6560 43673 6561
rect 43357 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43673 6560
rect 43357 6495 43673 6496
rect 14365 6490 14431 6493
rect 18413 6490 18479 6493
rect 14365 6488 18479 6490
rect 14365 6432 14370 6488
rect 14426 6432 18418 6488
rect 18474 6432 18479 6488
rect 14365 6430 18479 6432
rect 14365 6427 14431 6430
rect 18413 6427 18479 6430
rect 15193 6354 15259 6357
rect 33777 6354 33843 6357
rect 15193 6352 33843 6354
rect 15193 6296 15198 6352
rect 15254 6296 33782 6352
rect 33838 6296 33843 6352
rect 15193 6294 33843 6296
rect 15193 6291 15259 6294
rect 33777 6291 33843 6294
rect 5809 6218 5875 6221
rect 24025 6218 24091 6221
rect 5809 6216 24091 6218
rect 5809 6160 5814 6216
rect 5870 6160 24030 6216
rect 24086 6160 24091 6216
rect 5809 6158 24091 6160
rect 5809 6155 5875 6158
rect 24025 6155 24091 6158
rect 6247 6016 6563 6017
rect 6247 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6563 6016
rect 6247 5951 6563 5952
rect 16850 6016 17166 6017
rect 16850 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17166 6016
rect 16850 5951 17166 5952
rect 27453 6016 27769 6017
rect 27453 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27769 6016
rect 27453 5951 27769 5952
rect 38056 6016 38372 6017
rect 38056 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38372 6016
rect 38056 5951 38372 5952
rect 15285 5810 15351 5813
rect 24761 5810 24827 5813
rect 15285 5808 24827 5810
rect 15285 5752 15290 5808
rect 15346 5752 24766 5808
rect 24822 5752 24827 5808
rect 15285 5750 24827 5752
rect 15285 5747 15351 5750
rect 24761 5747 24827 5750
rect 9673 5674 9739 5677
rect 23381 5674 23447 5677
rect 9673 5672 23447 5674
rect 9673 5616 9678 5672
rect 9734 5616 23386 5672
rect 23442 5616 23447 5672
rect 9673 5614 23447 5616
rect 9673 5611 9739 5614
rect 23381 5611 23447 5614
rect 12341 5538 12407 5541
rect 20621 5538 20687 5541
rect 12341 5536 20687 5538
rect 12341 5480 12346 5536
rect 12402 5480 20626 5536
rect 20682 5480 20687 5536
rect 12341 5478 20687 5480
rect 12341 5475 12407 5478
rect 20621 5475 20687 5478
rect 11548 5472 11864 5473
rect 11548 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11864 5472
rect 11548 5407 11864 5408
rect 22151 5472 22467 5473
rect 22151 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22467 5472
rect 22151 5407 22467 5408
rect 32754 5472 33070 5473
rect 32754 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33070 5472
rect 32754 5407 33070 5408
rect 43357 5472 43673 5473
rect 43357 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43673 5472
rect 43357 5407 43673 5408
rect 10593 5266 10659 5269
rect 23197 5266 23263 5269
rect 10593 5264 23263 5266
rect 10593 5208 10598 5264
rect 10654 5208 23202 5264
rect 23258 5208 23263 5264
rect 10593 5206 23263 5208
rect 10593 5203 10659 5206
rect 23197 5203 23263 5206
rect 14917 5130 14983 5133
rect 33501 5130 33567 5133
rect 14917 5128 33567 5130
rect 14917 5072 14922 5128
rect 14978 5072 33506 5128
rect 33562 5072 33567 5128
rect 14917 5070 33567 5072
rect 14917 5067 14983 5070
rect 33501 5067 33567 5070
rect 6247 4928 6563 4929
rect 6247 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6563 4928
rect 6247 4863 6563 4864
rect 16850 4928 17166 4929
rect 16850 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17166 4928
rect 16850 4863 17166 4864
rect 27453 4928 27769 4929
rect 27453 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27769 4928
rect 27453 4863 27769 4864
rect 38056 4928 38372 4929
rect 38056 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38372 4928
rect 38056 4863 38372 4864
rect 14181 4722 14247 4725
rect 27061 4722 27127 4725
rect 14181 4720 27127 4722
rect 14181 4664 14186 4720
rect 14242 4664 27066 4720
rect 27122 4664 27127 4720
rect 14181 4662 27127 4664
rect 14181 4659 14247 4662
rect 27061 4659 27127 4662
rect 11548 4384 11864 4385
rect 11548 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11864 4384
rect 11548 4319 11864 4320
rect 22151 4384 22467 4385
rect 22151 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22467 4384
rect 22151 4319 22467 4320
rect 32754 4384 33070 4385
rect 32754 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33070 4384
rect 32754 4319 33070 4320
rect 43357 4384 43673 4385
rect 43357 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43673 4384
rect 43357 4319 43673 4320
rect 6247 3840 6563 3841
rect 6247 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6563 3840
rect 6247 3775 6563 3776
rect 16850 3840 17166 3841
rect 16850 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17166 3840
rect 16850 3775 17166 3776
rect 27453 3840 27769 3841
rect 27453 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27769 3840
rect 27453 3775 27769 3776
rect 38056 3840 38372 3841
rect 38056 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38372 3840
rect 38056 3775 38372 3776
rect 11548 3296 11864 3297
rect 11548 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11864 3296
rect 11548 3231 11864 3232
rect 22151 3296 22467 3297
rect 22151 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22467 3296
rect 22151 3231 22467 3232
rect 32754 3296 33070 3297
rect 32754 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33070 3296
rect 32754 3231 33070 3232
rect 43357 3296 43673 3297
rect 43357 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43673 3296
rect 43357 3231 43673 3232
rect 6247 2752 6563 2753
rect 6247 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6563 2752
rect 6247 2687 6563 2688
rect 16850 2752 17166 2753
rect 16850 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17166 2752
rect 16850 2687 17166 2688
rect 27453 2752 27769 2753
rect 27453 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27769 2752
rect 27453 2687 27769 2688
rect 38056 2752 38372 2753
rect 38056 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38372 2752
rect 38056 2687 38372 2688
rect 11548 2208 11864 2209
rect 11548 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11864 2208
rect 11548 2143 11864 2144
rect 22151 2208 22467 2209
rect 22151 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22467 2208
rect 22151 2143 22467 2144
rect 32754 2208 33070 2209
rect 32754 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33070 2208
rect 32754 2143 33070 2144
rect 43357 2208 43673 2209
rect 43357 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43673 2208
rect 43357 2143 43673 2144
<< via3 >>
rect 11554 7644 11618 7648
rect 11554 7588 11558 7644
rect 11558 7588 11614 7644
rect 11614 7588 11618 7644
rect 11554 7584 11618 7588
rect 11634 7644 11698 7648
rect 11634 7588 11638 7644
rect 11638 7588 11694 7644
rect 11694 7588 11698 7644
rect 11634 7584 11698 7588
rect 11714 7644 11778 7648
rect 11714 7588 11718 7644
rect 11718 7588 11774 7644
rect 11774 7588 11778 7644
rect 11714 7584 11778 7588
rect 11794 7644 11858 7648
rect 11794 7588 11798 7644
rect 11798 7588 11854 7644
rect 11854 7588 11858 7644
rect 11794 7584 11858 7588
rect 22157 7644 22221 7648
rect 22157 7588 22161 7644
rect 22161 7588 22217 7644
rect 22217 7588 22221 7644
rect 22157 7584 22221 7588
rect 22237 7644 22301 7648
rect 22237 7588 22241 7644
rect 22241 7588 22297 7644
rect 22297 7588 22301 7644
rect 22237 7584 22301 7588
rect 22317 7644 22381 7648
rect 22317 7588 22321 7644
rect 22321 7588 22377 7644
rect 22377 7588 22381 7644
rect 22317 7584 22381 7588
rect 22397 7644 22461 7648
rect 22397 7588 22401 7644
rect 22401 7588 22457 7644
rect 22457 7588 22461 7644
rect 22397 7584 22461 7588
rect 32760 7644 32824 7648
rect 32760 7588 32764 7644
rect 32764 7588 32820 7644
rect 32820 7588 32824 7644
rect 32760 7584 32824 7588
rect 32840 7644 32904 7648
rect 32840 7588 32844 7644
rect 32844 7588 32900 7644
rect 32900 7588 32904 7644
rect 32840 7584 32904 7588
rect 32920 7644 32984 7648
rect 32920 7588 32924 7644
rect 32924 7588 32980 7644
rect 32980 7588 32984 7644
rect 32920 7584 32984 7588
rect 33000 7644 33064 7648
rect 33000 7588 33004 7644
rect 33004 7588 33060 7644
rect 33060 7588 33064 7644
rect 33000 7584 33064 7588
rect 43363 7644 43427 7648
rect 43363 7588 43367 7644
rect 43367 7588 43423 7644
rect 43423 7588 43427 7644
rect 43363 7584 43427 7588
rect 43443 7644 43507 7648
rect 43443 7588 43447 7644
rect 43447 7588 43503 7644
rect 43503 7588 43507 7644
rect 43443 7584 43507 7588
rect 43523 7644 43587 7648
rect 43523 7588 43527 7644
rect 43527 7588 43583 7644
rect 43583 7588 43587 7644
rect 43523 7584 43587 7588
rect 43603 7644 43667 7648
rect 43603 7588 43607 7644
rect 43607 7588 43663 7644
rect 43663 7588 43667 7644
rect 43603 7584 43667 7588
rect 6253 7100 6317 7104
rect 6253 7044 6257 7100
rect 6257 7044 6313 7100
rect 6313 7044 6317 7100
rect 6253 7040 6317 7044
rect 6333 7100 6397 7104
rect 6333 7044 6337 7100
rect 6337 7044 6393 7100
rect 6393 7044 6397 7100
rect 6333 7040 6397 7044
rect 6413 7100 6477 7104
rect 6413 7044 6417 7100
rect 6417 7044 6473 7100
rect 6473 7044 6477 7100
rect 6413 7040 6477 7044
rect 6493 7100 6557 7104
rect 6493 7044 6497 7100
rect 6497 7044 6553 7100
rect 6553 7044 6557 7100
rect 6493 7040 6557 7044
rect 16856 7100 16920 7104
rect 16856 7044 16860 7100
rect 16860 7044 16916 7100
rect 16916 7044 16920 7100
rect 16856 7040 16920 7044
rect 16936 7100 17000 7104
rect 16936 7044 16940 7100
rect 16940 7044 16996 7100
rect 16996 7044 17000 7100
rect 16936 7040 17000 7044
rect 17016 7100 17080 7104
rect 17016 7044 17020 7100
rect 17020 7044 17076 7100
rect 17076 7044 17080 7100
rect 17016 7040 17080 7044
rect 17096 7100 17160 7104
rect 17096 7044 17100 7100
rect 17100 7044 17156 7100
rect 17156 7044 17160 7100
rect 17096 7040 17160 7044
rect 27459 7100 27523 7104
rect 27459 7044 27463 7100
rect 27463 7044 27519 7100
rect 27519 7044 27523 7100
rect 27459 7040 27523 7044
rect 27539 7100 27603 7104
rect 27539 7044 27543 7100
rect 27543 7044 27599 7100
rect 27599 7044 27603 7100
rect 27539 7040 27603 7044
rect 27619 7100 27683 7104
rect 27619 7044 27623 7100
rect 27623 7044 27679 7100
rect 27679 7044 27683 7100
rect 27619 7040 27683 7044
rect 27699 7100 27763 7104
rect 27699 7044 27703 7100
rect 27703 7044 27759 7100
rect 27759 7044 27763 7100
rect 27699 7040 27763 7044
rect 38062 7100 38126 7104
rect 38062 7044 38066 7100
rect 38066 7044 38122 7100
rect 38122 7044 38126 7100
rect 38062 7040 38126 7044
rect 38142 7100 38206 7104
rect 38142 7044 38146 7100
rect 38146 7044 38202 7100
rect 38202 7044 38206 7100
rect 38142 7040 38206 7044
rect 38222 7100 38286 7104
rect 38222 7044 38226 7100
rect 38226 7044 38282 7100
rect 38282 7044 38286 7100
rect 38222 7040 38286 7044
rect 38302 7100 38366 7104
rect 38302 7044 38306 7100
rect 38306 7044 38362 7100
rect 38362 7044 38366 7100
rect 38302 7040 38366 7044
rect 11554 6556 11618 6560
rect 11554 6500 11558 6556
rect 11558 6500 11614 6556
rect 11614 6500 11618 6556
rect 11554 6496 11618 6500
rect 11634 6556 11698 6560
rect 11634 6500 11638 6556
rect 11638 6500 11694 6556
rect 11694 6500 11698 6556
rect 11634 6496 11698 6500
rect 11714 6556 11778 6560
rect 11714 6500 11718 6556
rect 11718 6500 11774 6556
rect 11774 6500 11778 6556
rect 11714 6496 11778 6500
rect 11794 6556 11858 6560
rect 11794 6500 11798 6556
rect 11798 6500 11854 6556
rect 11854 6500 11858 6556
rect 11794 6496 11858 6500
rect 22157 6556 22221 6560
rect 22157 6500 22161 6556
rect 22161 6500 22217 6556
rect 22217 6500 22221 6556
rect 22157 6496 22221 6500
rect 22237 6556 22301 6560
rect 22237 6500 22241 6556
rect 22241 6500 22297 6556
rect 22297 6500 22301 6556
rect 22237 6496 22301 6500
rect 22317 6556 22381 6560
rect 22317 6500 22321 6556
rect 22321 6500 22377 6556
rect 22377 6500 22381 6556
rect 22317 6496 22381 6500
rect 22397 6556 22461 6560
rect 22397 6500 22401 6556
rect 22401 6500 22457 6556
rect 22457 6500 22461 6556
rect 22397 6496 22461 6500
rect 32760 6556 32824 6560
rect 32760 6500 32764 6556
rect 32764 6500 32820 6556
rect 32820 6500 32824 6556
rect 32760 6496 32824 6500
rect 32840 6556 32904 6560
rect 32840 6500 32844 6556
rect 32844 6500 32900 6556
rect 32900 6500 32904 6556
rect 32840 6496 32904 6500
rect 32920 6556 32984 6560
rect 32920 6500 32924 6556
rect 32924 6500 32980 6556
rect 32980 6500 32984 6556
rect 32920 6496 32984 6500
rect 33000 6556 33064 6560
rect 33000 6500 33004 6556
rect 33004 6500 33060 6556
rect 33060 6500 33064 6556
rect 33000 6496 33064 6500
rect 43363 6556 43427 6560
rect 43363 6500 43367 6556
rect 43367 6500 43423 6556
rect 43423 6500 43427 6556
rect 43363 6496 43427 6500
rect 43443 6556 43507 6560
rect 43443 6500 43447 6556
rect 43447 6500 43503 6556
rect 43503 6500 43507 6556
rect 43443 6496 43507 6500
rect 43523 6556 43587 6560
rect 43523 6500 43527 6556
rect 43527 6500 43583 6556
rect 43583 6500 43587 6556
rect 43523 6496 43587 6500
rect 43603 6556 43667 6560
rect 43603 6500 43607 6556
rect 43607 6500 43663 6556
rect 43663 6500 43667 6556
rect 43603 6496 43667 6500
rect 6253 6012 6317 6016
rect 6253 5956 6257 6012
rect 6257 5956 6313 6012
rect 6313 5956 6317 6012
rect 6253 5952 6317 5956
rect 6333 6012 6397 6016
rect 6333 5956 6337 6012
rect 6337 5956 6393 6012
rect 6393 5956 6397 6012
rect 6333 5952 6397 5956
rect 6413 6012 6477 6016
rect 6413 5956 6417 6012
rect 6417 5956 6473 6012
rect 6473 5956 6477 6012
rect 6413 5952 6477 5956
rect 6493 6012 6557 6016
rect 6493 5956 6497 6012
rect 6497 5956 6553 6012
rect 6553 5956 6557 6012
rect 6493 5952 6557 5956
rect 16856 6012 16920 6016
rect 16856 5956 16860 6012
rect 16860 5956 16916 6012
rect 16916 5956 16920 6012
rect 16856 5952 16920 5956
rect 16936 6012 17000 6016
rect 16936 5956 16940 6012
rect 16940 5956 16996 6012
rect 16996 5956 17000 6012
rect 16936 5952 17000 5956
rect 17016 6012 17080 6016
rect 17016 5956 17020 6012
rect 17020 5956 17076 6012
rect 17076 5956 17080 6012
rect 17016 5952 17080 5956
rect 17096 6012 17160 6016
rect 17096 5956 17100 6012
rect 17100 5956 17156 6012
rect 17156 5956 17160 6012
rect 17096 5952 17160 5956
rect 27459 6012 27523 6016
rect 27459 5956 27463 6012
rect 27463 5956 27519 6012
rect 27519 5956 27523 6012
rect 27459 5952 27523 5956
rect 27539 6012 27603 6016
rect 27539 5956 27543 6012
rect 27543 5956 27599 6012
rect 27599 5956 27603 6012
rect 27539 5952 27603 5956
rect 27619 6012 27683 6016
rect 27619 5956 27623 6012
rect 27623 5956 27679 6012
rect 27679 5956 27683 6012
rect 27619 5952 27683 5956
rect 27699 6012 27763 6016
rect 27699 5956 27703 6012
rect 27703 5956 27759 6012
rect 27759 5956 27763 6012
rect 27699 5952 27763 5956
rect 38062 6012 38126 6016
rect 38062 5956 38066 6012
rect 38066 5956 38122 6012
rect 38122 5956 38126 6012
rect 38062 5952 38126 5956
rect 38142 6012 38206 6016
rect 38142 5956 38146 6012
rect 38146 5956 38202 6012
rect 38202 5956 38206 6012
rect 38142 5952 38206 5956
rect 38222 6012 38286 6016
rect 38222 5956 38226 6012
rect 38226 5956 38282 6012
rect 38282 5956 38286 6012
rect 38222 5952 38286 5956
rect 38302 6012 38366 6016
rect 38302 5956 38306 6012
rect 38306 5956 38362 6012
rect 38362 5956 38366 6012
rect 38302 5952 38366 5956
rect 11554 5468 11618 5472
rect 11554 5412 11558 5468
rect 11558 5412 11614 5468
rect 11614 5412 11618 5468
rect 11554 5408 11618 5412
rect 11634 5468 11698 5472
rect 11634 5412 11638 5468
rect 11638 5412 11694 5468
rect 11694 5412 11698 5468
rect 11634 5408 11698 5412
rect 11714 5468 11778 5472
rect 11714 5412 11718 5468
rect 11718 5412 11774 5468
rect 11774 5412 11778 5468
rect 11714 5408 11778 5412
rect 11794 5468 11858 5472
rect 11794 5412 11798 5468
rect 11798 5412 11854 5468
rect 11854 5412 11858 5468
rect 11794 5408 11858 5412
rect 22157 5468 22221 5472
rect 22157 5412 22161 5468
rect 22161 5412 22217 5468
rect 22217 5412 22221 5468
rect 22157 5408 22221 5412
rect 22237 5468 22301 5472
rect 22237 5412 22241 5468
rect 22241 5412 22297 5468
rect 22297 5412 22301 5468
rect 22237 5408 22301 5412
rect 22317 5468 22381 5472
rect 22317 5412 22321 5468
rect 22321 5412 22377 5468
rect 22377 5412 22381 5468
rect 22317 5408 22381 5412
rect 22397 5468 22461 5472
rect 22397 5412 22401 5468
rect 22401 5412 22457 5468
rect 22457 5412 22461 5468
rect 22397 5408 22461 5412
rect 32760 5468 32824 5472
rect 32760 5412 32764 5468
rect 32764 5412 32820 5468
rect 32820 5412 32824 5468
rect 32760 5408 32824 5412
rect 32840 5468 32904 5472
rect 32840 5412 32844 5468
rect 32844 5412 32900 5468
rect 32900 5412 32904 5468
rect 32840 5408 32904 5412
rect 32920 5468 32984 5472
rect 32920 5412 32924 5468
rect 32924 5412 32980 5468
rect 32980 5412 32984 5468
rect 32920 5408 32984 5412
rect 33000 5468 33064 5472
rect 33000 5412 33004 5468
rect 33004 5412 33060 5468
rect 33060 5412 33064 5468
rect 33000 5408 33064 5412
rect 43363 5468 43427 5472
rect 43363 5412 43367 5468
rect 43367 5412 43423 5468
rect 43423 5412 43427 5468
rect 43363 5408 43427 5412
rect 43443 5468 43507 5472
rect 43443 5412 43447 5468
rect 43447 5412 43503 5468
rect 43503 5412 43507 5468
rect 43443 5408 43507 5412
rect 43523 5468 43587 5472
rect 43523 5412 43527 5468
rect 43527 5412 43583 5468
rect 43583 5412 43587 5468
rect 43523 5408 43587 5412
rect 43603 5468 43667 5472
rect 43603 5412 43607 5468
rect 43607 5412 43663 5468
rect 43663 5412 43667 5468
rect 43603 5408 43667 5412
rect 6253 4924 6317 4928
rect 6253 4868 6257 4924
rect 6257 4868 6313 4924
rect 6313 4868 6317 4924
rect 6253 4864 6317 4868
rect 6333 4924 6397 4928
rect 6333 4868 6337 4924
rect 6337 4868 6393 4924
rect 6393 4868 6397 4924
rect 6333 4864 6397 4868
rect 6413 4924 6477 4928
rect 6413 4868 6417 4924
rect 6417 4868 6473 4924
rect 6473 4868 6477 4924
rect 6413 4864 6477 4868
rect 6493 4924 6557 4928
rect 6493 4868 6497 4924
rect 6497 4868 6553 4924
rect 6553 4868 6557 4924
rect 6493 4864 6557 4868
rect 16856 4924 16920 4928
rect 16856 4868 16860 4924
rect 16860 4868 16916 4924
rect 16916 4868 16920 4924
rect 16856 4864 16920 4868
rect 16936 4924 17000 4928
rect 16936 4868 16940 4924
rect 16940 4868 16996 4924
rect 16996 4868 17000 4924
rect 16936 4864 17000 4868
rect 17016 4924 17080 4928
rect 17016 4868 17020 4924
rect 17020 4868 17076 4924
rect 17076 4868 17080 4924
rect 17016 4864 17080 4868
rect 17096 4924 17160 4928
rect 17096 4868 17100 4924
rect 17100 4868 17156 4924
rect 17156 4868 17160 4924
rect 17096 4864 17160 4868
rect 27459 4924 27523 4928
rect 27459 4868 27463 4924
rect 27463 4868 27519 4924
rect 27519 4868 27523 4924
rect 27459 4864 27523 4868
rect 27539 4924 27603 4928
rect 27539 4868 27543 4924
rect 27543 4868 27599 4924
rect 27599 4868 27603 4924
rect 27539 4864 27603 4868
rect 27619 4924 27683 4928
rect 27619 4868 27623 4924
rect 27623 4868 27679 4924
rect 27679 4868 27683 4924
rect 27619 4864 27683 4868
rect 27699 4924 27763 4928
rect 27699 4868 27703 4924
rect 27703 4868 27759 4924
rect 27759 4868 27763 4924
rect 27699 4864 27763 4868
rect 38062 4924 38126 4928
rect 38062 4868 38066 4924
rect 38066 4868 38122 4924
rect 38122 4868 38126 4924
rect 38062 4864 38126 4868
rect 38142 4924 38206 4928
rect 38142 4868 38146 4924
rect 38146 4868 38202 4924
rect 38202 4868 38206 4924
rect 38142 4864 38206 4868
rect 38222 4924 38286 4928
rect 38222 4868 38226 4924
rect 38226 4868 38282 4924
rect 38282 4868 38286 4924
rect 38222 4864 38286 4868
rect 38302 4924 38366 4928
rect 38302 4868 38306 4924
rect 38306 4868 38362 4924
rect 38362 4868 38366 4924
rect 38302 4864 38366 4868
rect 11554 4380 11618 4384
rect 11554 4324 11558 4380
rect 11558 4324 11614 4380
rect 11614 4324 11618 4380
rect 11554 4320 11618 4324
rect 11634 4380 11698 4384
rect 11634 4324 11638 4380
rect 11638 4324 11694 4380
rect 11694 4324 11698 4380
rect 11634 4320 11698 4324
rect 11714 4380 11778 4384
rect 11714 4324 11718 4380
rect 11718 4324 11774 4380
rect 11774 4324 11778 4380
rect 11714 4320 11778 4324
rect 11794 4380 11858 4384
rect 11794 4324 11798 4380
rect 11798 4324 11854 4380
rect 11854 4324 11858 4380
rect 11794 4320 11858 4324
rect 22157 4380 22221 4384
rect 22157 4324 22161 4380
rect 22161 4324 22217 4380
rect 22217 4324 22221 4380
rect 22157 4320 22221 4324
rect 22237 4380 22301 4384
rect 22237 4324 22241 4380
rect 22241 4324 22297 4380
rect 22297 4324 22301 4380
rect 22237 4320 22301 4324
rect 22317 4380 22381 4384
rect 22317 4324 22321 4380
rect 22321 4324 22377 4380
rect 22377 4324 22381 4380
rect 22317 4320 22381 4324
rect 22397 4380 22461 4384
rect 22397 4324 22401 4380
rect 22401 4324 22457 4380
rect 22457 4324 22461 4380
rect 22397 4320 22461 4324
rect 32760 4380 32824 4384
rect 32760 4324 32764 4380
rect 32764 4324 32820 4380
rect 32820 4324 32824 4380
rect 32760 4320 32824 4324
rect 32840 4380 32904 4384
rect 32840 4324 32844 4380
rect 32844 4324 32900 4380
rect 32900 4324 32904 4380
rect 32840 4320 32904 4324
rect 32920 4380 32984 4384
rect 32920 4324 32924 4380
rect 32924 4324 32980 4380
rect 32980 4324 32984 4380
rect 32920 4320 32984 4324
rect 33000 4380 33064 4384
rect 33000 4324 33004 4380
rect 33004 4324 33060 4380
rect 33060 4324 33064 4380
rect 33000 4320 33064 4324
rect 43363 4380 43427 4384
rect 43363 4324 43367 4380
rect 43367 4324 43423 4380
rect 43423 4324 43427 4380
rect 43363 4320 43427 4324
rect 43443 4380 43507 4384
rect 43443 4324 43447 4380
rect 43447 4324 43503 4380
rect 43503 4324 43507 4380
rect 43443 4320 43507 4324
rect 43523 4380 43587 4384
rect 43523 4324 43527 4380
rect 43527 4324 43583 4380
rect 43583 4324 43587 4380
rect 43523 4320 43587 4324
rect 43603 4380 43667 4384
rect 43603 4324 43607 4380
rect 43607 4324 43663 4380
rect 43663 4324 43667 4380
rect 43603 4320 43667 4324
rect 6253 3836 6317 3840
rect 6253 3780 6257 3836
rect 6257 3780 6313 3836
rect 6313 3780 6317 3836
rect 6253 3776 6317 3780
rect 6333 3836 6397 3840
rect 6333 3780 6337 3836
rect 6337 3780 6393 3836
rect 6393 3780 6397 3836
rect 6333 3776 6397 3780
rect 6413 3836 6477 3840
rect 6413 3780 6417 3836
rect 6417 3780 6473 3836
rect 6473 3780 6477 3836
rect 6413 3776 6477 3780
rect 6493 3836 6557 3840
rect 6493 3780 6497 3836
rect 6497 3780 6553 3836
rect 6553 3780 6557 3836
rect 6493 3776 6557 3780
rect 16856 3836 16920 3840
rect 16856 3780 16860 3836
rect 16860 3780 16916 3836
rect 16916 3780 16920 3836
rect 16856 3776 16920 3780
rect 16936 3836 17000 3840
rect 16936 3780 16940 3836
rect 16940 3780 16996 3836
rect 16996 3780 17000 3836
rect 16936 3776 17000 3780
rect 17016 3836 17080 3840
rect 17016 3780 17020 3836
rect 17020 3780 17076 3836
rect 17076 3780 17080 3836
rect 17016 3776 17080 3780
rect 17096 3836 17160 3840
rect 17096 3780 17100 3836
rect 17100 3780 17156 3836
rect 17156 3780 17160 3836
rect 17096 3776 17160 3780
rect 27459 3836 27523 3840
rect 27459 3780 27463 3836
rect 27463 3780 27519 3836
rect 27519 3780 27523 3836
rect 27459 3776 27523 3780
rect 27539 3836 27603 3840
rect 27539 3780 27543 3836
rect 27543 3780 27599 3836
rect 27599 3780 27603 3836
rect 27539 3776 27603 3780
rect 27619 3836 27683 3840
rect 27619 3780 27623 3836
rect 27623 3780 27679 3836
rect 27679 3780 27683 3836
rect 27619 3776 27683 3780
rect 27699 3836 27763 3840
rect 27699 3780 27703 3836
rect 27703 3780 27759 3836
rect 27759 3780 27763 3836
rect 27699 3776 27763 3780
rect 38062 3836 38126 3840
rect 38062 3780 38066 3836
rect 38066 3780 38122 3836
rect 38122 3780 38126 3836
rect 38062 3776 38126 3780
rect 38142 3836 38206 3840
rect 38142 3780 38146 3836
rect 38146 3780 38202 3836
rect 38202 3780 38206 3836
rect 38142 3776 38206 3780
rect 38222 3836 38286 3840
rect 38222 3780 38226 3836
rect 38226 3780 38282 3836
rect 38282 3780 38286 3836
rect 38222 3776 38286 3780
rect 38302 3836 38366 3840
rect 38302 3780 38306 3836
rect 38306 3780 38362 3836
rect 38362 3780 38366 3836
rect 38302 3776 38366 3780
rect 11554 3292 11618 3296
rect 11554 3236 11558 3292
rect 11558 3236 11614 3292
rect 11614 3236 11618 3292
rect 11554 3232 11618 3236
rect 11634 3292 11698 3296
rect 11634 3236 11638 3292
rect 11638 3236 11694 3292
rect 11694 3236 11698 3292
rect 11634 3232 11698 3236
rect 11714 3292 11778 3296
rect 11714 3236 11718 3292
rect 11718 3236 11774 3292
rect 11774 3236 11778 3292
rect 11714 3232 11778 3236
rect 11794 3292 11858 3296
rect 11794 3236 11798 3292
rect 11798 3236 11854 3292
rect 11854 3236 11858 3292
rect 11794 3232 11858 3236
rect 22157 3292 22221 3296
rect 22157 3236 22161 3292
rect 22161 3236 22217 3292
rect 22217 3236 22221 3292
rect 22157 3232 22221 3236
rect 22237 3292 22301 3296
rect 22237 3236 22241 3292
rect 22241 3236 22297 3292
rect 22297 3236 22301 3292
rect 22237 3232 22301 3236
rect 22317 3292 22381 3296
rect 22317 3236 22321 3292
rect 22321 3236 22377 3292
rect 22377 3236 22381 3292
rect 22317 3232 22381 3236
rect 22397 3292 22461 3296
rect 22397 3236 22401 3292
rect 22401 3236 22457 3292
rect 22457 3236 22461 3292
rect 22397 3232 22461 3236
rect 32760 3292 32824 3296
rect 32760 3236 32764 3292
rect 32764 3236 32820 3292
rect 32820 3236 32824 3292
rect 32760 3232 32824 3236
rect 32840 3292 32904 3296
rect 32840 3236 32844 3292
rect 32844 3236 32900 3292
rect 32900 3236 32904 3292
rect 32840 3232 32904 3236
rect 32920 3292 32984 3296
rect 32920 3236 32924 3292
rect 32924 3236 32980 3292
rect 32980 3236 32984 3292
rect 32920 3232 32984 3236
rect 33000 3292 33064 3296
rect 33000 3236 33004 3292
rect 33004 3236 33060 3292
rect 33060 3236 33064 3292
rect 33000 3232 33064 3236
rect 43363 3292 43427 3296
rect 43363 3236 43367 3292
rect 43367 3236 43423 3292
rect 43423 3236 43427 3292
rect 43363 3232 43427 3236
rect 43443 3292 43507 3296
rect 43443 3236 43447 3292
rect 43447 3236 43503 3292
rect 43503 3236 43507 3292
rect 43443 3232 43507 3236
rect 43523 3292 43587 3296
rect 43523 3236 43527 3292
rect 43527 3236 43583 3292
rect 43583 3236 43587 3292
rect 43523 3232 43587 3236
rect 43603 3292 43667 3296
rect 43603 3236 43607 3292
rect 43607 3236 43663 3292
rect 43663 3236 43667 3292
rect 43603 3232 43667 3236
rect 6253 2748 6317 2752
rect 6253 2692 6257 2748
rect 6257 2692 6313 2748
rect 6313 2692 6317 2748
rect 6253 2688 6317 2692
rect 6333 2748 6397 2752
rect 6333 2692 6337 2748
rect 6337 2692 6393 2748
rect 6393 2692 6397 2748
rect 6333 2688 6397 2692
rect 6413 2748 6477 2752
rect 6413 2692 6417 2748
rect 6417 2692 6473 2748
rect 6473 2692 6477 2748
rect 6413 2688 6477 2692
rect 6493 2748 6557 2752
rect 6493 2692 6497 2748
rect 6497 2692 6553 2748
rect 6553 2692 6557 2748
rect 6493 2688 6557 2692
rect 16856 2748 16920 2752
rect 16856 2692 16860 2748
rect 16860 2692 16916 2748
rect 16916 2692 16920 2748
rect 16856 2688 16920 2692
rect 16936 2748 17000 2752
rect 16936 2692 16940 2748
rect 16940 2692 16996 2748
rect 16996 2692 17000 2748
rect 16936 2688 17000 2692
rect 17016 2748 17080 2752
rect 17016 2692 17020 2748
rect 17020 2692 17076 2748
rect 17076 2692 17080 2748
rect 17016 2688 17080 2692
rect 17096 2748 17160 2752
rect 17096 2692 17100 2748
rect 17100 2692 17156 2748
rect 17156 2692 17160 2748
rect 17096 2688 17160 2692
rect 27459 2748 27523 2752
rect 27459 2692 27463 2748
rect 27463 2692 27519 2748
rect 27519 2692 27523 2748
rect 27459 2688 27523 2692
rect 27539 2748 27603 2752
rect 27539 2692 27543 2748
rect 27543 2692 27599 2748
rect 27599 2692 27603 2748
rect 27539 2688 27603 2692
rect 27619 2748 27683 2752
rect 27619 2692 27623 2748
rect 27623 2692 27679 2748
rect 27679 2692 27683 2748
rect 27619 2688 27683 2692
rect 27699 2748 27763 2752
rect 27699 2692 27703 2748
rect 27703 2692 27759 2748
rect 27759 2692 27763 2748
rect 27699 2688 27763 2692
rect 38062 2748 38126 2752
rect 38062 2692 38066 2748
rect 38066 2692 38122 2748
rect 38122 2692 38126 2748
rect 38062 2688 38126 2692
rect 38142 2748 38206 2752
rect 38142 2692 38146 2748
rect 38146 2692 38202 2748
rect 38202 2692 38206 2748
rect 38142 2688 38206 2692
rect 38222 2748 38286 2752
rect 38222 2692 38226 2748
rect 38226 2692 38282 2748
rect 38282 2692 38286 2748
rect 38222 2688 38286 2692
rect 38302 2748 38366 2752
rect 38302 2692 38306 2748
rect 38306 2692 38362 2748
rect 38362 2692 38366 2748
rect 38302 2688 38366 2692
rect 11554 2204 11618 2208
rect 11554 2148 11558 2204
rect 11558 2148 11614 2204
rect 11614 2148 11618 2204
rect 11554 2144 11618 2148
rect 11634 2204 11698 2208
rect 11634 2148 11638 2204
rect 11638 2148 11694 2204
rect 11694 2148 11698 2204
rect 11634 2144 11698 2148
rect 11714 2204 11778 2208
rect 11714 2148 11718 2204
rect 11718 2148 11774 2204
rect 11774 2148 11778 2204
rect 11714 2144 11778 2148
rect 11794 2204 11858 2208
rect 11794 2148 11798 2204
rect 11798 2148 11854 2204
rect 11854 2148 11858 2204
rect 11794 2144 11858 2148
rect 22157 2204 22221 2208
rect 22157 2148 22161 2204
rect 22161 2148 22217 2204
rect 22217 2148 22221 2204
rect 22157 2144 22221 2148
rect 22237 2204 22301 2208
rect 22237 2148 22241 2204
rect 22241 2148 22297 2204
rect 22297 2148 22301 2204
rect 22237 2144 22301 2148
rect 22317 2204 22381 2208
rect 22317 2148 22321 2204
rect 22321 2148 22377 2204
rect 22377 2148 22381 2204
rect 22317 2144 22381 2148
rect 22397 2204 22461 2208
rect 22397 2148 22401 2204
rect 22401 2148 22457 2204
rect 22457 2148 22461 2204
rect 22397 2144 22461 2148
rect 32760 2204 32824 2208
rect 32760 2148 32764 2204
rect 32764 2148 32820 2204
rect 32820 2148 32824 2204
rect 32760 2144 32824 2148
rect 32840 2204 32904 2208
rect 32840 2148 32844 2204
rect 32844 2148 32900 2204
rect 32900 2148 32904 2204
rect 32840 2144 32904 2148
rect 32920 2204 32984 2208
rect 32920 2148 32924 2204
rect 32924 2148 32980 2204
rect 32980 2148 32984 2204
rect 32920 2144 32984 2148
rect 33000 2204 33064 2208
rect 33000 2148 33004 2204
rect 33004 2148 33060 2204
rect 33060 2148 33064 2204
rect 33000 2144 33064 2148
rect 43363 2204 43427 2208
rect 43363 2148 43367 2204
rect 43367 2148 43423 2204
rect 43423 2148 43427 2204
rect 43363 2144 43427 2148
rect 43443 2204 43507 2208
rect 43443 2148 43447 2204
rect 43447 2148 43503 2204
rect 43503 2148 43507 2204
rect 43443 2144 43507 2148
rect 43523 2204 43587 2208
rect 43523 2148 43527 2204
rect 43527 2148 43583 2204
rect 43583 2148 43587 2204
rect 43523 2144 43587 2148
rect 43603 2204 43667 2208
rect 43603 2148 43607 2204
rect 43607 2148 43663 2204
rect 43663 2148 43667 2204
rect 43603 2144 43667 2148
<< metal4 >>
rect 6245 7104 6565 7664
rect 6245 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6565 7104
rect 6245 6016 6565 7040
rect 6245 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6565 6016
rect 6245 4928 6565 5952
rect 6245 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6565 4928
rect 6245 3840 6565 4864
rect 6245 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6565 3840
rect 6245 2752 6565 3776
rect 6245 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6565 2752
rect 6245 2128 6565 2688
rect 11546 7648 11866 7664
rect 11546 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11866 7648
rect 11546 6560 11866 7584
rect 11546 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11866 6560
rect 11546 5472 11866 6496
rect 11546 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11866 5472
rect 11546 4384 11866 5408
rect 11546 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11866 4384
rect 11546 3296 11866 4320
rect 11546 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11866 3296
rect 11546 2208 11866 3232
rect 11546 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11866 2208
rect 11546 2128 11866 2144
rect 16848 7104 17168 7664
rect 16848 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17168 7104
rect 16848 6016 17168 7040
rect 16848 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17168 6016
rect 16848 4928 17168 5952
rect 16848 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17168 4928
rect 16848 3840 17168 4864
rect 16848 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17168 3840
rect 16848 2752 17168 3776
rect 16848 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17168 2752
rect 16848 2128 17168 2688
rect 22149 7648 22469 7664
rect 22149 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22469 7648
rect 22149 6560 22469 7584
rect 22149 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22469 6560
rect 22149 5472 22469 6496
rect 22149 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22469 5472
rect 22149 4384 22469 5408
rect 22149 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22469 4384
rect 22149 3296 22469 4320
rect 22149 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22469 3296
rect 22149 2208 22469 3232
rect 22149 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22469 2208
rect 22149 2128 22469 2144
rect 27451 7104 27771 7664
rect 27451 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27771 7104
rect 27451 6016 27771 7040
rect 27451 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27771 6016
rect 27451 4928 27771 5952
rect 27451 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27771 4928
rect 27451 3840 27771 4864
rect 27451 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27771 3840
rect 27451 2752 27771 3776
rect 27451 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27771 2752
rect 27451 2128 27771 2688
rect 32752 7648 33072 7664
rect 32752 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33072 7648
rect 32752 6560 33072 7584
rect 32752 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33072 6560
rect 32752 5472 33072 6496
rect 32752 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33072 5472
rect 32752 4384 33072 5408
rect 32752 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33072 4384
rect 32752 3296 33072 4320
rect 32752 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33072 3296
rect 32752 2208 33072 3232
rect 32752 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33072 2208
rect 32752 2128 33072 2144
rect 38054 7104 38374 7664
rect 38054 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38374 7104
rect 38054 6016 38374 7040
rect 38054 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38374 6016
rect 38054 4928 38374 5952
rect 38054 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38374 4928
rect 38054 3840 38374 4864
rect 38054 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38374 3840
rect 38054 2752 38374 3776
rect 38054 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38374 2752
rect 38054 2128 38374 2688
rect 43355 7648 43675 7664
rect 43355 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43675 7648
rect 43355 6560 43675 7584
rect 43355 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43675 6560
rect 43355 5472 43675 6496
rect 43355 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43675 5472
rect 43355 4384 43675 5408
rect 43355 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43675 4384
rect 43355 3296 43675 4320
rect 43355 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43675 3296
rect 43355 2208 43675 3232
rect 43355 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43675 2208
rect 43355 2128 43675 2144
use sky130_fd_sc_hd__clkbuf_2  _01_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _02_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _03_
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _05_
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _06_
timestamp 1688980957
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 35512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 37812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _20_
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _21_
timestamp 1688980957
transform 1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _22_
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp 1688980957
transform 1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _24_
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _25_
timestamp 1688980957
transform 1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _26_
timestamp 1688980957
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _27_
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _30_
timestamp 1688980957
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 10672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1688980957
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1688980957
transform 1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _38_
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _39_
timestamp 1688980957
transform 1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _40_
timestamp 1688980957
transform 1 0 28336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _41_
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _42_
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _43_
timestamp 1688980957
transform 1 0 27232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _44_
timestamp 1688980957
transform 1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _45_
timestamp 1688980957
transform 1 0 26496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _46_
timestamp 1688980957
transform 1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _47_
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _48_
timestamp 1688980957
transform 1 0 25300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _49_
timestamp 1688980957
transform 1 0 25024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _50_
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _51_
timestamp 1688980957
transform 1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 14720 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1688980957
transform 1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1688980957
transform 1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1688980957
transform 1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1688980957
transform 1 0 33120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _73_
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform -1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform -1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_73
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_96
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_124
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_188
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_211
timestamp 1688980957
transform 1 0 20516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_234
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_246
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_257
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_321 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_326
timestamp 1688980957
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_334
timestamp 1688980957
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_354
timestamp 1688980957
transform 1 0 33672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_358
timestamp 1688980957
transform 1 0 34040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_368
timestamp 1688980957
transform 1 0 34960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_372
timestamp 1688980957
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_402
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_410
timestamp 1688980957
transform 1 0 38824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418
timestamp 1688980957
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_427
timestamp 1688980957
transform 1 0 40388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_435
timestamp 1688980957
transform 1 0 41124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_441
timestamp 1688980957
transform 1 0 41676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_452
timestamp 1688980957
transform 1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_172
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_184
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_233
timestamp 1688980957
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_257
timestamp 1688980957
transform 1 0 24748 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_262
timestamp 1688980957
transform 1 0 25208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_274
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_353
timestamp 1688980957
transform 1 0 33580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_365
timestamp 1688980957
transform 1 0 34684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_377
timestamp 1688980957
transform 1 0 35788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_389
timestamp 1688980957
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_402
timestamp 1688980957
transform 1 0 38088 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_414
timestamp 1688980957
transform 1 0 39192 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_426
timestamp 1688980957
transform 1 0 40296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_438
timestamp 1688980957
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_360
timestamp 1688980957
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_457
timestamp 1688980957
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_457
timestamp 1688980957
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_91
timestamp 1688980957
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_98
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_110
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_122
timestamp 1688980957
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_134
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_80
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_107
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_131
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_139
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_146
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_154
timestamp 1688980957
transform 1 0 15272 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_159
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_177
timestamp 1688980957
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_182
timestamp 1688980957
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_187
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_191
timestamp 1688980957
transform 1 0 18676 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_195
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_199
timestamp 1688980957
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_203
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_215
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_243
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_250
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_254
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_266
timestamp 1688980957
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1688980957
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_100
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_191
timestamp 1688980957
transform 1 0 18676 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_224
timestamp 1688980957
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_240
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_259
timestamp 1688980957
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_266
timestamp 1688980957
transform 1 0 25576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_271
timestamp 1688980957
transform 1 0 26036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_275
timestamp 1688980957
transform 1 0 26404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_279
timestamp 1688980957
transform 1 0 26772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_283
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_293
timestamp 1688980957
transform 1 0 28060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 1688980957
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_318
timestamp 1688980957
transform 1 0 30360 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_330
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_342
timestamp 1688980957
transform 1 0 32568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_346
timestamp 1688980957
transform 1 0 32936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_356
timestamp 1688980957
transform 1 0 33856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_362
timestamp 1688980957
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_88
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_94
timestamp 1688980957
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_98
timestamp 1688980957
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_122
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_126
timestamp 1688980957
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_251
timestamp 1688980957
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_355
timestamp 1688980957
transform 1 0 33764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_362
timestamp 1688980957
transform 1 0 34408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_433
timestamp 1688980957
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_445
timestamp 1688980957
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_457
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 24472 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 33396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 42964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 28612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 29808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 26036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 32936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 33488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 33028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform 1 0 31188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform 1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 37444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 38916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 38548 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 40388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 40388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 35236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 35788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 35236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 36340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 36340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 37812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 4968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 5520 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 9568 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 13432 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 14260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 14812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 10672 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform -1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 11408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform -1 0 12328 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 12880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 15364 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 15916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 16468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 33856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_term_single_147 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 34058 9840 34114 10300 0 FreeSans 224 90 0 0 Co
port 0 nsew signal tristate
flabel metal2 s 3238 -300 3294 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 26514 -300 26570 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 28630 -300 28686 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 30746 -300 30802 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 32862 -300 32918 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 34978 -300 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 37094 -300 37150 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 39210 -300 39266 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 41326 -300 41382 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 43442 -300 43498 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 7470 -300 7526 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 9586 -300 9642 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 11702 -300 11758 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 13818 -300 13874 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 15934 -300 15990 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 20166 -300 20222 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 22282 -300 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 34334 9840 34390 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 37094 9840 37150 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 37370 9840 37426 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 37646 9840 37702 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 37922 9840 37978 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 38198 9840 38254 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 38474 9840 38530 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 38750 9840 38806 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 39026 9840 39082 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 39302 9840 39358 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 39578 9840 39634 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 34610 9840 34666 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 34886 9840 34942 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 35162 9840 35218 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 35438 9840 35494 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 35714 9840 35770 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 35990 9840 36046 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 36266 9840 36322 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 36542 9840 36598 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 36818 9840 36874 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5078 9840 5134 10300 0 FreeSans 224 90 0 0 N1BEG[0]
port 41 nsew signal tristate
flabel metal2 s 5354 9840 5410 10300 0 FreeSans 224 90 0 0 N1BEG[1]
port 42 nsew signal tristate
flabel metal2 s 5630 9840 5686 10300 0 FreeSans 224 90 0 0 N1BEG[2]
port 43 nsew signal tristate
flabel metal2 s 5906 9840 5962 10300 0 FreeSans 224 90 0 0 N1BEG[3]
port 44 nsew signal tristate
flabel metal2 s 6182 9840 6238 10300 0 FreeSans 224 90 0 0 N2BEG[0]
port 45 nsew signal tristate
flabel metal2 s 6458 9840 6514 10300 0 FreeSans 224 90 0 0 N2BEG[1]
port 46 nsew signal tristate
flabel metal2 s 6734 9840 6790 10300 0 FreeSans 224 90 0 0 N2BEG[2]
port 47 nsew signal tristate
flabel metal2 s 7010 9840 7066 10300 0 FreeSans 224 90 0 0 N2BEG[3]
port 48 nsew signal tristate
flabel metal2 s 7286 9840 7342 10300 0 FreeSans 224 90 0 0 N2BEG[4]
port 49 nsew signal tristate
flabel metal2 s 7562 9840 7618 10300 0 FreeSans 224 90 0 0 N2BEG[5]
port 50 nsew signal tristate
flabel metal2 s 7838 9840 7894 10300 0 FreeSans 224 90 0 0 N2BEG[6]
port 51 nsew signal tristate
flabel metal2 s 8114 9840 8170 10300 0 FreeSans 224 90 0 0 N2BEG[7]
port 52 nsew signal tristate
flabel metal2 s 8390 9840 8446 10300 0 FreeSans 224 90 0 0 N2BEGb[0]
port 53 nsew signal tristate
flabel metal2 s 8666 9840 8722 10300 0 FreeSans 224 90 0 0 N2BEGb[1]
port 54 nsew signal tristate
flabel metal2 s 8942 9840 8998 10300 0 FreeSans 224 90 0 0 N2BEGb[2]
port 55 nsew signal tristate
flabel metal2 s 9218 9840 9274 10300 0 FreeSans 224 90 0 0 N2BEGb[3]
port 56 nsew signal tristate
flabel metal2 s 9494 9840 9550 10300 0 FreeSans 224 90 0 0 N2BEGb[4]
port 57 nsew signal tristate
flabel metal2 s 9770 9840 9826 10300 0 FreeSans 224 90 0 0 N2BEGb[5]
port 58 nsew signal tristate
flabel metal2 s 10046 9840 10102 10300 0 FreeSans 224 90 0 0 N2BEGb[6]
port 59 nsew signal tristate
flabel metal2 s 10322 9840 10378 10300 0 FreeSans 224 90 0 0 N2BEGb[7]
port 60 nsew signal tristate
flabel metal2 s 10598 9840 10654 10300 0 FreeSans 224 90 0 0 N4BEG[0]
port 61 nsew signal tristate
flabel metal2 s 13358 9840 13414 10300 0 FreeSans 224 90 0 0 N4BEG[10]
port 62 nsew signal tristate
flabel metal2 s 13634 9840 13690 10300 0 FreeSans 224 90 0 0 N4BEG[11]
port 63 nsew signal tristate
flabel metal2 s 13910 9840 13966 10300 0 FreeSans 224 90 0 0 N4BEG[12]
port 64 nsew signal tristate
flabel metal2 s 14186 9840 14242 10300 0 FreeSans 224 90 0 0 N4BEG[13]
port 65 nsew signal tristate
flabel metal2 s 14462 9840 14518 10300 0 FreeSans 224 90 0 0 N4BEG[14]
port 66 nsew signal tristate
flabel metal2 s 14738 9840 14794 10300 0 FreeSans 224 90 0 0 N4BEG[15]
port 67 nsew signal tristate
flabel metal2 s 10874 9840 10930 10300 0 FreeSans 224 90 0 0 N4BEG[1]
port 68 nsew signal tristate
flabel metal2 s 11150 9840 11206 10300 0 FreeSans 224 90 0 0 N4BEG[2]
port 69 nsew signal tristate
flabel metal2 s 11426 9840 11482 10300 0 FreeSans 224 90 0 0 N4BEG[3]
port 70 nsew signal tristate
flabel metal2 s 11702 9840 11758 10300 0 FreeSans 224 90 0 0 N4BEG[4]
port 71 nsew signal tristate
flabel metal2 s 11978 9840 12034 10300 0 FreeSans 224 90 0 0 N4BEG[5]
port 72 nsew signal tristate
flabel metal2 s 12254 9840 12310 10300 0 FreeSans 224 90 0 0 N4BEG[6]
port 73 nsew signal tristate
flabel metal2 s 12530 9840 12586 10300 0 FreeSans 224 90 0 0 N4BEG[7]
port 74 nsew signal tristate
flabel metal2 s 12806 9840 12862 10300 0 FreeSans 224 90 0 0 N4BEG[8]
port 75 nsew signal tristate
flabel metal2 s 13082 9840 13138 10300 0 FreeSans 224 90 0 0 N4BEG[9]
port 76 nsew signal tristate
flabel metal2 s 15014 9840 15070 10300 0 FreeSans 224 90 0 0 NN4BEG[0]
port 77 nsew signal tristate
flabel metal2 s 17774 9840 17830 10300 0 FreeSans 224 90 0 0 NN4BEG[10]
port 78 nsew signal tristate
flabel metal2 s 18050 9840 18106 10300 0 FreeSans 224 90 0 0 NN4BEG[11]
port 79 nsew signal tristate
flabel metal2 s 18326 9840 18382 10300 0 FreeSans 224 90 0 0 NN4BEG[12]
port 80 nsew signal tristate
flabel metal2 s 18602 9840 18658 10300 0 FreeSans 224 90 0 0 NN4BEG[13]
port 81 nsew signal tristate
flabel metal2 s 18878 9840 18934 10300 0 FreeSans 224 90 0 0 NN4BEG[14]
port 82 nsew signal tristate
flabel metal2 s 19154 9840 19210 10300 0 FreeSans 224 90 0 0 NN4BEG[15]
port 83 nsew signal tristate
flabel metal2 s 15290 9840 15346 10300 0 FreeSans 224 90 0 0 NN4BEG[1]
port 84 nsew signal tristate
flabel metal2 s 15566 9840 15622 10300 0 FreeSans 224 90 0 0 NN4BEG[2]
port 85 nsew signal tristate
flabel metal2 s 15842 9840 15898 10300 0 FreeSans 224 90 0 0 NN4BEG[3]
port 86 nsew signal tristate
flabel metal2 s 16118 9840 16174 10300 0 FreeSans 224 90 0 0 NN4BEG[4]
port 87 nsew signal tristate
flabel metal2 s 16394 9840 16450 10300 0 FreeSans 224 90 0 0 NN4BEG[5]
port 88 nsew signal tristate
flabel metal2 s 16670 9840 16726 10300 0 FreeSans 224 90 0 0 NN4BEG[6]
port 89 nsew signal tristate
flabel metal2 s 16946 9840 17002 10300 0 FreeSans 224 90 0 0 NN4BEG[7]
port 90 nsew signal tristate
flabel metal2 s 17222 9840 17278 10300 0 FreeSans 224 90 0 0 NN4BEG[8]
port 91 nsew signal tristate
flabel metal2 s 17498 9840 17554 10300 0 FreeSans 224 90 0 0 NN4BEG[9]
port 92 nsew signal tristate
flabel metal2 s 19430 9840 19486 10300 0 FreeSans 224 90 0 0 S1END[0]
port 93 nsew signal input
flabel metal2 s 19706 9840 19762 10300 0 FreeSans 224 90 0 0 S1END[1]
port 94 nsew signal input
flabel metal2 s 19982 9840 20038 10300 0 FreeSans 224 90 0 0 S1END[2]
port 95 nsew signal input
flabel metal2 s 20258 9840 20314 10300 0 FreeSans 224 90 0 0 S1END[3]
port 96 nsew signal input
flabel metal2 s 20534 9840 20590 10300 0 FreeSans 224 90 0 0 S2END[0]
port 97 nsew signal input
flabel metal2 s 20810 9840 20866 10300 0 FreeSans 224 90 0 0 S2END[1]
port 98 nsew signal input
flabel metal2 s 21086 9840 21142 10300 0 FreeSans 224 90 0 0 S2END[2]
port 99 nsew signal input
flabel metal2 s 21362 9840 21418 10300 0 FreeSans 224 90 0 0 S2END[3]
port 100 nsew signal input
flabel metal2 s 21638 9840 21694 10300 0 FreeSans 224 90 0 0 S2END[4]
port 101 nsew signal input
flabel metal2 s 21914 9840 21970 10300 0 FreeSans 224 90 0 0 S2END[5]
port 102 nsew signal input
flabel metal2 s 22190 9840 22246 10300 0 FreeSans 224 90 0 0 S2END[6]
port 103 nsew signal input
flabel metal2 s 22466 9840 22522 10300 0 FreeSans 224 90 0 0 S2END[7]
port 104 nsew signal input
flabel metal2 s 22742 9840 22798 10300 0 FreeSans 224 90 0 0 S2MID[0]
port 105 nsew signal input
flabel metal2 s 23018 9840 23074 10300 0 FreeSans 224 90 0 0 S2MID[1]
port 106 nsew signal input
flabel metal2 s 23294 9840 23350 10300 0 FreeSans 224 90 0 0 S2MID[2]
port 107 nsew signal input
flabel metal2 s 23570 9840 23626 10300 0 FreeSans 224 90 0 0 S2MID[3]
port 108 nsew signal input
flabel metal2 s 23846 9840 23902 10300 0 FreeSans 224 90 0 0 S2MID[4]
port 109 nsew signal input
flabel metal2 s 24122 9840 24178 10300 0 FreeSans 224 90 0 0 S2MID[5]
port 110 nsew signal input
flabel metal2 s 24398 9840 24454 10300 0 FreeSans 224 90 0 0 S2MID[6]
port 111 nsew signal input
flabel metal2 s 24674 9840 24730 10300 0 FreeSans 224 90 0 0 S2MID[7]
port 112 nsew signal input
flabel metal2 s 24950 9840 25006 10300 0 FreeSans 224 90 0 0 S4END[0]
port 113 nsew signal input
flabel metal2 s 27710 9840 27766 10300 0 FreeSans 224 90 0 0 S4END[10]
port 114 nsew signal input
flabel metal2 s 27986 9840 28042 10300 0 FreeSans 224 90 0 0 S4END[11]
port 115 nsew signal input
flabel metal2 s 28262 9840 28318 10300 0 FreeSans 224 90 0 0 S4END[12]
port 116 nsew signal input
flabel metal2 s 28538 9840 28594 10300 0 FreeSans 224 90 0 0 S4END[13]
port 117 nsew signal input
flabel metal2 s 28814 9840 28870 10300 0 FreeSans 224 90 0 0 S4END[14]
port 118 nsew signal input
flabel metal2 s 29090 9840 29146 10300 0 FreeSans 224 90 0 0 S4END[15]
port 119 nsew signal input
flabel metal2 s 25226 9840 25282 10300 0 FreeSans 224 90 0 0 S4END[1]
port 120 nsew signal input
flabel metal2 s 25502 9840 25558 10300 0 FreeSans 224 90 0 0 S4END[2]
port 121 nsew signal input
flabel metal2 s 25778 9840 25834 10300 0 FreeSans 224 90 0 0 S4END[3]
port 122 nsew signal input
flabel metal2 s 26054 9840 26110 10300 0 FreeSans 224 90 0 0 S4END[4]
port 123 nsew signal input
flabel metal2 s 26330 9840 26386 10300 0 FreeSans 224 90 0 0 S4END[5]
port 124 nsew signal input
flabel metal2 s 26606 9840 26662 10300 0 FreeSans 224 90 0 0 S4END[6]
port 125 nsew signal input
flabel metal2 s 26882 9840 26938 10300 0 FreeSans 224 90 0 0 S4END[7]
port 126 nsew signal input
flabel metal2 s 27158 9840 27214 10300 0 FreeSans 224 90 0 0 S4END[8]
port 127 nsew signal input
flabel metal2 s 27434 9840 27490 10300 0 FreeSans 224 90 0 0 S4END[9]
port 128 nsew signal input
flabel metal2 s 29366 9840 29422 10300 0 FreeSans 224 90 0 0 SS4END[0]
port 129 nsew signal input
flabel metal2 s 32126 9840 32182 10300 0 FreeSans 224 90 0 0 SS4END[10]
port 130 nsew signal input
flabel metal2 s 32402 9840 32458 10300 0 FreeSans 224 90 0 0 SS4END[11]
port 131 nsew signal input
flabel metal2 s 32678 9840 32734 10300 0 FreeSans 224 90 0 0 SS4END[12]
port 132 nsew signal input
flabel metal2 s 32954 9840 33010 10300 0 FreeSans 224 90 0 0 SS4END[13]
port 133 nsew signal input
flabel metal2 s 33230 9840 33286 10300 0 FreeSans 224 90 0 0 SS4END[14]
port 134 nsew signal input
flabel metal2 s 33506 9840 33562 10300 0 FreeSans 224 90 0 0 SS4END[15]
port 135 nsew signal input
flabel metal2 s 29642 9840 29698 10300 0 FreeSans 224 90 0 0 SS4END[1]
port 136 nsew signal input
flabel metal2 s 29918 9840 29974 10300 0 FreeSans 224 90 0 0 SS4END[2]
port 137 nsew signal input
flabel metal2 s 30194 9840 30250 10300 0 FreeSans 224 90 0 0 SS4END[3]
port 138 nsew signal input
flabel metal2 s 30470 9840 30526 10300 0 FreeSans 224 90 0 0 SS4END[4]
port 139 nsew signal input
flabel metal2 s 30746 9840 30802 10300 0 FreeSans 224 90 0 0 SS4END[5]
port 140 nsew signal input
flabel metal2 s 31022 9840 31078 10300 0 FreeSans 224 90 0 0 SS4END[6]
port 141 nsew signal input
flabel metal2 s 31298 9840 31354 10300 0 FreeSans 224 90 0 0 SS4END[7]
port 142 nsew signal input
flabel metal2 s 31574 9840 31630 10300 0 FreeSans 224 90 0 0 SS4END[8]
port 143 nsew signal input
flabel metal2 s 31850 9840 31906 10300 0 FreeSans 224 90 0 0 SS4END[9]
port 144 nsew signal input
flabel metal2 s 1122 -300 1178 160 0 FreeSans 224 90 0 0 UserCLK
port 145 nsew signal input
flabel metal2 s 33782 9840 33838 10300 0 FreeSans 224 90 0 0 UserCLKo
port 146 nsew signal tristate
flabel metal4 s 6245 2128 6565 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 16848 2128 17168 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 27451 2128 27771 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 38054 2128 38374 7664 0 FreeSans 1920 90 0 0 vccd1
port 147 nsew power bidirectional
flabel metal4 s 11546 2128 11866 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 22149 2128 22469 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 32752 2128 33072 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
flabel metal4 s 43355 2128 43675 7664 0 FreeSans 1920 90 0 0 vssd1
port 148 nsew ground bidirectional
rlabel metal1 22310 7072 22310 7072 0 vccd1
rlabel via1 22389 7616 22389 7616 0 vssd1
rlabel metal2 3266 1248 3266 1248 0 FrameStrobe[0]
rlabel metal2 24571 68 24571 68 0 FrameStrobe[10]
rlabel metal2 26542 687 26542 687 0 FrameStrobe[11]
rlabel metal2 28711 68 28711 68 0 FrameStrobe[12]
rlabel metal2 30919 68 30919 68 0 FrameStrobe[13]
rlabel metal2 32890 738 32890 738 0 FrameStrobe[14]
rlabel metal2 35151 68 35151 68 0 FrameStrobe[15]
rlabel metal2 37122 1299 37122 1299 0 FrameStrobe[16]
rlabel metal2 39238 143 39238 143 0 FrameStrobe[17]
rlabel metal2 41354 755 41354 755 0 FrameStrobe[18]
rlabel metal2 43325 68 43325 68 0 FrameStrobe[19]
rlabel metal2 5435 68 5435 68 0 FrameStrobe[1]
rlabel metal2 7551 68 7551 68 0 FrameStrobe[2]
rlabel metal2 9614 755 9614 755 0 FrameStrobe[3]
rlabel metal2 11875 68 11875 68 0 FrameStrobe[4]
rlabel metal2 13846 1248 13846 1248 0 FrameStrobe[5]
rlabel metal2 16107 68 16107 68 0 FrameStrobe[6]
rlabel metal2 18223 68 18223 68 0 FrameStrobe[7]
rlabel metal2 20339 68 20339 68 0 FrameStrobe[8]
rlabel metal2 22310 143 22310 143 0 FrameStrobe[9]
rlabel metal2 34362 8680 34362 8680 0 FrameStrobe_O[0]
rlabel metal1 37490 6834 37490 6834 0 FrameStrobe_O[10]
rlabel metal1 38134 6834 38134 6834 0 FrameStrobe_O[11]
rlabel metal1 37950 6630 37950 6630 0 FrameStrobe_O[12]
rlabel metal1 38548 6426 38548 6426 0 FrameStrobe_O[13]
rlabel metal1 38594 6630 38594 6630 0 FrameStrobe_O[14]
rlabel metal1 38686 6698 38686 6698 0 FrameStrobe_O[15]
rlabel metal2 38778 9173 38778 9173 0 FrameStrobe_O[16]
rlabel metal1 39560 6766 39560 6766 0 FrameStrobe_O[17]
rlabel metal2 39330 8680 39330 8680 0 FrameStrobe_O[18]
rlabel metal1 40204 6834 40204 6834 0 FrameStrobe_O[19]
rlabel metal2 34638 8646 34638 8646 0 FrameStrobe_O[1]
rlabel metal2 34914 9173 34914 9173 0 FrameStrobe_O[2]
rlabel metal1 35420 6834 35420 6834 0 FrameStrobe_O[3]
rlabel metal2 35466 9241 35466 9241 0 FrameStrobe_O[4]
rlabel metal1 35972 6834 35972 6834 0 FrameStrobe_O[5]
rlabel metal1 36294 6630 36294 6630 0 FrameStrobe_O[6]
rlabel metal2 36294 9173 36294 9173 0 FrameStrobe_O[7]
rlabel metal1 36892 6630 36892 6630 0 FrameStrobe_O[8]
rlabel metal2 36846 9173 36846 9173 0 FrameStrobe_O[9]
rlabel metal2 5106 9037 5106 9037 0 N1BEG[0]
rlabel metal1 5198 7514 5198 7514 0 N1BEG[1]
rlabel metal2 5658 9037 5658 9037 0 N1BEG[2]
rlabel metal1 5750 7514 5750 7514 0 N1BEG[3]
rlabel metal2 6210 9037 6210 9037 0 N2BEG[0]
rlabel metal1 6302 7310 6302 7310 0 N2BEG[1]
rlabel metal2 6762 8136 6762 8136 0 N2BEG[2]
rlabel metal2 7038 8340 7038 8340 0 N2BEG[3]
rlabel metal1 7176 7514 7176 7514 0 N2BEG[4]
rlabel metal2 7590 8340 7590 8340 0 N2BEG[5]
rlabel metal1 7728 7514 7728 7514 0 N2BEG[6]
rlabel metal2 8142 8340 8142 8340 0 N2BEG[7]
rlabel metal1 8280 7514 8280 7514 0 N2BEGb[0]
rlabel metal2 8694 8340 8694 8340 0 N2BEGb[1]
rlabel metal1 8832 7514 8832 7514 0 N2BEGb[2]
rlabel metal2 9246 8136 9246 8136 0 N2BEGb[3]
rlabel metal2 9522 7864 9522 7864 0 N2BEGb[4]
rlabel metal2 9798 8136 9798 8136 0 N2BEGb[5]
rlabel metal1 9844 6834 9844 6834 0 N2BEGb[6]
rlabel metal2 10350 8136 10350 8136 0 N2BEGb[7]
rlabel metal1 10396 6834 10396 6834 0 N4BEG[0]
rlabel metal2 13386 8340 13386 8340 0 N4BEG[10]
rlabel metal1 13478 7514 13478 7514 0 N4BEG[11]
rlabel metal2 13938 8136 13938 8136 0 N4BEG[12]
rlabel metal1 14030 7514 14030 7514 0 N4BEG[13]
rlabel metal2 14490 9037 14490 9037 0 N4BEG[14]
rlabel metal2 14766 8340 14766 8340 0 N4BEG[15]
rlabel metal2 10902 8408 10902 8408 0 N4BEG[1]
rlabel metal1 10902 7514 10902 7514 0 N4BEG[2]
rlabel metal2 11454 8408 11454 8408 0 N4BEG[3]
rlabel metal1 11454 7310 11454 7310 0 N4BEG[4]
rlabel metal2 12006 8408 12006 8408 0 N4BEG[5]
rlabel metal2 12282 8136 12282 8136 0 N4BEG[6]
rlabel metal2 12558 8680 12558 8680 0 N4BEG[7]
rlabel metal2 12834 8340 12834 8340 0 N4BEG[8]
rlabel metal1 12834 6732 12834 6732 0 N4BEG[9]
rlabel metal1 14904 7514 14904 7514 0 NN4BEG[0]
rlabel metal2 17802 9173 17802 9173 0 NN4BEG[10]
rlabel metal2 18078 8340 18078 8340 0 NN4BEG[11]
rlabel metal2 18354 9173 18354 9173 0 NN4BEG[12]
rlabel metal2 18630 9173 18630 9173 0 NN4BEG[13]
rlabel metal2 18906 8646 18906 8646 0 NN4BEG[14]
rlabel metal2 19182 8680 19182 8680 0 NN4BEG[15]
rlabel metal2 15318 8340 15318 8340 0 NN4BEG[1]
rlabel metal1 15456 7514 15456 7514 0 NN4BEG[2]
rlabel metal2 15870 8340 15870 8340 0 NN4BEG[3]
rlabel metal1 15962 7514 15962 7514 0 NN4BEG[4]
rlabel metal2 16422 8340 16422 8340 0 NN4BEG[5]
rlabel metal1 16606 7378 16606 7378 0 NN4BEG[6]
rlabel metal2 16974 9037 16974 9037 0 NN4BEG[7]
rlabel metal2 17250 9173 17250 9173 0 NN4BEG[8]
rlabel metal2 17526 8340 17526 8340 0 NN4BEG[9]
rlabel metal2 19458 8306 19458 8306 0 S1END[0]
rlabel metal2 19734 9105 19734 9105 0 S1END[1]
rlabel metal2 20010 9105 20010 9105 0 S1END[2]
rlabel metal2 20286 9785 20286 9785 0 S1END[3]
rlabel metal2 20562 9105 20562 9105 0 S2END[0]
rlabel metal2 20838 9105 20838 9105 0 S2END[1]
rlabel metal2 21114 8612 21114 8612 0 S2END[2]
rlabel metal2 21390 9105 21390 9105 0 S2END[3]
rlabel metal2 21666 8612 21666 8612 0 S2END[4]
rlabel metal2 21942 8306 21942 8306 0 S2END[5]
rlabel metal2 22218 9241 22218 9241 0 S2END[6]
rlabel metal2 22494 9309 22494 9309 0 S2END[7]
rlabel metal2 22770 8612 22770 8612 0 S2MID[0]
rlabel metal2 23046 8612 23046 8612 0 S2MID[1]
rlabel metal2 23322 8612 23322 8612 0 S2MID[2]
rlabel metal2 23598 8833 23598 8833 0 S2MID[3]
rlabel metal2 23874 9241 23874 9241 0 S2MID[4]
rlabel metal2 24150 9241 24150 9241 0 S2MID[5]
rlabel metal2 24426 8646 24426 8646 0 S2MID[6]
rlabel metal2 24702 8680 24702 8680 0 S2MID[7]
rlabel metal2 24978 9054 24978 9054 0 S4END[0]
rlabel metal2 27738 8918 27738 8918 0 S4END[10]
rlabel metal2 28014 9241 28014 9241 0 S4END[11]
rlabel metal2 28290 9309 28290 9309 0 S4END[12]
rlabel metal2 28566 9105 28566 9105 0 S4END[13]
rlabel metal2 28842 9241 28842 9241 0 S4END[14]
rlabel metal2 29118 8544 29118 8544 0 S4END[15]
rlabel metal2 25254 9020 25254 9020 0 S4END[1]
rlabel metal2 25530 8612 25530 8612 0 S4END[2]
rlabel metal2 25806 9241 25806 9241 0 S4END[3]
rlabel metal2 26082 9309 26082 9309 0 S4END[4]
rlabel metal2 26358 9241 26358 9241 0 S4END[5]
rlabel metal2 26634 9241 26634 9241 0 S4END[6]
rlabel metal2 26910 9309 26910 9309 0 S4END[7]
rlabel metal2 27186 9377 27186 9377 0 S4END[8]
rlabel metal2 27462 9445 27462 9445 0 S4END[9]
rlabel metal2 29394 9241 29394 9241 0 SS4END[0]
rlabel metal2 32154 9173 32154 9173 0 SS4END[10]
rlabel metal2 32430 9241 32430 9241 0 SS4END[11]
rlabel metal2 32706 8629 32706 8629 0 SS4END[12]
rlabel metal2 32982 8782 32982 8782 0 SS4END[13]
rlabel metal2 33350 6833 33350 6833 0 SS4END[14]
rlabel metal2 33626 6833 33626 6833 0 SS4END[15]
rlabel metal2 29670 8969 29670 8969 0 SS4END[1]
rlabel metal2 29946 9173 29946 9173 0 SS4END[2]
rlabel metal2 30222 9241 30222 9241 0 SS4END[3]
rlabel metal2 30498 8680 30498 8680 0 SS4END[4]
rlabel metal2 30774 8578 30774 8578 0 SS4END[5]
rlabel metal1 31786 7412 31786 7412 0 SS4END[6]
rlabel metal1 32016 7378 32016 7378 0 SS4END[7]
rlabel metal1 32430 7446 32430 7446 0 SS4END[8]
rlabel metal2 31878 9241 31878 9241 0 SS4END[9]
rlabel metal2 1150 1248 1150 1248 0 UserCLK
rlabel metal2 33810 8680 33810 8680 0 UserCLKo
rlabel metal2 4094 2244 4094 2244 0 net1
rlabel metal1 40894 2414 40894 2414 0 net10
rlabel metal2 9706 5899 9706 5899 0 net100
rlabel metal2 7222 7480 7222 7480 0 net101
rlabel metal2 19826 5542 19826 5542 0 net102
rlabel metal3 16284 8092 16284 8092 0 net103
rlabel metal2 15134 8211 15134 8211 0 net104
rlabel metal2 13754 6987 13754 6987 0 net105
rlabel metal1 20746 7174 20746 7174 0 net106
rlabel metal1 8418 6732 8418 6732 0 net107
rlabel metal1 21344 6630 21344 6630 0 net108
rlabel via2 20010 6613 20010 6613 0 net109
rlabel metal1 42826 2414 42826 2414 0 net11
rlabel metal1 10396 5678 10396 5678 0 net110
rlabel metal1 12926 6324 12926 6324 0 net111
rlabel metal2 10718 6528 10718 6528 0 net112
rlabel metal1 10074 6290 10074 6290 0 net113
rlabel metal2 10626 5967 10626 5967 0 net114
rlabel metal2 16790 5780 16790 5780 0 net115
rlabel metal2 16514 7633 16514 7633 0 net116
rlabel metal2 15410 5814 15410 5814 0 net117
rlabel metal2 15962 7633 15962 7633 0 net118
rlabel metal2 14398 7378 14398 7378 0 net119
rlabel metal2 5658 3060 5658 3060 0 net12
rlabel metal2 18446 6885 18446 6885 0 net120
rlabel metal2 10810 5848 10810 5848 0 net121
rlabel metal1 10304 7514 10304 7514 0 net122
rlabel metal2 12650 5916 12650 5916 0 net123
rlabel metal1 12558 8058 12558 8058 0 net124
rlabel metal2 15134 5406 15134 5406 0 net125
rlabel metal2 12466 5542 12466 5542 0 net126
rlabel metal2 12650 7786 12650 7786 0 net127
rlabel metal2 14214 5729 14214 5729 0 net128
rlabel metal2 17250 5542 17250 5542 0 net129
rlabel metal1 7774 1972 7774 1972 0 net13
rlabel metal1 14766 6154 14766 6154 0 net130
rlabel metal1 17986 6426 17986 6426 0 net131
rlabel metal1 18354 6426 18354 6426 0 net132
rlabel metal1 18676 6426 18676 6426 0 net133
rlabel metal1 18814 6970 18814 6970 0 net134
rlabel metal1 19550 6086 19550 6086 0 net135
rlabel metal1 19458 6426 19458 6426 0 net136
rlabel metal1 14950 6426 14950 6426 0 net137
rlabel metal1 14812 7378 14812 7378 0 net138
rlabel metal1 15502 6392 15502 6392 0 net139
rlabel metal2 9890 2176 9890 2176 0 net14
rlabel metal1 15778 6426 15778 6426 0 net140
rlabel metal1 16468 6426 16468 6426 0 net141
rlabel metal1 16422 7446 16422 7446 0 net142
rlabel metal1 17020 6426 17020 6426 0 net143
rlabel metal1 17204 6154 17204 6154 0 net144
rlabel metal1 17664 6426 17664 6426 0 net145
rlabel metal1 33166 2584 33166 2584 0 net146
rlabel metal1 34224 6834 34224 6834 0 net147
rlabel metal1 12282 2312 12282 2312 0 net15
rlabel metal1 14582 2312 14582 2312 0 net16
rlabel metal1 16376 2618 16376 2618 0 net17
rlabel metal1 18400 2618 18400 2618 0 net18
rlabel metal1 20516 2618 20516 2618 0 net19
rlabel metal1 24748 2618 24748 2618 0 net2
rlabel metal1 22540 2618 22540 2618 0 net20
rlabel metal1 16192 6902 16192 6902 0 net21
rlabel metal1 6578 6188 6578 6188 0 net22
rlabel metal1 17342 5848 17342 5848 0 net23
rlabel metal1 16514 5678 16514 5678 0 net24
rlabel metal2 20654 6069 20654 6069 0 net25
rlabel metal1 18354 6664 18354 6664 0 net26
rlabel metal1 13110 6324 13110 6324 0 net27
rlabel metal1 21666 6664 21666 6664 0 net28
rlabel metal1 19826 6732 19826 6732 0 net29
rlabel metal1 37030 7378 37030 7378 0 net3
rlabel metal1 21206 6800 21206 6800 0 net30
rlabel metal1 20378 7412 20378 7412 0 net31
rlabel metal1 21114 7276 21114 7276 0 net32
rlabel metal1 21206 7344 21206 7344 0 net33
rlabel metal1 22310 6834 22310 6834 0 net34
rlabel metal1 22678 6732 22678 6732 0 net35
rlabel metal1 22954 6800 22954 6800 0 net36
rlabel metal1 22862 7412 22862 7412 0 net37
rlabel viali 23230 6292 23230 6292 0 net38
rlabel metal1 23874 6324 23874 6324 0 net39
rlabel metal1 37490 2006 37490 2006 0 net4
rlabel metal1 24748 6290 24748 6290 0 net40
rlabel metal1 24978 7344 24978 7344 0 net41
rlabel metal1 27830 6800 27830 6800 0 net42
rlabel metal1 28566 6766 28566 6766 0 net43
rlabel metal1 29072 6766 29072 6766 0 net44
rlabel metal1 29578 6732 29578 6732 0 net45
rlabel metal1 29808 6766 29808 6766 0 net46
rlabel metal1 30084 6766 30084 6766 0 net47
rlabel metal1 25530 7412 25530 7412 0 net48
rlabel metal1 25070 6834 25070 6834 0 net49
rlabel metal1 36846 2040 36846 2040 0 net5
rlabel metal1 25346 6800 25346 6800 0 net50
rlabel metal1 25806 6732 25806 6732 0 net51
rlabel metal1 26174 6800 26174 6800 0 net52
rlabel metal1 26542 6732 26542 6732 0 net53
rlabel metal1 27048 6766 27048 6766 0 net54
rlabel metal1 27278 6800 27278 6800 0 net55
rlabel metal1 27554 6732 27554 6732 0 net56
rlabel metal1 23138 6324 23138 6324 0 net57
rlabel metal1 33258 7242 33258 7242 0 net58
rlabel metal1 33534 7174 33534 7174 0 net59
rlabel metal1 33488 2618 33488 2618 0 net6
rlabel metal2 33718 7956 33718 7956 0 net60
rlabel metal2 33258 6681 33258 6681 0 net61
rlabel metal2 33534 5865 33534 5865 0 net62
rlabel metal2 33810 6477 33810 6477 0 net63
rlabel metal2 19366 5916 19366 5916 0 net64
rlabel metal1 21022 6902 21022 6902 0 net65
rlabel metal1 19274 6222 19274 6222 0 net66
rlabel metal2 18630 6018 18630 6018 0 net67
rlabel metal2 18354 6868 18354 6868 0 net68
rlabel metal1 32062 7174 32062 7174 0 net69
rlabel metal1 35742 2380 35742 2380 0 net7
rlabel metal2 32338 6664 32338 6664 0 net70
rlabel via2 31786 7259 31786 7259 0 net71
rlabel metal1 32660 7174 32660 7174 0 net72
rlabel metal1 1702 1904 1702 1904 0 net73
rlabel metal1 33994 2618 33994 2618 0 net74
rlabel metal2 36754 6596 36754 6596 0 net75
rlabel metal1 38502 7480 38502 7480 0 net76
rlabel metal1 37536 2618 37536 2618 0 net77
rlabel metal1 38180 2550 38180 2550 0 net78
rlabel metal1 37214 3128 37214 3128 0 net79
rlabel metal2 37858 2822 37858 2822 0 net8
rlabel metal1 38962 2312 38962 2312 0 net80
rlabel metal1 38226 3162 38226 3162 0 net81
rlabel metal1 39514 2618 39514 2618 0 net82
rlabel metal1 40342 2618 40342 2618 0 net83
rlabel metal1 41906 2618 41906 2618 0 net84
rlabel metal1 34224 3706 34224 3706 0 net85
rlabel metal1 35926 7310 35926 7310 0 net86
rlabel metal1 35052 2618 35052 2618 0 net87
rlabel metal1 36294 7378 36294 7378 0 net88
rlabel metal2 35926 5304 35926 5304 0 net89
rlabel metal1 39284 2414 39284 2414 0 net9
rlabel metal2 33718 4828 33718 4828 0 net90
rlabel metal2 37306 4963 37306 4963 0 net91
rlabel metal1 37030 6392 37030 6392 0 net92
rlabel metal2 37950 3077 37950 3077 0 net93
rlabel metal1 4738 6766 4738 6766 0 net94
rlabel metal1 5658 6154 5658 6154 0 net95
rlabel metal1 6026 6426 6026 6426 0 net96
rlabel metal1 5842 7446 5842 7446 0 net97
rlabel metal3 12420 6800 12420 6800 0 net98
rlabel metal2 5842 6783 5842 6783 0 net99
<< properties >>
string FIXED_BBOX 0 0 44700 10000
<< end >>
