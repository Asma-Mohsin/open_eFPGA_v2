VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BlockRAM_1KB
  CLASS BLOCK ;
  FOREIGN BlockRAM_1KB ;
  ORIGIN 0.000 0.000 ;
  SIZE 575.000 BY 450.000 ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.790 4.000 99.090 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 4.000 103.850 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 4.000 108.610 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.070 4.000 113.370 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.230 4.000 308.530 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.990 4.000 313.290 ;
    END
  END C5
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 287.200 0.000 287.340 4.000 ;
    END
  END clk
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.830 4.000 118.130 ;
    END
  END rd_addr[0]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.590 4.000 122.890 ;
    END
  END rd_addr[1]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.350 4.000 127.650 ;
    END
  END rd_addr[2]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.110 4.000 132.410 ;
    END
  END rd_addr[3]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.870 4.000 137.170 ;
    END
  END rd_addr[4]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 4.000 141.930 ;
    END
  END rd_addr[5]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.390 4.000 146.690 ;
    END
  END rd_addr[6]
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.150 4.000 151.450 ;
    END
  END rd_addr[7]
  PIN rd_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.630 4.000 22.930 ;
    END
  END rd_data[0]
  PIN rd_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 4.000 70.530 ;
    END
  END rd_data[10]
  PIN rd_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.990 4.000 75.290 ;
    END
  END rd_data[11]
  PIN rd_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.750 4.000 80.050 ;
    END
  END rd_data[12]
  PIN rd_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 4.000 84.810 ;
    END
  END rd_data[13]
  PIN rd_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 4.000 89.570 ;
    END
  END rd_data[14]
  PIN rd_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.030 4.000 94.330 ;
    END
  END rd_data[15]
  PIN rd_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.070 4.000 232.370 ;
    END
  END rd_data[16]
  PIN rd_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.830 4.000 237.130 ;
    END
  END rd_data[17]
  PIN rd_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.590 4.000 241.890 ;
    END
  END rd_data[18]
  PIN rd_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.350 4.000 246.650 ;
    END
  END rd_data[19]
  PIN rd_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.390 4.000 27.690 ;
    END
  END rd_data[1]
  PIN rd_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.110 4.000 251.410 ;
    END
  END rd_data[20]
  PIN rd_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.870 4.000 256.170 ;
    END
  END rd_data[21]
  PIN rd_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.630 4.000 260.930 ;
    END
  END rd_data[22]
  PIN rd_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.390 4.000 265.690 ;
    END
  END rd_data[23]
  PIN rd_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.150 4.000 270.450 ;
    END
  END rd_data[24]
  PIN rd_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.910 4.000 275.210 ;
    END
  END rd_data[25]
  PIN rd_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.670 4.000 279.970 ;
    END
  END rd_data[26]
  PIN rd_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.430 4.000 284.730 ;
    END
  END rd_data[27]
  PIN rd_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.190 4.000 289.490 ;
    END
  END rd_data[28]
  PIN rd_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.950 4.000 294.250 ;
    END
  END rd_data[29]
  PIN rd_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.150 4.000 32.450 ;
    END
  END rd_data[2]
  PIN rd_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.710 4.000 299.010 ;
    END
  END rd_data[30]
  PIN rd_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.470 4.000 303.770 ;
    END
  END rd_data[31]
  PIN rd_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.910 4.000 37.210 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.670 4.000 41.970 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.430 4.000 46.730 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.190 4.000 51.490 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.950 4.000 56.250 ;
    END
  END rd_data[7]
  PIN rd_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.710 4.000 61.010 ;
    END
  END rd_data[8]
  PIN rd_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.470 4.000 65.770 ;
    END
  END rd_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 -2.160 -0.480 450.960 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 -2.160 577.080 -0.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 449.360 577.080 450.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.480 -2.160 577.080 450.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.020 -5.460 19.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 -5.460 39.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 -5.460 59.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.020 -5.460 79.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.020 432.480 79.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.020 -5.460 99.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.020 432.480 99.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.020 -5.460 119.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.020 432.480 119.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 -5.460 139.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 432.480 139.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.020 -5.460 159.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.020 432.480 159.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 178.020 -5.460 179.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 178.020 432.480 179.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 198.020 -5.460 199.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 198.020 432.480 199.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.020 -5.460 219.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.020 433.100 219.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 -5.460 239.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 432.480 239.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.020 -5.460 259.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.020 432.480 259.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.020 -5.460 279.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.020 433.100 279.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 298.020 -5.460 299.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 298.020 433.100 299.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.020 -5.460 319.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.020 433.100 319.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 -5.460 339.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 432.480 339.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.020 -5.460 359.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.020 432.480 359.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.020 -5.460 379.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.020 433.100 379.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 398.020 -5.460 399.620 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 398.020 433.100 399.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.020 -5.460 419.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.020 432.480 419.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.020 -5.460 439.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 438.020 432.480 439.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.020 -5.460 459.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.020 432.480 459.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 478.020 -5.460 479.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 478.020 432.480 479.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.020 -5.460 499.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.020 432.480 499.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.020 -5.460 519.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 518.020 433.100 519.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 538.020 -5.460 539.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 538.020 432.480 539.620 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.020 -5.460 559.620 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.020 432.480 559.620 454.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 27.940 580.380 29.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 417.940 580.380 419.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 561.780 10.640 563.380 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -5.460 -3.780 454.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -5.460 580.380 -3.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 452.660 580.380 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 578.780 -5.460 580.380 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.720 -5.460 16.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 -5.460 36.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.720 -5.460 56.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.720 -5.460 76.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.720 432.480 76.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.720 -5.460 96.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.720 432.480 96.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 -5.460 116.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 432.480 116.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 -5.460 136.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 432.480 136.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.720 -5.460 156.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.720 432.480 156.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.720 -5.460 176.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.720 432.480 176.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 194.720 -5.460 196.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 194.720 432.480 196.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.720 -5.460 216.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.720 432.480 216.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 -5.460 236.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 433.100 236.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.720 -5.460 256.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.720 433.100 256.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.720 -5.460 276.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.720 432.480 276.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.720 -5.460 296.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.720 432.480 296.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.720 -5.460 316.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.720 432.480 316.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 -5.460 336.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 433.100 336.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.720 -5.460 356.320 14.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.720 433.100 356.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.720 -5.460 376.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.720 432.480 376.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.720 -5.460 396.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.720 432.480 396.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.720 -5.460 416.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.720 432.480 416.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.720 -5.460 436.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.720 432.480 436.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.720 -5.460 456.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.720 432.480 456.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.720 -5.460 476.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.720 432.480 476.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.720 -5.460 496.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.720 432.480 496.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.720 -5.460 516.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.720 432.480 516.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.720 -5.460 536.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.720 432.480 536.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.720 -5.460 556.320 15.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.720 432.480 556.320 454.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 24.640 580.380 26.240 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 414.640 580.380 416.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.460 10.640 567.060 438.160 ;
    END
  END vssd1
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.750 4.000 318.050 ;
    END
  END wr_addr[0]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.510 4.000 322.810 ;
    END
  END wr_addr[1]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.270 4.000 327.570 ;
    END
  END wr_addr[2]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.030 4.000 332.330 ;
    END
  END wr_addr[3]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.790 4.000 337.090 ;
    END
  END wr_addr[4]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.550 4.000 341.850 ;
    END
  END wr_addr[5]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.310 4.000 346.610 ;
    END
  END wr_addr[6]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.070 4.000 351.370 ;
    END
  END wr_addr[7]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 4.000 156.210 ;
    END
  END wr_data[0]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.510 4.000 203.810 ;
    END
  END wr_data[10]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.270 4.000 208.570 ;
    END
  END wr_data[11]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 4.000 213.330 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.790 4.000 218.090 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.550 4.000 222.850 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.310 4.000 227.610 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.830 4.000 356.130 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.590 4.000 360.890 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.350 4.000 365.650 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.110 4.000 370.410 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.670 4.000 160.970 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.870 4.000 375.170 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.630 4.000 379.930 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.390 4.000 384.690 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.150 4.000 389.450 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.910 4.000 394.210 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.670 4.000 398.970 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.430 4.000 403.730 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.190 4.000 408.490 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.950 4.000 413.250 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.710 4.000 418.010 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.430 4.000 165.730 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.470 4.000 422.770 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.230 4.000 427.530 ;
    END
  END wr_data[31]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.190 4.000 170.490 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.950 4.000 175.250 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.710 4.000 180.010 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.470 4.000 184.770 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.230 4.000 189.530 ;
    END
  END wr_data[7]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.990 4.000 194.290 ;
    END
  END wr_data[8]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.750 4.000 199.050 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 569.480 443.445 ;
      LAYER met1 ;
        RECT 4.670 2.420 569.480 443.600 ;
      LAYER met2 ;
        RECT 4.690 4.280 567.030 443.545 ;
        RECT 4.690 2.390 286.920 4.280 ;
        RECT 287.620 2.390 567.030 4.280 ;
      LAYER met3 ;
        RECT 3.070 427.930 567.050 443.525 ;
        RECT 4.400 426.830 567.050 427.930 ;
        RECT 3.070 423.170 567.050 426.830 ;
        RECT 4.400 422.070 567.050 423.170 ;
        RECT 3.070 418.410 567.050 422.070 ;
        RECT 4.400 417.310 567.050 418.410 ;
        RECT 3.070 413.650 567.050 417.310 ;
        RECT 4.400 412.550 567.050 413.650 ;
        RECT 3.070 408.890 567.050 412.550 ;
        RECT 4.400 407.790 567.050 408.890 ;
        RECT 3.070 404.130 567.050 407.790 ;
        RECT 4.400 403.030 567.050 404.130 ;
        RECT 3.070 399.370 567.050 403.030 ;
        RECT 4.400 398.270 567.050 399.370 ;
        RECT 3.070 394.610 567.050 398.270 ;
        RECT 4.400 393.510 567.050 394.610 ;
        RECT 3.070 389.850 567.050 393.510 ;
        RECT 4.400 388.750 567.050 389.850 ;
        RECT 3.070 385.090 567.050 388.750 ;
        RECT 4.400 383.990 567.050 385.090 ;
        RECT 3.070 380.330 567.050 383.990 ;
        RECT 4.400 379.230 567.050 380.330 ;
        RECT 3.070 375.570 567.050 379.230 ;
        RECT 4.400 374.470 567.050 375.570 ;
        RECT 3.070 370.810 567.050 374.470 ;
        RECT 4.400 369.710 567.050 370.810 ;
        RECT 3.070 366.050 567.050 369.710 ;
        RECT 4.400 364.950 567.050 366.050 ;
        RECT 3.070 361.290 567.050 364.950 ;
        RECT 4.400 360.190 567.050 361.290 ;
        RECT 3.070 356.530 567.050 360.190 ;
        RECT 4.400 355.430 567.050 356.530 ;
        RECT 3.070 351.770 567.050 355.430 ;
        RECT 4.400 350.670 567.050 351.770 ;
        RECT 3.070 347.010 567.050 350.670 ;
        RECT 4.400 345.910 567.050 347.010 ;
        RECT 3.070 342.250 567.050 345.910 ;
        RECT 4.400 341.150 567.050 342.250 ;
        RECT 3.070 337.490 567.050 341.150 ;
        RECT 4.400 336.390 567.050 337.490 ;
        RECT 3.070 332.730 567.050 336.390 ;
        RECT 4.400 331.630 567.050 332.730 ;
        RECT 3.070 327.970 567.050 331.630 ;
        RECT 4.400 326.870 567.050 327.970 ;
        RECT 3.070 323.210 567.050 326.870 ;
        RECT 4.400 322.110 567.050 323.210 ;
        RECT 3.070 318.450 567.050 322.110 ;
        RECT 4.400 317.350 567.050 318.450 ;
        RECT 3.070 313.690 567.050 317.350 ;
        RECT 4.400 312.590 567.050 313.690 ;
        RECT 3.070 308.930 567.050 312.590 ;
        RECT 4.400 307.830 567.050 308.930 ;
        RECT 3.070 304.170 567.050 307.830 ;
        RECT 4.400 303.070 567.050 304.170 ;
        RECT 3.070 299.410 567.050 303.070 ;
        RECT 4.400 298.310 567.050 299.410 ;
        RECT 3.070 294.650 567.050 298.310 ;
        RECT 4.400 293.550 567.050 294.650 ;
        RECT 3.070 289.890 567.050 293.550 ;
        RECT 4.400 288.790 567.050 289.890 ;
        RECT 3.070 285.130 567.050 288.790 ;
        RECT 4.400 284.030 567.050 285.130 ;
        RECT 3.070 280.370 567.050 284.030 ;
        RECT 4.400 279.270 567.050 280.370 ;
        RECT 3.070 275.610 567.050 279.270 ;
        RECT 4.400 274.510 567.050 275.610 ;
        RECT 3.070 270.850 567.050 274.510 ;
        RECT 4.400 269.750 567.050 270.850 ;
        RECT 3.070 266.090 567.050 269.750 ;
        RECT 4.400 264.990 567.050 266.090 ;
        RECT 3.070 261.330 567.050 264.990 ;
        RECT 4.400 260.230 567.050 261.330 ;
        RECT 3.070 256.570 567.050 260.230 ;
        RECT 4.400 255.470 567.050 256.570 ;
        RECT 3.070 251.810 567.050 255.470 ;
        RECT 4.400 250.710 567.050 251.810 ;
        RECT 3.070 247.050 567.050 250.710 ;
        RECT 4.400 245.950 567.050 247.050 ;
        RECT 3.070 242.290 567.050 245.950 ;
        RECT 4.400 241.190 567.050 242.290 ;
        RECT 3.070 237.530 567.050 241.190 ;
        RECT 4.400 236.430 567.050 237.530 ;
        RECT 3.070 232.770 567.050 236.430 ;
        RECT 4.400 231.670 567.050 232.770 ;
        RECT 3.070 228.010 567.050 231.670 ;
        RECT 4.400 226.910 567.050 228.010 ;
        RECT 3.070 223.250 567.050 226.910 ;
        RECT 4.400 222.150 567.050 223.250 ;
        RECT 3.070 218.490 567.050 222.150 ;
        RECT 4.400 217.390 567.050 218.490 ;
        RECT 3.070 213.730 567.050 217.390 ;
        RECT 4.400 212.630 567.050 213.730 ;
        RECT 3.070 208.970 567.050 212.630 ;
        RECT 4.400 207.870 567.050 208.970 ;
        RECT 3.070 204.210 567.050 207.870 ;
        RECT 4.400 203.110 567.050 204.210 ;
        RECT 3.070 199.450 567.050 203.110 ;
        RECT 4.400 198.350 567.050 199.450 ;
        RECT 3.070 194.690 567.050 198.350 ;
        RECT 4.400 193.590 567.050 194.690 ;
        RECT 3.070 189.930 567.050 193.590 ;
        RECT 4.400 188.830 567.050 189.930 ;
        RECT 3.070 185.170 567.050 188.830 ;
        RECT 4.400 184.070 567.050 185.170 ;
        RECT 3.070 180.410 567.050 184.070 ;
        RECT 4.400 179.310 567.050 180.410 ;
        RECT 3.070 175.650 567.050 179.310 ;
        RECT 4.400 174.550 567.050 175.650 ;
        RECT 3.070 170.890 567.050 174.550 ;
        RECT 4.400 169.790 567.050 170.890 ;
        RECT 3.070 166.130 567.050 169.790 ;
        RECT 4.400 165.030 567.050 166.130 ;
        RECT 3.070 161.370 567.050 165.030 ;
        RECT 4.400 160.270 567.050 161.370 ;
        RECT 3.070 156.610 567.050 160.270 ;
        RECT 4.400 155.510 567.050 156.610 ;
        RECT 3.070 151.850 567.050 155.510 ;
        RECT 4.400 150.750 567.050 151.850 ;
        RECT 3.070 147.090 567.050 150.750 ;
        RECT 4.400 145.990 567.050 147.090 ;
        RECT 3.070 142.330 567.050 145.990 ;
        RECT 4.400 141.230 567.050 142.330 ;
        RECT 3.070 137.570 567.050 141.230 ;
        RECT 4.400 136.470 567.050 137.570 ;
        RECT 3.070 132.810 567.050 136.470 ;
        RECT 4.400 131.710 567.050 132.810 ;
        RECT 3.070 128.050 567.050 131.710 ;
        RECT 4.400 126.950 567.050 128.050 ;
        RECT 3.070 123.290 567.050 126.950 ;
        RECT 4.400 122.190 567.050 123.290 ;
        RECT 3.070 118.530 567.050 122.190 ;
        RECT 4.400 117.430 567.050 118.530 ;
        RECT 3.070 113.770 567.050 117.430 ;
        RECT 4.400 112.670 567.050 113.770 ;
        RECT 3.070 109.010 567.050 112.670 ;
        RECT 4.400 107.910 567.050 109.010 ;
        RECT 3.070 104.250 567.050 107.910 ;
        RECT 4.400 103.150 567.050 104.250 ;
        RECT 3.070 99.490 567.050 103.150 ;
        RECT 4.400 98.390 567.050 99.490 ;
        RECT 3.070 94.730 567.050 98.390 ;
        RECT 4.400 93.630 567.050 94.730 ;
        RECT 3.070 89.970 567.050 93.630 ;
        RECT 4.400 88.870 567.050 89.970 ;
        RECT 3.070 85.210 567.050 88.870 ;
        RECT 4.400 84.110 567.050 85.210 ;
        RECT 3.070 80.450 567.050 84.110 ;
        RECT 4.400 79.350 567.050 80.450 ;
        RECT 3.070 75.690 567.050 79.350 ;
        RECT 4.400 74.590 567.050 75.690 ;
        RECT 3.070 70.930 567.050 74.590 ;
        RECT 4.400 69.830 567.050 70.930 ;
        RECT 3.070 66.170 567.050 69.830 ;
        RECT 4.400 65.070 567.050 66.170 ;
        RECT 3.070 61.410 567.050 65.070 ;
        RECT 4.400 60.310 567.050 61.410 ;
        RECT 3.070 56.650 567.050 60.310 ;
        RECT 4.400 55.550 567.050 56.650 ;
        RECT 3.070 51.890 567.050 55.550 ;
        RECT 4.400 50.790 567.050 51.890 ;
        RECT 3.070 47.130 567.050 50.790 ;
        RECT 4.400 46.030 567.050 47.130 ;
        RECT 3.070 42.370 567.050 46.030 ;
        RECT 4.400 41.270 567.050 42.370 ;
        RECT 3.070 37.610 567.050 41.270 ;
        RECT 4.400 36.510 567.050 37.610 ;
        RECT 3.070 32.850 567.050 36.510 ;
        RECT 4.400 31.750 567.050 32.850 ;
        RECT 3.070 28.090 567.050 31.750 ;
        RECT 4.400 26.990 567.050 28.090 ;
        RECT 3.070 23.330 567.050 26.990 ;
        RECT 4.400 22.230 567.050 23.330 ;
        RECT 3.070 5.275 567.050 22.230 ;
      LAYER met4 ;
        RECT 52.735 6.295 54.320 439.105 ;
        RECT 56.720 6.295 57.620 439.105 ;
        RECT 60.020 432.080 74.320 439.105 ;
        RECT 76.720 432.080 77.620 439.105 ;
        RECT 80.020 432.080 94.320 439.105 ;
        RECT 96.720 432.080 97.620 439.105 ;
        RECT 100.020 432.080 114.320 439.105 ;
        RECT 116.720 432.080 117.620 439.105 ;
        RECT 120.020 432.080 134.320 439.105 ;
        RECT 136.720 432.080 137.620 439.105 ;
        RECT 140.020 432.080 154.320 439.105 ;
        RECT 156.720 432.080 157.620 439.105 ;
        RECT 160.020 432.080 174.320 439.105 ;
        RECT 176.720 432.080 177.620 439.105 ;
        RECT 180.020 432.080 194.320 439.105 ;
        RECT 196.720 432.080 197.620 439.105 ;
        RECT 200.020 432.080 214.320 439.105 ;
        RECT 216.720 432.700 217.620 439.105 ;
        RECT 220.020 432.700 234.320 439.105 ;
        RECT 236.720 432.700 237.620 439.105 ;
        RECT 216.720 432.080 237.620 432.700 ;
        RECT 240.020 432.700 254.320 439.105 ;
        RECT 256.720 432.700 257.620 439.105 ;
        RECT 240.020 432.080 257.620 432.700 ;
        RECT 260.020 432.080 274.320 439.105 ;
        RECT 276.720 432.700 277.620 439.105 ;
        RECT 280.020 432.700 294.320 439.105 ;
        RECT 276.720 432.080 294.320 432.700 ;
        RECT 296.720 432.700 297.620 439.105 ;
        RECT 300.020 432.700 314.320 439.105 ;
        RECT 296.720 432.080 314.320 432.700 ;
        RECT 316.720 432.700 317.620 439.105 ;
        RECT 320.020 432.700 334.320 439.105 ;
        RECT 336.720 432.700 337.620 439.105 ;
        RECT 316.720 432.080 337.620 432.700 ;
        RECT 340.020 432.700 354.320 439.105 ;
        RECT 356.720 432.700 357.620 439.105 ;
        RECT 340.020 432.080 357.620 432.700 ;
        RECT 360.020 432.080 374.320 439.105 ;
        RECT 376.720 432.700 377.620 439.105 ;
        RECT 380.020 432.700 394.320 439.105 ;
        RECT 376.720 432.080 394.320 432.700 ;
        RECT 396.720 432.700 397.620 439.105 ;
        RECT 400.020 432.700 414.320 439.105 ;
        RECT 396.720 432.080 414.320 432.700 ;
        RECT 416.720 432.080 417.620 439.105 ;
        RECT 420.020 432.080 434.320 439.105 ;
        RECT 436.720 432.080 437.620 439.105 ;
        RECT 440.020 432.080 454.320 439.105 ;
        RECT 456.720 432.080 457.620 439.105 ;
        RECT 460.020 432.080 474.320 439.105 ;
        RECT 476.720 432.080 477.620 439.105 ;
        RECT 480.020 432.080 494.320 439.105 ;
        RECT 496.720 432.080 497.620 439.105 ;
        RECT 500.020 432.080 514.320 439.105 ;
        RECT 516.720 432.700 517.620 439.105 ;
        RECT 520.020 432.700 534.320 439.105 ;
        RECT 516.720 432.080 534.320 432.700 ;
        RECT 536.720 432.080 537.620 439.105 ;
        RECT 540.020 432.080 549.160 439.105 ;
        RECT 60.020 15.420 549.160 432.080 ;
        RECT 60.020 6.295 74.320 15.420 ;
        RECT 76.720 6.295 77.620 15.420 ;
        RECT 80.020 6.295 94.320 15.420 ;
        RECT 96.720 14.800 114.320 15.420 ;
        RECT 96.720 6.295 97.620 14.800 ;
        RECT 100.020 6.295 114.320 14.800 ;
        RECT 116.720 6.295 117.620 15.420 ;
        RECT 120.020 6.295 134.320 15.420 ;
        RECT 136.720 6.295 137.620 15.420 ;
        RECT 140.020 6.295 154.320 15.420 ;
        RECT 156.720 14.800 177.620 15.420 ;
        RECT 156.720 6.295 157.620 14.800 ;
        RECT 160.020 6.295 174.320 14.800 ;
        RECT 176.720 6.295 177.620 14.800 ;
        RECT 180.020 14.800 197.620 15.420 ;
        RECT 180.020 6.295 194.320 14.800 ;
        RECT 196.720 6.295 197.620 14.800 ;
        RECT 200.020 14.800 237.620 15.420 ;
        RECT 200.020 6.295 214.320 14.800 ;
        RECT 216.720 6.295 217.620 14.800 ;
        RECT 220.020 6.295 234.320 14.800 ;
        RECT 236.720 6.295 237.620 14.800 ;
        RECT 240.020 14.800 317.620 15.420 ;
        RECT 240.020 6.295 254.320 14.800 ;
        RECT 256.720 6.295 257.620 14.800 ;
        RECT 260.020 6.295 274.320 14.800 ;
        RECT 276.720 6.295 277.620 14.800 ;
        RECT 280.020 6.295 294.320 14.800 ;
        RECT 296.720 6.295 297.620 14.800 ;
        RECT 300.020 6.295 314.320 14.800 ;
        RECT 316.720 6.295 317.620 14.800 ;
        RECT 320.020 14.800 374.320 15.420 ;
        RECT 320.020 6.295 334.320 14.800 ;
        RECT 336.720 6.295 337.620 14.800 ;
        RECT 340.020 6.295 354.320 14.800 ;
        RECT 356.720 6.295 357.620 14.800 ;
        RECT 360.020 6.295 374.320 14.800 ;
        RECT 376.720 14.800 394.320 15.420 ;
        RECT 376.720 6.295 377.620 14.800 ;
        RECT 380.020 6.295 394.320 14.800 ;
        RECT 396.720 14.800 414.320 15.420 ;
        RECT 396.720 6.295 397.620 14.800 ;
        RECT 400.020 6.295 414.320 14.800 ;
        RECT 416.720 6.295 417.620 15.420 ;
        RECT 420.020 6.295 434.320 15.420 ;
        RECT 436.720 6.295 437.620 15.420 ;
        RECT 440.020 6.295 454.320 15.420 ;
        RECT 456.720 6.295 457.620 15.420 ;
        RECT 460.020 6.295 474.320 15.420 ;
        RECT 476.720 6.295 477.620 15.420 ;
        RECT 480.020 6.295 494.320 15.420 ;
        RECT 496.720 6.295 497.620 15.420 ;
        RECT 500.020 6.295 514.320 15.420 ;
        RECT 516.720 6.295 517.620 15.420 ;
        RECT 520.020 6.295 534.320 15.420 ;
        RECT 536.720 6.295 537.620 15.420 ;
        RECT 540.020 6.295 549.160 15.420 ;
  END
END BlockRAM_1KB
END LIBRARY

