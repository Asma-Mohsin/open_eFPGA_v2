* NGSPICE file created from eFPGA_Config.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt eFPGA_Config CLK ComActive ConfigWriteData[0] ConfigWriteData[10] ConfigWriteData[11]
+ ConfigWriteData[12] ConfigWriteData[13] ConfigWriteData[14] ConfigWriteData[15]
+ ConfigWriteData[16] ConfigWriteData[17] ConfigWriteData[18] ConfigWriteData[19]
+ ConfigWriteData[1] ConfigWriteData[20] ConfigWriteData[21] ConfigWriteData[22] ConfigWriteData[23]
+ ConfigWriteData[24] ConfigWriteData[25] ConfigWriteData[26] ConfigWriteData[27]
+ ConfigWriteData[28] ConfigWriteData[29] ConfigWriteData[2] ConfigWriteData[30] ConfigWriteData[31]
+ ConfigWriteData[3] ConfigWriteData[4] ConfigWriteData[5] ConfigWriteData[6] ConfigWriteData[7]
+ ConfigWriteData[8] ConfigWriteData[9] ConfigWriteStrobe FrameAddressRegister[0]
+ FrameAddressRegister[10] FrameAddressRegister[11] FrameAddressRegister[12] FrameAddressRegister[13]
+ FrameAddressRegister[14] FrameAddressRegister[15] FrameAddressRegister[16] FrameAddressRegister[17]
+ FrameAddressRegister[18] FrameAddressRegister[19] FrameAddressRegister[1] FrameAddressRegister[20]
+ FrameAddressRegister[21] FrameAddressRegister[22] FrameAddressRegister[23] FrameAddressRegister[24]
+ FrameAddressRegister[25] FrameAddressRegister[26] FrameAddressRegister[27] FrameAddressRegister[28]
+ FrameAddressRegister[29] FrameAddressRegister[2] FrameAddressRegister[30] FrameAddressRegister[31]
+ FrameAddressRegister[3] FrameAddressRegister[4] FrameAddressRegister[5] FrameAddressRegister[6]
+ FrameAddressRegister[7] FrameAddressRegister[8] FrameAddressRegister[9] LongFrameStrobe
+ ReceiveLED RowSelect[0] RowSelect[1] RowSelect[2] RowSelect[3] RowSelect[4] Rx SelfWriteData[0]
+ SelfWriteData[10] SelfWriteData[11] SelfWriteData[12] SelfWriteData[13] SelfWriteData[14]
+ SelfWriteData[15] SelfWriteData[16] SelfWriteData[17] SelfWriteData[18] SelfWriteData[19]
+ SelfWriteData[1] SelfWriteData[20] SelfWriteData[21] SelfWriteData[22] SelfWriteData[23]
+ SelfWriteData[24] SelfWriteData[25] SelfWriteData[26] SelfWriteData[27] SelfWriteData[28]
+ SelfWriteData[29] SelfWriteData[2] SelfWriteData[30] SelfWriteData[31] SelfWriteData[3]
+ SelfWriteData[4] SelfWriteData[5] SelfWriteData[6] SelfWriteData[7] SelfWriteData[8]
+ SelfWriteData[9] SelfWriteStrobe resetn s_clk s_data vccd1 vssd1
XINST_config_UART._1187_ net1 INST_config_UART._0056_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._345_ Inst_bitbang._172_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._074_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1335__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._414_ net1 Inst_bitbang._051_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._276_ Inst_bitbang.serial_data\[6\] Inst_bitbang.serial_data\[7\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1041_ INST_config_UART.CRCReg\[6\] INST_config_UART._0499_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0500_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1110_ INST_config_UART.ID_Reg\[0\] INST_config_UART._0223_ INST_config_UART._0553_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0756_ INST_config_UART.blink\[22\] INST_config_UART._0304_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0825_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[10\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0348_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0687_ INST_config_UART._0266_ INST_config_UART._0267_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0007_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1308_ net1 INST_config_UART._0143_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[5\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1239_ net1 INST_config_UART._0101_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HighReg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1251__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._328_ Inst_bitbang.s_clk_sample\[2\] Inst_bitbang.s_clk_sample\[3\]
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._163_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_bitbang._259_ Inst_bitbang._126_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._034_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINST_config_UART._0610_ INST_config_UART._0203_ INST_config_UART._0204_ INST_config_UART._0206_
+ INST_config_UART._0209_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0210_ sky130_fd_sc_hd__and4_1
XANTENNA_INST_config_UART._1257__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1024_ INST_config_UART._0483_ INST_config_UART._0485_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0486_ sky130_fd_sc_hd__xnor2_1
XINST_config_UART._0739_ INST_config_UART.blink\[14\] INST_config_UART._0294_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0297_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0808_ INST_config_UART._0243_ INST_config_UART.WriteData\[8\] INST_config_UART._0215_
+ INST_config_UART._0338_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0072_ sky130_fd_sc_hd__a31o_1
XANTENNA_INST_config_UART._1274__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__209__A ConfigFSM_inst.WriteData\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_200_ ConfigFSM_inst.WriteData\[19\] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1350__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_131_ _039_ INST_config_UART.WriteData\[17\] _023_ vssd1 vssd1 vccd1 vccd1 _040_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1297__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0655__B1 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._142_ ConfigFSM_inst._061_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._062_
+ sky130_fd_sc_hd__buf_4
XConfigFSM_inst._211_ ConfigFSM_inst._102_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._024_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1007_ INST_config_UART._0312_ INST_config_UART._0393_ INST_config_UART._0470_
+ INST_config_UART.CRCReg\[1\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0471_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1144__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._448__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_114_ _028_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[11\] sky130_fd_sc_hd__buf_2
XFILLER_0_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._266__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1272__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1201__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1312__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._125_ ConfigFSM_inst.WriteData\[17\] ConfigFSM_inst.WriteData\[16\]
+ ConfigFSM_inst.WriteData\[19\] ConfigFSM_inst.WriteData\[14\] vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._046_ sky130_fd_sc_hd__or4b_1
XFILLER_0_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1335__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._0623__C_N INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1341_ net1 INST_config_UART._0004_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[1\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1272_ net1 INST_config_UART._0130_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._366__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0987_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0322_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0456_ sky130_fd_sc_hd__and3_1
XInst_bitbang._430_ net1 net38 net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.s_data_sample\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._361_ Inst_bitbang._180_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._082_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1208__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._292_ Inst_bitbang._144_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._049_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1194__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1358__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[31] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[21] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[11] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_bitbang._389__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[3] sky130_fd_sc_hd__buf_2
XINST_config_UART._0772_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[2\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0317_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0910_ INST_config_UART._0407_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0408_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._0841_ INST_config_UART._0359_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0084_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1324_ net1 INST_config_UART._0159_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1186_ net1 INST_config_UART._0055_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[2\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1255_ net1 INST_config_UART._0116_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._237__A0 ConfigFSM_inst.WriteData\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._275_ Inst_bitbang._135_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._041_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1304__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._413_ net1 Inst_bitbang._050_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._344_ Inst_bitbang.serial_control\[6\] Inst_bitbang.serial_control\[7\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1180__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1040_ INST_config_UART.ReceivedWord\[6\] INST_config_UART.HighReg\[2\]
+ INST_config_UART.Command\[7\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._404__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0755_ INST_config_UART._0304_ INST_config_UART._0305_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0044_ sky130_fd_sc_hd__nand2_1
XANTENNA_ConfigFSM_inst._257__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0824_ INST_config_UART.ComTick vssd1 vssd1 vccd1 vccd1 INST_config_UART._0347_
+ sky130_fd_sc_hd__clkbuf_2
XINST_config_UART._1307_ net1 INST_config_UART._0142_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[4\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0686_ INST_config_UART.ComCount\[4\] INST_config_UART._0253_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1238_ net1 INST_config_UART._0016_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceiveState sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._385__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1169_ INST_config_UART.ComState\[5\] INST_config_UART.ComState\[8\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._327_ Inst_bitbang._162_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._066_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._258_ Inst_bitbang.serial_data\[31\] Inst_bitbang.data\[31\] Inst_bitbang._087_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._126_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._198__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XInst_bitbang._189_ Inst_bitbang._089_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._001_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1297__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._427__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1226__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1023_ INST_config_UART._0484_ INST_config_UART._0478_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0485_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0738_ INST_config_UART.blink\[14\] INST_config_UART._0294_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0296_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0807_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0314_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0338_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0669_ INST_config_UART.ComCount\[6\] INST_config_UART._0254_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0255_ sky130_fd_sc_hd__or2_1
XConfigFSM_inst._287_ net1 ConfigFSM_inst.FSM_Reset net112 vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst.old_reset sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_130_ net11 Inst_bitbang.data\[17\] _021_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._210_ ConfigFSM_inst.WriteData\[14\] ConfigFSM_inst.FrameAddressRegister\[14\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._141_ ConfigFSM_inst.WriteData\[20\] ConfigFSM_inst._041_ ConfigFSM_inst._043_
+ ConfigFSM_inst.state\[2\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._061_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1241__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1006_ INST_config_UART._0222_ INST_config_UART._0246_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0470_ sky130_fd_sc_hd__or2_1
XANTENNA_ConfigFSM_inst._272__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1144__B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_113_ _027_ INST_config_UART.WriteData\[11\] _023_ vssd1 vssd1 vccd1 vccd1 _028_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._417__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1264__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0876__A1 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1241__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._131__C_N ConfigFSM_inst.WriteData\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._124_ ConfigFSM_inst.WriteData\[18\] ConfigFSM_inst.WriteData\[22\]
+ ConfigFSM_inst.WriteData\[23\] ConfigFSM_inst.WriteData\[21\] vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._045_ sky130_fd_sc_hd__or4bb_1
XANTENNA_INST_config_UART._1329__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1287__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1340_ net1 INST_config_UART._0001_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1271_ net1 INST_config_UART._0129_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.ReceiveLED
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0986_ INST_config_UART._0242_ INST_config_UART.WriteData\[27\]
+ INST_config_UART._0234_ INST_config_UART._0455_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0133_
+ sky130_fd_sc_hd__a31o_1
XInst_bitbang._291_ Inst_bitbang.serial_data\[13\] Inst_bitbang.serial_data\[14\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._144_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._360_ Inst_bitbang.serial_control\[14\] Inst_bitbang.serial_control\[15\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[22] sky130_fd_sc_hd__buf_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[12] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[3] sky130_fd_sc_hd__buf_2
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[23] sky130_fd_sc_hd__buf_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[4] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[12] sky130_fd_sc_hd__clkbuf_4
XANTENNA_ConfigFSM_inst._256__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._191__A0 ConfigFSM_inst.WriteData\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1302__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._432__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0771_ INST_config_UART.WriteData\[1\] INST_config_UART._0240_ INST_config_UART._0316_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0840_ INST_config_UART.ID_Reg\[18\] INST_config_UART._0221_ INST_config_UART._0356_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1323_ net1 INST_config_UART._0158_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1185_ net1 INST_config_UART._0030_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[6\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1254_ net1 INST_config_UART._0115_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0969_ INST_config_UART.CRCReg\[15\] INST_config_UART._0442_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0443_ sky130_fd_sc_hd__nand2_1
XInst_bitbang._412_ net1 Inst_bitbang._049_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._274_ Inst_bitbang.serial_data\[5\] Inst_bitbang.serial_data\[6\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._135_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1325__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._343_ Inst_bitbang._171_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._073_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._279__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1344__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__138__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0754_ INST_config_UART.blink\[20\] INST_config_UART._0302_ INST_config_UART.blink\[21\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0305_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._0823_ INST_config_UART._0339_ INST_config_UART.WriteData\[15\]
+ INST_config_UART._0215_ INST_config_UART._0346_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0079_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0685_ INST_config_UART.ComCount\[4\] INST_config_UART._0253_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0266_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1306_ net1 INST_config_UART._0141_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[3\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1237_ net1 INST_config_UART._0100_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1348__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1099_ INST_config_UART._0539_ INST_config_UART._0544_ INST_config_UART.CRCReg\[18\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0546_ sky130_fd_sc_hd__a21o_1
XINST_config_UART._1168_ INST_config_UART._0350_ INST_config_UART.ComState\[1\] INST_config_UART._0306_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0186_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_bitbang._379__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._188_ Inst_bitbang.old_local_strobe Inst_bitbang.local_strobe vssd1
+ vssd1 vccd1 vccd1 Inst_bitbang._089_ sky130_fd_sc_hd__and2b_1
XInst_bitbang._326_ Inst_bitbang.serial_data\[30\] Inst_bitbang.serial_data\[31\]
+ Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._162_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._257_ Inst_bitbang._125_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._033_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1266__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1022_ INST_config_UART.CRCReg\[2\] INST_config_UART._0476_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0806_ INST_config_UART._0243_ INST_config_UART.WriteData\[23\]
+ INST_config_UART._0236_ INST_config_UART._0337_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0071_
+ sky130_fd_sc_hd__a31o_1
XINST_config_UART._0737_ INST_config_UART._0294_ INST_config_UART._0295_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0035_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._286_ net1 ConfigFSM_inst._000_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameStrobe
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0668_ INST_config_UART.ComCount\[5\] INST_config_UART.ComCount\[4\]
+ INST_config_UART._0253_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0254_ sky130_fd_sc_hd__or3_1
XINST_config_UART._0599_ INST_config_UART._0198_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0199_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._309_ Inst_bitbang._153_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._057_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1193__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_189_ ConfigFSM_inst.WriteData\[8\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._140_ ConfigFSM_inst.FrameShiftState\[1\] ConfigFSM_inst._059_ ConfigFSM_inst._043_
+ ConfigFSM_inst.FrameShiftState\[0\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._060_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA_ConfigFSM_inst._129__D_N ConfigFSM_inst.WriteData\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1005_ INST_config_UART._0461_ INST_config_UART._0462_ INST_config_UART._0466_
+ INST_config_UART._0469_ INST_config_UART.CRCReg\[0\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0138_
+ sky130_fd_sc_hd__a32o_1
XANTENNA_INST_config_UART._1188__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._269_ net1 ConfigFSM_inst._024_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._417__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_112_ net5 Inst_bitbang.data\[11\] _021_ vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._123_ ConfigFSM_inst._043_ ConfigFSM_inst._041_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._044_ sky130_fd_sc_hd__nor2_1
XANTENNA_INST_config_UART._1210__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1281__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1369__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1231__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1270_ net1 INST_config_UART._0000_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ByteWriteStrobe sky130_fd_sc_hd__dfrtp_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0985_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0320_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0455_ sky130_fd_sc_hd__and3_1
XANTENNA_Inst_bitbang._379__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._290_ Inst_bitbang._143_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._048_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1254__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[23] sky130_fd_sc_hd__clkbuf_4
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[13] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[4] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[24] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[5] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[13] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._0770_ INST_config_UART._0312_ INST_config_UART.HexData\[1\] INST_config_UART._0315_
+ INST_config_UART._0242_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0316_ sky130_fd_sc_hd__o211a_1
XANTENNA_Inst_bitbang._401__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1322_ net1 INST_config_UART._0157_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1253_ net1 INST_config_UART._0114_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1184_ net1 INST_config_UART._0018_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0968_ INST_config_UART.CRCReg\[12\] INST_config_UART.CRCReg\[13\]
+ INST_config_UART.CRCReg\[14\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0442_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1277__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._411_ net1 Inst_bitbang._048_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._342_ Inst_bitbang.serial_control\[5\] Inst_bitbang.serial_control\[6\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._171_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0899_ INST_config_UART._0397_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0104_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._273_ Inst_bitbang._134_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._040_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1313__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0822_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0328_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0346_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0753_ INST_config_UART.blink\[20\] INST_config_UART.blink\[21\]
+ INST_config_UART._0302_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0304_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0684_ INST_config_UART._0253_ INST_config_UART._0265_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1305_ net1 INST_config_UART._0140_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[2\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1236_ net1 INST_config_UART._0099_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._450__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._266__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1098_ INST_config_UART.CRCReg\[18\] INST_config_UART._0539_ INST_config_UART._0544_
+ INST_config_UART._0497_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0545_ sky130_fd_sc_hd__a31oi_1
XINST_config_UART._1167_ INST_config_UART._0584_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0185_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._246__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._394__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._325_ Inst_bitbang._161_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._065_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1156__A1 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._187_ Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._000_
+ sky130_fd_sc_hd__inv_2
XInst_bitbang._256_ Inst_bitbang.serial_data\[30\] Inst_bitbang.data\[30\] Inst_bitbang._087_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._125_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1021_ INST_config_UART._0481_ INST_config_UART._0482_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0483_ sky130_fd_sc_hd__or2b_1
XANTENNA_INST_config_UART._1235__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1315__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0736_ INST_config_UART.blink\[11\] INST_config_UART.blink\[12\]
+ INST_config_UART._0290_ INST_config_UART.blink\[13\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0295_
+ sky130_fd_sc_hd__o31ai_1
XINST_config_UART._0805_ INST_config_UART._0335_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0328_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0337_ sky130_fd_sc_hd__and3_1
XConfigFSM_inst._285_ net1 ConfigFSM_inst._040_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._269__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0598_ INST_config_UART._0197_ INST_config_UART.ComState\[6\] INST_config_UART._0198_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0667_ INST_config_UART.ComCount\[3\] INST_config_UART._0252_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0253_ sky130_fd_sc_hd__or2_1
XANTENNA_INST_config_UART._1138__A1 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1219_ net1 INST_config_UART._0082_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._308_ Inst_bitbang.serial_data\[21\] Inst_bitbang.serial_data\[22\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._153_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._239_ Inst_bitbang._116_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._024_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1338__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_188_ ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1004_ INST_config_UART._0468_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0469_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._369__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0719_ INST_config_UART.blink\[5\] INST_config_UART._0284_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0049_ sky130_fd_sc_hd__xnor2_1
XANTENNA_ConfigFSM_inst._281__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._268_ net1 ConfigFSM_inst._023_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._199_ ConfigFSM_inst._061_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._096_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_111_ _026_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[10\] sky130_fd_sc_hd__buf_2
XFILLER_0_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1179__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._426__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._122_ net72 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._043_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_INST_config_UART._1250__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_ConfigFSM_inst._200__A0 ConfigFSM_inst.WriteData\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1338__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1183__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._407__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0984_ INST_config_UART._0339_ INST_config_UART.WriteData\[26\]
+ INST_config_UART._0234_ INST_config_UART._0454_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0132_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[24] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[14] sky130_fd_sc_hd__clkbuf_4
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[5] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[25] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[14] sky130_fd_sc_hd__buf_2
XINST_config_UART._1321_ net1 INST_config_UART._0156_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[18\] sky130_fd_sc_hd__dfstp_1
XANTENNA_Inst_bitbang._441__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1252_ net1 INST_config_UART._0113_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1183_ net1 INST_config_UART._0029_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0898_ INST_config_UART._0232_ INST_config_UART.HighReg\[3\] INST_config_UART._0389_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0397_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0967_ INST_config_UART.TimeToSendCounter\[14\] INST_config_UART._0440_
+ INST_config_UART._0399_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0128_ sky130_fd_sc_hd__a21o_1
XInst_bitbang._410_ net1 Inst_bitbang._047_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._341_ Inst_bitbang._170_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._072_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._272_ Inst_bitbang.serial_data\[4\] Inst_bitbang.serial_data\[5\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1221__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0752_ INST_config_UART.blink\[20\] INST_config_UART._0302_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0043_ sky130_fd_sc_hd__xnor2_1
XINST_config_UART._0821_ INST_config_UART._0339_ INST_config_UART.WriteData\[14\]
+ INST_config_UART._0215_ INST_config_UART._0345_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0078_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0683_ INST_config_UART.ComCount\[3\] INST_config_UART._0252_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0265_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1304_ net1 INST_config_UART._0139_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[1\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1235_ net1 INST_config_UART._0098_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1244__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1166_ INST_config_UART.ComState\[8\] INST_config_UART.ComState\[2\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0584_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1097_ INST_config_UART.CRCReg\[16\] INST_config_UART.CRCReg\[17\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0544_ sky130_fd_sc_hd__and2_1
XANTENNA_Inst_bitbang._363__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._255_ Inst_bitbang._124_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._032_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._324_ Inst_bitbang.serial_data\[29\] Inst_bitbang.serial_data\[30\]
+ Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._161_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._186_ Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._088_
+ sky130_fd_sc_hd__buf_4
XINST_config_UART._1020_ INST_config_UART.CRCReg\[3\] INST_config_UART._0480_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0482_ sky130_fd_sc_hd__nand2_1
XANTENNA_INST_config_UART._1267__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1275__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1204__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0735_ INST_config_UART.blink\[11\] INST_config_UART.blink\[12\]
+ INST_config_UART.blink\[13\] INST_config_UART._0290_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0294_
+ sky130_fd_sc_hd__or4_2
XConfigFSM_inst._284_ net1 ConfigFSM_inst._039_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0804_ INST_config_UART._0243_ INST_config_UART.WriteData\[22\]
+ INST_config_UART._0236_ INST_config_UART._0336_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0070_
+ sky130_fd_sc_hd__a31o_1
XINST_config_UART._0597_ INST_config_UART.RxLocal INST_config_UART.ComState\[0\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0198_ sky130_fd_sc_hd__and2b_1
XINST_config_UART._0666_ INST_config_UART.ComCount\[1\] INST_config_UART.ComCount\[0\]
+ INST_config_UART.ComCount\[2\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0252_ sky130_fd_sc_hd__or3_1
XANTENNA_INST_config_UART._0624__A INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._1149_ INST_config_UART._0575_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0176_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1218_ net1 INST_config_UART._0081_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._238_ Inst_bitbang.serial_data\[21\] Inst_bitbang.data\[21\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._116_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._307_ Inst_bitbang._152_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._056_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._440__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_187_ ConfigFSM_inst.WriteData\[6\] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1003_ INST_config_UART._0192_ INST_config_UART._0467_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0468_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0718_ INST_config_UART._0284_ INST_config_UART._0285_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0048_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0649_ INST_config_UART._0214_ INST_config_UART._0238_ INST_config_UART._0240_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._267_ net1 ConfigFSM_inst._022_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._198_ ConfigFSM_inst._095_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._018_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1197__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_110_ _025_ INST_config_UART.WriteData\[10\] _023_ vssd1 vssd1 vccd1 vccd1 _026_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1305__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._259__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_239_ ConfigFSM_inst.FrameAddressRegister\[26\] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._121_ net72 ConfigFSM_inst.state\[2\] ConfigFSM_inst.WriteData\[20\]
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._042_ sky130_fd_sc_hd__and3_1
XANTENNA_Inst_bitbang._204__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1290__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1307__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1328__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0983_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0318_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0454_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._185__A0 ConfigFSM_inst.WriteData\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__112__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._388__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[25] sky130_fd_sc_hd__buf_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[15] sky130_fd_sc_hd__buf_2
XFILLER_0_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[15] sky130_fd_sc_hd__buf_2
XINST_config_UART._1320_ net1 INST_config_UART._0155_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[17\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1251_ net1 INST_config_UART._0112_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1182_ net1 INST_config_UART._0028_ net112 vssd1 vssd1 vccd1 vccd1
+ net39 sky130_fd_sc_hd__dfrtp_4
XANTENNA_INST_config_UART._1229__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._410__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0897_ INST_config_UART._0396_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0103_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0966_ INST_config_UART._0440_ INST_config_UART._0441_ INST_config_UART._0418_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0127_ sky130_fd_sc_hd__a21oi_1
XInst_bitbang._271_ Inst_bitbang._133_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._039_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._340_ Inst_bitbang.serial_control\[4\] Inst_bitbang.serial_control\[5\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1322__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0751_ INST_config_UART._0302_ INST_config_UART._0303_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0041_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0820_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0326_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0345_ sky130_fd_sc_hd__and3_1
XANTENNA_INST_config_UART._1196__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0682_ INST_config_UART._0259_ INST_config_UART._0264_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0005_ sky130_fd_sc_hd__a21o_1
XINST_config_UART._1303_ net1 INST_config_UART._0138_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1096_ INST_config_UART._0543_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0155_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1234_ net1 INST_config_UART._0097_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[12\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1165_ INST_config_UART._0583_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0184_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._275__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0949_ INST_config_UART.TimeToSendCounter\[7\] INST_config_UART._0401_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0431_ sky130_fd_sc_hd__nor2_1
XANTENNA_INST_config_UART._1314__SET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._185_ Inst_bitbang._083_ Inst_bitbang._084_ Inst_bitbang._085_ Inst_bitbang._086_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._087_ sky130_fd_sc_hd__nand4_4
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._254_ Inst_bitbang.serial_data\[29\] Inst_bitbang.data\[29\] Inst_bitbang._087_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._124_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._323_ Inst_bitbang._160_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._064_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0734_ INST_config_UART.blink\[12\] INST_config_UART._0292_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0034_ sky130_fd_sc_hd__xnor2_1
XINST_config_UART._0803_ INST_config_UART._0335_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0326_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0336_ sky130_fd_sc_hd__and3_1
XConfigFSM_inst._283_ net1 ConfigFSM_inst._038_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0665_ INST_config_UART._0250_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0251_
+ sky130_fd_sc_hd__buf_2
XANTENNA__181__A ConfigFSM_inst.WriteData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0596_ INST_config_UART.ComTick vssd1 vssd1 vccd1 vccd1 INST_config_UART._0197_
+ sky130_fd_sc_hd__inv_2
XANTENNA_INST_config_UART._1211__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1217_ net1 INST_config_UART._0020_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1079_ INST_config_UART.CRCReg\[12\] INST_config_UART._0529_ INST_config_UART._0497_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0532_ sky130_fd_sc_hd__a21oi_1
XANTENNA_INST_config_UART._1361__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1148_ INST_config_UART.Data_Reg\[1\] INST_config_UART._0222_ INST_config_UART._0573_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._392__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._237_ Inst_bitbang._115_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._023_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._306_ Inst_bitbang.serial_data\[20\] Inst_bitbang.serial_data\[21\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1234__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_186_ ConfigFSM_inst.WriteData\[5\] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1002_ INST_config_UART._0464_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0467_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__115__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0717_ INST_config_UART.blink\[4\] INST_config_UART._0282_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0285_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0648_ INST_config_UART.PresentState\[5\] INST_config_UART._0017_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0240_ sky130_fd_sc_hd__nor2_4
XConfigFSM_inst._266_ net1 ConfigFSM_inst._021_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._197_ ConfigFSM_inst.WriteData\[8\] ConfigFSM_inst.FrameAddressRegister\[8\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1257__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._124__C_N ConfigFSM_inst.WriteData\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._435__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_169_ _065_ INST_config_UART.WriteData\[29\] net39 vssd1 vssd1 vccd1 vccd1 _066_
+ sky130_fd_sc_hd__mux2_1
X_238_ ConfigFSM_inst.FrameAddressRegister\[25\] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._120_ ConfigFSM_inst.old_reset ConfigFSM_inst.FSM_Reset vssd1 vssd1
+ vccd1 vccd1 ConfigFSM_inst._041_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._249_ net1 ConfigFSM_inst._009_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameShiftState\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._430__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._191__A Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1347__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0982_ INST_config_UART._0339_ INST_config_UART.WriteData\[25\]
+ INST_config_UART._0234_ INST_config_UART._0453_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0131_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._453__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0632__B INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._249__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._186__A Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[26] sky130_fd_sc_hd__clkbuf_4
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[16] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[7] sky130_fd_sc_hd__buf_2
XFILLER_0_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1181__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1250_ net1 INST_config_UART._0111_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1181_ net1 INST_config_UART._0027_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1269__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._450__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0965_ INST_config_UART.TimeToSendCounter\[13\] INST_config_UART._0405_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0441_ sky130_fd_sc_hd__nand2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__184__A ConfigFSM_inst.WriteData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0896_ INST_config_UART._0395_ INST_config_UART.HighReg\[2\] INST_config_UART._0389_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0396_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1318__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._270_ Inst_bitbang.serial_data\[3\] Inst_bitbang.serial_data\[4\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._399_ net1 Inst_bitbang._036_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1362__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0750_ INST_config_UART.blink\[19\] INST_config_UART._0300_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0681_ INST_config_UART._0252_ INST_config_UART._0263_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0264_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1302_ net1 INST_config_UART._0045_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[22\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1233_ net1 INST_config_UART._0096_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._0629__C_N INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1095_ INST_config_UART._0542_ INST_config_UART._0540_ INST_config_UART.CRCReg\[17\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0543_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1164_ INST_config_UART.ComState\[9\] INST_config_UART.ComState\[3\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0583_ sky130_fd_sc_hd__mux2_1
XANTENNA__118__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0948_ INST_config_UART._0401_ INST_config_UART._0430_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1290__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0879_ INST_config_UART._0382_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0099_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._322_ Inst_bitbang.serial_data\[28\] Inst_bitbang.serial_data\[29\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._160_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._184_ Inst_bitbang.serial_control\[3\] Inst_bitbang.serial_control\[2\]
+ Inst_bitbang.serial_control\[1\] Inst_bitbang.serial_control\[0\] vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang._086_ sky130_fd_sc_hd__nor4b_2
XInst_bitbang._253_ Inst_bitbang._123_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._031_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._372__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0802_ INST_config_UART.ByteWriteStrobe vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0335_ sky130_fd_sc_hd__clkbuf_2
XConfigFSM_inst._282_ net1 ConfigFSM_inst._037_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0733_ INST_config_UART._0292_ INST_config_UART._0293_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0033_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0595_ INST_config_UART._0192_ INST_config_UART._0194_ INST_config_UART._0196_
+ INST_config_UART.PresentState\[6\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0026_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_INST_config_UART._1284__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0664_ INST_config_UART.ComState\[0\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0250_
+ sky130_fd_sc_hd__clkbuf_2
XINST_config_UART._1216_ net1 INST_config_UART._0019_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1213__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1078_ INST_config_UART._0466_ INST_config_UART._0526_ INST_config_UART._0530_
+ INST_config_UART._0531_ INST_config_UART.CRCReg\[11\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0149_
+ sky130_fd_sc_hd__a32o_1
XINST_config_UART._1147_ INST_config_UART._0574_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0175_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1186__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._221__A0 ConfigFSM_inst.WriteData\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._305_ Inst_bitbang._151_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._055_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._236_ Inst_bitbang.serial_data\[20\] Inst_bitbang.data\[20\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._115_ sky130_fd_sc_hd__mux2_1
X_185_ ConfigFSM_inst.WriteData\[4\] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._212__A0 ConfigFSM_inst.WriteData\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1001_ INST_config_UART._0465_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0466_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._282__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._265_ net1 ConfigFSM_inst._020_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__192__A ConfigFSM_inst.WriteData\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0716_ INST_config_UART.blink\[4\] INST_config_UART._0282_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0284_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0647_ INST_config_UART._0239_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0017_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._196_ ConfigFSM_inst._094_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._017_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._219_ Inst_bitbang.serial_data\[12\] Inst_bitbang.data\[12\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._106_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1201__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._404__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_237_ ConfigFSM_inst.FrameAddressRegister\[24\] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
X_168_ net24 Inst_bitbang.data\[29\] Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _065_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1351__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_099_ _017_ INST_config_UART.WriteData\[7\] _001_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__mux2_1
XANTENNA__187__A ConfigFSM_inst.WriteData\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._382__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._248_ net1 ConfigFSM_inst._008_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameShiftState\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XConfigFSM_inst._179_ ConfigFSM_inst.FrameShiftState\[3\] ConfigFSM_inst._074_ ConfigFSM_inst._079_
+ ConfigFSM_inst.FrameShiftState\[4\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._086_
+ sky130_fd_sc_hd__o31a_1
XANTENNA_INST_config_UART._1224__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0981_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0316_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0453_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1247__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._269__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._397__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[27] sky130_fd_sc_hd__buf_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1180_ net1 INST_config_UART._0026_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0964_ INST_config_UART.TimeToSendCounter\[13\] INST_config_UART._0405_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0440_ sky130_fd_sc_hd__or2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0895_ INST_config_UART._0219_ INST_config_UART._0229_ INST_config_UART._0231_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0395_ sky130_fd_sc_hd__o21ai_2
XANTENNA_Inst_bitbang._420__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._398_ net1 Inst_bitbang._035_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1331__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0842__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._443__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0680_ INST_config_UART.ComCount\[2\] INST_config_UART._0260_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._1301_ net1 INST_config_UART._0044_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[21\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1232_ net1 INST_config_UART._0095_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[10\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1163_ INST_config_UART._0582_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0183_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._1094_ INST_config_UART.CRCReg\[16\] INST_config_UART._0465_ INST_config_UART._0539_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0542_ sky130_fd_sc_hd__and3_1
XANTENNA__195__A ConfigFSM_inst.WriteData\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0878_ INST_config_UART.ID_Reg\[14\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART._0375_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0382_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._0833__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._0947_ INST_config_UART.TimeToSendCounter\[6\] INST_config_UART._0428_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0430_ sky130_fd_sc_hd__nand2_1
XANTENNA_ConfigFSM_inst._284__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._321_ Inst_bitbang._159_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._063_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._183_ Inst_bitbang.serial_control\[6\] Inst_bitbang.serial_control\[7\]
+ Inst_bitbang.serial_control\[5\] Inst_bitbang.serial_control\[4\] vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang._085_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._252_ Inst_bitbang.serial_data\[28\] Inst_bitbang.data\[28\] Inst_bitbang._087_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._123_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1308__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._429__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0732_ INST_config_UART.blink\[11\] INST_config_UART._0290_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._281_ net1 ConfigFSM_inst._036_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0801_ INST_config_UART._0243_ INST_config_UART.WriteData\[21\]
+ INST_config_UART._0236_ INST_config_UART._0334_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0069_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0663_ INST_config_UART._0249_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0015_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0594_ INST_config_UART.TimeToSend INST_config_UART._0195_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1146_ INST_config_UART.Data_Reg\[0\] INST_config_UART._0223_ INST_config_UART._0573_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0574_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1253__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1215_ net1 INST_config_UART._0080_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[5\] sky130_fd_sc_hd__dfrtp_4
XINST_config_UART._1077_ INST_config_UART._0467_ INST_config_UART._0529_ INST_config_UART._0192_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0531_ sky130_fd_sc_hd__a21oi_1
XANTENNA_ConfigFSM_inst._183__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._235_ Inst_bitbang._114_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._022_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._304_ Inst_bitbang.serial_data\[19\] Inst_bitbang.serial_data\[20\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._151_ sky130_fd_sc_hd__mux2_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_184_ ConfigFSM_inst.WriteData\[3\] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._122__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1000_ INST_config_UART._0192_ INST_config_UART._0464_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0465_ sky130_fd_sc_hd__nor2_1
XANTENNA_INST_config_UART._1280__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._324__S Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0715_ INST_config_UART._0282_ INST_config_UART._0283_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0047_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._195_ ConfigFSM_inst.WriteData\[7\] ConfigFSM_inst.FrameAddressRegister\[7\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._094_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._264_ net1 ConfigFSM_inst._019_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0646_ INST_config_UART.ByteWriteStrobe INST_config_UART.GetWordState\[3\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0239_ sky130_fd_sc_hd__and2_1
XINST_config_UART._1129_ INST_config_UART._0564_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0167_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._218_ Inst_bitbang._105_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._014_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_098_ net32 Inst_bitbang.data\[7\] _000_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_236_ ConfigFSM_inst.FrameAddressRegister\[23\] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._197__A0 ConfigFSM_inst.WriteData\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_167_ _064_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[28\] sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_Inst_bitbang._444__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0629_ INST_config_UART.ReceivedWord\[4\] INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART.ReceivedWord\[6\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0225_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._247_ net1 ConfigFSM_inst._007_ net36 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameShiftState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._178_ ConfigFSM_inst._074_ ConfigFSM_inst._084_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0662__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._272__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0980_ INST_config_UART._0339_ INST_config_UART.WriteData\[24\]
+ INST_config_UART._0234_ INST_config_UART._0452_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0130_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_INST_config_UART._1199__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_219_ ConfigFSM_inst.FrameAddressRegister\[6\] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XANTENNA__198__A ConfigFSM_inst.WriteData\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._191__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._366__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[18] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1341__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1190__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._372__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._130__A ConfigFSM_inst.WriteData\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._0894_ INST_config_UART._0394_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0102_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1207__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0963_ INST_config_UART._0405_ INST_config_UART._0439_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0126_ sky130_fd_sc_hd__a21oi_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1278__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1214__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1364__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._397_ net1 Inst_bitbang._034_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._395__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1300__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1237__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._125__A ConfigFSM_inst.WriteData\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1300_ net1 INST_config_UART._0043_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[20\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1231_ net1 INST_config_UART._0094_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[9\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1093_ INST_config_UART.CRCReg\[16\] INST_config_UART._0540_ INST_config_UART._0541_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0154_ sky130_fd_sc_hd__a21o_1
XINST_config_UART._1162_ INST_config_UART.ComState\[10\] INST_config_UART.ComState\[5\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0582_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0877_ INST_config_UART._0381_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0098_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0946_ INST_config_UART._0428_ INST_config_UART._0429_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._251_ Inst_bitbang._122_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._030_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._320_ Inst_bitbang.serial_data\[27\] Inst_bitbang.serial_data\[28\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._159_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._182_ Inst_bitbang.serial_control\[8\] Inst_bitbang.serial_control\[10\]
+ Inst_bitbang.serial_control\[11\] Inst_bitbang.serial_control\[9\] vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang._084_ sky130_fd_sc_hd__and4bb_1
XANTENNA_ConfigFSM_inst._253__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_bitbang._381__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._449_ net1 Inst_bitbang._078_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._410__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0731_ INST_config_UART.blink\[11\] INST_config_UART._0290_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0292_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0662_ net39 INST_config_UART._0242_ INST_config_UART._0193_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0249_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0800_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0324_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0334_ sky130_fd_sc_hd__and3_1
XConfigFSM_inst._280_ net1 ConfigFSM_inst._035_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0593_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0195_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1076_ INST_config_UART._0529_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0530_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._1145_ INST_config_UART._0572_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0573_
+ sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._1214_ net1 INST_config_UART._0024_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.GetWordState\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1293__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1222__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0929_ INST_config_UART._0399_ INST_config_UART._0406_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0418_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._433__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._234_ Inst_bitbang.serial_data\[19\] Inst_bitbang.data\[19\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._114_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._303_ Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._150_
+ sky130_fd_sc_hd__clkbuf_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ ConfigFSM_inst.WriteData\[2\] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0645_ INST_config_UART.GetWordState\[0\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0238_ sky130_fd_sc_hd__inv_2
XINST_config_UART._0714_ INST_config_UART.blink\[3\] INST_config_UART._0280_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0283_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._194_ ConfigFSM_inst._093_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._016_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._263_ net1 ConfigFSM_inst._018_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1059_ INST_config_UART._0502_ INST_config_UART._0505_ INST_config_UART._0513_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0516_ sky130_fd_sc_hd__or3_1
XINST_config_UART._1128_ INST_config_UART.Command\[0\] INST_config_UART._0223_ INST_config_UART._0563_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._217_ Inst_bitbang.serial_data\[11\] Inst_bitbang.data\[11\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._105_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1140__A1 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_235_ ConfigFSM_inst.FrameAddressRegister\[22\] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
X_097_ _016_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[6\] sky130_fd_sc_hd__buf_2
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_166_ _063_ INST_config_UART.WriteData\[28\] _045_ vssd1 vssd1 vccd1 vccd1 _064_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._413__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0628_ INST_config_UART._0222_ INST_config_UART._0223_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0224_ sky130_fd_sc_hd__nor2_1
XConfigFSM_inst._177_ ConfigFSM_inst.FrameShiftState\[3\] ConfigFSM_inst.FrameShiftState\[4\]
+ ConfigFSM_inst._079_ ConfigFSM_inst.state\[1\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._084_
+ sky130_fd_sc_hd__o31a_1
XConfigFSM_inst._246_ net1 ConfigFSM_inst._006_ net36 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameShiftState\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_ConfigFSM_inst._189__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1122__A1 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1270__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1325__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_218_ ConfigFSM_inst.FrameAddressRegister\[5\] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
X_149_ _052_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[22\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_INST_config_UART._1293__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._278__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 ComActive sky130_fd_sc_hd__clkbuf_4
XANTENNA_INST_config_UART._1040__A0 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._229_ ConfigFSM_inst.WriteData\[24\] ConfigFSM_inst.FrameAddressRegister\[24\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._130__B ConfigFSM_inst.WriteData\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0893_ INST_config_UART._0393_ INST_config_UART.HighReg\[1\] INST_config_UART._0389_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0394_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0962_ INST_config_UART.TimeToSendCounter\[12\] INST_config_UART._0404_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0439_ sky130_fd_sc_hd__nand2_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1247__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._262__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1189__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1013__A0 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_bitbang._396_ net1 Inst_bitbang._033_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._125__B ConfigFSM_inst.WriteData\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._1230_ net1 INST_config_UART._0093_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._141__A ConfigFSM_inst.WriteData\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1340__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1161_ INST_config_UART._0581_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0182_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1092_ INST_config_UART.CRCReg\[16\] INST_config_UART._0465_ INST_config_UART._0539_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0541_ sky130_fd_sc_hd__and3b_1
XINST_config_UART._0945_ INST_config_UART.TimeToSendCounter\[4\] INST_config_UART._0400_
+ INST_config_UART.TimeToSendCounter\[5\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0429_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_INST_config_UART._1331__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0876_ INST_config_UART.ID_Reg\[13\] INST_config_UART.ReceivedWord\[5\]
+ INST_config_UART._0375_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0381_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._285__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._233__A0 ConfigFSM_inst.WriteData\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1359_ net1 INST_config_UART._0180_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_bitbang._181_ Inst_bitbang.serial_control\[13\] Inst_bitbang.serial_control\[12\]
+ Inst_bitbang.serial_control\[15\] Inst_bitbang.serial_control\[14\] vssd1 vssd1
+ vccd1 vccd1 Inst_bitbang._083_ sky130_fd_sc_hd__and4_1
XInst_bitbang._250_ Inst_bitbang.serial_data\[27\] Inst_bitbang.data\[27\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._122_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._197__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._362__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._379_ net1 Inst_bitbang._016_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._448_ net1 Inst_bitbang._077_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1204__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._438__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0730_ INST_config_UART._0290_ INST_config_UART._0291_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0032_ sky130_fd_sc_hd__nand2_1
XANTENNA_INST_config_UART._1354__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0592_ INST_config_UART.TimeToSend INST_config_UART._0193_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0194_ sky130_fd_sc_hd__nor2_1
XINST_config_UART._0661_ INST_config_UART._0248_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0000_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1213_ net1 INST_config_UART._0023_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.GetWordState\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1075_ INST_config_UART._0517_ INST_config_UART._0519_ INST_config_UART._0528_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0529_ sky130_fd_sc_hd__a21oi_4
XINST_config_UART._1144_ net39 net112 INST_config_UART._0193_ vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0572_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0928_ INST_config_UART._0417_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0113_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._206__A0 ConfigFSM_inst.WriteData\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._385__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1262__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._302_ Inst_bitbang._149_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._054_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0859_ INST_config_UART.RxLocal INST_config_UART._0369_ INST_config_UART._0370_
+ INST_config_UART.ReceivedWord\[4\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0091_
+ sky130_fd_sc_hd__o22a_1
XInst_bitbang._233_ Inst_bitbang._113_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._021_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1227__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ ConfigFSM_inst.WriteData\[1\] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._262_ net1 ConfigFSM_inst._017_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0644_ INST_config_UART._0236_ INST_config_UART._0237_ INST_config_UART.PresentState\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0022_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._0713_ INST_config_UART.blink\[0\] INST_config_UART.blink\[1\] INST_config_UART.blink\[2\]
+ INST_config_UART.blink\[3\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0282_ sky130_fd_sc_hd__or4_2
XConfigFSM_inst._193_ ConfigFSM_inst.WriteData\[6\] ConfigFSM_inst.FrameAddressRegister\[6\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._093_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1058_ INST_config_UART._0514_ INST_config_UART._0515_ INST_config_UART.CRCReg\[7\]
+ INST_config_UART._0469_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0145_ sky130_fd_sc_hd__a2bb2o_1
XINST_config_UART._1127_ INST_config_UART._0562_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0563_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._400__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._216_ Inst_bitbang._104_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._013_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1184__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_234_ ConfigFSM_inst.FrameAddressRegister\[21\] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
X_165_ net23 Inst_bitbang.data\[28\] _043_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__mux2_1
X_096_ _015_ INST_config_UART.WriteData\[6\] _001_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._453__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._245_ net1 ConfigFSM_inst._005_ net36 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameShiftState\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_Inst_bitbang._423__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0627_ INST_config_UART.ReceivedWord\[0\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0223_ sky130_fd_sc_hd__clkbuf_4
XConfigFSM_inst._176_ ConfigFSM_inst.FrameShiftState\[3\] ConfigFSM_inst._082_ ConfigFSM_inst._083_
+ ConfigFSM_inst._076_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._008_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1365__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._0872__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._446__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_217_ ConfigFSM_inst.FrameAddressRegister\[4\] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
X_148_ _051_ INST_config_UART.WriteData\[22\] _045_ vssd1 vssd1 vccd1 vccd1 _052_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_079_ _004_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[0\] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._0863__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._228_ ConfigFSM_inst._111_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._032_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._247__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._256__S Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._159_ ConfigFSM_inst._071_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.RowSelect\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._375__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0961_ INST_config_UART._0404_ INST_config_UART._0438_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0125_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0892_ INST_config_UART._0227_ INST_config_UART._0392_ INST_config_UART._0218_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0393_ sky130_fd_sc_hd__a21oi_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1287__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1260__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._395_ net1 Inst_bitbang._032_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._125__C ConfigFSM_inst.WriteData\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0763__A0 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._1091_ INST_config_UART.CRCReg\[16\] INST_config_UART._0467_ INST_config_UART._0539_
+ INST_config_UART._0192_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0540_ sky130_fd_sc_hd__a31oi_2
XINST_config_UART._1160_ INST_config_UART.Data_Reg\[7\] INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART._0573_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0581_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1283__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0944_ INST_config_UART.TimeToSendCounter\[5\] INST_config_UART._0426_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0428_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0875_ INST_config_UART._0380_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0097_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1358_ net1 INST_config_UART._0179_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XINST_config_UART._1289_ net1 INST_config_UART._0053_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._262__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._447_ net1 Inst_bitbang._076_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._378_ net1 Inst_bitbang._015_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._390__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0660_ INST_config_UART.LocalWriteStrobe INST_config_UART.HexWriteStrobe
+ INST_config_UART._0247_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0248_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0591_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0193_ sky130_fd_sc_hd__and2_1
XANTENNA_Inst_bitbang._407__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1143_ INST_config_UART._0571_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0174_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1212_ net1 INST_config_UART._0022_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.GetWordState\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1074_ INST_config_UART.CRCReg\[10\] INST_config_UART.CRCReg\[11\]
+ INST_config_UART._0445_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0528_ sky130_fd_sc_hd__nand3_2
XANTENNA_ConfigFSM_inst._252__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0927_ INST_config_UART.HexData\[7\] INST_config_UART.HighReg\[3\]
+ INST_config_UART._0014_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0417_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1179__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0858_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0370_ sky130_fd_sc_hd__and3b_1
XFILLER_0_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0789_ INST_config_UART.WriteData\[7\] INST_config_UART._0240_ INST_config_UART._0328_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0063_ sky130_fd_sc_hd__a22o_1
XANTENNA_INST_config_UART._1231__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._301_ Inst_bitbang.serial_data\[18\] Inst_bitbang.serial_data\[19\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._149_ sky130_fd_sc_hd__mux2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._232_ Inst_bitbang.serial_data\[18\] Inst_bitbang.data\[18\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._113_ sky130_fd_sc_hd__mux2_1
X_181_ ConfigFSM_inst.WriteData\[0\] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1319__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._275__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1321__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0712_ INST_config_UART._0280_ INST_config_UART._0281_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0046_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._261_ net1 ConfigFSM_inst._016_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0643_ INST_config_UART.ByteWriteStrobe INST_config_UART.GetWordState\[1\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0237_ sky130_fd_sc_hd__or2b_1
XConfigFSM_inst._192_ ConfigFSM_inst._092_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._015_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1126_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] INST_config_UART.PresentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0562_ sky130_fd_sc_hd__and3_1
XINST_config_UART._1057_ INST_config_UART._0501_ INST_config_UART._0509_ INST_config_UART._0513_
+ INST_config_UART._0497_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0515_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._215_ Inst_bitbang.serial_data\[10\] Inst_bitbang.data\[10\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._104_ sky130_fd_sc_hd__mux2_1
XANTENNA__172__S net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__201__A ConfigFSM_inst.WriteData\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1344__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_095_ net31 Inst_bitbang.data\[6\] _000_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_233_ net113 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[20] sky130_fd_sc_hd__buf_2
X_164_ _062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[27\] sky130_fd_sc_hd__buf_1
XANTENNA_Inst_bitbang._375__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._244_ ConfigFSM_inst._119_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._040_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._175_ ConfigFSM_inst._070_ ConfigFSM_inst._079_ ConfigFSM_inst._057_
+ ConfigFSM_inst.state\[1\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._083_ sky130_fd_sc_hd__o211a_1
XANTENNA_INST_config_UART._1217__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0626_ INST_config_UART.ReceivedWord\[1\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0222_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._422__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1367__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1109_ INST_config_UART._0552_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0553_
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_bitbang._398__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1334__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_078_ _003_ INST_config_UART.WriteData\[0\] _001_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__mux2_1
XANTENNA__106__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_147_ net17 Inst_bitbang.data\[22\] _043_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__mux2_1
X_216_ ConfigFSM_inst.FrameAddressRegister\[3\] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._158_ ConfigFSM_inst.FrameShiftState\[4\] ConfigFSM_inst._043_ vssd1
+ vssd1 vccd1 vccd1 ConfigFSM_inst._071_ sky130_fd_sc_hd__or2b_1
XConfigFSM_inst._227_ ConfigFSM_inst.WriteData\[23\] ConfigFSM_inst.FrameAddressRegister\[23\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0609_ INST_config_UART._0207_ INST_config_UART._0208_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0209_ sky130_fd_sc_hd__nor2_1
XANTENNA_ConfigFSM_inst._287__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._125__D_N ConfigFSM_inst.WriteData\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._413__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0891_ INST_config_UART._0391_ INST_config_UART._0219_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0392_ sky130_fd_sc_hd__or2_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0960_ INST_config_UART.TimeToSendCounter\[10\] INST_config_UART._0403_
+ INST_config_UART.TimeToSendCounter\[11\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0438_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1256__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._394_ net1 Inst_bitbang._031_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._436__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._0763__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1090_ INST_config_UART._0517_ INST_config_UART._0519_ INST_config_UART._0528_
+ INST_config_UART._0443_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0539_ sky130_fd_sc_hd__a211oi_4
XINST_config_UART._0874_ INST_config_UART.ID_Reg\[12\] INST_config_UART.ReceivedWord\[4\]
+ INST_config_UART._0375_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0380_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0943_ INST_config_UART._0426_ INST_config_UART._0427_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0118_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1357_ net1 INST_config_UART._0178_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XINST_config_UART._1288_ net1 INST_config_UART._0052_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__175__S net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__204__A ConfigFSM_inst.WriteData\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._377_ net1 Inst_bitbang._014_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._446_ net1 Inst_bitbang._075_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1178__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1250__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0590_ INST_config_UART.PresentState\[1\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0192_ sky130_fd_sc_hd__buf_2
XINST_config_UART._1073_ INST_config_UART._0497_ INST_config_UART._0525_ INST_config_UART._0526_
+ INST_config_UART._0527_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0148_ sky130_fd_sc_hd__o31ai_1
XINST_config_UART._1142_ INST_config_UART._0247_ INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART._0563_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0571_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._447__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1211_ net1 INST_config_UART._0021_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.GetWordState\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0926_ INST_config_UART._0416_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0112_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0857_ INST_config_UART._0368_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0369_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0788_ INST_config_UART._0312_ INST_config_UART.HexData\[7\] INST_config_UART._0327_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0328_ sky130_fd_sc_hd__o211a_1
XInst_bitbang._300_ Inst_bitbang._148_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._053_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._231_ Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._112_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1152__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1200__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_180_ Inst_bitbang.strobe INST_config_UART.ReceiveLED vssd1 vssd1 vccd1 vccd1 net105
+ sky130_fd_sc_hd__xor2_1
XANTENNA_INST_config_UART._1273__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XInst_bitbang._429_ net1 Inst_bitbang._066_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0711_ INST_config_UART.blink\[0\] INST_config_UART.blink\[1\] INST_config_UART.blink\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0281_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._0642_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0236_ sky130_fd_sc_hd__nand2_4
XConfigFSM_inst._260_ net1 ConfigFSM_inst._015_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._191_ ConfigFSM_inst.WriteData\[5\] ConfigFSM_inst.FrameAddressRegister\[5\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._092_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1056_ INST_config_UART._0501_ INST_config_UART._0509_ INST_config_UART._0513_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0514_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._1125_ INST_config_UART._0561_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0166_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1134__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1296__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0909_ INST_config_UART._0399_ INST_config_UART._0406_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0407_ sky130_fd_sc_hd__or2_2
XANTENNA_Inst_bitbang._369__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._214_ Inst_bitbang._103_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._012_
+ sky130_fd_sc_hd__clkbuf_1
X_232_ ConfigFSM_inst.FrameAddressRegister\[19\] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1315__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_094_ _014_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[5\] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1193__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_163_ _061_ INST_config_UART.WriteData\[27\] _045_ vssd1 vssd1 vccd1 vccd1 _062_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1116__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0625_ INST_config_UART.ReceivedWord\[2\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0221_ sky130_fd_sc_hd__clkbuf_4
XConfigFSM_inst._243_ ConfigFSM_inst.WriteData\[31\] ConfigFSM_inst.FrameAddressRegister\[31\]
+ ConfigFSM_inst._061_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._119_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._174_ ConfigFSM_inst._076_ ConfigFSM_inst._079_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1039_ INST_config_UART._0496_ INST_config_UART._0498_ INST_config_UART.CRCReg\[5\]
+ INST_config_UART._0469_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0143_ sky130_fd_sc_hd__a2bb2o_1
XINST_config_UART._1108_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] INST_config_UART.PresentState\[6\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0552_ sky130_fd_sc_hd__and3_1
XANTENNA_INST_config_UART._1107__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1107__B2 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._265__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1311__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__212__A ConfigFSM_inst.WriteData\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1034__A0 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1303__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_215_ ConfigFSM_inst.FrameAddressRegister\[2\] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
X_077_ net3 Inst_bitbang.data\[0\] _000_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__mux2_1
X_146_ _050_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[21\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0608_ INST_config_UART.ID_Reg\[14\] INST_config_UART.ID_Reg\[17\]
+ INST_config_UART.ID_Reg\[16\] INST_config_UART.ID_Reg\[15\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0208_ sky130_fd_sc_hd__or4b_1
XANTENNA_INST_config_UART._1334__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._226_ ConfigFSM_inst._110_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._031_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._157_ ConfigFSM_inst._043_ ConfigFSM_inst._070_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst.RowSelect\[3\] sky130_fd_sc_hd__nand2_1
XFILLER_0_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._256__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__178__S net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__207__A ConfigFSM_inst.WriteData\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._365__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._384__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1207__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0890_ INST_config_UART.ReceivedWord\[1\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0391_ sky130_fd_sc_hd__inv_2
XANTENNA_INST_config_UART._1357__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_129_ _038_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[16\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1296__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._388__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1225__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._209_ ConfigFSM_inst._101_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._023_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._393_ net1 Inst_bitbang._030_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._227__A0 ConfigFSM_inst.WriteData\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0873_ INST_config_UART._0379_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0096_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._218__A0 ConfigFSM_inst.WriteData\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0942_ INST_config_UART.TimeToSendCounter\[4\] INST_config_UART._0400_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0427_ sky130_fd_sc_hd__nand2_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1356_ net1 INST_config_UART._0177_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XINST_config_UART._1287_ net1 INST_config_UART._0051_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._403__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0976__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._250__SET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._376_ net1 Inst_bitbang._013_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._445_ net1 Inst_bitbang._074_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._271__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINST_config_UART._1210_ net1 INST_config_UART._0079_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[15\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1072_ INST_config_UART.CRCReg\[10\] INST_config_UART._0468_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0527_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1141_ INST_config_UART._0570_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0173_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0925_ INST_config_UART.HexData\[6\] INST_config_UART.HighReg\[2\]
+ INST_config_UART._0014_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0416_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._416__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0787_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[7\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0327_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0856_ INST_config_UART.ComState\[0\] INST_config_UART._0347_ INST_config_UART.ComState\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_bitbang._426__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1339_ net1 INST_config_UART._0174_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[7\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._230_ Inst_bitbang._111_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._020_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1240__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._359_ Inst_bitbang._179_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._081_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1328__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._428_ net1 Inst_bitbang._065_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._449__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0710_ INST_config_UART.blink\[0\] INST_config_UART.blink\[1\] INST_config_UART.blink\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0280_ sky130_fd_sc_hd__or3_1
XINST_config_UART._0641_ INST_config_UART._0234_ INST_config_UART._0235_ INST_config_UART.PresentState\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0023_ sky130_fd_sc_hd__a21oi_1
XConfigFSM_inst._190_ ConfigFSM_inst._091_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._014_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1055_ INST_config_UART._0511_ INST_config_UART._0512_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0513_ sky130_fd_sc_hd__or2b_1
XINST_config_UART._1124_ INST_config_UART.ID_Reg\[7\] INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART._0553_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0561_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0908_ INST_config_UART.TimeToSendCounter\[13\] INST_config_UART.TimeToSendCounter\[14\]
+ INST_config_UART._0405_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0406_ sky130_fd_sc_hd__or3_1
XINST_config_UART._0839_ INST_config_UART._0358_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0083_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._213_ Inst_bitbang.serial_data\[9\] Inst_bitbang.data\[9\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1240__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0636__A1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_231_ ConfigFSM_inst.FrameAddressRegister\[18\] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
X_162_ net22 Inst_bitbang.data\[27\] _043_ vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__mux2_1
X_093_ _013_ INST_config_UART.WriteData\[5\] _001_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0624_ INST_config_UART._0218_ INST_config_UART._0219_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0220_ sky130_fd_sc_hd__nor2_1
XConfigFSM_inst._242_ ConfigFSM_inst._118_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._039_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._173_ ConfigFSM_inst.FrameShiftState\[2\] ConfigFSM_inst._076_ ConfigFSM_inst._075_
+ ConfigFSM_inst._081_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._007_ sky130_fd_sc_hd__a22o_1
XANTENNA_INST_config_UART._1263__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1038_ INST_config_UART._0490_ INST_config_UART._0493_ INST_config_UART._0495_
+ INST_config_UART._0497_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0498_ sky130_fd_sc_hd__a31o_1
XANTENNA_Inst_bitbang._431__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1107_ INST_config_UART.RxLocal INST_config_UART._0550_ INST_config_UART._0551_
+ INST_config_UART.ReceivedWord\[6\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0158_
+ sky130_fd_sc_hd__o22a_1
Xinput1 CLK vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_16
XANTENNA_INST_config_UART._1321__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_ConfigFSM_inst._130__C_N ConfigFSM_inst.WriteData\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._196__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_214_ ConfigFSM_inst.FrameAddressRegister\[1\] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
X_145_ _049_ INST_config_UART.WriteData\[21\] _045_ vssd1 vssd1 vccd1 vccd1 _050_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1286__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1343__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_076_ _002_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FSM_Reset sky130_fd_sc_hd__buf_1
XANTENNA_INST_config_UART._0848__A1 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._225_ ConfigFSM_inst.WriteData\[22\] ConfigFSM_inst.FrameAddressRegister\[22\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0607_ INST_config_UART.ID_Reg\[19\] INST_config_UART.ID_Reg\[18\]
+ INST_config_UART.ID_Reg\[21\] INST_config_UART.ID_Reg\[20\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0207_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._156_ ConfigFSM_inst.FrameShiftState\[3\] vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst._070_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_128_ _037_ INST_config_UART.WriteData\[16\] _023_ vssd1 vssd1 vccd1 vccd1 _038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._255__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._181__A0 ConfigFSM_inst.WriteData\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1301__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1265__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._208_ ConfigFSM_inst.WriteData\[13\] ConfigFSM_inst.FrameAddressRegister\[13\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._101_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._392_ net1 Inst_bitbang._029_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._139_ ConfigFSM_inst.FrameShiftState\[3\] ConfigFSM_inst.FrameShiftState\[2\]
+ ConfigFSM_inst.FrameShiftState\[4\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._059_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1324__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._278__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0941_ INST_config_UART.TimeToSendCounter\[4\] INST_config_UART._0400_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0426_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0872_ INST_config_UART.ID_Reg\[11\] INST_config_UART._0218_ INST_config_UART._0375_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1355_ net1 INST_config_UART._0176_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1286_ net1 INST_config_UART._0050_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[6\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._444_ net1 Inst_bitbang._073_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._375_ net1 Inst_bitbang._012_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1347__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1187__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._378__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1071_ INST_config_UART.CRCReg\[10\] INST_config_UART._0445_ INST_config_UART._0520_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0526_ sky130_fd_sc_hd__and3_1
XINST_config_UART._1140_ INST_config_UART.Command\[6\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART._0563_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0924_ INST_config_UART._0415_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0111_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0786_ INST_config_UART.WriteData\[6\] INST_config_UART._0240_ INST_config_UART._0326_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0062_ sky130_fd_sc_hd__a22o_1
XINST_config_UART._0855_ INST_config_UART.RxLocal INST_config_UART._0366_ INST_config_UART._0367_
+ INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0090_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1338_ net1 INST_config_UART._0173_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[6\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1269_ net1 INST_config_UART._0015_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.LocalWriteStrobe sky130_fd_sc_hd__dfrtp_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1280__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._427_ net1 Inst_bitbang._064_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._289_ Inst_bitbang.serial_data\[12\] Inst_bitbang.serial_data\[13\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._143_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._358_ Inst_bitbang.serial_control\[13\] Inst_bitbang.serial_control\[14\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._179_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1368__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0640_ INST_config_UART._0216_ INST_config_UART.GetWordState\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0235_ sky130_fd_sc_hd__or2b_1
XINST_config_UART._1123_ INST_config_UART._0560_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0165_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1054_ INST_config_UART.CRCReg\[7\] INST_config_UART._0510_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0512_ sky130_fd_sc_hd__nand2_1
XANTENNA_INST_config_UART._1192__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0838_ INST_config_UART.ID_Reg\[17\] INST_config_UART._0222_ INST_config_UART._0356_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0358_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0907_ INST_config_UART.TimeToSendCounter\[12\] INST_config_UART._0404_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0405_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0769_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[1\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0315_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._212_ Inst_bitbang._102_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._011_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._378__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0636__A2 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_230_ ConfigFSM_inst.FrameAddressRegister\[17\] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
X_161_ _060_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[26\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_092_ net30 Inst_bitbang.data\[5\] _000_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._416__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._241_ ConfigFSM_inst.WriteData\[30\] ConfigFSM_inst.FrameAddressRegister\[30\]
+ ConfigFSM_inst._061_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._118_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0623_ INST_config_UART.ReceivedWord\[7\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART.ReceivedWord\[5\] INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0219_ sky130_fd_sc_hd__or4bb_2
XConfigFSM_inst._172_ ConfigFSM_inst._079_ ConfigFSM_inst._080_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._081_ sky130_fd_sc_hd__nand2_1
XANTENNA__136__A Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1219__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1106_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[1\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0551_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._400__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1037_ INST_config_UART._0192_ INST_config_UART._0464_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0497_ sky130_fd_sc_hd__or2_2
Xinput2 Rx vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._439__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_075_ _000_ _001_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_213_ ConfigFSM_inst.FrameAddressRegister\[0\] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
X_144_ net16 Inst_bitbang.data\[21\] _043_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._155_ ConfigFSM_inst._069_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.RowSelect\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._224_ ConfigFSM_inst._109_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._030_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1230__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0606_ INST_config_UART.ID_Reg\[1\] INST_config_UART.ID_Reg\[0\]
+ INST_config_UART._0205_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0206_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._265__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._393__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1253__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_127_ net10 Inst_bitbang.data\[16\] _021_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._138_ ConfigFSM_inst.state\[1\] ConfigFSM_inst._057_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._058_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._207_ ConfigFSM_inst._100_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._022_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1234__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._391_ net1 Inst_bitbang._028_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1276__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0871_ INST_config_UART._0378_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0095_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0940_ INST_config_UART._0399_ INST_config_UART._0424_ INST_config_UART._0425_
+ INST_config_UART._0407_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0117_ sky130_fd_sc_hd__o31a_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1354_ net1 INST_config_UART._0175_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XINST_config_UART._1285_ net1 INST_config_UART._0049_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1299__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0978__B2 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0978__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._374_ net1 Inst_bitbang._011_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._443_ net1 Inst_bitbang._072_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._280__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._245__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1070_ INST_config_UART._0445_ INST_config_UART._0520_ INST_config_UART.CRCReg\[10\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0525_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._0923_ INST_config_UART.HexData\[5\] INST_config_UART.HighReg\[1\]
+ INST_config_UART._0014_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0415_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0854_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[8\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0367_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0785_ INST_config_UART._0312_ INST_config_UART.HexData\[6\] INST_config_UART._0325_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0326_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._425__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1337_ net1 INST_config_UART._0172_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1268_ net1 INST_config_UART._0017_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteStrobe sky130_fd_sc_hd__dfrtp_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1199_ net1 INST_config_UART._0068_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1314__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._268__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._357_ Inst_bitbang._178_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._080_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._426_ net1 Inst_bitbang._063_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._288_ Inst_bitbang._142_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._047_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1337__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1122_ INST_config_UART.ID_Reg\[6\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART._0553_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0560_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1053_ INST_config_UART.CRCReg\[7\] INST_config_UART._0510_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_INST_config_UART._1337__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0837_ INST_config_UART._0357_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0082_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0906_ INST_config_UART.TimeToSendCounter\[11\] INST_config_UART.TimeToSendCounter\[10\]
+ INST_config_UART._0403_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0404_ sky130_fd_sc_hd__or3_1
XInst_bitbang._211_ Inst_bitbang.serial_data\[8\] Inst_bitbang.data\[8\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._102_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0768_ INST_config_UART.WriteData\[0\] INST_config_UART._0240_ INST_config_UART._0314_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0056_ sky130_fd_sc_hd__a22o_1
XINST_config_UART._0699_ INST_config_UART._0257_ INST_config_UART._0274_ INST_config_UART._0262_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0012_ sky130_fd_sc_hd__a21oi_1
XANTENNA_Inst_bitbang._368__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_091_ _012_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[4\] sky130_fd_sc_hd__buf_2
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_160_ _059_ INST_config_UART.WriteData\[26\] _045_ vssd1 vssd1 vccd1 vccd1 _060_
+ sky130_fd_sc_hd__mux2_1
XInst_bitbang._409_ net1 Inst_bitbang._046_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0622_ INST_config_UART.ReceivedWord\[3\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0218_ sky130_fd_sc_hd__buf_4
XConfigFSM_inst._171_ ConfigFSM_inst.FrameShiftState\[0\] ConfigFSM_inst.FrameShiftState\[1\]
+ ConfigFSM_inst.FrameShiftState\[2\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._080_
+ sky130_fd_sc_hd__o21ai_1
XConfigFSM_inst._240_ ConfigFSM_inst._117_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._038_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1036_ INST_config_UART._0490_ INST_config_UART._0493_ INST_config_UART._0495_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0496_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._1105_ INST_config_UART._0549_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0550_
+ sky130_fd_sc_hd__inv_2
Xinput3 SelfWriteData[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1259__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._440__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_212_ ConfigFSM_inst.WriteData\[31\] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
X_074_ net39 vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_143_ _048_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[20\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_INST_config_UART._1182__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1352__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0605_ INST_config_UART.ID_Reg\[3\] INST_config_UART.ID_Reg\[2\]
+ INST_config_UART.ID_Reg\[5\] INST_config_UART.ID_Reg\[4\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0205_ sky130_fd_sc_hd__and4_1
XConfigFSM_inst._154_ ConfigFSM_inst.FrameShiftState\[2\] ConfigFSM_inst._043_ vssd1
+ vssd1 vccd1 vccd1 ConfigFSM_inst._069_ sky130_fd_sc_hd__or2b_1
XConfigFSM_inst._223_ ConfigFSM_inst.WriteData\[21\] ConfigFSM_inst.FrameAddressRegister\[21\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1019_ INST_config_UART.CRCReg\[3\] INST_config_UART._0480_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0481_ sky130_fd_sc_hd__nor2_1
XANTENNA_Inst_bitbang._406__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._362__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_126_ _036_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[15\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1370_ net1 INST_config_UART._0191_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._429__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._390_ net1 Inst_bitbang._027_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._206_ ConfigFSM_inst.WriteData\[12\] ConfigFSM_inst.FrameAddressRegister\[12\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._137_ ConfigFSM_inst.old_reset ConfigFSM_inst.FSM_Reset vssd1 vssd1
+ vccd1 vccd1 ConfigFSM_inst._057_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1203__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1274__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0870_ INST_config_UART.ID_Reg\[10\] INST_config_UART._0221_ INST_config_UART._0375_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0378_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1220__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1370__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ net4 Inst_bitbang.data\[10\] _021_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1353_ net1 net2 net36 vssd1 vssd1 vccd1 vccd1 INST_config_UART.RxLocal
+ sky130_fd_sc_hd__dfstp_4
XINST_config_UART._1284_ net1 INST_config_UART._0048_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0999_ INST_config_UART._0014_ INST_config_UART._0463_ net39 vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0464_ sky130_fd_sc_hd__o21ai_2
XInst_bitbang._373_ net1 Inst_bitbang._010_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._442_ net1 Inst_bitbang._071_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1243__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1196__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0784_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[6\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0325_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0922_ INST_config_UART._0414_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0110_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0853_ INST_config_UART._0365_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0366_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1336_ net1 INST_config_UART._0171_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1267_ net1 INST_config_UART._0128_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1198_ net1 INST_config_UART._0067_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1266__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._287_ Inst_bitbang.serial_data\[11\] Inst_bitbang.serial_data\[12\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._142_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._356_ Inst_bitbang.serial_control\[12\] Inst_bitbang.serial_control\[13\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._425_ net1 Inst_bitbang._062_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1306__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1289__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1121_ INST_config_UART._0559_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0164_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1052_ INST_config_UART.ReceivedWord\[7\] INST_config_UART.HighReg\[3\]
+ INST_config_UART._0246_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0510_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._0878__A1 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0767_ INST_config_UART._0312_ INST_config_UART.HexData\[0\] INST_config_UART._0313_
+ INST_config_UART._0242_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0314_ sky130_fd_sc_hd__o211a_1
XINST_config_UART._0836_ INST_config_UART.ID_Reg\[16\] INST_config_UART._0223_ INST_config_UART._0356_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0357_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0905_ INST_config_UART.TimeToSendCounter\[9\] INST_config_UART._0402_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0403_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1319_ net1 INST_config_UART._0154_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[16\] sky130_fd_sc_hd__dfrtp_2
XInst_bitbang._210_ Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._101_
+ sky130_fd_sc_hd__buf_4
XINST_config_UART._0698_ INST_config_UART.ComCount\[9\] INST_config_UART._0256_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0274_ sky130_fd_sc_hd__nand2_1
XANTENNA_ConfigFSM_inst._259__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_090_ _011_ INST_config_UART.WriteData\[4\] _001_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._387__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._408_ net1 Inst_bitbang._045_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._339_ Inst_bitbang._169_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._071_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0621_ INST_config_UART.PresentState\[6\] INST_config_UART._0194_
+ INST_config_UART._0196_ INST_config_UART.PresentState\[2\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0030_ sky130_fd_sc_hd__a22o_1
XConfigFSM_inst._170_ ConfigFSM_inst.FrameShiftState\[0\] ConfigFSM_inst.FrameShiftState\[1\]
+ ConfigFSM_inst.FrameShiftState\[2\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._079_
+ sky130_fd_sc_hd__or3_2
XANTENNA_ConfigFSM_inst._258__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput4 SelfWriteData[10] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1035_ INST_config_UART.CRCReg\[5\] INST_config_UART._0494_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0495_ sky130_fd_sc_hd__xnor2_1
XANTENNA_INST_config_UART._1304__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1104_ INST_config_UART.ComState\[0\] INST_config_UART.ComTick INST_config_UART.ComState\[1\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1299__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1228__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0819_ INST_config_UART._0339_ INST_config_UART.WriteData\[13\]
+ INST_config_UART._0215_ INST_config_UART._0344_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0077_
+ sky130_fd_sc_hd__a31o_1
X_211_ ConfigFSM_inst.WriteData\[30\] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_142_ _047_ INST_config_UART.WriteData\[20\] _045_ vssd1 vssd1 vccd1 vccd1 _048_
+ sky130_fd_sc_hd__mux2_1
X_073_ Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_ConfigFSM_inst._193__A0 ConfigFSM_inst.WriteData\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1327__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0604_ INST_config_UART.ID_Reg\[10\] INST_config_UART.ID_Reg\[12\]
+ INST_config_UART.ID_Reg\[13\] INST_config_UART.ID_Reg\[11\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0204_ sky130_fd_sc_hd__and4bb_1
XConfigFSM_inst._153_ ConfigFSM_inst._068_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.RowSelect\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._222_ ConfigFSM_inst._108_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._029_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1018_ INST_config_UART._0218_ INST_config_UART._0232_ INST_config_UART._0246_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0480_ sky130_fd_sc_hd__mux2_1
XANTENNA__073__A Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._274__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0999__B1 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_125_ _035_ INST_config_UART.WriteData\[15\] _023_ vssd1 vssd1 vccd1 vccd1 _036_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._419__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._205_ ConfigFSM_inst._099_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._021_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._136_ ConfigFSM_inst._056_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._002_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1243__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0597__A_N INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_108_ _024_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[9\] sky130_fd_sc_hd__buf_2
XINST_config_UART._1352_ net1 INST_config_UART._0013_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComTick sky130_fd_sc_hd__dfrtp_4
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1283_ net1 INST_config_UART._0047_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._202__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0998_ INST_config_UART._0246_ INST_config_UART._0195_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0463_ sky130_fd_sc_hd__nor2_1
XANTENNA_INST_config_UART._1195__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._372_ net1 Inst_bitbang._009_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._441_ net1 Inst_bitbang._070_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._419__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0921_ INST_config_UART.HexData\[4\] INST_config_UART.HighReg\[0\]
+ INST_config_UART._0014_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0414_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0783_ INST_config_UART.WriteData\[5\] INST_config_UART._0240_ INST_config_UART._0324_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0061_ sky130_fd_sc_hd__a22o_1
XINST_config_UART._0852_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[8\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0365_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1335_ net1 INST_config_UART._0170_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._434__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1266_ net1 INST_config_UART._0127_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1197_ net1 INST_config_UART._0066_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._424_ net1 Inst_bitbang._061_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._286_ Inst_bitbang._141_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._046_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1210__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._355_ Inst_bitbang._177_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._079_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1360__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1346__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1051_ INST_config_UART._0504_ INST_config_UART._0506_ INST_config_UART._0502_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0509_ sky130_fd_sc_hd__a21o_1
XINST_config_UART._1120_ INST_config_UART.ID_Reg\[5\] INST_config_UART.ReceivedWord\[5\]
+ INST_config_UART._0553_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0559_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._391__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0904_ INST_config_UART.TimeToSendCounter\[8\] INST_config_UART.TimeToSendCounter\[7\]
+ INST_config_UART._0401_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0402_ sky130_fd_sc_hd__or3_2
XFILLER_0_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1233__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0766_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[0\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0313_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0835_ INST_config_UART._0355_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0356_
+ sky130_fd_sc_hd__buf_2
XINST_config_UART._0697_ INST_config_UART._0256_ INST_config_UART._0273_ INST_config_UART._0262_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0011_ sky130_fd_sc_hd__a21oi_1
XANTENNA__105__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1318_ net1 INST_config_UART._0153_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[15\] sky130_fd_sc_hd__dfstp_1
XINST_config_UART._1249_ net1 INST_config_UART._0110_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._407_ net1 Inst_bitbang._044_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._269_ Inst_bitbang._132_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._038_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._338_ Inst_bitbang.serial_control\[3\] Inst_bitbang.serial_control\[4\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0620_ INST_config_UART.PresentState\[2\] INST_config_UART._0194_
+ INST_config_UART._0196_ INST_config_UART.PresentState\[4\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0027_ sky130_fd_sc_hd__a22o_1
XANTENNA_INST_config_UART._1256__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1103_ INST_config_UART._0547_ INST_config_UART._0468_ INST_config_UART._0545_
+ INST_config_UART._0548_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0157_ sky130_fd_sc_hd__o31a_1
XANTENNA_INST_config_UART._1180__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 SelfWriteData[11] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1034_ INST_config_UART.ReceivedWord\[5\] INST_config_UART.HighReg\[1\]
+ INST_config_UART.Command\[7\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0494_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0818_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0324_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0344_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0749_ INST_config_UART.blink\[19\] INST_config_UART._0300_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0302_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1268__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1279__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_210_ ConfigFSM_inst.WriteData\[29\] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_141_ net15 Inst_bitbang.data\[20\] _043_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._221_ ConfigFSM_inst.WriteData\[19\] ConfigFSM_inst.FrameAddressRegister\[19\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0603_ INST_config_UART.ID_Reg\[8\] INST_config_UART.ID_Reg\[9\]
+ INST_config_UART.ID_Reg\[7\] INST_config_UART.ID_Reg\[6\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0203_ sky130_fd_sc_hd__and4b_1
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._152_ ConfigFSM_inst.FrameShiftState\[1\] ConfigFSM_inst._043_ vssd1
+ vssd1 vccd1 vccd1 ConfigFSM_inst._068_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1017_ INST_config_UART._0466_ INST_config_UART._0478_ INST_config_UART._0479_
+ INST_config_UART._0469_ INST_config_UART.CRCReg\[2\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0140_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_bitbang._452__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._248__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._371__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_124_ net9 Inst_bitbang.data\[15\] _021_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._204_ ConfigFSM_inst.WriteData\[11\] ConfigFSM_inst.FrameAddressRegister\[11\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._099_ sky130_fd_sc_hd__mux2_1
Xinput30 SelfWriteData[5] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._135_ ConfigFSM_inst._041_ ConfigFSM_inst._042_ ConfigFSM_inst._055_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._056_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1283__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1317__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1212__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1158__A1 INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_107_ _022_ INST_config_UART.WriteData\[9\] _023_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1282_ net1 INST_config_UART._0046_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[2\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1351_ net1 INST_config_UART._0003_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0623__D_N INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_load_slew111_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0997_ INST_config_UART.CRCReg\[0\] INST_config_UART._0460_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0462_ sky130_fd_sc_hd__nand2_1
XInst_bitbang._440_ net1 Inst_bitbang._069_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._371_ net1 Inst_bitbang._008_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0920_ INST_config_UART._0413_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0109_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0851_ INST_config_UART._0364_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0089_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0782_ INST_config_UART._0312_ INST_config_UART.HexData\[5\] INST_config_UART._0323_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0324_ sky130_fd_sc_hd__o211a_1
XINST_config_UART._1334_ net1 INST_config_UART._0169_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1265_ net1 INST_config_UART._0126_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1196_ net1 INST_config_UART._0065_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._403__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._423_ net1 Inst_bitbang._060_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._285_ Inst_bitbang.serial_data\[10\] Inst_bitbang.serial_data\[11\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._141_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._354_ Inst_bitbang.serial_control\[11\] Inst_bitbang.serial_control\[12\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1185__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1050_ INST_config_UART.CRCReg\[6\] INST_config_UART._0469_ INST_config_UART._0466_
+ INST_config_UART._0508_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0834_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] INST_config_UART.PresentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0355_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0903_ INST_config_UART.TimeToSendCounter\[6\] INST_config_UART.TimeToSendCounter\[5\]
+ INST_config_UART.TimeToSendCounter\[4\] INST_config_UART._0400_ vssd1 vssd1 vccd1
+ vccd1 INST_config_UART._0401_ sky130_fd_sc_hd__or4_2
XANTENNA__182__A ConfigFSM_inst.WriteData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._208__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0765_ INST_config_UART._0246_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0312_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_ConfigFSM_inst._202__A0 ConfigFSM_inst.WriteData\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0696_ INST_config_UART.ComCount\[7\] INST_config_UART._0255_ INST_config_UART.ComCount\[8\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0273_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._1317_ net1 INST_config_UART._0152_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[14\] sky130_fd_sc_hd__dfstp_1
XINST_config_UART._1248_ net1 INST_config_UART._0109_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__121__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1179_ net1 INST_config_UART._0025_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.PresentState\[0\] sky130_fd_sc_hd__dfstp_1
XANTENNA_Inst_bitbang._409__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._281__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._268__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._406_ net1 Inst_bitbang._043_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._337_ Inst_bitbang._168_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._070_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._199_ Inst_bitbang._095_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._005_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._268_ Inst_bitbang.serial_data\[2\] Inst_bitbang.serial_data\[3\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._132_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._396__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1102_ INST_config_UART.CRCReg\[18\] INST_config_UART._0465_ INST_config_UART._0539_
+ INST_config_UART._0544_ INST_config_UART.CRCReg\[19\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0548_
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 SelfWriteData[12] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1033_ INST_config_UART._0466_ INST_config_UART._0492_ INST_config_UART._0493_
+ INST_config_UART._0469_ INST_config_UART.CRCReg\[4\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0142_
+ sky130_fd_sc_hd__a32o_1
XINST_config_UART._0817_ INST_config_UART._0339_ INST_config_UART.WriteData\[12\]
+ INST_config_UART._0215_ INST_config_UART._0343_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0076_
+ sky130_fd_sc_hd__a31o_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1200__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1350__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0748_ INST_config_UART._0300_ INST_config_UART._0301_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1237__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0679_ INST_config_UART._0260_ INST_config_UART._0261_ INST_config_UART._0262_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._381__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_140_ _046_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[19\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1223__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0602_ INST_config_UART.Command\[5\] INST_config_UART.Command\[4\]
+ INST_config_UART.Command\[6\] INST_config_UART._0201_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0202_
+ sky130_fd_sc_hd__or4_1
XConfigFSM_inst._151_ ConfigFSM_inst._067_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.RowSelect\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._220_ ConfigFSM_inst._061_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._107_
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_bitbang._282__A Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1330__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1016_ INST_config_UART._0471_ INST_config_UART._0474_ INST_config_UART._0477_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0479_ sky130_fd_sc_hd__nand3_1
XFILLER_0_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1246__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._283__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_123_ _034_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[14\] sky130_fd_sc_hd__buf_2
XFILLER_0_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 SelfWriteData[6] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1316__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput20 SelfWriteData[25] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._203_ ConfigFSM_inst._098_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._020_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._134_ ConfigFSM_inst._044_ ConfigFSM_inst._049_ ConfigFSM_inst._054_
+ ConfigFSM_inst.state\[0\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._055_ sky130_fd_sc_hd__o31a_1
XANTENNA__190__A ConfigFSM_inst.WriteData\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._131__D_N ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1269__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._428__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._187__A Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1252__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ net39 vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._1281_ net1 INST_config_UART._0042_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1350_ net1 INST_config_UART._0002_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__185__A ConfigFSM_inst.WriteData\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0996_ INST_config_UART.CRCReg\[0\] INST_config_UART._0460_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0461_ sky130_fd_sc_hd__or2_1
XInst_bitbang._370_ net1 Inst_bitbang._007_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._442__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__124__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0781_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[5\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0323_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0850_ INST_config_UART.ID_Reg\[23\] INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART._0356_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1307__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1333_ net1 INST_config_UART._0168_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1195_ net1 INST_config_UART._0064_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[16\] sky130_fd_sc_hd__dfrtp_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1264_ net1 INST_config_UART._0125_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._443__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0979_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0314_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0452_ sky130_fd_sc_hd__and3_1
XInst_bitbang._353_ Inst_bitbang._176_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._078_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._422_ net1 Inst_bitbang._059_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._284_ Inst_bitbang._140_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._045_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0764_ INST_config_UART._0311_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0055_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0833_ INST_config_UART.RxLocal INST_config_UART._0353_ INST_config_UART._0354_
+ INST_config_UART._0222_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0081_ sky130_fd_sc_hd__o22a_1
XINST_config_UART._0902_ INST_config_UART.TimeToSendCounter\[3\] INST_config_UART.TimeToSendCounter\[2\]
+ INST_config_UART.TimeToSendCounter\[1\] INST_config_UART.TimeToSendCounter\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0400_ sky130_fd_sc_hd__or4_2
XINST_config_UART._0695_ INST_config_UART._0271_ INST_config_UART._0272_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0010_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._1316_ net1 INST_config_UART._0151_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[13\] sky130_fd_sc_hd__dfstp_1
XINST_config_UART._1247_ net1 INST_config_UART._0108_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[2\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1178_ net1 INST_config_UART._0054_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._405_ net1 Inst_bitbang._042_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._267_ Inst_bitbang._131_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._037_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._336_ Inst_bitbang.serial_control\[2\] Inst_bitbang.serial_control\[3\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._168_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._198_ Inst_bitbang.serial_data\[2\] Inst_bitbang.data\[2\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._095_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._365__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINST_config_UART._1032_ INST_config_UART._0487_ INST_config_UART._0491_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0493_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1101_ INST_config_UART.CRCReg\[19\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0547_
+ sky130_fd_sc_hd__inv_2
Xinput7 SelfWriteData[13] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__193__A ConfigFSM_inst.WriteData\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0747_ INST_config_UART.blink\[17\] INST_config_UART._0298_ INST_config_UART.blink\[18\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0301_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._0816_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0322_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0343_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._187__A0 ConfigFSM_inst.WriteData\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._0678_ INST_config_UART._0250_ INST_config_UART._0259_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0262_ sky130_fd_sc_hd__nand2b_1
XANTENNA_INST_config_UART._1206__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1277__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._319_ Inst_bitbang._158_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._062_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0601_ INST_config_UART.ID_Reg\[23\] INST_config_UART.ID_Reg\[22\]
+ INST_config_UART.Command\[3\] INST_config_UART.Command\[2\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0201_ sky130_fd_sc_hd__or4_1
XConfigFSM_inst._150_ ConfigFSM_inst.FrameShiftState\[0\] ConfigFSM_inst._043_ vssd1
+ vssd1 vccd1 vccd1 ConfigFSM_inst._067_ sky130_fd_sc_hd__or2b_1
X_199_ ConfigFSM_inst.WriteData\[18\] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__188__A ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1015_ INST_config_UART._0471_ INST_config_UART._0474_ INST_config_UART._0477_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0478_ sky130_fd_sc_hd__a21o_1
XANTENNA_ConfigFSM_inst._271__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1370__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1198__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__127__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._279_ net1 ConfigFSM_inst._034_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._181__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_122_ _033_ INST_config_UART.WriteData\[14\] _023_ vssd1 vssd1 vccd1 vccd1 _034_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._252__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1199__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._380__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1340__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 SelfWriteData[7] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput21 SelfWriteData[26] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 SelfWriteData[16] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._202_ ConfigFSM_inst.WriteData\[10\] ConfigFSM_inst.FrameAddressRegister\[10\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._098_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._133_ ConfigFSM_inst._050_ ConfigFSM_inst._051_ ConfigFSM_inst._052_
+ ConfigFSM_inst._053_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._054_ sky130_fd_sc_hd__or4b_1
XANTENNA_Inst_bitbang._371__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0633__B_N INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1292__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1213__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1221__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1363__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_105_ net34 Inst_bitbang.data\[9\] _021_ vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__mux2_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1309__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1280_ net1 INST_config_UART._0031_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_Inst_bitbang._394__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0995_ INST_config_UART._0223_ INST_config_UART._0387_ INST_config_UART._0246_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0460_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1236__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0780_ INST_config_UART.WriteData\[4\] INST_config_UART._0240_ INST_config_UART._0322_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0060_ sky130_fd_sc_hd__a22o_1
XANTENNA_INST_config_UART._1259__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1332_ net1 INST_config_UART._0167_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.Command\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1194_ net1 INST_config_UART._0063_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1263_ net1 INST_config_UART._0124_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__196__A ConfigFSM_inst.WriteData\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0978_ net111 INST_config_UART.ReceiveLED INST_config_UART._0451_
+ net39 vssd1 vssd1 vccd1 vccd1 INST_config_UART._0129_ sky130_fd_sc_hd__o22a_1
XInst_bitbang._283_ Inst_bitbang.serial_data\[9\] Inst_bitbang.serial_data\[10\] Inst_bitbang._139_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._140_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._412__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._352_ Inst_bitbang.serial_control\[10\] Inst_bitbang.serial_control\[11\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._176_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._421_ net1 Inst_bitbang._058_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._432__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0901_ INST_config_UART._0398_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0399_
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1324__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0763_ INST_config_UART._0221_ INST_config_UART.RxLocal INST_config_UART._0310_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0311_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0832_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[9\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0354_ sky130_fd_sc_hd__and3b_1
XINST_config_UART._0694_ INST_config_UART.ComCount\[7\] INST_config_UART._0255_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0272_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1315_ net1 INST_config_UART._0150_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[12\] sky130_fd_sc_hd__dfstp_1
XINST_config_UART._1246_ net1 INST_config_UART._0107_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[1\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1177_ INST_config_UART._0588_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0191_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._404_ net1 Inst_bitbang._041_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._266_ Inst_bitbang.serial_data\[1\] Inst_bitbang.serial_data\[2\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._131_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._335_ Inst_bitbang._167_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._069_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._277__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._197_ Inst_bitbang._094_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._004_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 SelfWriteData[14] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1031_ INST_config_UART._0487_ INST_config_UART._0491_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0492_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1100_ INST_config_UART.CRCReg\[18\] INST_config_UART._0469_ INST_config_UART._0545_
+ INST_config_UART._0546_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0815_ INST_config_UART._0339_ INST_config_UART.WriteData\[11\]
+ INST_config_UART._0215_ INST_config_UART._0342_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0075_
+ sky130_fd_sc_hd__a31o_1
XINST_config_UART._0746_ INST_config_UART.blink\[17\] INST_config_UART.blink\[18\]
+ INST_config_UART._0298_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0300_ sky130_fd_sc_hd__or3_1
XINST_config_UART._0677_ INST_config_UART.ComCount\[1\] INST_config_UART.ComCount\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0261_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1229_ net1 INST_config_UART._0092_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1246__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._249_ Inst_bitbang._121_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._029_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._318_ Inst_bitbang.serial_data\[26\] Inst_bitbang.serial_data\[27\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0600_ INST_config_UART.Command\[1\] INST_config_UART.Command\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0200_ sky130_fd_sc_hd__xnor2_1
X_198_ ConfigFSM_inst.WriteData\[17\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1014_ INST_config_UART.CRCReg\[2\] INST_config_UART._0476_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0729_ INST_config_UART.blink\[9\] INST_config_UART._0288_ INST_config_UART.blink\[10\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0291_ sky130_fd_sc_hd__o21ai_1
XConfigFSM_inst._278_ net1 ConfigFSM_inst._033_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1292__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_121_ net8 Inst_bitbang.data\[14\] _021_ vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._201_ ConfigFSM_inst._097_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._019_
+ sky130_fd_sc_hd__clkbuf_1
Xinput33 SelfWriteData[8] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput22 SelfWriteData[27] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 SelfWriteData[17] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._132_ ConfigFSM_inst.WriteData\[11\] ConfigFSM_inst.WriteData\[13\]
+ ConfigFSM_inst.WriteData\[12\] ConfigFSM_inst.WriteData\[15\] vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._053_ sky130_fd_sc_hd__and4_1
XANTENNA__199__A ConfigFSM_inst.WriteData\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._437__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1261__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_104_ Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__buf_4
XANTENNA_ConfigFSM_inst._241__A0 ConfigFSM_inst.WriteData\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._131__A ConfigFSM_inst.WriteData\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._261__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1188__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_233__113 vssd1 vssd1 vccd1 vccd1 _233__113/HI net113 sky130_fd_sc_hd__conb_1
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1349__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0994_ INST_config_UART._0242_ INST_config_UART.WriteData\[31\]
+ INST_config_UART._0234_ INST_config_UART._0459_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0137_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._187__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1330__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._284__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._223__A0 ConfigFSM_inst.WriteData\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._126__A ConfigFSM_inst.WriteData\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._214__A0 ConfigFSM_inst.WriteData\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1331_ net1 INST_config_UART._0166_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1183__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1262_ net1 INST_config_UART._0123_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[9\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1193_ net1 INST_config_UART._0062_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1203__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0977_ INST_config_UART.PresentState\[0\] INST_config_UART.blink\[22\]
+ INST_config_UART._0449_ INST_config_UART._0450_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0451_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1353__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._420_ net1 Inst_bitbang._057_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._282_ Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._139_
+ sky130_fd_sc_hd__clkbuf_4
XInst_bitbang._351_ Inst_bitbang._175_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._077_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._452__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._384__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1226__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0831_ INST_config_UART._0352_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0353_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._0900_ INST_config_UART.ComState\[4\] INST_config_UART.PresentState\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0398_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0762_ INST_config_UART.ComState\[0\] INST_config_UART.ComState\[2\]
+ INST_config_UART._0245_ INST_config_UART._0309_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0310_
+ sky130_fd_sc_hd__o211a_1
XINST_config_UART._0693_ INST_config_UART.ComCount\[7\] INST_config_UART._0255_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0271_ sky130_fd_sc_hd__or2_1
XANTENNA_INST_config_UART._1364__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1314_ net1 INST_config_UART._0149_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[11\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1245_ net1 INST_config_UART._0106_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexData\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1176_ INST_config_UART.ComState\[1\] INST_config_UART.ComState\[10\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0588_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._403_ net1 Inst_bitbang._040_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._265_ Inst_bitbang._130_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._036_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._196_ Inst_bitbang.serial_data\[1\] Inst_bitbang.data\[1\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._094_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1249__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._334_ Inst_bitbang.serial_control\[1\] Inst_bitbang.serial_control\[2\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._167_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._246__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._374__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 SelfWriteData[15] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1030_ INST_config_UART._0489_ INST_config_UART._0490_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0491_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0814_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0320_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0342_ sky130_fd_sc_hd__and3_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0745_ INST_config_UART.blink\[17\] INST_config_UART._0298_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0676_ INST_config_UART.ComCount\[1\] INST_config_UART.ComCount\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0260_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1228_ net1 INST_config_UART._0091_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[4\] sky130_fd_sc_hd__dfrtp_4
XINST_config_UART._1159_ INST_config_UART._0580_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0181_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._195__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1286__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._422__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1215__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._317_ Inst_bitbang._157_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._061_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._248_ Inst_bitbang.serial_data\[26\] Inst_bitbang.data\[26\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._121_ sky130_fd_sc_hd__mux2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_197_ ConfigFSM_inst.WriteData\[16\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1013_ INST_config_UART._0221_ INST_config_UART._0395_ INST_config_UART._0246_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0476_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._445__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._277_ net1 ConfigFSM_inst._032_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0659_ INST_config_UART._0246_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0247_
+ sky130_fd_sc_hd__buf_2
XINST_config_UART._0728_ INST_config_UART.blink\[9\] INST_config_UART.blink\[10\]
+ INST_config_UART._0288_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0290_ sky130_fd_sc_hd__or3_2
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 RowSelect[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_120_ _032_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[13\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._129__A ConfigFSM_inst.WriteData\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._261__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0844__A1 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._200_ ConfigFSM_inst.WriteData\[9\] ConfigFSM_inst.FrameAddressRegister\[9\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._097_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._131_ ConfigFSM_inst.WriteData\[8\] ConfigFSM_inst.WriteData\[10\]
+ ConfigFSM_inst.WriteData\[9\] ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst._052_ sky130_fd_sc_hd__or4bb_1
Xinput34 SelfWriteData[9] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 SelfWriteData[28] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 SelfWriteData[18] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_249_ ConfigFSM_inst.RowSelect\[4\] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._406__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1230__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_103_ _020_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[8\] sky130_fd_sc_hd__buf_2
XANTENNA_ConfigFSM_inst._131__B ConfigFSM_inst.WriteData\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0993_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0328_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0459_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1282__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._399__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._126__B ConfigFSM_inst.WriteData\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1330_ net1 INST_config_UART._0165_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[6\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1261_ net1 INST_config_UART._0122_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1192_ net1 INST_config_UART._0061_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0976_ net111 vssd1 vssd1 vccd1 vccd1 INST_config_UART._0450_ sky130_fd_sc_hd__inv_2
XInst_bitbang._350_ Inst_bitbang.serial_control\[9\] Inst_bitbang.serial_control\[10\]
+ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._281_ Inst_bitbang._138_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._044_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._254__S Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._421__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._251__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1178__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0830_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[9\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0352_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0761_ INST_config_UART._0197_ INST_config_UART.ComState\[2\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0309_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0692_ INST_config_UART._0255_ INST_config_UART._0270_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0009_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1313_ net1 INST_config_UART._0148_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1333__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1244_ net1 INST_config_UART._0105_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.TimeToSend
+ sky130_fd_sc_hd__dfxtp_1
XINST_config_UART._1175_ INST_config_UART._0350_ INST_config_UART.ComState\[9\] INST_config_UART._0309_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0190_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._274__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1320__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0959_ INST_config_UART._0436_ INST_config_UART._0437_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0124_ sky130_fd_sc_hd__a21oi_1
XInst_bitbang._402_ net1 Inst_bitbang._039_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._333_ Inst_bitbang._166_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._068_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._264_ Inst_bitbang.serial_data\[0\] Inst_bitbang.serial_data\[1\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._130_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._195_ Inst_bitbang._093_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._003_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._286__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1343__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0813_ INST_config_UART._0339_ INST_config_UART.WriteData\[10\]
+ INST_config_UART._0215_ INST_config_UART._0341_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0074_
+ sky130_fd_sc_hd__a31o_1
XINST_config_UART._0744_ INST_config_UART._0298_ INST_config_UART._0299_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0038_ sky130_fd_sc_hd__nand2_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0675_ INST_config_UART._0251_ INST_config_UART.ComCount\[0\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0001_ sky130_fd_sc_hd__nor2_1
XANTENNA_Inst_bitbang._374__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1158_ INST_config_UART.Data_Reg\[6\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART._0573_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0580_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1227_ net1 INST_config_UART._0090_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ReceivedWord\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1089_ INST_config_UART._0538_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0153_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1216__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1255__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._247_ Inst_bitbang._120_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._028_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._316_ Inst_bitbang.serial_data\[25\] Inst_bitbang.serial_data\[26\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._157_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1366__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_196_ ConfigFSM_inst.WriteData\[15\] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._397__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1012_ INST_config_UART._0466_ INST_config_UART._0474_ INST_config_UART._0475_
+ INST_config_UART._0469_ INST_config_UART.CRCReg\[1\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0139_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1239__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0727_ INST_config_UART.blink\[9\] INST_config_UART._0288_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._276_ net1 ConfigFSM_inst._031_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0658_ INST_config_UART.Command\[7\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0246_
+ sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._0589_ INST_config_UART.blink\[0\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0031_
+ sky130_fd_sc_hd__inv_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[6] sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1311__SET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._129__B ConfigFSM_inst.WriteData\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._124__D_N ConfigFSM_inst.WriteData\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput13 SelfWriteData[19] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._130_ ConfigFSM_inst.WriteData\[1\] ConfigFSM_inst.WriteData\[3\]
+ ConfigFSM_inst.WriteData\[20\] ConfigFSM_inst.WriteData\[0\] vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst._051_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_179_ _072_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlymetal6s2s_1
X_248_ ConfigFSM_inst.RowSelect\[3\] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
Xinput24 SelfWriteData[29] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 SelfWriteStrobe vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
XFILLER_0_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._412__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._129__C_N ConfigFSM_inst.WriteData\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._446__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._259_ net1 ConfigFSM_inst._014_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1270__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_102_ _019_ INST_config_UART.WriteData\[8\] _001_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._435__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0992_ INST_config_UART._0242_ INST_config_UART.WriteData\[30\]
+ INST_config_UART._0234_ INST_config_UART._0458_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0136_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._368__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._1191_ net1 INST_config_UART._0060_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1260_ net1 INST_config_UART._0121_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__104__A Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0975_ INST_config_UART._0443_ INST_config_UART._0446_ INST_config_UART._0447_
+ INST_config_UART._0448_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0449_ sky130_fd_sc_hd__or4_1
XANTENNA_INST_config_UART._1192__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._280_ Inst_bitbang.serial_data\[8\] Inst_bitbang.serial_data\[9\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1209__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0760_ INST_config_UART._0308_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0054_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1272__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1312_ net1 INST_config_UART._0147_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[9\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0691_ INST_config_UART.ComCount\[6\] INST_config_UART._0254_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0270_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._1243_ net1 INST_config_UART._0014_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HexWriteStrobe sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1174_ INST_config_UART._0587_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0189_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1302__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0892__B1 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._0889_ INST_config_UART._0390_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0101_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0958_ INST_config_UART.TimeToSendCounter\[10\] INST_config_UART._0403_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0437_ sky130_fd_sc_hd__nand2_1
XInst_bitbang._401_ net1 Inst_bitbang._038_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._263_ Inst_bitbang._129_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._035_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._332_ Inst_bitbang.serial_control\[0\] Inst_bitbang.serial_control\[1\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._194_ Inst_bitbang.serial_data\[0\] Inst_bitbang.data\[0\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._093_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1295__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._255__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._383__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0812_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0318_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0341_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0743_ INST_config_UART.blink\[15\] INST_config_UART._0296_ INST_config_UART.blink\[16\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0299_ sky130_fd_sc_hd__o21ai_1
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0674_ INST_config_UART._0251_ INST_config_UART._0259_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1157_ INST_config_UART._0579_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0180_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1088_ INST_config_UART._0537_ INST_config_UART._0535_ INST_config_UART.CRCReg\[15\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0538_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1226_ net1 INST_config_UART._0089_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__202__A ConfigFSM_inst.WriteData\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1295__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1224__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._315_ Inst_bitbang._156_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._060_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._246_ Inst_bitbang.serial_data\[25\] Inst_bitbang.data\[25\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_ConfigFSM_inst._264__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_195_ ConfigFSM_inst.WriteData\[14\] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1310__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1011_ INST_config_UART.CRCReg\[0\] INST_config_UART._0460_ INST_config_UART._0471_
+ INST_config_UART._0473_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0726_ INST_config_UART._0288_ INST_config_UART._0289_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0052_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0657_ INST_config_UART._0195_ INST_config_UART._0245_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._275_ net1 ConfigFSM_inst._030_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1209_ net1 INST_config_UART._0078_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__168__S Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1333__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_ConfigFSM_inst._287__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._229_ Inst_bitbang.serial_data\[17\] Inst_bitbang.data\[17\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 SelfWriteData[1] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 SelfWriteData[2] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._364__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput36 resetn vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_16
X_247_ ConfigFSM_inst.RowSelect\[2\] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._270__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_178_ _071_ INST_config_UART.WriteStrobe net39 vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1206__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1356__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0709_ INST_config_UART.blink\[0\] INST_config_UART.blink\[1\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0042_ sky130_fd_sc_hd__xnor2_1
XConfigFSM_inst._258_ net1 ConfigFSM_inst._013_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._189_ ConfigFSM_inst.WriteData\[4\] ConfigFSM_inst.FrameAddressRegister\[4\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._091_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._415__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._387__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_101_ net33 Inst_bitbang.data\[8\] _000_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1229__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0991_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0326_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0458_ sky130_fd_sc_hd__and3_1
XANTENNA_INST_config_UART._1327__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1238__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._208__A0 ConfigFSM_inst.WriteData\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._402__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1190_ net1 INST_config_UART._0059_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0974_ INST_config_UART.CRCReg\[16\] INST_config_UART.CRCReg\[17\]
+ INST_config_UART.CRCReg\[19\] INST_config_UART.CRCReg\[18\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0448_ sky130_fd_sc_hd__or4b_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1249__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._430__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._425__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__205__A ConfigFSM_inst.WriteData\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0690_ INST_config_UART._0259_ INST_config_UART._0269_ INST_config_UART._0251_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0008_ sky130_fd_sc_hd__a21o_1
XINST_config_UART._1311_ net1 INST_config_UART._0146_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[8\] sky130_fd_sc_hd__dfstp_1
XINST_config_UART._1242_ net1 INST_config_UART._0104_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HighReg\[3\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1173_ INST_config_UART.ComState\[3\] INST_config_UART.ComState\[6\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0587_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._448__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1342__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._400_ net1 Inst_bitbang._037_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0888_ INST_config_UART._0387_ INST_config_UART.HighReg\[0\] INST_config_UART._0389_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0390_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0957_ INST_config_UART.TimeToSendCounter\[10\] INST_config_UART._0403_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0436_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._262_ Inst_bitbang.s_data_sample\[3\] Inst_bitbang.serial_data\[0\]
+ Inst_bitbang._128_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._129_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._331_ Inst_bitbang._165_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._067_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._193_ Inst_bitbang._088_ Inst_bitbang._092_ vssd1 vssd1 vccd1 vccd1
+ Inst_bitbang._002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._0811_ INST_config_UART._0339_ INST_config_UART.WriteData\[9\] INST_config_UART._0215_
+ INST_config_UART._0340_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0073_ sky130_fd_sc_hd__a31o_1
XANTENNA_INST_config_UART._0874__A1 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0742_ INST_config_UART.blink\[14\] INST_config_UART.blink\[15\]
+ INST_config_UART.blink\[16\] INST_config_UART._0294_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0298_
+ sky130_fd_sc_hd__or4_2
XFILLER_0_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0673_ INST_config_UART.ComCount\[11\] INST_config_UART._0258_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0259_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1225_ net1 INST_config_UART._0088_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[22\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1156_ INST_config_UART.Data_Reg\[5\] INST_config_UART.ReceivedWord\[5\]
+ INST_config_UART._0573_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0579_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1087_ INST_config_UART._0442_ INST_config_UART._0465_ INST_config_UART._0529_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0537_ sky130_fd_sc_hd__and3_1
XANTENNA_INST_config_UART._1262__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._314_ Inst_bitbang.serial_data\[24\] Inst_bitbang.serial_data\[25\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._156_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._245_ Inst_bitbang._119_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._027_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1264__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_194_ ConfigFSM_inst.WriteData\[13\] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1010_ INST_config_UART.CRCReg\[0\] INST_config_UART._0460_ INST_config_UART._0471_
+ INST_config_UART._0473_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0474_ sky130_fd_sc_hd__nand4_1
XINST_config_UART._0725_ INST_config_UART.blink\[7\] INST_config_UART._0286_ INST_config_UART.blink\[8\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0289_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._0656_ INST_config_UART.RxLocal INST_config_UART.ComState\[0\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0245_ sky130_fd_sc_hd__nand2_1
XConfigFSM_inst._274_ net1 ConfigFSM_inst._029_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1208_ net1 INST_config_UART._0077_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1285__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[8] sky130_fd_sc_hd__buf_2
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1139_ INST_config_UART._0569_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0172_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._228_ Inst_bitbang._110_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._019_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._0829__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._0829__B2 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 s_clk vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
X_177_ net35 Inst_bitbang.strobe Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _071_
+ sky130_fd_sc_hd__mux2_1
Xinput15 SelfWriteData[20] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 SelfWriteData[30] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_246_ ConfigFSM_inst.RowSelect\[1\] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1186__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._257_ net1 ConfigFSM_inst._012_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0708_ INST_config_UART._0279_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0018_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0639_ INST_config_UART._0214_ INST_config_UART.GetWordState\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0234_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._188_ ConfigFSM_inst._090_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._013_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._254__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1300__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_100_ _018_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[7\] sky130_fd_sc_hd__buf_2
XFILLER_0_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0990_ INST_config_UART._0242_ INST_config_UART.WriteData\[29\]
+ INST_config_UART._0234_ INST_config_UART._0457_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0135_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_INST_config_UART._1367__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_229_ ConfigFSM_inst.FrameAddressRegister\[16\] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._277__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1323__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._249__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_bitbang._194__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._377__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1346__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0973_ INST_config_UART.CRCReg\[6\] INST_config_UART.CRCReg\[7\]
+ INST_config_UART.CRCReg\[10\] INST_config_UART.CRCReg\[11\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0447_ sky130_fd_sc_hd__or4b_1
XANTENNA_Inst_bitbang._377__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1219__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1317__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1289__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1218__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1369__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1310_ net1 INST_config_UART._0145_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[7\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1241_ net1 INST_config_UART._0103_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HighReg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1172_ INST_config_UART._0586_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0188_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0956_ INST_config_UART._0403_ INST_config_UART._0435_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0123_ sky130_fd_sc_hd__a21oi_1
XInst_bitbang._330_ Inst_bitbang.s_data_sample\[3\] Inst_bitbang.serial_control\[0\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._165_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0887_ INST_config_UART._0388_ INST_config_UART._0233_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0389_ sky130_fd_sc_hd__or2_2
XInst_bitbang._261_ Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._128_
+ sky130_fd_sc_hd__buf_4
XInst_bitbang._192_ Inst_bitbang._083_ Inst_bitbang._084_ Inst_bitbang._085_ Inst_bitbang._090_
+ Inst_bitbang._091_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._092_ sky130_fd_sc_hd__a41o_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1191__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._264__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0810_ INST_config_UART._0335_ INST_config_UART.GetWordState\[1\]
+ INST_config_UART._0316_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0340_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0741_ INST_config_UART.blink\[15\] INST_config_UART._0296_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._392__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0672_ INST_config_UART.ComCount\[10\] INST_config_UART._0257_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0258_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1155_ INST_config_UART._0578_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0179_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1224_ net1 INST_config_UART._0087_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._415__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1086_ INST_config_UART.CRCReg\[14\] INST_config_UART._0535_ INST_config_UART._0536_
+ INST_config_UART.CRCReg\[13\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0152_ sky130_fd_sc_hd__a22o_1
XANTENNA_Inst_bitbang._409__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0939_ INST_config_UART.TimeToSendCounter\[3\] INST_config_UART._0422_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0425_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._313_ Inst_bitbang._155_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._059_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._244_ Inst_bitbang.serial_data\[24\] Inst_bitbang.data\[24\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._119_ sky130_fd_sc_hd__mux2_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1233__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_193_ ConfigFSM_inst.WriteData\[12\] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._438__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output39_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._231__A Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0724_ INST_config_UART.blink\[7\] INST_config_UART.blink\[8\] INST_config_UART._0286_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0288_ sky130_fd_sc_hd__or3_2
XConfigFSM_inst._273_ net1 ConfigFSM_inst._028_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0655_ INST_config_UART._0243_ INST_config_UART._0211_ net39 INST_config_UART._0244_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0028_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[9] sky130_fd_sc_hd__buf_2
XFILLER_0_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1207_ net1 INST_config_UART._0076_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[12\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1138_ INST_config_UART.Command\[5\] INST_config_UART.ReceivedWord\[5\]
+ INST_config_UART._0563_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1069_ INST_config_UART._0466_ INST_config_UART._0523_ INST_config_UART._0524_
+ INST_config_UART._0468_ INST_config_UART.CRCReg\[9\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0147_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._227_ Inst_bitbang.serial_data\[16\] Inst_bitbang.data\[16\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._110_ sky130_fd_sc_hd__mux2_1
Xinput38 s_data vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 SelfWriteData[31] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 SelfWriteData[21] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_245_ ConfigFSM_inst.RowSelect\[0\] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
X_176_ _070_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[31\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1252__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0707_ INST_config_UART._0244_ INST_config_UART._0192_ INST_config_UART._0193_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0279_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._256_ net1 ConfigFSM_inst._011_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0638_ INST_config_UART.ReceiveState INST_config_UART._0233_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0014_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._187_ ConfigFSM_inst.WriteData\[3\] ConfigFSM_inst.FrameAddressRegister\[3\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._424__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1275__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_228_ ConfigFSM_inst.FrameAddressRegister\[15\] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
X_159_ net21 Inst_bitbang.data\[26\] _043_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1336__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._239_ ConfigFSM_inst.WriteData\[29\] ConfigFSM_inst.FrameAddressRegister\[29\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._117_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1154__A1 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1298__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._0972_ INST_config_UART.CRCReg\[0\] INST_config_UART.CRCReg\[1\]
+ INST_config_UART._0444_ INST_config_UART._0445_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0446_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_INST_config_UART._1136__A1 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1258__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1313__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._267__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1240_ net1 INST_config_UART._0102_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.HighReg\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1118__A1 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1171_ INST_config_UART.ComState\[4\] INST_config_UART.ComState\[7\]
+ INST_config_UART._0350_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0586_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0886_ INST_config_UART.ReceiveState vssd1 vssd1 vccd1 vccd1 INST_config_UART._0388_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._0955_ INST_config_UART.TimeToSendCounter\[9\] INST_config_UART._0402_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._260_ Inst_bitbang.s_clk_sample\[3\] Inst_bitbang.s_clk_sample\[2\]
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._127_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1351__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._191_ Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 Inst_bitbang._091_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._1369_ net1 INST_config_UART._0190_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1336__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._389_ net1 Inst_bitbang._026_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._367__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0740_ INST_config_UART._0296_ INST_config_UART._0297_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0671_ INST_config_UART.ComCount\[9\] INST_config_UART._0256_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0257_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1154_ INST_config_UART.Data_Reg\[4\] INST_config_UART.ReceivedWord\[4\]
+ INST_config_UART._0573_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0578_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1209__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1223_ net1 INST_config_UART._0086_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[20\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1085_ INST_config_UART._0442_ INST_config_UART._0465_ INST_config_UART._0529_
+ INST_config_UART.CRCReg\[12\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0536_ sky130_fd_sc_hd__and4b_1
XANTENNA_INST_config_UART._1359__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1027__A0 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0869_ INST_config_UART._0377_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0094_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0938_ INST_config_UART._0400_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0424_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._449__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._243_ Inst_bitbang._118_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._026_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._312_ Inst_bitbang.serial_data\[23\] Inst_bitbang.serial_data\[24\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1018__A0 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_192_ ConfigFSM_inst.WriteData\[11\] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1273__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1202__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0723_ INST_config_UART.blink\[7\] INST_config_UART._0286_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0051_ sky130_fd_sc_hd__xnor2_1
XConfigFSM_inst._272_ net1 ConfigFSM_inst._027_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0654_ INST_config_UART.TimeToSend vssd1 vssd1 vccd1 vccd1 INST_config_UART._0244_
+ sky130_fd_sc_hd__inv_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 LongFrameStrobe sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1068_ INST_config_UART._0445_ INST_config_UART._0520_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0524_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1206_ net1 INST_config_UART._0075_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1181__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1137_ INST_config_UART._0568_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0171_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._226_ Inst_bitbang._109_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._018_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._229__A0 ConfigFSM_inst.WriteData\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._405__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_244_ ConfigFSM_inst.FrameAddressRegister\[31\] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
Xinput28 SelfWriteData[3] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 SelfWriteData[22] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_175_ _069_ INST_config_UART.WriteData\[31\] net39 vssd1 vssd1 vccd1 vccd1 _070_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1195__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0706_ INST_config_UART._0278_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0016_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0637_ INST_config_UART._0220_ INST_config_UART._0232_ INST_config_UART._0193_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0233_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._186_ ConfigFSM_inst._089_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._012_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._255_ net1 ConfigFSM_inst._010_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._428__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._209_ Inst_bitbang._100_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._010_
+ sky130_fd_sc_hd__clkbuf_1
X_227_ ConfigFSM_inst.FrameAddressRegister\[14\] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_089_ net29 Inst_bitbang.data\[4\] _000_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__mux2_1
X_158_ _058_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[25\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_INST_config_UART._1305__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._169_ ConfigFSM_inst.FrameShiftState\[1\] ConfigFSM_inst._076_ ConfigFSM_inst._075_
+ ConfigFSM_inst._078_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._006_ sky130_fd_sc_hd__a22o_1
XConfigFSM_inst._238_ ConfigFSM_inst._116_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._037_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._258__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1242__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0971_ INST_config_UART.CRCReg\[8\] INST_config_UART.CRCReg\[9\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0445_ sky130_fd_sc_hd__and2_1
XANTENNA_Inst_bitbang._386__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1298__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1265__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1227__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1170_ INST_config_UART._0585_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0187_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0885_ INST_config_UART._0223_ INST_config_UART._0385_ INST_config_UART._0386_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0387_ sky130_fd_sc_hd__a21bo_1
XINST_config_UART._0954_ INST_config_UART._0399_ INST_config_UART._0433_ INST_config_UART._0434_
+ INST_config_UART._0407_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0122_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1288__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1299_ net1 INST_config_UART._0041_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[19\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._190_ Inst_bitbang.serial_control\[3\] Inst_bitbang.serial_control\[2\]
+ Inst_bitbang.serial_control\[1\] vssd1 vssd1 vccd1 vccd1 Inst_bitbang._090_ sky130_fd_sc_hd__nor3_1
XANTENNA_INST_config_UART._1320__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1368_ net1 INST_config_UART._0189_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._388_ net1 Inst_bitbang._025_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._0859__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0859__B2 INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_ConfigFSM_inst._273__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0670_ INST_config_UART.ComCount\[7\] INST_config_UART.ComCount\[8\]
+ INST_config_UART._0255_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0256_ sky130_fd_sc_hd__or3_1
XINST_config_UART._1084_ INST_config_UART._0442_ INST_config_UART._0467_ INST_config_UART._0529_
+ INST_config_UART._0192_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0535_ sky130_fd_sc_hd__a31oi_1
XINST_config_UART._1153_ INST_config_UART._0577_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0178_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1222_ net1 INST_config_UART._0085_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0868_ INST_config_UART.ID_Reg\[9\] INST_config_UART._0222_ INST_config_UART._0375_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0377_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0937_ INST_config_UART._0422_ INST_config_UART._0423_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0116_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0799_ INST_config_UART._0243_ INST_config_UART.WriteData\[20\]
+ INST_config_UART._0236_ INST_config_UART._0333_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0068_
+ sky130_fd_sc_hd__a31o_1
XInst_bitbang._242_ Inst_bitbang.serial_data\[23\] Inst_bitbang.data\[23\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._118_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._311_ Inst_bitbang._154_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._058_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._257__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1303__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._418__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_191_ ConfigFSM_inst.WriteData\[10\] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1242__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0722_ INST_config_UART._0286_ INST_config_UART._0287_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0050_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0653_ INST_config_UART._0242_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0243_
+ sky130_fd_sc_hd__clkbuf_4
XConfigFSM_inst._271_ net1 ConfigFSM_inst._026_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1205_ net1 INST_config_UART._0074_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ReceiveLED sky130_fd_sc_hd__buf_2
XANTENNA_ConfigFSM_inst._183__A0 ConfigFSM_inst.WriteData\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1067_ INST_config_UART.CRCReg\[8\] INST_config_UART._0520_ INST_config_UART.CRCReg\[9\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0523_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1326__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1136_ INST_config_UART.Command\[4\] INST_config_UART.ReceivedWord\[4\]
+ INST_config_UART._0563_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0568_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._0612__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._225_ Inst_bitbang.serial_data\[15\] Inst_bitbang.data\[15\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_243_ ConfigFSM_inst.FrameAddressRegister\[30\] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
Xinput18 SelfWriteData[23] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 SelfWriteData[4] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1349__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_174_ net27 Inst_bitbang.data\[31\] Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _069_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0705_ INST_config_UART.PresentState\[6\] INST_config_UART._0192_
+ INST_config_UART._0233_ INST_config_UART._0277_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0278_
+ sky130_fd_sc_hd__or4_1
XINST_config_UART._0636_ INST_config_UART._0218_ INST_config_UART._0221_ INST_config_UART._0227_
+ INST_config_UART._0228_ INST_config_UART._0231_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0232_
+ sky130_fd_sc_hd__o311ai_4
XConfigFSM_inst._185_ ConfigFSM_inst.WriteData\[2\] ConfigFSM_inst.FrameAddressRegister\[2\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._089_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._254_ net1 ConfigFSM_inst.FrameStrobe net112 vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst.oldFrameStrobe sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1119_ INST_config_UART._0558_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0163_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._433__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._208_ Inst_bitbang.serial_data\[7\] Inst_bitbang.data\[7\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._100_ sky130_fd_sc_hd__mux2_1
X_226_ ConfigFSM_inst.FrameAddressRegister\[13\] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
X_157_ _057_ INST_config_UART.WriteData\[25\] _045_ vssd1 vssd1 vccd1 vccd1 _058_
+ sky130_fd_sc_hd__mux2_1
X_088_ _010_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[3\] sky130_fd_sc_hd__buf_2
XFILLER_0_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1345__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._237_ ConfigFSM_inst.WriteData\[28\] ConfigFSM_inst.FrameAddressRegister\[28\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._116_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0619_ INST_config_UART._0215_ INST_config_UART._0217_ INST_config_UART.PresentState\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0024_ sky130_fd_sc_hd__a21oi_1
XConfigFSM_inst._168_ ConfigFSM_inst.FrameShiftState\[0\] ConfigFSM_inst.FrameShiftState\[1\]
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1194__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINST_config_UART._0970_ INST_config_UART.CRCReg\[2\] INST_config_UART.CRCReg\[3\]
+ INST_config_UART.CRCReg\[4\] INST_config_UART.CRCReg\[5\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0444_ sky130_fd_sc_hd__or4_1
X_209_ ConfigFSM_inst.WriteData\[28\] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._418__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1267__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._0953_ INST_config_UART.TimeToSendCounter\[7\] INST_config_UART._0401_
+ INST_config_UART.TimeToSendCounter\[8\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0434_
+ sky130_fd_sc_hd__o21a_1
XINST_config_UART._0884_ INST_config_UART.ReceivedWord\[0\] INST_config_UART.ReceivedWord\[3\]
+ INST_config_UART._0225_ INST_config_UART._0384_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0386_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1367_ net1 INST_config_UART._0188_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[4\] sky130_fd_sc_hd__dfrtp_2
XINST_config_UART._1298_ net1 INST_config_UART._0040_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_bitbang._390__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1232__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._387_ net1 Inst_bitbang._024_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1221_ net1 INST_config_UART._0084_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[18\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1189__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._261__A Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1083_ INST_config_UART._0533_ INST_config_UART._0468_ INST_config_UART._0532_
+ INST_config_UART._0534_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0151_ sky130_fd_sc_hd__o31a_1
XINST_config_UART._1152_ INST_config_UART.Data_Reg\[3\] INST_config_UART._0218_ INST_config_UART._0573_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0577_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._370__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._200__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0936_ INST_config_UART.TimeToSendCounter\[2\] INST_config_UART._0420_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0423_ sky130_fd_sc_hd__nand2_1
XANTENNA_INST_config_UART._1255__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0867_ INST_config_UART._0376_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0093_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0798_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0322_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0333_ sky130_fd_sc_hd__and3_1
XInst_bitbang._310_ Inst_bitbang.serial_data\[22\] Inst_bitbang.serial_data\[23\]
+ Inst_bitbang._150_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._154_ sky130_fd_sc_hd__mux2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_bitbang._241_ Inst_bitbang._117_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._025_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_190_ ConfigFSM_inst.WriteData\[9\] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._439_ net1 Inst_bitbang._068_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1282__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._270_ net1 ConfigFSM_inst._025_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.FrameAddressRegister\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1278__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0652_ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0242_
+ sky130_fd_sc_hd__buf_2
XINST_config_UART._0721_ INST_config_UART.blink\[5\] INST_config_UART._0284_ INST_config_UART.blink\[6\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0287_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1204_ net1 INST_config_UART._0073_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1135_ INST_config_UART._0567_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0170_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 RowSelect[0] sky130_fd_sc_hd__buf_2
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1066_ INST_config_UART._0466_ INST_config_UART._0521_ INST_config_UART._0522_
+ INST_config_UART._0469_ INST_config_UART.CRCReg\[8\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0146_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0919_ INST_config_UART.HexData\[3\] INST_config_UART._0232_ INST_config_UART._0014_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0759__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_bitbang._224_ Inst_bitbang._108_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._017_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 SelfWriteData[24] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_242_ ConfigFSM_inst.FrameAddressRegister\[29\] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
X_173_ _068_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[30\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._451__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0704_ INST_config_UART.PresentState\[2\] INST_config_UART.PresentState\[4\]
+ INST_config_UART.PresentState\[5\] INST_config_UART.PresentState\[0\] vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0277_ sky130_fd_sc_hd__or4_1
XConfigFSM_inst._253_ net1 ConfigFSM_inst._001_ net112 vssd1 vssd1 vccd1 vccd1 net104
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._247__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0635_ INST_config_UART._0226_ INST_config_UART._0229_ INST_config_UART._0230_
+ INST_config_UART._0225_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0231_ sky130_fd_sc_hd__a211o_1
XConfigFSM_inst._184_ ConfigFSM_inst._088_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._011_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1118_ INST_config_UART.ID_Reg\[4\] INST_config_UART.ReceivedWord\[4\]
+ INST_config_UART._0553_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1049_ INST_config_UART._0502_ INST_config_UART._0507_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__074__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._207_ Inst_bitbang._099_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._009_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._402__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1316__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_087_ _009_ INST_config_UART.WriteData\[3\] _001_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__mux2_1
X_225_ ConfigFSM_inst.FrameAddressRegister\[12\] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
X_156_ net20 Inst_bitbang.data\[25\] _043_ vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._236_ ConfigFSM_inst._115_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._036_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0618_ INST_config_UART._0216_ INST_config_UART.GetWordState\[3\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._167_ ConfigFSM_inst._077_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._005_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1339__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1312__SET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._267__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_208_ ConfigFSM_inst.WriteData\[27\] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_139_ _044_ INST_config_UART.WriteData\[19\] _045_ vssd1 vssd1 vccd1 vccd1 _046_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._395__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._219_ ConfigFSM_inst._106_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._028_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1236__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._210__A0 ConfigFSM_inst.WriteData\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0883_ INST_config_UART.ReceivedWord\[3\] INST_config_UART._0384_
+ INST_config_UART._0219_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0385_ sky130_fd_sc_hd__a21oi_1
XINST_config_UART._0952_ INST_config_UART._0402_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0433_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1297_ net1 INST_config_UART._0039_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1184__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1366_ net1 INST_config_UART._0187_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._386_ net1 Inst_bitbang._023_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._408__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._280__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1151_ INST_config_UART._0576_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0177_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1220_ net1 INST_config_UART._0083_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[17\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1082_ INST_config_UART.CRCReg\[12\] INST_config_UART._0466_ INST_config_UART._0529_
+ INST_config_UART.CRCReg\[13\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0534_ sky130_fd_sc_hd__a31o_1
XANTENNA_ConfigFSM_inst._282__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0866_ INST_config_UART.ID_Reg\[8\] INST_config_UART._0223_ INST_config_UART._0375_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0376_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0935_ INST_config_UART.TimeToSendCounter\[2\] INST_config_UART._0420_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0422_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._240_ Inst_bitbang.serial_data\[22\] Inst_bitbang.data\[22\] Inst_bitbang._112_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0797_ INST_config_UART._0243_ INST_config_UART.WriteData\[19\]
+ INST_config_UART._0236_ INST_config_UART._0332_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0067_
+ sky130_fd_sc_hd__a31o_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1349_ net1 INST_config_UART._0012_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1216__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._427__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._369_ net1 Inst_bitbang._006_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._438_ net1 Inst_bitbang._067_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1251__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._380__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0720_ INST_config_UART.blink\[4\] INST_config_UART.blink\[5\] INST_config_UART.blink\[6\]
+ INST_config_UART._0282_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0286_ sky130_fd_sc_hd__or4_2
XINST_config_UART._0651_ INST_config_UART.PresentState\[5\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0241_ sky130_fd_sc_hd__inv_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 RowSelect[1] sky130_fd_sc_hd__buf_2
XINST_config_UART._1203_ net1 INST_config_UART._0072_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[8\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1134_ INST_config_UART.Command\[3\] INST_config_UART._0218_ INST_config_UART._0563_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1065_ INST_config_UART.CRCReg\[8\] INST_config_UART._0520_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1339__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1222__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0918_ INST_config_UART._0412_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0108_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._0849_ INST_config_UART._0363_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0088_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._223_ Inst_bitbang.serial_data\[14\] Inst_bitbang.data\[14\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ ConfigFSM_inst.FrameAddressRegister\[28\] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
X_172_ _067_ INST_config_UART.WriteData\[30\] net39 vssd1 vssd1 vccd1 vccd1 _068_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1245__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0703_ INST_config_UART._0276_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0003_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._183_ ConfigFSM_inst.WriteData\[1\] ConfigFSM_inst.FrameAddressRegister\[1\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._088_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._252_ net1 ConfigFSM_inst._004_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._206__S Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0634_ INST_config_UART.ReceivedWord\[3\] INST_config_UART.ReceivedWord\[2\]
+ INST_config_UART.ReceivedWord\[1\] INST_config_UART.ReceivedWord\[0\] vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0230_ sky130_fd_sc_hd__o211a_1
XINST_config_UART._1048_ INST_config_UART._0504_ INST_config_UART._0506_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0507_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1117_ INST_config_UART._0557_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0162_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._0623__B INST_config_UART.ReceivedWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._206_ Inst_bitbang.serial_data\[6\] Inst_bitbang.data\[6\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._099_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1268__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._130__D_N ConfigFSM_inst.WriteData\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._442__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0840__A1 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_224_ ConfigFSM_inst.FrameAddressRegister\[11\] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
X_086_ net28 Inst_bitbang.data\[3\] _000_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_155_ _056_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[24\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0617_ INST_config_UART.ByteWriteStrobe vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0216_ sky130_fd_sc_hd__buf_2
XConfigFSM_inst._166_ ConfigFSM_inst._075_ ConfigFSM_inst._076_ ConfigFSM_inst.FrameShiftState\[0\]
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._077_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._235_ ConfigFSM_inst.WriteData\[27\] ConfigFSM_inst.FrameAddressRegister\[27\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._441__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_207_ ConfigFSM_inst.WriteData\[26\] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_138_ net39 vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._364__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__109__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._0629__A INST_config_UART.ReceivedWord\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._149_ ConfigFSM_inst._066_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._001_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._218_ ConfigFSM_inst.WriteData\[18\] ConfigFSM_inst.FrameAddressRegister\[18\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1306__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1205__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1276__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0882_ INST_config_UART.ReceivedWord\[1\] INST_config_UART.ReceivedWord\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0384_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0951_ INST_config_UART._0399_ INST_config_UART._0431_ INST_config_UART._0432_
+ INST_config_UART._0407_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0121_ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_INST_config_UART._1329__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1296_ net1 INST_config_UART._0038_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[16\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1365_ net1 INST_config_UART._0186_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_bitbang._385_ net1 Inst_bitbang._022_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._195__A0 ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XINST_config_UART._1081_ INST_config_UART.CRCReg\[13\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0533_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._1150_ INST_config_UART.Data_Reg\[2\] INST_config_UART._0221_ INST_config_UART._0573_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0576_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._251__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__183__A ConfigFSM_inst.WriteData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0865_ INST_config_UART._0374_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0375_
+ sky130_fd_sc_hd__buf_2
XINST_config_UART._0796_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0320_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0332_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0934_ INST_config_UART._0420_ INST_config_UART._0421_ INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0115_ sky130_fd_sc_hd__a21oi_1
XANTENNA_INST_config_UART._1198__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1279_ net1 INST_config_UART._0137_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[31\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1348_ net1 INST_config_UART._0011_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._368_ net1 Inst_bitbang._005_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._437_ net1 Inst_bitbang.s_clk_sample\[2\] net111 vssd1 vssd1 vccd1 vccd1
+ Inst_bitbang.s_clk_sample\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._299_ Inst_bitbang.serial_data\[17\] Inst_bitbang.serial_data\[18\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._148_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1291__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1220__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0650_ INST_config_UART.PresentState\[4\] INST_config_UART._0194_
+ INST_config_UART._0198_ INST_config_UART.PresentState\[0\] vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 RowSelect[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1064_ INST_config_UART.CRCReg\[8\] INST_config_UART._0520_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0521_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1133_ INST_config_UART._0566_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0169_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[26] sky130_fd_sc_hd__buf_2
XINST_config_UART._1202_ net1 INST_config_UART._0071_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[23\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1308__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0779_ INST_config_UART._0312_ INST_config_UART.HexData\[4\] INST_config_UART._0321_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0322_ sky130_fd_sc_hd__o211a_1
XINST_config_UART._0917_ INST_config_UART.HexData\[2\] INST_config_UART._0395_ INST_config_UART._0014_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0848_ INST_config_UART.ID_Reg\[22\] INST_config_UART.ReceivedWord\[6\]
+ INST_config_UART._0356_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._222_ Inst_bitbang._107_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._016_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._270__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1197__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_240_ ConfigFSM_inst.FrameAddressRegister\[27\] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_171_ net26 Inst_bitbang.data\[30\] Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _067_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0633_ INST_config_UART.ReceivedWord\[3\] INST_config_UART._0221_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0229_ sky130_fd_sc_hd__or2b_1
XANTENNA_Inst_bitbang._389__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._251_ net1 ConfigFSM_inst._003_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XConfigFSM_inst._182_ ConfigFSM_inst._087_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._010_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0702_ INST_config_UART._0251_ INST_config_UART.ComCount\[11\] INST_config_UART._0258_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0276_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1047_ INST_config_UART._0484_ INST_config_UART._0478_ INST_config_UART._0482_
+ INST_config_UART._0505_ INST_config_UART._0481_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0506_
+ sky130_fd_sc_hd__a311o_1
XINST_config_UART._1116_ INST_config_UART.ID_Reg\[3\] INST_config_UART._0218_ INST_config_UART._0553_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0557_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._193__A Inst_bitbang._088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._370__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._205_ Inst_bitbang._098_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._008_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._411__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_223_ ConfigFSM_inst.FrameAddressRegister\[10\] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
X_085_ _008_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[2\] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1212__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_154_ _055_ INST_config_UART.WriteData\[24\] _045_ vssd1 vssd1 vccd1 vccd1 _056_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1362__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__191__A ConfigFSM_inst.WriteData\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0616_ INST_config_UART._0214_ INST_config_UART.GetWordState\[1\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0215_ sky130_fd_sc_hd__nand2_4
XConfigFSM_inst._165_ ConfigFSM_inst._042_ ConfigFSM_inst._073_ ConfigFSM_inst._057_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._076_ sky130_fd_sc_hd__o21a_1
XConfigFSM_inst._234_ ConfigFSM_inst._114_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._035_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._393__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__130__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1323__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1235__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_206_ ConfigFSM_inst.WriteData\[25\] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._276__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_137_ net13 Inst_bitbang.data\[19\] _043_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__186__A ConfigFSM_inst.WriteData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._217_ ConfigFSM_inst._105_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._027_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1258__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._148_ ConfigFSM_inst.oldFrameStrobe ConfigFSM_inst.FrameStrobe vssd1
+ vssd1 vccd1 vccd1 ConfigFSM_inst._066_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1245__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0881_ INST_config_UART._0383_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0100_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0950_ INST_config_UART.TimeToSendCounter\[7\] INST_config_UART._0401_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0432_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1364_ net1 INST_config_UART._0185_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._431__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1295_ net1 INST_config_UART._0037_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._453_ net1 Inst_bitbang._082_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._384_ net1 Inst_bitbang._021_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1080_ INST_config_UART.CRCReg\[12\] INST_config_UART._0531_ INST_config_UART._0532_
+ INST_config_UART._0529_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0933_ INST_config_UART.TimeToSendCounter\[1\] INST_config_UART.TimeToSendCounter\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0421_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._0864_ INST_config_UART.ComTick INST_config_UART.ComState\[4\] INST_config_UART.PresentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0374_ sky130_fd_sc_hd__and3_1
XINST_config_UART._0795_ INST_config_UART._0243_ INST_config_UART.WriteData\[18\]
+ INST_config_UART._0236_ INST_config_UART._0331_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0066_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1347_ net1 INST_config_UART._0010_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1278_ net1 INST_config_UART._0136_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[30\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1120__A1 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._436_ net1 Inst_bitbang.s_clk_sample\[1\] net111 vssd1 vssd1 vccd1 vccd1
+ Inst_bitbang.s_clk_sample\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._367_ net1 Inst_bitbang._004_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._436__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._298_ Inst_bitbang._147_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._052_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1318__SET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1319__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1260__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 RowSelect[3] sky130_fd_sc_hd__buf_2
XINST_config_UART._1201_ net1 INST_config_UART._0070_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output72_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1063_ INST_config_UART._0517_ INST_config_UART._0519_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0520_ sky130_fd_sc_hd__nand2_2
XINST_config_UART._1132_ INST_config_UART.Command\[2\] INST_config_UART._0221_ INST_config_UART._0563_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0566_ sky130_fd_sc_hd__mux2_1
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[27] sky130_fd_sc_hd__clkbuf_4
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[16] sky130_fd_sc_hd__buf_2
XANTENNA__194__A ConfigFSM_inst.WriteData\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0916_ INST_config_UART._0411_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0107_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0778_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[4\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0321_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0847_ INST_config_UART._0362_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0087_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1348__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._221_ Inst_bitbang.serial_data\[13\] Inst_bitbang.data\[13\] Inst_bitbang._101_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._107_ sky130_fd_sc_hd__mux2_1
XANTENNA__133__S _021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_170_ _066_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[29\] sky130_fd_sc_hd__buf_1
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._419_ net1 Inst_bitbang._056_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._250_ net1 ConfigFSM_inst._002_ net112 vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_INST_config_UART._1291__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._0632_ INST_config_UART._0222_ INST_config_UART._0221_ INST_config_UART._0219_
+ INST_config_UART.ReceivedWord\[3\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0228_
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._181_ ConfigFSM_inst.WriteData\[0\] ConfigFSM_inst.FrameAddressRegister\[0\]
+ ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._087_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0701_ INST_config_UART._0258_ INST_config_UART._0275_ INST_config_UART._0262_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0002_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__189__A ConfigFSM_inst.WriteData\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1046_ INST_config_UART._0491_ INST_config_UART._0495_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0505_ sky130_fd_sc_hd__or2_1
XINST_config_UART._1115_ INST_config_UART._0556_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0161_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1182__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._204_ Inst_bitbang.serial_data\[5\] Inst_bitbang.data\[5\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._451__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_153_ net19 Inst_bitbang.data\[24\] _043_ vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__mux2_1
X_222_ ConfigFSM_inst.FrameAddressRegister\[9\] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
X_084_ _007_ INST_config_UART.WriteData\[2\] _001_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._121__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._233_ ConfigFSM_inst.WriteData\[26\] ConfigFSM_inst.FrameAddressRegister\[26\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._114_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0615_ INST_config_UART.ByteWriteStrobe vssd1 vssd1 vccd1 vccd1
+ INST_config_UART._0214_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_ConfigFSM_inst._231__A0 ConfigFSM_inst.WriteData\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._164_ ConfigFSM_inst._058_ ConfigFSM_inst._074_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._075_ sky130_fd_sc_hd__nor2_1
XANTENNA_ConfigFSM_inst._260__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1187__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1029_ INST_config_UART.CRCReg\[4\] INST_config_UART._0488_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0490_ sky130_fd_sc_hd__nand2_1
XANTENNA_INST_config_UART._1363__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._283__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_205_ ConfigFSM_inst.WriteData\[24\] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_136_ Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_ConfigFSM_inst._245__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._373__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._216_ ConfigFSM_inst.WriteData\[17\] ConfigFSM_inst.FrameAddressRegister\[17\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._105_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._204__A0 ConfigFSM_inst.WriteData\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XConfigFSM_inst._147_ ConfigFSM_inst._063_ ConfigFSM_inst._064_ ConfigFSM_inst._065_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._004_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1202__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1352__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1214__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1285__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0880_ INST_config_UART.ID_Reg\[15\] INST_config_UART.ReceivedWord\[7\]
+ INST_config_UART._0375_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0383_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._383__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_119_ _031_ INST_config_UART.WriteData\[13\] _023_ vssd1 vssd1 vccd1 vccd1 _032_
+ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1363_ net1 INST_config_UART._0184_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1294_ net1 INST_config_UART._0036_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1225__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xload_slew111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__197__A ConfigFSM_inst.WriteData\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._452_ net1 Inst_bitbang._081_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._383_ net1 Inst_bitbang._020_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._0656__A INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1248__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0863_ INST_config_UART.RxLocal INST_config_UART._0372_ INST_config_UART._0373_
+ INST_config_UART._0223_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0092_ sky130_fd_sc_hd__o22a_1
XINST_config_UART._0932_ INST_config_UART.TimeToSendCounter\[1\] INST_config_UART.TimeToSendCounter\[0\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0420_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0794_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0318_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0331_ sky130_fd_sc_hd__and3_1
XANTENNA_ConfigFSM_inst._260__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1346_ net1 INST_config_UART._0009_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[6\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1277_ net1 INST_config_UART._0135_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._185__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._435_ net1 Inst_bitbang.s_clk_sample\[0\] net111 vssd1 vssd1 vccd1 vccd1
+ Inst_bitbang.s_clk_sample\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._366_ net1 Inst_bitbang._003_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._297_ Inst_bitbang.serial_data\[16\] Inst_bitbang.serial_data\[17\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._147_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._405__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0870__A1 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._421__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._124__A ConfigFSM_inst.WriteData\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[8] sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._1131_ INST_config_UART._0565_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0168_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._326__S Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1200_ net1 INST_config_UART._0069_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1062_ INST_config_UART._0501_ INST_config_UART._0511_ INST_config_UART._0512_
+ INST_config_UART._0518_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0519_ sky130_fd_sc_hd__o211a_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[28] sky130_fd_sc_hd__clkbuf_4
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[17] sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._0915_ INST_config_UART.HexData\[1\] INST_config_UART._0393_ INST_config_UART._0014_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0411_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0846_ INST_config_UART.ID_Reg\[21\] INST_config_UART.ReceivedWord\[5\]
+ INST_config_UART._0356_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0362_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0777_ INST_config_UART.WriteData\[3\] INST_config_UART._0240_ INST_config_UART._0320_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._220_ Inst_bitbang._106_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._015_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1329_ net1 INST_config_UART._0164_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._444__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._349_ Inst_bitbang._174_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._076_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._418_ net1 Inst_bitbang._055_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._0700_ INST_config_UART.ComCount\[10\] INST_config_UART._0257_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0631_ INST_config_UART._0224_ INST_config_UART._0225_ INST_config_UART._0226_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0227_ sky130_fd_sc_hd__or3b_2
XConfigFSM_inst._180_ ConfigFSM_inst._085_ ConfigFSM_inst._086_ ConfigFSM_inst._057_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._009_ sky130_fd_sc_hd__o21a_1
XANTENNA_Inst_bitbang._398__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1114_ INST_config_UART.ID_Reg\[2\] INST_config_UART._0221_ INST_config_UART._0553_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0556_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1045_ INST_config_UART.CRCReg\[5\] INST_config_UART._0494_ INST_config_UART._0503_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0504_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINST_config_UART._0829_ INST_config_UART.RxLocal INST_config_UART._0349_ INST_config_UART._0351_
+ INST_config_UART.ReceivedWord\[5\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0080_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._203_ Inst_bitbang._097_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._007_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._1309__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_083_ net25 Inst_bitbang.data\[2\] _000_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1239__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_221_ ConfigFSM_inst.FrameAddressRegister\[8\] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_152_ _054_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[23\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._420__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._232_ ConfigFSM_inst._113_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._034_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._163_ ConfigFSM_inst._042_ ConfigFSM_inst._073_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._074_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0614_ INST_config_UART.PresentState\[0\] INST_config_UART._0199_
+ INST_config_UART._0211_ INST_config_UART.PresentState\[5\] INST_config_UART._0213_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1028_ INST_config_UART.CRCReg\[4\] INST_config_UART._0488_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0489_ sky130_fd_sc_hd__or2_1
XANTENNA_ConfigFSM_inst._193__S ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1332__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1281__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_204_ ConfigFSM_inst.WriteData\[23\] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_ConfigFSM_inst._132__A ConfigFSM_inst.WriteData\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_135_ _042_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[18\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_ConfigFSM_inst._285__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XConfigFSM_inst._215_ ConfigFSM_inst._104_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._026_
+ sky130_fd_sc_hd__clkbuf_1
XConfigFSM_inst._146_ ConfigFSM_inst.state\[1\] ConfigFSM_inst._057_ ConfigFSM_inst._060_
+ ConfigFSM_inst._044_ ConfigFSM_inst.state\[2\] vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._065_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1254__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._250__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_118_ net7 Inst_bitbang.data\[13\] _021_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1293_ net1 INST_config_UART._0035_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xload_slew112 net36 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1362_ net1 INST_config_UART._0183_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComState\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._451_ net1 Inst_bitbang._080_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._382_ net1 Inst_bitbang._019_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_ConfigFSM_inst._189__A0 ConfigFSM_inst.WriteData\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XConfigFSM_inst._129_ ConfigFSM_inst.WriteData\[2\] ConfigFSM_inst.WriteData\[6\]
+ ConfigFSM_inst.WriteData\[5\] ConfigFSM_inst.WriteData\[4\] vssd1 vssd1 vccd1 vccd1
+ ConfigFSM_inst._050_ sky130_fd_sc_hd__or4bb_1
XANTENNA_ConfigFSM_inst._273__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1211__SET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0862_ INST_config_UART._0250_ INST_config_UART._0347_ INST_config_UART.ComState\[3\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0373_ sky130_fd_sc_hd__and3b_1
XINST_config_UART._0931_ INST_config_UART.TimeToSendCounter\[0\] INST_config_UART._0419_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0793_ INST_config_UART._0243_ INST_config_UART.WriteData\[17\]
+ INST_config_UART._0236_ INST_config_UART._0330_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0065_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_1 ConfigFSM_inst.WriteData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1345_ net1 INST_config_UART._0008_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1342__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1276_ net1 INST_config_UART._0134_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._434_ net1 net37 net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.s_clk_sample\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._365_ net1 Inst_bitbang.local_strobe net111 vssd1 vssd1 vccd1 vccd1
+ Inst_bitbang.old_local_strobe sky130_fd_sc_hd__dfrtp_1
XANTENNA_Inst_bitbang._373__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._296_ Inst_bitbang._146_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._051_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._445__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._124__B ConfigFSM_inst.WriteData\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1215__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[9] sky130_fd_sc_hd__buf_2
XINST_config_UART._1061_ INST_config_UART._0502_ INST_config_UART._0504_ INST_config_UART._0513_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0518_ sky130_fd_sc_hd__or3_1
XINST_config_UART._1130_ INST_config_UART.Command\[1\] INST_config_UART._0222_ INST_config_UART._0563_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0565_ sky130_fd_sc_hd__mux2_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[29] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[18] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1365__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._0914_ INST_config_UART._0410_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0106_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0776_ INST_config_UART._0312_ INST_config_UART.HexData\[3\] INST_config_UART._0319_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0845_ INST_config_UART._0361_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0086_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._396__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1328_ net1 INST_config_UART._0163_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_bitbang._252__S Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1259_ net1 INST_config_UART._0120_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1238__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._348_ Inst_bitbang.serial_control\[8\] Inst_bitbang.serial_control\[9\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._174_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._417_ net1 Inst_bitbang._054_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._279_ Inst_bitbang._137_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._043_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0630_ INST_config_UART._0222_ INST_config_UART._0223_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0226_ sky130_fd_sc_hd__nand2_1
XANTENNA_Inst_bitbang._367__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1044_ INST_config_UART.CRCReg\[5\] INST_config_UART._0494_ INST_config_UART._0488_
+ INST_config_UART.CRCReg\[4\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0503_ sky130_fd_sc_hd__o211a_1
XINST_config_UART._1113_ INST_config_UART._0555_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0160_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0759_ INST_config_UART.ReceivedWord\[7\] INST_config_UART.RxLocal
+ INST_config_UART._0307_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0308_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0828_ INST_config_UART._0251_ INST_config_UART._0350_ INST_config_UART.ComState\[10\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0351_ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._202_ Inst_bitbang.serial_data\[4\] Inst_bitbang.data\[4\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._097_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1191__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._411__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_220_ ConfigFSM_inst.FrameAddressRegister\[7\] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_082_ _006_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[1\] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1279__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_151_ _053_ INST_config_UART.WriteData\[23\] _045_ vssd1 vssd1 vccd1 vccd1 _054_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._121__C ConfigFSM_inst.WriteData\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1208__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._0613_ INST_config_UART.PresentState\[6\] INST_config_UART._0212_
+ INST_config_UART.TimeToSend vssd1 vssd1 vccd1 vccd1 INST_config_UART._0213_ sky130_fd_sc_hd__o21a_1
XConfigFSM_inst._231_ ConfigFSM_inst.WriteData\[25\] ConfigFSM_inst.FrameAddressRegister\[25\]
+ ConfigFSM_inst._107_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._113_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._162_ ConfigFSM_inst.state\[2\] ConfigFSM_inst.state\[1\] ConfigFSM_inst._043_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._073_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1027_ INST_config_UART.ReceivedWord\[4\] INST_config_UART.HighReg\[0\]
+ INST_config_UART.Command\[7\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0488_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._434__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1301__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_203_ ConfigFSM_inst.WriteData\[22\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_134_ _041_ INST_config_UART.WriteData\[18\] _023_ vssd1 vssd1 vccd1 vccd1 _042_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._132__B ConfigFSM_inst.WriteData\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._254__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XConfigFSM_inst._214_ ConfigFSM_inst.WriteData\[16\] ConfigFSM_inst.FrameAddressRegister\[16\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._104_ sky130_fd_sc_hd__mux2_1
XConfigFSM_inst._145_ ConfigFSM_inst._043_ ConfigFSM_inst.state\[0\] ConfigFSM_inst._057_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._064_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._382__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1150__A1 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_ConfigFSM_inst._127__B ConfigFSM_inst.WriteData\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_117_ _030_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[12\] sky130_fd_sc_hd__buf_2
XANTENNA_INST_config_UART._1294__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1223__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1292_ net1 INST_config_UART._0034_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[12\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1361_ net1 INST_config_UART._0182_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_load_slew112_A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1132__A1 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1271__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._381_ net1 Inst_bitbang._018_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._450_ net1 Inst_bitbang._079_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_control\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XConfigFSM_inst._128_ ConfigFSM_inst._045_ ConfigFSM_inst._046_ ConfigFSM_inst._047_
+ ConfigFSM_inst._048_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._049_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1114__A1 INST_config_UART._0221_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1294__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0930_ INST_config_UART._0418_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0419_
+ sky130_fd_sc_hd__buf_2
XINST_config_UART._0861_ INST_config_UART._0371_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0372_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._0792_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0316_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0330_ sky130_fd_sc_hd__and3_1
XINST_config_UART._1344_ net1 INST_config_UART._0007_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 ConfigFSM_inst.WriteData\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINST_config_UART._1275_ net1 INST_config_UART._0133_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[27\] sky130_fd_sc_hd__dfrtp_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._433_ net1 Inst_bitbang.s_data_sample\[2\] net111 vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang.s_data_sample\[3\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._364_ net1 Inst_bitbang._000_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.local_strobe
+ sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._295_ Inst_bitbang.serial_data\[15\] Inst_bitbang.serial_data\[16\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._414__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 ConfigWriteStrobe sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[29] sky130_fd_sc_hd__clkbuf_4
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[19] sky130_fd_sc_hd__buf_2
XINST_config_UART._1060_ INST_config_UART._0484_ INST_config_UART._0478_ INST_config_UART._0482_
+ INST_config_UART._0516_ INST_config_UART._0481_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0517_
+ sky130_fd_sc_hd__a311o_2
XFILLER_0_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[19] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[2] sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._0913_ INST_config_UART.HexData\[0\] INST_config_UART._0387_ INST_config_UART._0014_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0410_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1353__SET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0775_ INST_config_UART._0247_ INST_config_UART.Data_Reg\[3\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0319_ sky130_fd_sc_hd__or2_1
XINST_config_UART._0844_ INST_config_UART.ID_Reg\[20\] INST_config_UART.ReceivedWord\[4\]
+ INST_config_UART._0356_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0361_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._263__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1327_ net1 INST_config_UART._0162_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1189_ net1 INST_config_UART._0058_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1258_ net1 INST_config_UART._0119_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1326__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._278_ Inst_bitbang.serial_data\[7\] Inst_bitbang.serial_data\[8\] Inst_bitbang._128_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._137_ sky130_fd_sc_hd__mux2_1
XInst_bitbang._347_ Inst_bitbang._173_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._075_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._416_ net1 Inst_bitbang._053_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1332__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._286__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._243__A0 ConfigFSM_inst.WriteData\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._279__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1043_ INST_config_UART._0500_ INST_config_UART._0501_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0502_ sky130_fd_sc_hd__nand2_1
XINST_config_UART._1112_ INST_config_UART.ID_Reg\[1\] INST_config_UART._0222_ INST_config_UART._0553_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0555_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._363__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0827_ INST_config_UART._0347_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0350_
+ sky130_fd_sc_hd__clkbuf_4
XINST_config_UART._0758_ INST_config_UART.ComState\[0\] INST_config_UART.ComState\[7\]
+ INST_config_UART._0245_ INST_config_UART._0306_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0307_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0689_ INST_config_UART._0254_ INST_config_UART._0268_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0269_ sky130_fd_sc_hd__nand2_1
XInst_bitbang._201_ Inst_bitbang._096_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._006_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_INST_config_UART._1205__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1355__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._225__A0 ConfigFSM_inst.WriteData\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_150_ net18 Inst_bitbang.data\[23\] _043_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__mux2_1
X_081_ _005_ INST_config_UART.WriteData\[1\] _001_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1248__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XConfigFSM_inst._230_ ConfigFSM_inst._112_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._033_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._386__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0612_ net39 INST_config_UART._0192_ INST_config_UART.PresentState\[2\]
+ INST_config_UART.PresentState\[4\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0212_
+ sky130_fd_sc_hd__or4_1
XConfigFSM_inst._161_ ConfigFSM_inst._072_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._000_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_ConfigFSM_inst._216__A0 ConfigFSM_inst.WriteData\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1228__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1026_ INST_config_UART._0484_ INST_config_UART._0478_ INST_config_UART._0482_
+ INST_config_UART._0481_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0487_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._258__S Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__171__S Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1341__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__200__A ConfigFSM_inst.WriteData\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_202_ ConfigFSM_inst.WriteData\[21\] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_133_ net12 Inst_bitbang.data\[18\] _021_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__mux2_1
XANTENNA_ConfigFSM_inst._132__C ConfigFSM_inst.WriteData\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XConfigFSM_inst._213_ ConfigFSM_inst._103_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._025_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_bitbang._401__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._144_ ConfigFSM_inst._049_ ConfigFSM_inst._054_ vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XINST_config_UART._1009_ INST_config_UART._0246_ INST_config_UART._0393_ INST_config_UART._0472_
+ INST_config_UART.CRCReg\[1\] vssd1 vssd1 vccd1 vccd1 INST_config_UART._0473_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._439__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_ConfigFSM_inst._127__C ConfigFSM_inst.WriteData\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._424__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_116_ _029_ INST_config_UART.WriteData\[12\] _023_ vssd1 vssd1 vccd1 vccd1 _030_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINST_config_UART._1360_ net1 INST_config_UART._0181_ vssd1 vssd1 vccd1 vccd1 INST_config_UART.Data_Reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_INST_config_UART._1263__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1291_ net1 INST_config_UART._0033_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[11\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._380_ net1 Inst_bitbang._017_ net36 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._127_ ConfigFSM_inst.WriteData\[29\] ConfigFSM_inst.WriteData\[28\]
+ ConfigFSM_inst.WriteData\[31\] ConfigFSM_inst.WriteData\[30\] vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._048_ sky130_fd_sc_hd__and4_1
XANTENNA_Inst_bitbang._447__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._0791_ INST_config_UART._0243_ INST_config_UART.WriteData\[16\]
+ INST_config_UART._0236_ INST_config_UART._0329_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0064_
+ sky130_fd_sc_hd__a31o_1
XINST_config_UART._0860_ INST_config_UART.ComState\[0\] INST_config_UART.ComTick INST_config_UART.ComState\[3\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0371_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._210__A Inst_bitbang._087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINST_config_UART._1343_ net1 INST_config_UART._0006_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1274_ net1 INST_config_UART._0132_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_bitbang._432_ net1 Inst_bitbang.s_data_sample\[1\] net111 vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang.s_data_sample\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1185__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0989_ INST_config_UART._0216_ INST_config_UART.GetWordState\[0\]
+ INST_config_UART._0324_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0457_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._294_ Inst_bitbang._145_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._050_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._363_ net1 Inst_bitbang._002_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.active
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_INST_config_UART._0855__A1 INST_config_UART.RxLocal vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0855__B2 INST_config_UART._0218_ vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[2] sky130_fd_sc_hd__clkbuf_4
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[1] sky130_fd_sc_hd__buf_2
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[0] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_INST_config_UART._1261__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[30] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[0] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[1] sky130_fd_sc_hd__buf_2
XINST_config_UART._0912_ INST_config_UART._0409_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0105_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_INST_config_UART._0846__A1 INST_config_UART.ReceivedWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0843_ INST_config_UART._0360_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0085_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._0774_ INST_config_UART.WriteData\[2\] INST_config_UART._0240_ INST_config_UART._0318_
+ INST_config_UART._0017_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0058_ sky130_fd_sc_hd__a22o_1
XINST_config_UART._1326_ net1 INST_config_UART._0161_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[2\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1257_ net1 INST_config_UART._0118_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINST_config_UART._1188_ net1 INST_config_UART._0057_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_INST_config_UART._1366__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__174__S Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_bitbang._415_ net1 Inst_bitbang._052_ net112 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.serial_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__203__A ConfigFSM_inst.WriteData\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_bitbang._277_ Inst_bitbang._136_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._042_
+ sky130_fd_sc_hd__clkbuf_1
XInst_bitbang._346_ Inst_bitbang.serial_control\[7\] Inst_bitbang.serial_control\[8\]
+ Inst_bitbang._164_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._173_ sky130_fd_sc_hd__mux2_1
XANTENNA_INST_config_UART._1284__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1111_ INST_config_UART._0554_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0159_
+ sky130_fd_sc_hd__clkbuf_1
XINST_config_UART._1042_ INST_config_UART.CRCReg\[6\] INST_config_UART._0499_ vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0501_ sky130_fd_sc_hd__nand2_1
XANTENNA_ConfigFSM_inst._248__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._376__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0826_ INST_config_UART._0348_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0349_
+ sky130_fd_sc_hd__inv_2
XINST_config_UART._0757_ INST_config_UART._0197_ INST_config_UART.ComState\[7\] vssd1
+ vssd1 vccd1 vccd1 INST_config_UART._0306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0688_ INST_config_UART.ComCount\[4\] INST_config_UART._0253_ INST_config_UART.ComCount\[5\]
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0268_ sky130_fd_sc_hd__o21ai_1
XINST_config_UART._1309_ net1 INST_config_UART._0144_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.CRCReg\[6\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._200_ Inst_bitbang.serial_data\[3\] Inst_bitbang.data\[3\] Inst_bitbang._088_
+ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__169__S net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_080_ net14 Inst_bitbang.data\[1\] _000_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._329_ Inst_bitbang._163_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._164_
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_INST_config_UART._1288__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._253__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_INST_config_UART._1217__RESET_B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._0611_ INST_config_UART._0200_ INST_config_UART._0202_ INST_config_UART._0210_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0211_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._160_ ConfigFSM_inst.state\[1\] ConfigFSM_inst._057_ ConfigFSM_inst._060_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._072_ sky130_fd_sc_hd__and3_1
XINST_config_UART._1025_ INST_config_UART.CRCReg\[3\] INST_config_UART._0469_ INST_config_UART._0466_
+ INST_config_UART._0486_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0809_ INST_config_UART._0242_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0339_
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1322__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._143__B1 ConfigFSM_inst._062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._276__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._303__A Inst_bitbang._127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1310__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._0911__S net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_201_ ConfigFSM_inst.WriteData\[20\] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_132_ _040_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst.WriteData\[17\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_ConfigFSM_inst._132__D ConfigFSM_inst.WriteData\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._143_ ConfigFSM_inst._058_ ConfigFSM_inst._060_ ConfigFSM_inst._062_
+ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._003_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._212_ ConfigFSM_inst.WriteData\[15\] ConfigFSM_inst.FrameAddressRegister\[15\]
+ ConfigFSM_inst._096_ vssd1 vssd1 vccd1 vccd1 ConfigFSM_inst._103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_ConfigFSM_inst._263__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1345__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1008_ INST_config_UART._0391_ INST_config_UART._0246_ vssd1 vssd1
+ vccd1 vccd1 INST_config_UART._0472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_bitbang._391__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_bitbang._376__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__211__A ConfigFSM_inst.WriteData\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_bitbang._408__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1218__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_ConfigFSM_inst._127__D ConfigFSM_inst.WriteData\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_115_ net6 Inst_bitbang.data\[12\] _021_ vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._1290_ net1 INST_config_UART._0032_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.blink\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_INST_config_UART._1368__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_INST_config_UART._1232__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._399__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XConfigFSM_inst._126_ ConfigFSM_inst.WriteData\[24\] ConfigFSM_inst.WriteData\[26\]
+ ConfigFSM_inst.WriteData\[27\] ConfigFSM_inst.WriteData\[25\] vssd1 vssd1 vccd1
+ vccd1 ConfigFSM_inst._047_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__177__S Inst_bitbang.active vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__206__A ConfigFSM_inst.WriteData\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_INST_config_UART._1190__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0790_ INST_config_UART._0214_ INST_config_UART.GetWordState\[2\]
+ INST_config_UART._0314_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0329_ sky130_fd_sc_hd__and3_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1273_ net1 INST_config_UART._0131_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.WriteData\[25\] sky130_fd_sc_hd__dfrtp_1
XINST_config_UART._1342_ net1 INST_config_UART._0005_ net112 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ComCount\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ConfigFSM_inst._126__D_N ConfigFSM_inst.WriteData\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._0988_ INST_config_UART._0242_ INST_config_UART.WriteData\[28\]
+ INST_config_UART._0234_ INST_config_UART._0456_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0134_
+ sky130_fd_sc_hd__a31o_1
XInst_bitbang._431_ net1 Inst_bitbang.s_data_sample\[0\] net111 vssd1 vssd1 vccd1
+ vccd1 Inst_bitbang.s_data_sample\[1\] sky130_fd_sc_hd__dfrtp_1
XInst_bitbang._362_ net1 Inst_bitbang._001_ net111 vssd1 vssd1 vccd1 vccd1 Inst_bitbang.strobe
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_bitbang._293_ Inst_bitbang.serial_data\[14\] Inst_bitbang.serial_data\[15\]
+ Inst_bitbang._139_ vssd1 vssd1 vccd1 vccd1 Inst_bitbang._145_ sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_bitbang._414__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[20] sky130_fd_sc_hd__clkbuf_4
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[10] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ConfigWriteData[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[31] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[21] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_bitbang._423__RESET_B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 FrameAddressRegister[10] sky130_fd_sc_hd__buf_2
XINST_config_UART._0842_ INST_config_UART.ID_Reg\[19\] INST_config_UART._0218_ INST_config_UART._0356_
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0360_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0911_ INST_config_UART.TimeToSend INST_config_UART._0408_ net111
+ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0409_ sky130_fd_sc_hd__mux2_1
XINST_config_UART._0773_ INST_config_UART._0312_ INST_config_UART.HexData\[2\] INST_config_UART._0317_
+ INST_config_UART._0241_ vssd1 vssd1 vccd1 vccd1 INST_config_UART._0318_ sky130_fd_sc_hd__o211a_2
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINST_config_UART._1325_ net1 INST_config_UART._0160_ net36 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.ID_Reg\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_bitbang._437__CLK net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINST_config_UART._1256_ net1 INST_config_UART._0117_ net111 vssd1 vssd1 vccd1 vccd1
+ INST_config_UART.TimeToSendCounter\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

