* NGSPICE file created from RAM_IO.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt RAM_IO Config_accessC_bit0 Config_accessC_bit1 Config_accessC_bit2 Config_accessC_bit3
+ E1END[0] E1END[1] E1END[2] E1END[3] E2END[0] E2END[1] E2END[2] E2END[3] E2END[4]
+ E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5]
+ E2MID[6] E2MID[7] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4]
+ E6END[5] E6END[6] E6END[7] E6END[8] E6END[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12]
+ EE4END[13] EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5]
+ EE4END[6] EE4END[7] EE4END[8] EE4END[9] FAB2RAM_A0_O0 FAB2RAM_A0_O1 FAB2RAM_A0_O2
+ FAB2RAM_A0_O3 FAB2RAM_A1_O0 FAB2RAM_A1_O1 FAB2RAM_A1_O2 FAB2RAM_A1_O3 FAB2RAM_C_O0
+ FAB2RAM_C_O1 FAB2RAM_C_O2 FAB2RAM_C_O3 FAB2RAM_D0_O0 FAB2RAM_D0_O1 FAB2RAM_D0_O2
+ FAB2RAM_D0_O3 FAB2RAM_D1_O0 FAB2RAM_D1_O1 FAB2RAM_D1_O2 FAB2RAM_D1_O3 FAB2RAM_D2_O0
+ FAB2RAM_D2_O1 FAB2RAM_D2_O2 FAB2RAM_D2_O3 FAB2RAM_D3_O0 FAB2RAM_D3_O1 FAB2RAM_D3_O2
+ FAB2RAM_D3_O3 FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] RAM2FAB_D0_I0 RAM2FAB_D0_I1 RAM2FAB_D0_I2
+ RAM2FAB_D0_I3 RAM2FAB_D1_I0 RAM2FAB_D1_I1 RAM2FAB_D1_I2 RAM2FAB_D1_I3 RAM2FAB_D2_I0
+ RAM2FAB_D2_I1 RAM2FAB_D2_I2 RAM2FAB_D2_I3 RAM2FAB_D3_I0 RAM2FAB_D3_I1 RAM2FAB_D3_I2
+ RAM2FAB_D3_I3 S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0]
+ S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1]
+ S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2]
+ S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12]
+ S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6]
+ S4BEG[7] S4BEG[8] S4BEG[9] S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14]
+ S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8]
+ S4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2] W1BEG[3] W2BEG[0]
+ W2BEG[1] W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1]
+ W2BEGb[2] W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W6BEG[0] W6BEG[10] W6BEG[11]
+ W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
XInst_FAB2RAM_D2_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0 net1 net27 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\] Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N1BEG0 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S4BEG2 sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame6_bit3 net74 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_12._0_ strobe_inbuf_12.X VGND VGND VPWR VPWR strobe_outbuf_12.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_7._0_ data_inbuf_7.X VGND VGND VPWR VPWR data_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3 net104 net130 net156 net182
+ Inst_RAM_IO_ConfigMem.ConfigBits\[278\] Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame2_bit18 net58 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit29 net70 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput264 net264 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput253 net253 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput286 net286 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput275 net275 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput242 net242 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput231 net231 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit6 net77 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput220 net220 VGND VGND VPWR VPWR FAB2RAM_D3_O3 sky130_fd_sc_hd__buf_2
Xoutput297 net297 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
X_062_ Inst_RAM_IO_switch_matrix.N2BEG6 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
X_131_ Inst_RAM_IO_switch_matrix.W2BEG3 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit17 net57 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit28 net69 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_045_ strobe_outbuf_13.X VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_1
X_114_ S4BEG_outbuf_6.X VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0 net17 net9 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
+ net399 Inst_RAM_IO_ConfigMem.ConfigBits\[256\] Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_2
XFILLER_0_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame0_bit9 net80 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame0_bit27 net68 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit16 net56 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit1 net60 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_028_ data_outbuf_28.X VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 Inst_RAM_IO_switch_matrix.S2BEG1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_7._0_ strobe_inbuf_7.X VGND VGND VPWR VPWR strobe_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame10_bit27 net68 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_1._0_ net60 VGND VGND VPWR VPWR data_inbuf_1.X sky130_fd_sc_hd__clkbuf_1
Xinput175 S4END[11] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xinput164 S2END[7] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xinput153 S1END[0] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_2
Xinput186 S4END[7] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xinput142 RAM2FAB_D1_I1 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_1
Xinput131 N4END[4] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xinput120 N2MID[7] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[136\] Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG4 sky130_fd_sc_hd__mux4_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux._2_ UserCLK net139 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1 net2 net28 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[50\] Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N1BEG1 sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[116\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit4 net75 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4 net101 net121 net153 net173
+ Inst_RAM_IO_ConfigMem.ConfigBits\[280\] Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG4 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit19 net59 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__o21ai_1
XN4END_inbuf_7._0_ net123 VGND VGND VPWR VPWR N4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput265 net265 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput276 net276 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput254 net254 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput298 net298 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
Xoutput221 net221 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput243 net243 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit7 net78 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput210 net210 VGND VGND VPWR VPWR FAB2RAM_D1_O1 sky130_fd_sc_hd__buf_2
XFILLER_0_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_130_ Inst_RAM_IO_switch_matrix.W2BEG2 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_1
X_061_ Inst_RAM_IO_switch_matrix.N2BEG5 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit18 net58 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit29 net70 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_113_ S4BEG_outbuf_5.X VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_1
X_044_ strobe_outbuf_12.X VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1 net18 net10 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
+ net400 Inst_RAM_IO_ConfigMem.ConfigBits\[258\] Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame0_bit17 net57 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit2 net71 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit28 net69 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ net143 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_10._0_ data_inbuf_10.X VGND VGND VPWR VPWR data_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 Inst_RAM_IO_switch_matrix.S2BEG3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_027_ data_outbuf_27.X VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame10_bit28 net69 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__o21ai_1
Xinput110 N2END[5] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput154 S1END[1] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xinput165 S2MID[0] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
Xinput176 S4END[12] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput187 S4END[8] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput143 RAM2FAB_D1_I2 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xinput132 N4END[5] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput121 N4END[0] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[138\] Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG5 sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2 net3 net29 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[52\] Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N1BEG2 sky130_fd_sc_hd__mux4_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux._1_ UserCLK net138 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0 net1 net21 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
+ net403 Inst_RAM_IO_ConfigMem.ConfigBits\[264\] Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0 net2 net37
+ net28 Inst_RAM_IO_switch_matrix.J_NS4_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[112\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_ConfigMem.Inst_frame6_bit5 net76 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5 net102 net128 net154 net180
+ Inst_RAM_IO_ConfigMem.ConfigBits\[282\] Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG5 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput200 net200 VGND VGND VPWR VPWR FAB2RAM_A1_O3 sky130_fd_sc_hd__clkbuf_4
Xoutput255 net255 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput299 net299 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput266 net266 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput244 net244 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__buf_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput222 net222 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame3_bit8 net79 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput211 net211 VGND VGND VPWR VPWR FAB2RAM_D1_O2 sky130_fd_sc_hd__clkbuf_4
X_060_ Inst_RAM_IO_switch_matrix.N2BEG4 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit19 net59 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_30._0_ net72 VGND VGND VPWR VPWR data_inbuf_30.X sky130_fd_sc_hd__clkbuf_1
X_043_ strobe_outbuf_11.X VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
X_112_ S4BEG_outbuf_4.X VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2 net19 net11 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
+ net401 Inst_RAM_IO_ConfigMem.ConfigBits\[260\] Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_21._0_ net62 VGND VGND VPWR VPWR data_inbuf_21.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame0_bit18 net58 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_0._0_ net81 VGND VGND VPWR VPWR strobe_inbuf_0.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_12._0_ net52 VGND VGND VPWR VPWR data_inbuf_12.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit3 net74 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit29 net70 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_026_ data_outbuf_26.X VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
XANTENNA_7 Inst_RAM_IO_switch_matrix.S2BEG3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame10_bit29 net70 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_8_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput144 RAM2FAB_D1_I3 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
Xinput133 N4END[6] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput122 N4END[10] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
Xinput100 FrameStrobe[9] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_8
Xinput111 N2END[6] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput166 S2MID[1] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
Xinput155 S1END[2] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xinput177 S4END[13] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput188 S4END[9] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_15._0_ strobe_inbuf_15.X VGND VGND VPWR VPWR strobe_outbuf_15.X sky130_fd_sc_hd__clkbuf_1
X_009_ data_outbuf_9.X VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[140\] Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG6 sky130_fd_sc_hd__mux4_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux._0_ UserCLK net137 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3 net4 net30 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[54\] Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N1BEG3 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1 net2 net24 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
+ net404 Inst_RAM_IO_ConfigMem.ConfigBits\[266\] Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG9 Inst_RAM_IO_switch_matrix.J_NS4_BEG13 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
+ Inst_RAM_IO_ConfigMem.ConfigBits\[111\] Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit6 net77 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_A0_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6 net103 net129 net155 net181
+ Inst_RAM_IO_ConfigMem.ConfigBits\[284\] Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput234 net234 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput223 net223 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput212 net212 VGND VGND VPWR VPWR FAB2RAM_D1_O3 sky130_fd_sc_hd__buf_2
Xoutput201 net201 VGND VGND VPWR VPWR FAB2RAM_C_O0 sky130_fd_sc_hd__buf_2
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput256 net256 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput289 net289 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput278 net278 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput245 net245 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit9 net80 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_inbuf_12._0_ net84 VGND VGND VPWR VPWR strobe_inbuf_12.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0 net43 net36 net27 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
+ Inst_RAM_IO_ConfigMem.ConfigBits\[224\] Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ net151 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_042_ strobe_outbuf_10.X VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_1
X_111_ S4BEG_outbuf_3.X VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3 net20 net12 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
+ net402 Inst_RAM_IO_ConfigMem.ConfigBits\[262\] Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS4_BEG5
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[180\] Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG10 sky130_fd_sc_hd__mux4_1
XFILLER_0_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit19 net59 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit4 net75 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_025_ data_outbuf_25.X VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_4._0_ net75 VGND VGND VPWR VPWR data_inbuf_4.X sky130_fd_sc_hd__clkbuf_1
XANTENNA_8 Inst_RAM_IO_switch_matrix.S2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_73_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput167 S2MID[2] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xinput156 S1END[3] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xinput178 S4END[14] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xinput145 RAM2FAB_D2_I0 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xinput123 N4END[11] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput134 N4END[7] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput112 N2END[7] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput101 N1END[0] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_008_ data_outbuf_8.X VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[142\] Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG7 sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__o21ai_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2 net3 net25 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
+ net405 Inst_RAM_IO_ConfigMem.ConfigBits\[268\] Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame6_bit7 net78 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ net137 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7 net104 net130 net156 net182
+ Inst_RAM_IO_ConfigMem.ConfigBits\[286\] Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG7 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4BEG_outbuf_2._0_ N4BEG_outbuf_2.A VGND VGND VPWR VPWR N4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput268 net268 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput257 net257 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput235 net235 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
Xoutput224 net224 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput246 net246 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput202 net202 VGND VGND VPWR VPWR FAB2RAM_C_O1 sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR FAB2RAM_D2_O0 sky130_fd_sc_hd__buf_2
Xoutput279 net279 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1 net44 net37 net28 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
+ Inst_RAM_IO_ConfigMem.ConfigBits\[226\] Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_36_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_31._0_ data_inbuf_31.X VGND VGND VPWR VPWR data_outbuf_31.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396/HI net396 sky130_fd_sc_hd__conb_1
XFILLER_0_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_22._0_ data_inbuf_22.X VGND VGND VPWR VPWR data_outbuf_22.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ S4BEG_outbuf_2.X VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_1
X_041_ strobe_outbuf_9.X VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_13._0_ data_inbuf_13.X VGND VGND VPWR VPWR data_outbuf_13.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_2._0_ S4BEG_outbuf_2.A VGND VGND VPWR VPWR S4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS4_BEG4
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[182\] Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG11 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame9_bit5 net76 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__o21ai_2
XS4END_inbuf_0._0_ net183 VGND VGND VPWR VPWR S4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_1
X_024_ data_outbuf_24.X VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 Inst_RAM_IO_switch_matrix.S2BEGb3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput168 S2MID[3] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
Xinput157 S2END[0] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xinput179 S4END[15] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
Xinput135 N4END[8] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput124 N4END[12] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
Xinput113 N2MID[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
Xinput102 N1END[1] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_2
Xinput146 RAM2FAB_D2_I1 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__o21ai_1
X_007_ data_outbuf_7.X VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3 net4 net26 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
+ net409 Inst_RAM_IO_ConfigMem.ConfigBits\[270\] Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_4_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__o21ai_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit8 net79 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8 net101 net121 net153 net173
+ Inst_RAM_IO_ConfigMem.ConfigBits\[288\] Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG8 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S4BEG1 sky130_fd_sc_hd__o21ai_4
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput258 net258 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput269 net269 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput236 net236 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput225 net225 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput203 net203 VGND VGND VPWR VPWR FAB2RAM_C_O2 sky130_fd_sc_hd__clkbuf_4
Xoutput214 net214 VGND VGND VPWR VPWR FAB2RAM_D2_O1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0 net20 net12 net31 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_ConfigMem.ConfigBits\[92\] Inst_RAM_IO_ConfigMem.ConfigBits\[93\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG0 sky130_fd_sc_hd__mux4_2
Xdata_outbuf_0._0_ data_inbuf_0.X VGND VGND VPWR VPWR data_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2 net45 net38 net29 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
+ Inst_RAM_IO_ConfigMem.ConfigBits\[228\] Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit0 net49 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_24._0_ net65 VGND VGND VPWR VPWR data_inbuf_24.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_3._0_ net94 VGND VGND VPWR VPWR strobe_inbuf_3.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_15._0_ net55 VGND VGND VPWR VPWR data_inbuf_15.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_040_ strobe_outbuf_8.X VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_169_ Inst_RAM_IO_switch_matrix.WW4BEG13 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS4_BEG3
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[184\] Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG12 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit6 net77 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
X_023_ data_outbuf_23.X VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_outbuf_18._0_ strobe_inbuf_18.X VGND VGND VPWR VPWR strobe_outbuf_18.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ net145 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput169 S2MID[4] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
Xinput158 S2END[1] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
Xinput125 N4END[13] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
Xinput136 N4END[9] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
Xinput147 RAM2FAB_D2_I2 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
Xinput103 N1END[2] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xinput114 N2MID[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_2
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_006_ data_outbuf_6.X VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit9 net80 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9 net102 net128 net154 net180
+ Inst_RAM_IO_ConfigMem.ConfigBits\[290\] Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG9 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[113\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xstrobe_outbuf_0._0_ strobe_inbuf_0.X VGND VGND VPWR VPWR strobe_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_15._0_ net87 VGND VGND VPWR VPWR strobe_inbuf_15.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput259 net259 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput237 net237 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput226 net226 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput248 net248 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput204 net204 VGND VGND VPWR VPWR FAB2RAM_C_O3 sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR FAB2RAM_D2_O2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1 net19 net11 net32 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_ConfigMem.ConfigBits\[94\] Inst_RAM_IO_ConfigMem.ConfigBits\[95\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix._47_ net172 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb7
+ sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3 net46 net39 net30 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
+ Inst_RAM_IO_ConfigMem.ConfigBits\[230\] Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame2_bit1 net60 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[83\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XN4END_inbuf_0._0_ net131 VGND VGND VPWR VPWR N4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406/HI
+ net406 sky130_fd_sc_hd__conb_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10 net103 net129 net155 net181
+ Inst_RAM_IO_ConfigMem.ConfigBits\[292\] Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG10 sky130_fd_sc_hd__mux4_2
Xdata_inbuf_7._0_ net78 VGND VGND VPWR VPWR data_inbuf_7.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_168_ Inst_RAM_IO_switch_matrix.WW4BEG12 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
X_099_ Inst_RAM_IO_switch_matrix.S2BEG7 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS4_BEG2
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[186\] Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG13 sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit7 net78 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
X_022_ data_outbuf_22.X VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput126 N4END[14] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xinput115 N2MID[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_1
Xinput104 N1END[3] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
Xinput159 S2END[2] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
Xinput148 RAM2FAB_D2_I3 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
Xinput137 RAM2FAB_D0_I0 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ data_outbuf_5.X VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XN4BEG_outbuf_5._0_ N4BEG_outbuf_5.A VGND VGND VPWR VPWR N4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\] sky130_fd_sc_hd__o21ai_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput205 net205 VGND VGND VPWR VPWR FAB2RAM_D0_O0 sky130_fd_sc_hd__clkbuf_4
Xoutput216 net216 VGND VGND VPWR VPWR FAB2RAM_D2_O3 sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput227 net227 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
Xoutput249 net249 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2 net18 net10 net22 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_ConfigMem.ConfigBits\[96\] Inst_RAM_IO_ConfigMem.ConfigBits\[97\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG2 sky130_fd_sc_hd__mux4_2
Xdata_outbuf_25._0_ data_inbuf_25.X VGND VGND VPWR VPWR data_outbuf_25.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix._46_ net171 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb6
+ sky130_fd_sc_hd__buf_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_16._0_ data_inbuf_16.X VGND VGND VPWR VPWR data_outbuf_16.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit2 net71 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_5._0_ S4BEG_outbuf_5.A VGND VGND VPWR VPWR S4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_35_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D1_InPass4_frame_config_mux._3_ UserCLK net144 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4END_inbuf_3._0_ net186 VGND VGND VPWR VPWR S4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11 net104 net130 net156 net182
+ Inst_RAM_IO_ConfigMem.ConfigBits\[294\] Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG11 sky130_fd_sc_hd__mux4_2
X_098_ Inst_RAM_IO_switch_matrix.S2BEG6 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
X_167_ Inst_RAM_IO_switch_matrix.WW4BEG11 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS4_BEG1
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[188\] Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG14 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame9_bit8 net79 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_021_ data_outbuf_21.X VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput149 RAM2FAB_D3_I0 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xinput116 N2MID[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 N2END[0] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput127 N4END[15] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput138 RAM2FAB_D0_I1 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_004_ data_outbuf_4.X VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0 net101 net153 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[121\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit0 net49 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XN4END_inbuf_11._0_ net127 VGND VGND VPWR VPWR N4BEG_outbuf_11.A sky130_fd_sc_hd__buf_2
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ net140 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_3._0_ data_inbuf_3.X VGND VGND VPWR VPWR data_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
Xoutput239 net239 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput228 net228 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput206 net206 VGND VGND VPWR VPWR FAB2RAM_D0_O1 sky130_fd_sc_hd__clkbuf_4
Xoutput217 net217 VGND VGND VPWR VPWR FAB2RAM_D3_O0 sky130_fd_sc_hd__clkbuf_4
Xdata_inbuf_27._0_ net68 VGND VGND VPWR VPWR data_inbuf_27.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3 net17 net9 net23 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_ConfigMem.ConfigBits\[98\] Inst_RAM_IO_ConfigMem.ConfigBits\[99\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG3 sky130_fd_sc_hd__mux4_2
Xdata_inbuf_18._0_ net58 VGND VGND VPWR VPWR data_inbuf_18.X sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_6._0_ net97 VGND VGND VPWR VPWR strobe_inbuf_6.X sky130_fd_sc_hd__buf_1
XInst_RAM_IO_switch_matrix._45_ net170 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb5
+ sky130_fd_sc_hd__clkbuf_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame2_bit3 net74 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0 net3 net38
+ net29 Inst_RAM_IO_switch_matrix.J_NS4_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[115\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux._2_ UserCLK net143 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404/HI net404 sky130_fd_sc_hd__conb_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12 net101 net121 net153 net173
+ Inst_RAM_IO_ConfigMem.ConfigBits\[296\] Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG12 sky130_fd_sc_hd__mux4_2
X_097_ Inst_RAM_IO_switch_matrix.S2BEG5 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
X_166_ Inst_RAM_IO_switch_matrix.WW4BEG10 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS4_BEG0
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\] Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG15 sky130_fd_sc_hd__mux4_1
XFILLER_0_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_11._0_ net179 VGND VGND VPWR VPWR S4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit9 net80 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_020_ data_outbuf_20.X VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_149_ Inst_RAM_IO_switch_matrix.W6BEG5 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput117 N2MID[4] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput128 N4END[1] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
Xinput106 N2END[1] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xinput139 RAM2FAB_D0_I2 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_003_ data_outbuf_3.X VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_3._0_ strobe_inbuf_3.X VGND VGND VPWR VPWR strobe_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1 net102 net154 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[123\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_18._0_ net90 VGND VGND VPWR VPWR strobe_inbuf_18.X sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit1 net60 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
Xoutput229 net229 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput207 net207 VGND VGND VPWR VPWR FAB2RAM_D0_O2 sky130_fd_sc_hd__buf_2
Xoutput218 net218 VGND VGND VPWR VPWR FAB2RAM_D3_O1 sky130_fd_sc_hd__buf_2
XN4END_inbuf_3._0_ net134 VGND VGND VPWR VPWR N4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4 net1 net16 net8 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
+ Inst_RAM_IO_ConfigMem.ConfigBits\[100\] Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG4 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix._44_ net169 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb4
+ sky130_fd_sc_hd__clkbuf_2
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit4 net75 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG10 Inst_RAM_IO_switch_matrix.J_NS4_BEG14 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
+ Inst_RAM_IO_ConfigMem.ConfigBits\[114\] Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM2FAB_D1_InPass4_frame_config_mux._1_ UserCLK net142 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13 net102 net128 net154 net180
+ Inst_RAM_IO_ConfigMem.ConfigBits\[298\] Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG13 sky130_fd_sc_hd__mux4_2
XFILLER_0_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_165_ Inst_RAM_IO_switch_matrix.WW4BEG9 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
X_096_ Inst_RAM_IO_switch_matrix.S2BEG4 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput390 net390 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_148_ Inst_RAM_IO_switch_matrix.W6BEG4 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_1
X_079_ N4BEG_outbuf_7.X VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_8._0_ N4BEG_outbuf_8.A VGND VGND VPWR VPWR N4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput107 N2END[2] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xinput118 N2MID[5] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_1
Xinput129 N4END[2] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
XS4BEG_outbuf_11._0_ S4BEG_outbuf_11.A VGND VGND VPWR VPWR S4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_002_ data_outbuf_2.X VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ net148 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2 net103 net155 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[125\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit2 net71 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__o21ai_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402/HI net402 sky130_fd_sc_hd__conb_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S4BEG0 sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_28._0_ data_inbuf_28.X VGND VGND VPWR VPWR data_outbuf_28.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_D0_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_19._0_ data_inbuf_19.X VGND VGND VPWR VPWR data_outbuf_19.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 net208 VGND VGND VPWR VPWR FAB2RAM_D0_O3 sky130_fd_sc_hd__clkbuf_4
Xoutput219 net219 VGND VGND VPWR VPWR FAB2RAM_D3_O2 sky130_fd_sc_hd__clkbuf_4
XS4BEG_outbuf_8._0_ S4BEG_outbuf_8.A VGND VGND VPWR VPWR S4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__o21ai_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5 net2 net15 net7 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
+ Inst_RAM_IO_ConfigMem.ConfigBits\[102\] Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG5 sky130_fd_sc_hd__mux4_2
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix._43_ net168 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb3
+ sky130_fd_sc_hd__clkbuf_2
XS4END_inbuf_6._0_ net174 VGND VGND VPWR VPWR S4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit5 net76 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux._0_ UserCLK net141 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N4BEG2 sky130_fd_sc_hd__o21ai_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14 net103 net129 net155 net181
+ Inst_RAM_IO_ConfigMem.ConfigBits\[300\] Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG14 sky130_fd_sc_hd__mux4_2
X_095_ Inst_RAM_IO_switch_matrix.S2BEG3 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
X_164_ Inst_RAM_IO_switch_matrix.WW4BEG8 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_1
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput380 net380 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput391 net391 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_078_ N4BEG_outbuf_6.X VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame8_bit0 net49 net99 VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
X_147_ Inst_RAM_IO_switch_matrix.W6BEG3 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_1
XFILLER_0_73_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 N2END[3] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
Xinput119 N2MID[6] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_001_ data_outbuf_1.X VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3 net104 net156 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[127\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 FrameStrobe[18] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_11._0_ strobe_inbuf_11.X VGND VGND VPWR VPWR strobe_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_6._0_ data_inbuf_6.X VGND VGND VPWR VPWR data_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit3 net74 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[110\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xstrobe_inbuf_9._0_ net100 VGND VGND VPWR VPWR strobe_inbuf_9.X sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput209 net209 VGND VGND VPWR VPWR FAB2RAM_D1_O0 sky130_fd_sc_hd__buf_2
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6 net3 net14 net6 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
+ Inst_RAM_IO_ConfigMem.ConfigBits\[104\] Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG6 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_switch_matrix._42_ net167 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame2_bit6 net77 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[80\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15 net104 net130 net156 net182
+ Inst_RAM_IO_ConfigMem.ConfigBits\[302\] Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG15 sky130_fd_sc_hd__mux4_2
X_094_ Inst_RAM_IO_switch_matrix.S2BEG2 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_163_ Inst_RAM_IO_switch_matrix.WW4BEG7 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput392 net392 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput381 net381 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput370 net370 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__clkbuf_4
X_077_ N4BEG_outbuf_5.X VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit1 net60 net99 VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
X_146_ Inst_RAM_IO_switch_matrix.W6BEG2 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_6._0_ strobe_inbuf_6.X VGND VGND VPWR VPWR strobe_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput109 N2END[4] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_000_ data_outbuf_0.X VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_0._0_ net49 VGND VGND VPWR VPWR data_inbuf_0.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_129_ Inst_RAM_IO_switch_matrix.W2BEG1 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 FrameData[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xinput91 FrameStrobe[19] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit4 net75 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4END_inbuf_6._0_ net122 VGND VGND VPWR VPWR N4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ net142 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7 net4 net13 net5 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
+ Inst_RAM_IO_ConfigMem.ConfigBits\[106\] Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEG7 sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix._41_ net166 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb1
+ sky130_fd_sc_hd__clkbuf_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame2_bit7 net78 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_51_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_162_ Inst_RAM_IO_switch_matrix.WW4BEG6 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
X_093_ Inst_RAM_IO_switch_matrix.S2BEG1 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput1 E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput360 net360 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput393 net393 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput371 net371 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput382 net382 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
X_145_ Inst_RAM_IO_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit2 net71 net99 VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
X_076_ N4BEG_outbuf_4.X VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput190 net190 VGND VGND VPWR VPWR Config_accessC_bit1 sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ Inst_RAM_IO_switch_matrix.W2BEG0 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_1
X_059_ Inst_RAM_IO_switch_matrix.N2BEG3 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0 net1 net33
+ net31 Inst_RAM_IO_switch_matrix.J_NS4_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[73\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput70 FrameData[29] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_4
Xinput92 FrameStrobe[1] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_8
Xinput81 FrameStrobe[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_8
XFILLER_0_66_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame5_bit5 net76 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_11._0_ N4BEG_outbuf_11.A VGND VGND VPWR VPWR N4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XS4END_inbuf_9._0_ net177 VGND VGND VPWR VPWR S4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix._40_ net165 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S2BEGb0
+ sky130_fd_sc_hd__clkbuf_2
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit8 net79 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_161_ Inst_RAM_IO_switch_matrix.WW4BEG5 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
X_092_ Inst_RAM_IO_switch_matrix.S2BEG0 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_20._0_ net61 VGND VGND VPWR VPWR data_inbuf_20.X sky130_fd_sc_hd__clkbuf_1
Xinput2 E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_11._0_ net51 VGND VGND VPWR VPWR data_inbuf_11.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput350 net350 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput361 net361 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput383 net383 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput372 net372 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__clkbuf_4
X_075_ N4BEG_outbuf_3.X VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit3 net74 net99 VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
X_144_ Inst_RAM_IO_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_1
XFILLER_0_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput191 net191 VGND VGND VPWR VPWR Config_accessC_bit2 sky130_fd_sc_hd__buf_2
Xstrobe_outbuf_14._0_ strobe_inbuf_14.X VGND VGND VPWR VPWR strobe_outbuf_14.X sky130_fd_sc_hd__clkbuf_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ Inst_RAM_IO_switch_matrix.N2BEG2 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_9._0_ data_inbuf_9.X VGND VGND VPWR VPWR data_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
X_127_ Inst_RAM_IO_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG8 Inst_RAM_IO_switch_matrix.J_NS4_BEG12 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_ConfigMem.ConfigBits\[72\] Inst_RAM_IO_ConfigMem.ConfigBits\[73\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput71 FrameData[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xinput60 FrameData[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
Xinput82 FrameStrobe[10] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput93 FrameStrobe[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_16
XInst_RAM_IO_ConfigMem.Inst_frame5_bit6 net77 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ net150 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit9 net80 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_11._0_ net83 VGND VGND VPWR VPWR strobe_inbuf_11.X sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395/HI net395 sky130_fd_sc_hd__conb_1
XFILLER_0_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_091_ Inst_RAM_IO_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
X_160_ Inst_RAM_IO_switch_matrix.WW4BEG4 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_9._0_ strobe_inbuf_9.X VGND VGND VPWR VPWR strobe_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
Xinput3 E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput351 net351 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput362 net362 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput340 net340 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput384 net384 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput373 net373 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__clkbuf_4
X_074_ N4BEG_outbuf_2.X VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_3._0_ net74 VGND VGND VPWR VPWR data_inbuf_3.X sky130_fd_sc_hd__clkbuf_1
X_143_ Inst_RAM_IO_switch_matrix.W2BEGb7 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit4 net75 net99 VGND VGND VPWR VPWR Inst_Config_accessConfig_access.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0 net4 net39
+ net30 Inst_RAM_IO_switch_matrix.J_NS4_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[118\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinst_clk_buf UserCLK VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_16
Xoutput192 net192 VGND VGND VPWR VPWR Config_accessC_bit3 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_057_ Inst_RAM_IO_switch_matrix.N2BEG1 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
X_126_ Inst_RAM_IO_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__o21ai_1
Xinput72 FrameData[30] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
Xinput61 FrameData[20] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_4
Xinput50 FrameData[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XN4END_inbuf_9._0_ net125 VGND VGND VPWR VPWR N4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput83 FrameStrobe[11] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 FrameStrobe[3] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D2_InPass4_frame_config_mux._3_ UserCLK net148 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit7 net78 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XN4BEG_outbuf_1._0_ N4BEG_outbuf_1.A VGND VGND VPWR VPWR N4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_C_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ S4BEG_outbuf_1.X VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_30._0_ data_inbuf_30.X VGND VGND VPWR VPWR data_outbuf_30.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_21._0_ data_inbuf_21.X VGND VGND VPWR VPWR data_outbuf_21.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ Inst_RAM_IO_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_12._0_ data_inbuf_12.X VGND VGND VPWR VPWR data_outbuf_12.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_1._0_ S4BEG_outbuf_1.A VGND VGND VPWR VPWR S4BEG_outbuf_1.X sky130_fd_sc_hd__buf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0 net33 net47 net31 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
+ Inst_RAM_IO_ConfigMem.ConfigBits\[232\] Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N4BEG1 sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_0_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__o21ai_2
Xoutput352 net352 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput330 net330 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput341 net341 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput363 net363 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput374 net374 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__clkbuf_4
X_142_ Inst_RAM_IO_switch_matrix.W2BEGb6 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
X_073_ N4BEG_outbuf_1.X VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit5 net76 net99 VGND VGND VPWR VPWR Inst_Config_accessConfig_access.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG11 Inst_RAM_IO_switch_matrix.J_NS4_BEG15 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
+ Inst_RAM_IO_ConfigMem.ConfigBits\[117\] Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_20 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_31 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput193 net193 VGND VGND VPWR VPWR FAB2RAM_A0_O0 sky130_fd_sc_hd__buf_2
XFILLER_0_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__o21ai_1
X_125_ Inst_RAM_IO_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_1
X_056_ Inst_RAM_IO_switch_matrix.N2BEG0 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
Xinput73 FrameData[31] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
Xinput62 FrameData[21] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_4
Xinput51 FrameData[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__o21ai_1
Xinput40 EE4END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
Xinput84 FrameStrobe[12] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 FrameStrobe[4] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_8
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux._2_ UserCLK net147 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit8 net79 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
X_108_ S4BEG_outbuf_0.X VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_039_ strobe_outbuf_7.X VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS4_BEG15
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[160\] Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0 net1 net31 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\] Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S1BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_35_185 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_23._0_ net64 VGND VGND VPWR VPWR data_inbuf_23.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame1_bit0 net49 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_2._0_ net93 VGND VGND VPWR VPWR strobe_inbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_14._0_ net54 VGND VGND VPWR VPWR data_inbuf_14.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1 net40 net48 net32 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
+ Inst_RAM_IO_ConfigMem.ConfigBits\[234\] Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[77\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
Xoutput364 net364 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput331 net331 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput320 net320 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput342 net342 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput353 net353 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput386 net386 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput375 net375 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_141_ Inst_RAM_IO_switch_matrix.W2BEGb5 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
X_072_ N4BEG_outbuf_0.X VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit6 net77 net99 VGND VGND VPWR VPWR Inst_Config_accessConfig_access.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_17._0_ strobe_inbuf_17.X VGND VGND VPWR VPWR strobe_outbuf_17.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_21 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_10 Inst_RAM_IO_switch_matrix.S2BEGb6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput194 net194 VGND VGND VPWR VPWR FAB2RAM_A0_O1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
X_055_ Inst_RAM_IO_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
X_124_ Inst_RAM_IO_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_75_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 FrameData[22] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_4
Xinput52 FrameData[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
Xinput74 FrameData[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
Xinput30 E6END[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
Xinput41 EE4END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput85 FrameStrobe[13] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput96 FrameStrobe[5] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_8
XFILLER_0_59_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux._1_ UserCLK net146 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit9 net80 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_C_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
X_038_ strobe_outbuf_6.X VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit30 net72 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
X_107_ Inst_RAM_IO_switch_matrix.S2BEGb7 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS4_BEG14
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[162\] Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_14._0_ net86 VGND VGND VPWR VPWR strobe_inbuf_14.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1 net2 net32 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[86\] Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S1BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame1_bit1 net60 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_6._0_ net77 VGND VGND VPWR VPWR data_inbuf_6.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2 net41 net34 net22 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
+ Inst_RAM_IO_ConfigMem.ConfigBits\[236\] Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
Xinput6 E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput321 net321 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput310 net310 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput343 net343 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
Xoutput365 net365 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput354 net354 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput387 net387 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput376 net376 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__clkbuf_4
X_071_ Inst_RAM_IO_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_1
X_140_ Inst_RAM_IO_switch_matrix.W2BEGb4 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit7 net78 net99 VGND VGND VPWR VPWR Inst_Config_accessConfig_access.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 N4BEG_outbuf_1.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput195 net195 VGND VGND VPWR VPWR FAB2RAM_A0_O2 sky130_fd_sc_hd__buf_2
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
X_054_ Inst_RAM_IO_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
X_123_ Inst_RAM_IO_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394/HI
+ net394 sky130_fd_sc_hd__conb_1
XFILLER_0_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XN4BEG_outbuf_4._0_ N4BEG_outbuf_4.A VGND VGND VPWR VPWR N4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
Xinput31 E6END[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
Xinput20 E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 FrameData[23] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
Xinput53 FrameData[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_4
Xinput75 FrameData[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
Xinput42 EE4END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 FrameStrobe[14] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 FrameStrobe[6] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_8
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM2FAB_D2_InPass4_frame_config_mux._0_ UserCLK net145 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\] sky130_fd_sc_hd__o21ai_4
XInst_RAM_IO_ConfigMem.Inst_frame9_bit31 net73 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit20 net61 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
X_037_ strobe_outbuf_5.X VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ Inst_RAM_IO_switch_matrix.S2BEGb6 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS4_BEG13
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[164\] Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_24._0_ data_inbuf_24.X VGND VGND VPWR VPWR data_outbuf_24.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2 net3 net22 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[88\] Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S1BEG2 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame8_bit30 net72 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_15._0_ data_inbuf_15.X VGND VGND VPWR VPWR data_outbuf_15.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_4._0_ S4BEG_outbuf_4.A VGND VGND VPWR VPWR S4BEG_outbuf_4.X sky130_fd_sc_hd__buf_2
XFILLER_0_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame1_bit2 net71 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403/HI net403 sky130_fd_sc_hd__conb_1
XFILLER_0_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XS4END_inbuf_2._0_ net185 VGND VGND VPWR VPWR S4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3 net42 net35 net23 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
+ Inst_RAM_IO_ConfigMem.ConfigBits\[238\] Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
Xoutput300 net300 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput344 net344 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput333 net333 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput311 net311 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput322 net322 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput355 net355 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput366 net366 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput377 net377 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput388 net388 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
X_070_ Inst_RAM_IO_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame8_bit8 net79 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ net139 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__o21ai_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 N4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 N4BEG_outbuf_3.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_34 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput196 net196 VGND VGND VPWR VPWR FAB2RAM_A0_O3 sky130_fd_sc_hd__buf_2
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_053_ Inst_RAM_IO_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
X_122_ Inst_RAM_IO_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput54 FrameData[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 E6END[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput21 E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput43 EE4END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput10 E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput65 FrameData[24] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
Xinput76 FrameData[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xinput87 FrameStrobe[15] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 FrameStrobe[7] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_8
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame9_bit21 net62 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit10 net50 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
X_105_ Inst_RAM_IO_switch_matrix.S2BEGb5 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_036_ strobe_outbuf_4.X VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XN4END_inbuf_10._0_ net126 VGND VGND VPWR VPWR N4BEG_outbuf_10.A sky130_fd_sc_hd__buf_2
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame4_bit0 net49 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS4_BEG12
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[166\] Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0 net113 net105 net165 net157
+ Inst_RAM_IO_ConfigMem.ConfigBits\[304\] Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG0 sky130_fd_sc_hd__mux4_2
Xdata_outbuf_2._0_ data_inbuf_2.X VGND VGND VPWR VPWR data_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_019_ data_outbuf_19.X VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_26._0_ net67 VGND VGND VPWR VPWR data_inbuf_26.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3 net4 net23 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
+ Inst_RAM_IO_switch_matrix.J_NS1_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[90\] Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S1BEG3 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame8_bit20 net61 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit31 net73 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_17._0_ net57 VGND VGND VPWR VPWR data_inbuf_17.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0 net2 net40
+ net32 Inst_RAM_IO_switch_matrix.J_NS4_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[76\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
Xstrobe_inbuf_5._0_ net96 VGND VGND VPWR VPWR strobe_inbuf_5.X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame1_bit3 net74 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XS4END_inbuf_10._0_ net178 VGND VGND VPWR VPWR S4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit30 net72 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput301 net301 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput345 net345 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput334 net334 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput323 net323 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput312 net312 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput356 net356 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput389 net389 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput378 net378 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput367 net367 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame8_bit9 net80 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_13 N4BEG_outbuf_11.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 N4BEG_outbuf_6.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_35 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput197 net197 VGND VGND VPWR VPWR FAB2RAM_A1_O0 sky130_fd_sc_hd__clkbuf_4
X_121_ Inst_RAM_IO_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_1
X_052_ Inst_RAM_IO_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_1
XFILLER_0_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_outbuf_2._0_ strobe_inbuf_2.X VGND VGND VPWR VPWR strobe_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xinput66 FrameData[25] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_4
Xinput55 FrameData[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_4
Xinput77 FrameData[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_4
Xinput22 E6END[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput44 EE4END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput88 FrameStrobe[16] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
Xinput11 E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
Xinput33 EE4END[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput99 FrameStrobe[8] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_8
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
X_035_ strobe_outbuf_3.X VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit11 net51 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_17._0_ net89 VGND VGND VPWR VPWR strobe_inbuf_17.X sky130_fd_sc_hd__clkbuf_2
X_104_ Inst_RAM_IO_switch_matrix.S2BEGb4 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit22 net63 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame4_bit1 net60 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401/HI net401 sky130_fd_sc_hd__conb_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS4_BEG11
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[168\] Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1 net114 net106 net166 net158
+ Inst_RAM_IO_ConfigMem.ConfigBits\[306\] Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_018_ data_outbuf_18.X VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XN4END_inbuf_2._0_ net133 VGND VGND VPWR VPWR N4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_2
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398/HI net398 sky130_fd_sc_hd__conb_1
XFILLER_0_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit10 net50 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit21 net62 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG9 Inst_RAM_IO_switch_matrix.J_NS4_BEG13 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_ConfigMem.ConfigBits\[75\] Inst_RAM_IO_ConfigMem.ConfigBits\[76\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
Xdata_inbuf_9._0_ net80 VGND VGND VPWR VPWR data_inbuf_9.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame1_bit4 net75 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ net147 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit31 net73 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit20 net61 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput302 net302 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput335 net335 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput346 net346 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput357 net357 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput324 net324 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput313 net313 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput379 net379 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput368 net368 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N4BEG0 sky130_fd_sc_hd__o21ai_2
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XN4BEG_outbuf_7._0_ N4BEG_outbuf_7.A VGND VGND VPWR VPWR N4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XANTENNA_14 N4BEG_outbuf_4.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput198 net198 VGND VGND VPWR VPWR FAB2RAM_A1_O1 sky130_fd_sc_hd__buf_2
XFILLER_0_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4BEG_outbuf_10._0_ S4BEG_outbuf_10.A VGND VGND VPWR VPWR S4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_2
X_051_ strobe_outbuf_19.X VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_1
X_120_ Inst_RAM_IO_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit30 net72 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput67 FrameData[26] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
Xinput56 FrameData[16] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_4
Xinput78 FrameData[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput23 E6END[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
Xinput34 EE4END[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 EE4END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
Xinput89 FrameStrobe[17] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
Xinput12 E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
X_034_ strobe_outbuf_2.X VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit23 net64 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
X_103_ Inst_RAM_IO_switch_matrix.S2BEGb3 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit12 net52 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__o21ai_2
XInst_RAM_IO_ConfigMem.Inst_frame4_bit2 net71 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS4_BEG10
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[170\] Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_0_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_27._0_ data_inbuf_27.X VGND VGND VPWR VPWR data_outbuf_27.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2 net115 net107 net167 net159
+ Inst_RAM_IO_ConfigMem.ConfigBits\[308\] Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_18._0_ data_inbuf_18.X VGND VGND VPWR VPWR data_outbuf_18.X sky130_fd_sc_hd__clkbuf_1
X_017_ data_outbuf_17.X VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XS4BEG_outbuf_7._0_ S4BEG_outbuf_7.A VGND VGND VPWR VPWR S4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_2
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame8_bit11 net51 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit22 net63 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XS4END_inbuf_5._0_ net188 VGND VGND VPWR VPWR S4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame1_bit5 net76 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput303 net303 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame7_bit10 net50 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput325 net325 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput314 net314 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame7_bit21 net62 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput347 net347 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput358 net358 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput336 net336 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput369 net369 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[74\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_26 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 RAM2FAB_D1_I0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 Inst_RAM_IO_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit0 net49 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput199 net199 VGND VGND VPWR VPWR FAB2RAM_A1_O2 sky130_fd_sc_hd__buf_2
X_050_ strobe_outbuf_18.X VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit31 net73 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit20 net61 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
Xinput68 FrameData[27] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput57 FrameData[17] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_4
Xinput79 FrameData[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
Xinput24 E6END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
Xinput35 EE4END[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
Xinput46 EE4END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
XFILLER_0_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit13 net53 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
X_033_ strobe_outbuf_1.X VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_10._0_ strobe_inbuf_10.X VGND VGND VPWR VPWR strobe_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
X_102_ Inst_RAM_IO_switch_matrix.S2BEGb2 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit24 net65 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_5._0_ data_inbuf_5.X VGND VGND VPWR VPWR data_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit3 net74 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_29._0_ net70 VGND VGND VPWR VPWR data_inbuf_29.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS4_BEG9
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG1 Inst_RAM_IO_ConfigMem.ConfigBits\[172\] Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG6 sky130_fd_sc_hd__mux4_1
XFILLER_0_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit30 net72 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_8._0_ net99 VGND VGND VPWR VPWR strobe_inbuf_8.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3 net116 net108 net168 net160
+ Inst_RAM_IO_ConfigMem.ConfigBits\[310\] Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG3 sky130_fd_sc_hd__mux4_2
X_016_ data_outbuf_16.X VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408/HI
+ net408 sky130_fd_sc_hd__conb_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame8_bit23 net64 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit12 net52 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame1_bit6 net77 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM2FAB_D3_InPass4_frame_config_mux._3_ UserCLK net152 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput304 net304 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame7_bit11 net51 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit22 net63 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput348 net348 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput326 net326 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput315 net315 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput337 net337 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput359 net359 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_5._0_ strobe_inbuf_5.X VGND VGND VPWR VPWR strobe_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 strobe_inbuf_12.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit1 net60 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput189 net189 VGND VGND VPWR VPWR Config_accessC_bit0 sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ net141 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame6_bit10 net50 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit21 net62 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 EE4END[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput25 E6END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 FrameData[28] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
Xinput58 FrameData[18] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
Xinput47 EE4END[8] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame9_bit25 net66 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit14 net54 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
X_101_ Inst_RAM_IO_switch_matrix.S2BEGb1 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
X_032_ strobe_outbuf_0.X VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XN4END_inbuf_5._0_ net136 VGND VGND VPWR VPWR N4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_ConfigMem.Inst_frame4_bit4 net75 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS4_BEG8
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\] Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG7 sky130_fd_sc_hd__mux4_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4 net117 net109 net169 net161
+ Inst_RAM_IO_ConfigMem.ConfigBits\[312\] Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG4 sky130_fd_sc_hd__mux4_2
XFILLER_0_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame5_bit20 net61 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit31 net73 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_015_ data_outbuf_15.X VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame8_bit24 net65 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit13 net53 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_ConfigMem.Inst_frame1_bit7 net78 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit30 net72 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux._2_ UserCLK net151 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit12 net52 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput305 net305 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit23 net64 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput349 net349 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput327 net327 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput338 net338 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_28 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit2 net71 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_17 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix._39_ net120 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit22 net63 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit11 net51 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput59 FrameData[19] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
Xinput26 E6END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 EE4END[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput48 EE4END[9] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput15 E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_031_ data_outbuf_31.X VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit15 net55 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
X_100_ Inst_RAM_IO_switch_matrix.S2BEGb0 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit26 net67 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame4_bit5 net76 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS4_BEG7
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[176\] Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG8 sky130_fd_sc_hd__mux4_1
XN4BEG_outbuf_10._0_ N4BEG_outbuf_10.A VGND VGND VPWR VPWR N4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit21 net62 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit10 net50 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5 net118 net110 net170 net162
+ Inst_RAM_IO_ConfigMem.ConfigBits\[314\] Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG5 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_014_ data_outbuf_14.X VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4END_inbuf_8._0_ net176 VGND VGND VPWR VPWR S4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 net13 net5 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ net395 Inst_RAM_IO_ConfigMem.ConfigBits\[248\] Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit25 net66 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit14 net54 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame1_bit8 net79 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame4_bit20 net61 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit31 net73 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM2FAB_D3_InPass4_frame_config_mux._1_ UserCLK net150 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit13 net53 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit24 net65 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput306 net306 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput339 net339 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput328 net328 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput317 net317 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_0_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0 net121 net173 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG15 Inst_RAM_IO_ConfigMem.ConfigBits\[192\] Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux4_1
Xdata_inbuf_10._0_ net50 VGND VGND VPWR VPWR data_inbuf_10.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ net149 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame3_bit30 net72 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_29 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit3 net74 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0 net20 net12 net30 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_ConfigMem.ConfigBits\[56\] Inst_RAM_IO_ConfigMem.ConfigBits\[57\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399/HI net399 sky130_fd_sc_hd__conb_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit12 net52 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit23 net64 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix._38_ net119 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_13._0_ strobe_inbuf_13.X VGND VGND VPWR VPWR strobe_outbuf_13.X sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_8._0_ data_inbuf_8.X VGND VGND VPWR VPWR data_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
Xinput49 FrameData[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
Xinput27 E6END[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput38 EE4END[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
Xinput16 E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_030_ data_outbuf_30.X VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit27 net68 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit16 net56 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_159_ Inst_RAM_IO_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit6 net77 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS4_BEG6
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[178\] Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.WW4BEG9 sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit11 net51 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6 net119 net111 net171 net163
+ Inst_RAM_IO_ConfigMem.ConfigBits\[316\] Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG6 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit22 net63 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
X_013_ data_outbuf_13.X VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1 net14 net6 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ net396 Inst_RAM_IO_ConfigMem.ConfigBits\[250\] Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame8_bit15 net55 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame8_bit26 net67 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_10._0_ net82 VGND VGND VPWR VPWR strobe_inbuf_10.X sky130_fd_sc_hd__clkbuf_2
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit9 net80 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit21 net62 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit10 net50 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM2FAB_D3_InPass4_frame_config_mux._0_ UserCLK net149 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput307 net307 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit14 net54 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit25 net66 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput318 net318 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xstrobe_outbuf_8._0_ strobe_inbuf_8.X VGND VGND VPWR VPWR strobe_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1 net128 net180 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG14 Inst_RAM_IO_ConfigMem.ConfigBits\[194\] Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_45_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame3_bit31 net73 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_2._0_ net71 VGND VGND VPWR VPWR data_inbuf_2.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit20 net61 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_19 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit4 net75 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0 net3 net41
+ net22 Inst_RAM_IO_switch_matrix.J_NS4_BEG2 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[79\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1 net19 net11 net29 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_ConfigMem.ConfigBits\[58\] Inst_RAM_IO_ConfigMem.ConfigBits\[59\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame6_bit13 net53 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit24 net65 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix._37_ net118 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb5
+ sky130_fd_sc_hd__clkbuf_2
Xinput39 EE4END[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
Xinput28 E6END[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
Xinput17 E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4END_inbuf_8._0_ net124 VGND VGND VPWR VPWR N4BEG_outbuf_8.A sky130_fd_sc_hd__buf_2
XFILLER_0_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame2_bit30 net72 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit17 net57 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit28 net69 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XN4BEG_outbuf_0._0_ N4BEG_outbuf_0.A VGND VGND VPWR VPWR N4BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
X_089_ Inst_RAM_IO_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_158_ Inst_RAM_IO_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit7 net78 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit12 net52 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit23 net64 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7 net120 net112 net172 net164
+ Inst_RAM_IO_ConfigMem.ConfigBits\[318\] Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS2_BEG7 sky130_fd_sc_hd__mux4_2
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
X_012_ data_outbuf_12.X VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2 net15 net7 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ net397 Inst_RAM_IO_ConfigMem.ConfigBits\[252\] Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame8_bit16 net56 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit27 net68 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit22 net63 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit11 net51 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_20._0_ data_inbuf_20.X VGND VGND VPWR VPWR data_outbuf_20.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_11._0_ data_inbuf_11.X VGND VGND VPWR VPWR data_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_0._0_ S4BEG_outbuf_0.A VGND VGND VPWR VPWR S4BEG_outbuf_0.X sky130_fd_sc_hd__buf_2
XFILLER_0_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput308 net308 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame7_bit15 net55 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit26 net67 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput319 net319 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__buf_2
XInst_Config_accessConfig_access._3_ Inst_Config_accessConfig_access.ConfigBits\[3\]
+ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2 net129 net181 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG13 Inst_RAM_IO_ConfigMem.ConfigBits\[196\] Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__o21ai_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit10 net50 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit21 net62 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit5 net76 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG10 Inst_RAM_IO_switch_matrix.J_NS4_BEG14 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_ConfigMem.ConfigBits\[78\] Inst_RAM_IO_ConfigMem.ConfigBits\[79\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2 net18 net10 net28 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_ConfigMem.ConfigBits\[60\] Inst_RAM_IO_ConfigMem.ConfigBits\[61\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_switch_matrix._36_ net117 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit14 net54 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit25 net66 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
Xinput29 E6END[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ net144 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit31 net73 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit29 net70 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit20 net61 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit18 net58 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[144\] Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb0 sky130_fd_sc_hd__mux4_1
XFILLER_0_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_157_ Inst_RAM_IO_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0 net33 net47 net21 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
+ Inst_RAM_IO_ConfigMem.ConfigBits\[216\] Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
X_088_ Inst_RAM_IO_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\] sky130_fd_sc_hd__o21ai_4
XInst_RAM_IO_ConfigMem.Inst_frame4_bit8 net79 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame5_bit13 net53 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit24 net65 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
X_011_ data_outbuf_11.X VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3 net16 net8 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ net398 Inst_RAM_IO_ConfigMem.ConfigBits\[254\] Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit30 net72 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit28 net69 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit17 net57 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409/HI net409 sky130_fd_sc_hd__conb_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_31._0_ net73 VGND VGND VPWR VPWR data_inbuf_31.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit12 net52 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit23 net64 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_22._0_ net63 VGND VGND VPWR VPWR data_inbuf_22.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_1._0_ net92 VGND VGND VPWR VPWR strobe_inbuf_1.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_13._0_ net53 VGND VGND VPWR VPWR data_inbuf_13.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame0_bit0 net49 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_Config_accessConfig_access._2_ Inst_Config_accessConfig_access.ConfigBits\[2\]
+ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit27 net68 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput309 net309 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame7_bit16 net56 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3 net130 net182 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG12 Inst_RAM_IO_ConfigMem.ConfigBits\[198\] Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG3 sky130_fd_sc_hd__mux4_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame3_bit22 net63 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit11 net51 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_16._0_ strobe_inbuf_16.X VGND VGND VPWR VPWR strobe_outbuf_16.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit6 net77 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0 net1 net43 net36 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
+ Inst_RAM_IO_ConfigMem.ConfigBits\[240\] Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3 net17 net9 net27 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_ConfigMem.ConfigBits\[62\] Inst_RAM_IO_ConfigMem.ConfigBits\[63\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix._35_ net116 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb3
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit15 net55 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit26 net67 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput19 E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit10 net50 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit21 net62 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame9_bit19 net59 net100 VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[146\] Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb1 sky130_fd_sc_hd__mux4_1
XFILLER_0_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1 net40 net48 net24 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
+ Inst_RAM_IO_ConfigMem.ConfigBits\[218\] Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_2
X_087_ Inst_RAM_IO_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_1
X_156_ Inst_RAM_IO_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit9 net80 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame5_bit14 net54 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit25 net66 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_010_ data_outbuf_10.X VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_13._0_ net85 VGND VGND VPWR VPWR strobe_inbuf_13.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_139_ Inst_RAM_IO_switch_matrix.W2BEGb3 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit29 net70 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit18 net58 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit31 net73 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit20 net61 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit13 net53 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame4_bit24 net65 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit1 net60 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit30 net72 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_5._0_ net76 VGND VGND VPWR VPWR data_inbuf_5.X sky130_fd_sc_hd__clkbuf_1
XInst_Config_accessConfig_access._1_ Inst_Config_accessConfig_access.ConfigBits\[1\]
+ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit17 net57 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit28 net69 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG7 Inst_RAM_IO_switch_matrix.J_NS4_BEG11 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_ConfigMem.ConfigBits\[200\] Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_0_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame10_bit30 net72 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame3_bit23 net64 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame3_bit12 net52 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1 net2 net44 net37 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
+ Inst_RAM_IO_ConfigMem.ConfigBits\[242\] Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\] sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit7 net78 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4 net16 net8 net26 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
+ Inst_RAM_IO_ConfigMem.ConfigBits\[64\] Inst_RAM_IO_ConfigMem.ConfigBits\[65\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG4 sky130_fd_sc_hd__mux4_1
XFILLER_0_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ net152 VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_switch_matrix._34_ net115 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb2
+ sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_ConfigMem.Inst_frame6_bit27 net68 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit16 net56 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XN4BEG_outbuf_3._0_ N4BEG_outbuf_3.A VGND VGND VPWR VPWR N4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame2_bit22 net63 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit11 net51 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\] sky130_fd_sc_hd__o21ai_4
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[148\] Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb2 sky130_fd_sc_hd__mux4_1
X_086_ Inst_RAM_IO_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2 net41 net34 net25 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
+ Inst_RAM_IO_ConfigMem.ConfigBits\[220\] Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
X_155_ Inst_RAM_IO_switch_matrix.W6BEG11 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit26 net67 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit15 net55 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 net290 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ Inst_RAM_IO_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit10 net50 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_138_ Inst_RAM_IO_switch_matrix.W2BEGb2 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit21 net62 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame8_bit19 net59 net99 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
+ Inst_RAM_IO_ConfigMem.Inst_frame8_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ net138 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_23._0_ data_inbuf_23.X VGND VGND VPWR VPWR data_outbuf_23.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_14._0_ data_inbuf_14.X VGND VGND VPWR VPWR data_outbuf_14.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_3._0_ S4BEG_outbuf_3.A VGND VGND VPWR VPWR S4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_ConfigMem.Inst_frame4_bit14 net54 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit25 net66 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XS4END_inbuf_1._0_ net184 VGND VGND VPWR VPWR S4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit2 net71 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit20 net61 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit18 net58 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit31 net73 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_Config_accessConfig_access._0_ Inst_Config_accessConfig_access.ConfigBits\[0\]
+ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit29 net70 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG6 Inst_RAM_IO_switch_matrix.J_NS4_BEG10 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_ConfigMem.ConfigBits\[202\] Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG5 sky130_fd_sc_hd__mux4_1
XFILLER_0_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame10_bit31 net73 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit13 net53 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit24 net65 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__o21ai_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2 net3 net45 net38 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
+ Inst_RAM_IO_ConfigMem.ConfigBits\[244\] Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\] sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame7_bit8 net79 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5 net15 net7 net25 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
+ Inst_RAM_IO_ConfigMem.ConfigBits\[66\] Inst_RAM_IO_ConfigMem.ConfigBits\[67\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG5 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix._33_ net114 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb1
+ sky130_fd_sc_hd__clkbuf_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit28 net69 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit17 net57 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
X_171_ Inst_RAM_IO_switch_matrix.WW4BEG15 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_1
XFILLER_0_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\] sky130_fd_sc_hd__o21ai_4
XFILLER_0_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit23 net64 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit12 net52 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\] VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\] sky130_fd_sc_hd__o21ai_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[150\] Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb3 sky130_fd_sc_hd__mux4_1
X_085_ Inst_RAM_IO_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3 net42 net35 net26 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
+ Inst_RAM_IO_ConfigMem.ConfigBits\[222\] Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
X_154_ Inst_RAM_IO_switch_matrix.W6BEG10 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame5_bit27 net68 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit16 net56 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400/HI net400 sky130_fd_sc_hd__conb_1
XFILLER_0_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_FAB2RAM_D3_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit0 net49 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput291 net291 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput280 net280 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xdata_outbuf_1._0_ data_inbuf_1.X VGND VGND VPWR VPWR data_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
X_137_ Inst_RAM_IO_switch_matrix.W2BEGb1 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
X_068_ Inst_RAM_IO_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit11 net51 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit22 net63 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0 net101 net21 net153 net406
+ Inst_RAM_IO_ConfigMem.ConfigBits\[320\] Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS1_BEG0 sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397/HI net397 sky130_fd_sc_hd__conb_1
Xdata_inbuf_25._0_ net66 VGND VGND VPWR VPWR data_inbuf_25.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_4._0_ net95 VGND VGND VPWR VPWR strobe_inbuf_4.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_16._0_ net56 VGND VGND VPWR VPWR data_inbuf_16.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame4_bit26 net67 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit15 net55 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame0_bit3 net74 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit21 net62 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit10 net50 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit19 net59 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_19._0_ strobe_inbuf_19.X VGND VGND VPWR VPWR strobe_outbuf_19.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG5 Inst_RAM_IO_switch_matrix.J_NS4_BEG9 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_ConfigMem.ConfigBits\[204\] Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG6 sky130_fd_sc_hd__mux4_1
XFILLER_0_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit14 net54 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit25 net66 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3 net4 net46 net39 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
+ Inst_RAM_IO_ConfigMem.ConfigBits\[246\] Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\] sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame7_bit9 net80 net98 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
+ Inst_RAM_IO_ConfigMem.Inst_frame7_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_ Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.S4BEG3 sky130_fd_sc_hd__o21ai_2
Xinput180 S4END[1] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6 net14 net6 net24 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
+ Inst_RAM_IO_ConfigMem.ConfigBits\[68\] Inst_RAM_IO_ConfigMem.ConfigBits\[69\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG6 sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix._32_ net113 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit29 net70 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit18 net58 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ Inst_RAM_IO_switch_matrix.WW4BEG14 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_1._0_ strobe_inbuf_1.X VGND VGND VPWR VPWR strobe_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\] sky130_fd_sc_hd__o21ai_2
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame2_bit13 net53 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit24 net65 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_ Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[152\] Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb4 sky130_fd_sc_hd__mux4_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_153_ Inst_RAM_IO_switch_matrix.W6BEG9 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
X_084_ Inst_RAM_IO_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_16._0_ net88 VGND VGND VPWR VPWR strobe_inbuf_16.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ net146 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame5_bit17 net57 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit28 net69 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
Xoutput270 net270 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit1 net60 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput292 net292 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput281 net281 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_136_ Inst_RAM_IO_switch_matrix.W2BEGb0 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
X_067_ Inst_RAM_IO_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1 net102 net24 net154 net407
+ Inst_RAM_IO_ConfigMem.ConfigBits\[322\] Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS1_BEG1 sky130_fd_sc_hd__mux4_2
XInst_RAM_IO_ConfigMem.Inst_frame1_bit23 net64 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit12 net52 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4END_inbuf_1._0_ net132 VGND VGND VPWR VPWR N4BEG_outbuf_1.A sky130_fd_sc_hd__buf_2
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0 net1 net36
+ net27 Inst_RAM_IO_switch_matrix.J_NS4_BEG0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[109\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit27 net68 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit16 net56 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_8._0_ net79 VGND VGND VPWR VPWR data_inbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_119_ S4BEG_outbuf_11.X VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG1 Inst_RAM_IO_switch_matrix.J_NS4_BEG5 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
+ Inst_RAM_IO_ConfigMem.ConfigBits\[212\] Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG10 sky130_fd_sc_hd__mux4_1
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame0_bit4 net75 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit22 net63 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit11 net51 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG4 Inst_RAM_IO_switch_matrix.J_NS4_BEG8 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_ConfigMem.ConfigBits\[206\] Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG7 sky130_fd_sc_hd__mux4_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame3_bit26 net67 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit15 net55 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[119\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput181 S4END[2] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_2
Xinput170 S2MID[5] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7 net13 net5 net21 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
+ Inst_RAM_IO_ConfigMem.ConfigBits\[70\] Inst_RAM_IO_ConfigMem.ConfigBits\[71\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.N2BEG7 sky130_fd_sc_hd__mux4_2
XN4BEG_outbuf_6._0_ N4BEG_outbuf_6.A VGND VGND VPWR VPWR N4BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit19 net59 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit14 net54 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit25 net66 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[154\] Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb5 sky130_fd_sc_hd__mux4_1
X_083_ N4BEG_outbuf_11.X VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
X_152_ Inst_RAM_IO_switch_matrix.W6BEG8 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_1
XFILLER_0_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit18 net58 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit29 net70 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux._1_ UserCLK Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\] sky130_fd_sc_hd__dfxtp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 net260 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput271 net271 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput282 net282 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput293 net293 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xdata_outbuf_26._0_ data_inbuf_26.X VGND VGND VPWR VPWR data_outbuf_26.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit2 net71 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0 net4 net42
+ net23 Inst_RAM_IO_switch_matrix.J_NS4_BEG3 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
+ Inst_RAM_IO_ConfigMem.ConfigBits\[82\] VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_066_ Inst_RAM_IO_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_1
X_135_ Inst_RAM_IO_switch_matrix.W2BEG7 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_1
XFILLER_0_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_17._0_ data_inbuf_17.X VGND VGND VPWR VPWR data_outbuf_17.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit24 net65 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit13 net53 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2 net103 net25 net155 net408
+ Inst_RAM_IO_ConfigMem.ConfigBits\[324\] Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS1_BEG2 sky130_fd_sc_hd__mux4_2
XS4BEG_outbuf_6._0_ S4BEG_outbuf_6.A VGND VGND VPWR VPWR S4BEG_outbuf_6.X sky130_fd_sc_hd__buf_2
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407 VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407/HI
+ net407 sky130_fd_sc_hd__conb_1
XFILLER_0_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4END_inbuf_4._0_ net187 VGND VGND VPWR VPWR S4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG8 Inst_RAM_IO_switch_matrix.J_NS4_BEG12 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
+ Inst_RAM_IO_ConfigMem.ConfigBits\[108\] Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit28 net69 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit17 net57 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_049_ strobe_outbuf_17.X VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
X_118_ S4BEG_outbuf_10.X VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
+ Inst_RAM_IO_ConfigMem.ConfigBits\[214\] Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG11 sky130_fd_sc_hd__mux4_1
XFILLER_0_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit5 net76 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit23 net64 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit12 net52 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_1 Inst_RAM_IO_switch_matrix.N2BEG7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG3 Inst_RAM_IO_switch_matrix.J_NS4_BEG7 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
+ Inst_RAM_IO_ConfigMem.ConfigBits\[208\] Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG8 sky130_fd_sc_hd__mux4_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame3_bit27 net68 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit16 net56 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
Xinput171 S2MID[6] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
Xinput182 S4END[3] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xinput160 S2END[3] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\] Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[128\] Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG0 sky130_fd_sc_hd__mux4_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit0 net49 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\] sky130_fd_sc_hd__o21ai_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0 net101 net121 net153 net173
+ Inst_RAM_IO_ConfigMem.ConfigBits\[272\] Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG0 sky130_fd_sc_hd__mux4_2
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_ Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame2_bit15 net55 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit26 net67 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\] VGND VGND VPWR VPWR Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[156\] Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb6 sky130_fd_sc_hd__mux4_1
XFILLER_0_64_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ N4BEG_outbuf_10.X VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
X_151_ Inst_RAM_IO_switch_matrix.W6BEG7 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_4._0_ data_inbuf_4.X VGND VGND VPWR VPWR data_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame5_bit19 net59 net96 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
+ Inst_RAM_IO_ConfigMem.Inst_frame5_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_28._0_ net69 VGND VGND VPWR VPWR data_inbuf_28.X sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux._0_ UserCLK Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput294 net294 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput261 net261 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput272 net272 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput283 net283 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput250 net250 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit3 net74 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_19._0_ net59 VGND VGND VPWR VPWR data_inbuf_19.X sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_7._0_ net98 VGND VGND VPWR VPWR strobe_inbuf_7.X sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG11 Inst_RAM_IO_switch_matrix.J_NS4_BEG15 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_ConfigMem.ConfigBits\[81\] Inst_RAM_IO_ConfigMem.ConfigBits\[82\] VGND
+ VGND VPWR VPWR Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_065_ Inst_RAM_IO_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit14 net54 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
X_134_ Inst_RAM_IO_switch_matrix.W2BEG6 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit25 net66 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3 net104 net26 net156 net394
+ Inst_RAM_IO_ConfigMem.ConfigBits\[326\] Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS1_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame4_bit18 net58 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit29 net70 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
X_117_ S4BEG_outbuf_9.X VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_048_ strobe_outbuf_16.X VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM_IO_ConfigMem.Inst_frame0_bit6 net77 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit13 net53 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit24 net65 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM_IO_switch_matrix.J_NS4_BEG2 Inst_RAM_IO_switch_matrix.J_NS4_BEG6 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
+ Inst_RAM_IO_ConfigMem.ConfigBits\[210\] Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W6BEG9 sky130_fd_sc_hd__mux4_1
XANTENNA_2 Inst_RAM_IO_switch_matrix.N4BEG0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame10_bit24 net65 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit28 net69 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit17 net57 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput183 S4END[4] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xinput172 S2MID[7] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
Xinput161 S2END[4] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput150 RAM2FAB_D3_I1 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_4._0_ strobe_inbuf_4.X VGND VGND VPWR VPWR strobe_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\] Inst_RAM_IO_switch_matrix.J_NS2_BEG1
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG6 Inst_RAM_IO_ConfigMem.ConfigBits\[130\] Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG1 sky130_fd_sc_hd__mux4_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame6_bit1 net60 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1 net102 net128 net154 net180
+ Inst_RAM_IO_ConfigMem.ConfigBits\[274\] Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG1 sky130_fd_sc_hd__mux4_2
Xstrobe_inbuf_19._0_ net91 VGND VGND VPWR VPWR strobe_inbuf_19.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_RAM_IO_ConfigMem.Inst_frame2_bit16 net56 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit27 net68 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS2_BEG0
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG7 Inst_RAM_IO_ConfigMem.ConfigBits\[158\] Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEGb7 sky130_fd_sc_hd__mux4_1
XFILLER_0_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_150_ Inst_RAM_IO_switch_matrix.W6BEG6 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_1
X_081_ N4BEG_outbuf_9.X VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XN4END_inbuf_4._0_ net135 VGND VGND VPWR VPWR N4BEG_outbuf_4.A sky130_fd_sc_hd__buf_2
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput295 net295 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput284 net284 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput273 net273 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput262 net262 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput240 net240 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput251 net251 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__buf_2
XInst_RAM_IO_ConfigMem.Inst_frame3_bit4 net75 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_133_ Inst_RAM_IO_switch_matrix.W2BEG5 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_064_ Inst_RAM_IO_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit26 net67 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit15 net55 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405 VGND VGND VPWR VPWR
+ Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405/HI net405 sky130_fd_sc_hd__conb_1
XInst_RAM_IO_ConfigMem.Inst_frame4_bit19 net59 net95 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
+ Inst_RAM_IO_ConfigMem.Inst_frame4_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
X_116_ S4BEG_outbuf_8.X VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_1
X_047_ strobe_outbuf_15.X VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit7 net78 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit14 net54 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit25 net66 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 Inst_RAM_IO_switch_matrix.S1BEG1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_9._0_ N4BEG_outbuf_9.A VGND VGND VPWR VPWR N4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_RAM_IO_ConfigMem.Inst_frame10_bit25 net66 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit18 net58 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame3_bit29 net70 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput162 S2END[5] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_1
Xinput151 RAM2FAB_D3_I2 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
Xinput140 RAM2FAB_D0_I3 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xinput184 S4END[5] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput173 S4END[0] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\] VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\] Inst_RAM_IO_switch_matrix.J_NS2_BEG2
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG5 Inst_RAM_IO_ConfigMem.ConfigBits\[132\] Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG2 sky130_fd_sc_hd__mux4_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux._3_ UserCLK Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_ConfigMem.Inst_frame6_bit2 net71 net97 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
+ Inst_RAM_IO_ConfigMem.Inst_frame6_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_ Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2 net103 net129 net155 net181
+ Inst_RAM_IO_ConfigMem.ConfigBits\[276\] Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.J_NS4_BEG2 sky130_fd_sc_hd__mux4_2
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_RAM_IO_ConfigMem.Inst_frame2_bit28 net69 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame2_bit17 net57 net93 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
+ Inst_RAM_IO_ConfigMem.Inst_frame2_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
+ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_ Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
+ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__o21ai_2
X_080_ N4BEG_outbuf_8.X VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_29._0_ data_inbuf_29.X VGND VGND VPWR VPWR data_outbuf_29.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XS4BEG_outbuf_9._0_ S4BEG_outbuf_9.A VGND VGND VPWR VPWR S4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput241 net241 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput230 net230 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput252 net252 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
XInst_RAM_IO_ConfigMem.Inst_frame3_bit5 net76 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput285 net285 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput263 net263 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput296 net296 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__clkbuf_4
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
+ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_063_ Inst_RAM_IO_switch_matrix.N2BEG7 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_132_ Inst_RAM_IO_switch_matrix.W2BEG4 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_1
XS4END_inbuf_7._0_ net175 VGND VGND VPWR VPWR S4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit27 net68 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame1_bit16 net56 net92 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
+ Inst_RAM_IO_ConfigMem.Inst_frame1_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_A1_OutPass4_frame_config_mux._2_ UserCLK Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
+ VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\] sky130_fd_sc_hd__dfxtp_1
XInst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_ Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
+ Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\] VGND VGND VPWR VPWR Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_046_ strobe_outbuf_14.X VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_1
X_115_ S4BEG_outbuf_7.X VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_RAM_IO_ConfigMem.Inst_frame0_bit8 net79 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit26 net67 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame0_bit15 net55 net81 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
+ Inst_RAM_IO_ConfigMem.Inst_frame0_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_RAM_IO_ConfigMem.Inst_frame9_bit0 net49 net100 VGND VGND VPWR VPWR Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
+ Inst_RAM_IO_ConfigMem.Inst_frame9_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_029_ data_outbuf_29.X VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 Inst_RAM_IO_switch_matrix.S1BEG3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM_IO_ConfigMem.Inst_frame10_bit26 net67 net82 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
+ Inst_RAM_IO_ConfigMem.Inst_frame10_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_ConfigMem.Inst_frame3_bit19 net59 net94 VGND VGND VPWR VPWR Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
+ Inst_RAM_IO_ConfigMem.Inst_frame3_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
+ Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\] VGND VGND VPWR VPWR Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput163 S2END[6] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xinput185 S4END[6] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput174 S4END[10] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xinput152 RAM2FAB_D3_I3 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
Xinput141 RAM2FAB_D1_I0 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_1
Xinput130 N4END[3] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
+ Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\] Inst_RAM_IO_switch_matrix.J_NS2_BEG3
+ Inst_RAM_IO_switch_matrix.J_NS2_BEG4 Inst_RAM_IO_ConfigMem.ConfigBits\[134\] Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
+ VGND VGND VPWR VPWR Inst_RAM_IO_switch_matrix.W2BEG3 sky130_fd_sc_hd__mux4_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_RAM2FAB_D0_InPass4_frame_config_mux._3_ UserCLK net140 VGND VGND VPWR VPWR Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
+ sky130_fd_sc_hd__dfxtp_1
.ends

